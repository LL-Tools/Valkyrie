

module b21_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10662;

  INV_X1 U4920 ( .A(n5863), .ZN(n6061) );
  XNOR2_X1 U4921 ( .A(n5770), .B(SI_12_), .ZN(n7706) );
  XNOR2_X1 U4922 ( .A(n5129), .B(n5561), .ZN(n5770) );
  INV_X4 U4923 ( .A(n8188), .ZN(n8197) );
  OR2_X2 U4924 ( .A1(n6411), .A2(n4976), .ZN(n7853) );
  INV_X1 U4925 ( .A(n8572), .ZN(n5956) );
  INV_X1 U4927 ( .A(n10662), .ZN(n4857) );
  BUF_X1 U4928 ( .A(n8719), .Z(n4860) );
  NAND2_X1 U4929 ( .A1(n9796), .A2(n8809), .ZN(n9776) );
  INV_X1 U4930 ( .A(n5991), .ZN(n8580) );
  INV_X2 U4931 ( .A(n8768), .ZN(n6870) );
  INV_X1 U4932 ( .A(n6724), .ZN(n6906) );
  INV_X1 U4933 ( .A(n5865), .ZN(n5757) );
  INV_X1 U4934 ( .A(n4865), .ZN(n8029) );
  INV_X4 U4936 ( .A(n4858), .ZN(n4862) );
  NOR2_X1 U4937 ( .A1(n9691), .A2(n9859), .ZN(n9669) );
  NAND2_X1 U4938 ( .A1(n8808), .A2(n8377), .ZN(n9812) );
  NAND2_X1 U4939 ( .A1(n5167), .A2(n5166), .ZN(n8932) );
  NAND2_X1 U4940 ( .A1(n6411), .A2(n8243), .ZN(n4858) );
  NAND2_X1 U4941 ( .A1(n9374), .A2(n5498), .ZN(n6030) );
  NOR3_X2 U4942 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n5483) );
  AOI21_X2 U4943 ( .B1(n9757), .B2(n8812), .A(n8811), .ZN(n9719) );
  CLKBUF_X2 U4944 ( .A(n6560), .Z(n4859) );
  NAND2_X2 U4945 ( .A1(n6723), .A2(n6722), .ZN(n10413) );
  INV_X2 U4946 ( .A(n6787), .ZN(n6746) );
  AOI21_X2 U4947 ( .B1(n9734), .B2(n8788), .A(n5322), .ZN(n9716) );
  NAND2_X2 U4948 ( .A1(n6411), .A2(n4976), .ZN(n6787) );
  XNOR2_X2 U4949 ( .A(n6404), .B(n9950), .ZN(n6411) );
  NOR2_X1 U4950 ( .A1(n8587), .A2(n8774), .ZN(n8719) );
  AOI21_X2 U4951 ( .B1(n9776), .B2(n9777), .A(n8810), .ZN(n9756) );
  NAND2_X1 U4952 ( .A1(n6098), .A2(n5582), .ZN(n6492) );
  XNOR2_X2 U4953 ( .A(n5512), .B(n5511), .ZN(n6098) );
  BUF_X4 U4954 ( .A(n6030), .Z(n4861) );
  OAI222_X1 U4955 ( .A1(n6411), .A2(P1_U3084), .B1(n8830), .B2(n9376), .C1(
        n8829), .C2(n9961), .ZN(P1_U3323) );
  XNOR2_X2 U4956 ( .A(n5139), .B(n6403), .ZN(n6386) );
  OAI21_X2 U4957 ( .B1(n6165), .B2(n5400), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5139) );
  XNOR2_X1 U4958 ( .A(n6004), .B(n6003), .ZN(n8876) );
  NAND2_X1 U4959 ( .A1(n5969), .A2(n5968), .ZN(n9305) );
  OR2_X1 U4960 ( .A1(n9892), .A2(n9790), .ZN(n9774) );
  NAND2_X1 U4961 ( .A1(n7770), .A2(n7769), .ZN(n9917) );
  NAND2_X1 U4962 ( .A1(n7377), .A2(n7281), .ZN(n7450) );
  NAND2_X1 U4963 ( .A1(n10391), .A2(n7102), .ZN(n8419) );
  INV_X1 U4964 ( .A(n8496), .ZN(n10405) );
  BUF_X2 U4966 ( .A(n8191), .Z(n8185) );
  INV_X1 U4967 ( .A(n10413), .ZN(n5013) );
  INV_X4 U4968 ( .A(n8199), .ZN(n8191) );
  BUF_X1 U4969 ( .A(n7101), .Z(n9544) );
  CLKBUF_X2 U4970 ( .A(n6724), .Z(n8184) );
  NAND4_X1 U4971 ( .A1(n6793), .A2(n6792), .A3(n6791), .A4(n6790), .ZN(n6954)
         );
  INV_X2 U4972 ( .A(n8719), .ZN(n8727) );
  CLKBUF_X2 U4973 ( .A(n6901), .Z(n4864) );
  NAND2_X1 U4974 ( .A1(n7049), .A2(n8253), .ZN(n6901) );
  INV_X4 U4975 ( .A(n6225), .ZN(n6197) );
  NAND2_X2 U4976 ( .A1(n6125), .A2(n9383), .ZN(n6225) );
  OR2_X1 U4977 ( .A1(n9840), .A2(n9684), .ZN(n5228) );
  AND2_X1 U4978 ( .A1(n5229), .A2(n5103), .ZN(n9840) );
  OAI21_X1 U4979 ( .B1(n4959), .B2(n9811), .A(n4957), .ZN(n9853) );
  AOI21_X1 U4980 ( .B1(n8362), .B2(n8476), .A(n8456), .ZN(n8365) );
  NOR2_X1 U4981 ( .A1(n9656), .A2(n4960), .ZN(n4959) );
  INV_X1 U4982 ( .A(n5116), .ZN(n9656) );
  OAI21_X2 U4983 ( .B1(n8876), .B2(n8874), .A(n4875), .ZN(n8865) );
  NAND2_X1 U4984 ( .A1(n8565), .A2(n8735), .ZN(n9055) );
  NAND2_X1 U4985 ( .A1(n5471), .A2(n9417), .ZN(n9474) );
  NAND2_X1 U4986 ( .A1(n9169), .A2(n9168), .ZN(n9167) );
  NAND2_X1 U4987 ( .A1(n8042), .A2(n8043), .ZN(n9493) );
  NAND2_X1 U4988 ( .A1(n5994), .A2(n5993), .ZN(n9298) );
  NAND2_X1 U4989 ( .A1(n4949), .A2(n6016), .ZN(n9294) );
  NAND2_X1 U4990 ( .A1(n8109), .A2(n8108), .ZN(n9869) );
  NAND3_X1 U4991 ( .A1(n5111), .A2(n5108), .A3(n9797), .ZN(n9796) );
  NAND2_X1 U4992 ( .A1(n8091), .A2(n8090), .ZN(n9874) );
  NAND2_X1 U4993 ( .A1(n5953), .A2(n5952), .ZN(n9311) );
  NAND2_X1 U4994 ( .A1(n5941), .A2(n5940), .ZN(n9316) );
  NAND2_X1 U4995 ( .A1(n8073), .A2(n8072), .ZN(n9881) );
  INV_X1 U4996 ( .A(n5142), .ZN(n4863) );
  AND2_X1 U4997 ( .A1(n5056), .A2(n5055), .ZN(n8014) );
  NAND2_X1 U4998 ( .A1(n5919), .A2(n5918), .ZN(n9321) );
  OAI21_X1 U4999 ( .B1(n7877), .B2(n4888), .A(n5057), .ZN(n5056) );
  OAI21_X1 U5000 ( .B1(n5069), .B2(n5068), .A(n4874), .ZN(n5799) );
  NAND2_X1 U5001 ( .A1(n5389), .A2(n5390), .ZN(n7877) );
  NAND2_X1 U5002 ( .A1(n8031), .A2(n8030), .ZN(n9895) );
  NAND2_X1 U5003 ( .A1(n8023), .A2(n8022), .ZN(n9901) );
  NAND2_X1 U5004 ( .A1(n5862), .A2(n5861), .ZN(n9337) );
  NOR2_X1 U5005 ( .A1(n7738), .A2(n7740), .ZN(n7555) );
  NOR2_X1 U5006 ( .A1(n7547), .A2(n7548), .ZN(n7738) );
  NAND2_X1 U5007 ( .A1(n4973), .A2(n4972), .ZN(n7646) );
  NAND2_X1 U5008 ( .A1(n5148), .A2(n5143), .ZN(n7813) );
  INV_X1 U5009 ( .A(n10591), .ZN(n4973) );
  NAND2_X1 U5010 ( .A1(n7529), .A2(n7528), .ZN(n9925) );
  AND2_X1 U5011 ( .A1(n8633), .A2(n10582), .ZN(n8751) );
  NAND2_X1 U5012 ( .A1(n5208), .A2(n4899), .ZN(n7201) );
  NAND2_X1 U5013 ( .A1(n5319), .A2(n7284), .ZN(n10534) );
  AND2_X2 U5014 ( .A1(n6579), .A2(n10628), .ZN(n8918) );
  NAND2_X1 U5015 ( .A1(n7401), .A2(n7400), .ZN(n10547) );
  AND2_X1 U5016 ( .A1(n7131), .A2(n7130), .ZN(n7392) );
  INV_X2 U5017 ( .A(n10605), .ZN(n10607) );
  NAND2_X2 U5018 ( .A1(n7390), .A2(n9819), .ZN(n9822) );
  XNOR2_X1 U5019 ( .A(n6802), .B(n8197), .ZN(n6890) );
  AND2_X1 U5020 ( .A1(n7053), .A2(n7052), .ZN(n10485) );
  INV_X1 U5021 ( .A(n7109), .ZN(n8490) );
  NAND2_X1 U5022 ( .A1(n8598), .A2(n8599), .ZN(n8741) );
  NOR2_X1 U5023 ( .A1(n10400), .A2(n10426), .ZN(n7223) );
  AND3_X1 U5024 ( .A1(n6799), .A2(n6798), .A3(n6797), .ZN(n10443) );
  NAND3_X1 U5025 ( .A1(n6647), .A2(n6646), .A3(n6645), .ZN(n6676) );
  NAND4_X1 U5026 ( .A1(n6433), .A2(n6432), .A3(n6431), .A4(n6430), .ZN(n7290)
         );
  AND3_X1 U5027 ( .A1(n6809), .A2(n6808), .A3(n6807), .ZN(n7225) );
  AND4_X1 U5028 ( .A1(n7152), .A2(n7151), .A3(n7150), .A4(n7149), .ZN(n7445)
         );
  AND2_X2 U5029 ( .A1(n6724), .A2(n6649), .ZN(n8155) );
  NAND2_X2 U5030 ( .A1(n6155), .A2(n6653), .ZN(n8199) );
  NAND4_X1 U5031 ( .A1(n6750), .A2(n6749), .A3(n6748), .A4(n6747), .ZN(n6813)
         );
  AND2_X1 U5032 ( .A1(n8934), .A2(n6568), .ZN(n6840) );
  CLKBUF_X1 U5033 ( .A(n6901), .Z(n4865) );
  BUF_X2 U5034 ( .A(n5651), .Z(n8581) );
  NAND2_X2 U5035 ( .A1(n6386), .A2(n6387), .ZN(n7049) );
  INV_X1 U5036 ( .A(n8243), .ZN(n4976) );
  INV_X1 U5037 ( .A(n9377), .ZN(n5498) );
  NAND2_X1 U5038 ( .A1(n5497), .A2(n9377), .ZN(n5865) );
  NAND2_X1 U5039 ( .A1(n5489), .A2(n4870), .ZN(n9377) );
  XNOR2_X1 U5040 ( .A(n6636), .B(n6635), .ZN(n9781) );
  NOR2_X1 U5041 ( .A1(n5009), .A2(n5223), .ZN(n6405) );
  OR2_X1 U5042 ( .A1(n5521), .A2(SI_1_), .ZN(n5522) );
  OAI21_X1 U5043 ( .B1(n5859), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5885) );
  NAND2_X1 U5044 ( .A1(n4870), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U5045 ( .A1(n5401), .A2(n6163), .ZN(n5400) );
  INV_X1 U5046 ( .A(n5402), .ZN(n5401) );
  NAND2_X1 U5047 ( .A1(n5482), .A2(n5503), .ZN(n5592) );
  NAND2_X1 U5048 ( .A1(n5463), .A2(n5403), .ZN(n5402) );
  NOR2_X1 U5049 ( .A1(n5399), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n5398) );
  INV_X1 U5050 ( .A(n6148), .ZN(n5403) );
  INV_X1 U5051 ( .A(n5455), .ZN(n5453) );
  AND2_X1 U5052 ( .A1(n5224), .A2(n5011), .ZN(n5010) );
  NAND2_X1 U5053 ( .A1(n6147), .A2(n6167), .ZN(n6148) );
  XNOR2_X1 U5054 ( .A(n5026), .B(P2_IR_REG_1__SCAN_IN), .ZN(n10316) );
  INV_X1 U5055 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6159) );
  INV_X1 U5056 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6339) );
  NOR2_X1 U5057 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n6139) );
  INV_X1 U5058 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6160) );
  INV_X1 U5059 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6158) );
  INV_X1 U5060 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5814) );
  NOR2_X1 U5061 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5478) );
  NOR2_X1 U5062 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5476) );
  NOR2_X1 U5063 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5603) );
  INV_X1 U5064 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6632) );
  INV_X1 U5065 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6141) );
  NOR2_X1 U5066 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5472) );
  NOR2_X1 U5067 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5473) );
  INV_X1 U5068 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5729) );
  INV_X1 U5069 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5733) );
  INV_X4 U5070 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  XNOR2_X2 U5071 ( .A(n5674), .B(n5467), .ZN(n6900) );
  OR2_X1 U5072 ( .A1(n9294), .A2(n8914), .ZN(n8707) );
  INV_X1 U5073 ( .A(n5388), .ZN(n5386) );
  INV_X1 U5074 ( .A(n6648), .ZN(n6667) );
  AND2_X1 U5075 ( .A1(n5583), .A2(n6877), .ZN(n5584) );
  INV_X1 U5076 ( .A(n8574), .ZN(n8567) );
  CLKBUF_X1 U5077 ( .A(n5757), .Z(n5738) );
  NAND2_X2 U5078 ( .A1(n9374), .A2(n9377), .ZN(n8574) );
  NAND3_X1 U5079 ( .A1(n8046), .A2(n9492), .A3(n5385), .ZN(n5030) );
  INV_X1 U5080 ( .A(n5962), .ZN(n5076) );
  NOR2_X1 U5081 ( .A1(n5435), .A2(n5082), .ZN(n5081) );
  NOR2_X1 U5082 ( .A1(n8902), .A2(n8900), .ZN(n5082) );
  NAND2_X1 U5083 ( .A1(n5436), .A2(n5437), .ZN(n5435) );
  NAND2_X1 U5084 ( .A1(n8731), .A2(n4911), .ZN(n5284) );
  INV_X1 U5085 ( .A(n8730), .ZN(n5283) );
  NAND2_X1 U5086 ( .A1(n5333), .A2(n9011), .ZN(n8760) );
  AND2_X1 U5087 ( .A1(n5334), .A2(n8723), .ZN(n8726) );
  OR2_X1 U5088 ( .A1(n8998), .A2(n8729), .ZN(n5334) );
  OR2_X1 U5089 ( .A1(n9278), .A2(n8923), .ZN(n8715) );
  OR2_X1 U5090 ( .A1(n9327), .A2(n8924), .ZN(n8668) );
  AOI21_X1 U5091 ( .B1(n4867), .B2(n7239), .A(n5266), .ZN(n5265) );
  NAND2_X1 U5092 ( .A1(n5297), .A2(n5506), .ZN(n5296) );
  INV_X1 U5093 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5506) );
  INV_X1 U5094 ( .A(n5505), .ZN(n5297) );
  AND2_X1 U5095 ( .A1(n7116), .A2(n6155), .ZN(n6724) );
  AOI21_X1 U5096 ( .B1(n8349), .B2(n8488), .A(n8351), .ZN(n4953) );
  OR2_X1 U5097 ( .A1(n9859), .A2(n9690), .ZN(n8816) );
  INV_X1 U5098 ( .A(n7753), .ZN(n5134) );
  OR2_X1 U5099 ( .A1(n7800), .A2(n7808), .ZN(n8392) );
  XNOR2_X1 U5100 ( .A(n7101), .B(n5013), .ZN(n8496) );
  NAND2_X1 U5101 ( .A1(n9843), .A2(n5107), .ZN(n5106) );
  OR2_X1 U5102 ( .A1(n9837), .A2(n8348), .ZN(n8488) );
  NAND2_X1 U5103 ( .A1(n8532), .A2(n10415), .ZN(n8351) );
  NAND2_X1 U5104 ( .A1(n8239), .A2(n8238), .ZN(n8245) );
  INV_X1 U5105 ( .A(SI_20_), .ZN(n10127) );
  INV_X1 U5106 ( .A(n5938), .ZN(n5936) );
  AND3_X1 U5107 ( .A1(n4980), .A2(n4979), .A3(n4978), .ZN(n6146) );
  INV_X1 U5108 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n4978) );
  NAND2_X1 U5109 ( .A1(n5571), .A2(n5570), .ZN(n5850) );
  NAND2_X1 U5110 ( .A1(n5813), .A2(n4935), .ZN(n5571) );
  INV_X1 U5111 ( .A(SI_16_), .ZN(n5572) );
  OR2_X1 U5112 ( .A1(n5920), .A2(n10187), .ZN(n5943) );
  AND2_X1 U5113 ( .A1(n4859), .A2(n8768), .ZN(n5405) );
  XNOR2_X1 U5114 ( .A(n5407), .B(n7009), .ZN(n5406) );
  AND2_X1 U5115 ( .A1(n6225), .A2(n6718), .ZN(n5651) );
  AND2_X1 U5116 ( .A1(n8998), .A2(n8729), .ZN(n8761) );
  AND2_X1 U5117 ( .A1(n6013), .A2(n6012), .ZN(n8914) );
  NAND2_X1 U5118 ( .A1(n9047), .A2(n9273), .ZN(n9038) );
  NAND2_X1 U5119 ( .A1(n5245), .A2(n5247), .ZN(n8565) );
  NOR2_X1 U5120 ( .A1(n5246), .A2(n8564), .ZN(n5245) );
  INV_X1 U5121 ( .A(n5248), .ZN(n5246) );
  OR2_X1 U5122 ( .A1(n9110), .A2(n9111), .ZN(n9108) );
  AND2_X1 U5123 ( .A1(n8697), .A2(n8692), .ZN(n9111) );
  NOR2_X1 U5124 ( .A1(n5458), .A2(n8756), .ZN(n5182) );
  NAND2_X1 U5125 ( .A1(n5162), .A2(n5161), .ZN(n9212) );
  INV_X1 U5126 ( .A(n9343), .ZN(n5161) );
  NAND2_X1 U5127 ( .A1(n5269), .A2(n5268), .ZN(n5267) );
  NAND2_X1 U5128 ( .A1(n10436), .A2(n7041), .ZN(n7040) );
  INV_X1 U5129 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5486) );
  INV_X1 U5130 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5503) );
  INV_X1 U5131 ( .A(n7116), .ZN(n6653) );
  NAND2_X1 U5132 ( .A1(n5030), .A2(n4900), .ZN(n5471) );
  INV_X1 U5133 ( .A(n9419), .ZN(n5031) );
  INV_X1 U5134 ( .A(n6411), .ZN(n4977) );
  AND2_X1 U5135 ( .A1(n8819), .A2(n8450), .ZN(n9624) );
  OAI21_X1 U5136 ( .B1(n9655), .B2(n8797), .A(n8798), .ZN(n9639) );
  OR2_X1 U5137 ( .A1(n7855), .A2(n7854), .ZN(n7907) );
  OAI21_X1 U5138 ( .B1(n7903), .B2(n7902), .A(n8394), .ZN(n7904) );
  INV_X1 U5139 ( .A(n6899), .ZN(n8355) );
  NAND2_X1 U5140 ( .A1(n7049), .A2(n6718), .ZN(n6899) );
  AND2_X1 U5141 ( .A1(n6376), .A2(n6378), .ZN(n6629) );
  INV_X1 U5142 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6137) );
  BUF_X1 U5143 ( .A(n5577), .Z(n8253) );
  XNOR2_X1 U5144 ( .A(n5406), .B(n5405), .ZN(n6696) );
  NAND2_X1 U5145 ( .A1(n6696), .A2(n6697), .ZN(n6695) );
  AOI21_X1 U5146 ( .B1(n9838), .B2(n9825), .A(n8825), .ZN(n5227) );
  OR2_X1 U5147 ( .A1(n8613), .A2(n5291), .ZN(n5290) );
  NAND2_X1 U5148 ( .A1(n5292), .A2(n4889), .ZN(n5291) );
  AOI21_X1 U5149 ( .B1(n8617), .B2(n8616), .A(n8747), .ZN(n5289) );
  AND2_X1 U5150 ( .A1(n8752), .A2(n5302), .ZN(n5301) );
  INV_X1 U5151 ( .A(n5303), .ZN(n5302) );
  OAI22_X1 U5152 ( .A1(n4869), .A2(n4860), .B1(n4866), .B2(n8727), .ZN(n5303)
         );
  NOR2_X1 U5153 ( .A1(n9137), .A2(n8680), .ZN(n5309) );
  OR2_X1 U5154 ( .A1(n8689), .A2(n8691), .ZN(n5307) );
  AOI21_X1 U5155 ( .B1(n5418), .B2(n5419), .A(n5417), .ZN(n5416) );
  INV_X1 U5156 ( .A(n8832), .ZN(n5417) );
  INV_X1 U5157 ( .A(n5421), .ZN(n5418) );
  INV_X1 U5158 ( .A(n8856), .ZN(n5436) );
  INV_X1 U5159 ( .A(n7533), .ZN(n7534) );
  INV_X1 U5160 ( .A(n9446), .ZN(n5381) );
  NAND2_X1 U5161 ( .A1(n4876), .A2(n9438), .ZN(n5378) );
  NOR2_X1 U5162 ( .A1(n8502), .A2(n5218), .ZN(n5217) );
  INV_X1 U5163 ( .A(n8387), .ZN(n5218) );
  AOI21_X1 U5164 ( .B1(n6021), .B2(n6025), .A(n5362), .ZN(n5361) );
  INV_X1 U5165 ( .A(n6039), .ZN(n5362) );
  INV_X1 U5166 ( .A(n6025), .ZN(n5359) );
  INV_X1 U5167 ( .A(SI_26_), .ZN(n10109) );
  AOI21_X1 U5168 ( .B1(n5345), .B2(n5346), .A(n5343), .ZN(n5342) );
  INV_X1 U5169 ( .A(n5590), .ZN(n5343) );
  INV_X1 U5170 ( .A(SI_8_), .ZN(n10093) );
  NOR2_X1 U5171 ( .A1(n5706), .A2(n5348), .ZN(n5347) );
  INV_X1 U5172 ( .A(n5548), .ZN(n5348) );
  INV_X1 U5173 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5048) );
  INV_X1 U5174 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5047) );
  OAI21_X1 U5175 ( .B1(n5083), .B2(n5076), .A(n4919), .ZN(n5073) );
  INV_X1 U5176 ( .A(n5414), .ZN(n5412) );
  AND2_X1 U5177 ( .A1(n5781), .A2(n5445), .ZN(n5444) );
  NAND2_X1 U5178 ( .A1(n7634), .A2(n5769), .ZN(n5445) );
  AND2_X1 U5179 ( .A1(n7792), .A2(n5780), .ZN(n5781) );
  NAND2_X1 U5180 ( .A1(n5081), .A2(n8902), .ZN(n5080) );
  NOR2_X1 U5181 ( .A1(n8699), .A2(n8708), .ZN(n8704) );
  AND2_X1 U5182 ( .A1(n8736), .A2(n8707), .ZN(n8709) );
  NAND2_X1 U5183 ( .A1(n8760), .A2(n5328), .ZN(n5327) );
  NOR2_X1 U5184 ( .A1(n9044), .A2(n5329), .ZN(n5328) );
  NAND2_X1 U5185 ( .A1(n5277), .A2(n5330), .ZN(n5329) );
  NOR2_X1 U5186 ( .A1(n9079), .A2(n5331), .ZN(n5330) );
  OR2_X1 U5187 ( .A1(n9289), .A2(n8867), .ZN(n8736) );
  INV_X1 U5188 ( .A(n9019), .ZN(n5181) );
  OAI21_X1 U5189 ( .B1(n4871), .B2(n5181), .A(n9137), .ZN(n5180) );
  OR2_X1 U5190 ( .A1(n9305), .A2(n8894), .ZN(n8693) );
  NOR2_X1 U5191 ( .A1(n9145), .A2(n9168), .ZN(n5241) );
  NOR2_X1 U5192 ( .A1(n9192), .A2(n5238), .ZN(n5237) );
  NOR2_X1 U5193 ( .A1(n8756), .A2(n5239), .ZN(n5238) );
  INV_X1 U5194 ( .A(n8662), .ZN(n5239) );
  OR2_X1 U5195 ( .A1(n8221), .A2(n7841), .ZN(n8650) );
  INV_X1 U5196 ( .A(n7333), .ZN(n5256) );
  INV_X1 U5197 ( .A(n10582), .ZN(n5255) );
  INV_X1 U5198 ( .A(n7468), .ZN(n5257) );
  AND2_X1 U5199 ( .A1(n8774), .A2(n8592), .ZN(n6129) );
  OR2_X1 U5200 ( .A1(n7225), .A2(n6906), .ZN(n6810) );
  OR2_X1 U5201 ( .A1(n7853), .A2(n10424), .ZN(n6639) );
  OR2_X1 U5202 ( .A1(n6787), .A2(n6638), .ZN(n6640) );
  NOR2_X1 U5203 ( .A1(n9837), .A2(n5153), .ZN(n5152) );
  INV_X1 U5204 ( .A(n5154), .ZN(n5153) );
  OR2_X1 U5205 ( .A1(n9848), .A2(n9659), .ZN(n8818) );
  NAND2_X1 U5206 ( .A1(n8781), .A2(n5118), .ZN(n5117) );
  INV_X1 U5207 ( .A(n7925), .ZN(n5118) );
  NAND2_X1 U5208 ( .A1(n8510), .A2(n5007), .ZN(n5006) );
  AND2_X1 U5209 ( .A1(n5120), .A2(n8781), .ZN(n5119) );
  INV_X1 U5210 ( .A(n7864), .ZN(n5007) );
  NAND2_X1 U5211 ( .A1(n8397), .A2(n8806), .ZN(n5233) );
  NOR2_X1 U5212 ( .A1(n7898), .A2(n5121), .ZN(n5120) );
  INV_X1 U5213 ( .A(n7892), .ZN(n5121) );
  OR2_X1 U5214 ( .A1(n7891), .A2(n9520), .ZN(n8394) );
  AND2_X1 U5215 ( .A1(n5315), .A2(n4997), .ZN(n4996) );
  NAND2_X1 U5216 ( .A1(n8505), .A2(n7612), .ZN(n4997) );
  NOR2_X1 U5217 ( .A1(n5316), .A2(n8506), .ZN(n5315) );
  INV_X1 U5218 ( .A(n7801), .ZN(n5316) );
  NAND2_X1 U5219 ( .A1(n5144), .A2(n7625), .ZN(n5146) );
  INV_X1 U5220 ( .A(n5149), .ZN(n5144) );
  INV_X1 U5221 ( .A(n7457), .ZN(n5148) );
  INV_X1 U5222 ( .A(n5217), .ZN(n5216) );
  NOR2_X1 U5223 ( .A1(n8284), .A2(n8276), .ZN(n7449) );
  NOR2_X1 U5224 ( .A1(n7118), .A2(n7206), .ZN(n5137) );
  INV_X1 U5225 ( .A(n8420), .ZN(n5211) );
  INV_X1 U5226 ( .A(n8415), .ZN(n5212) );
  OR2_X1 U5227 ( .A1(n6667), .A2(n8525), .ZN(n7116) );
  INV_X1 U5228 ( .A(n8531), .ZN(n6677) );
  AND2_X1 U5229 ( .A1(n8252), .A2(n8251), .ZN(n8353) );
  AND2_X1 U5230 ( .A1(n8246), .A2(n8242), .ZN(n8244) );
  NAND2_X1 U5231 ( .A1(n6015), .A2(n6014), .ZN(n6022) );
  INV_X1 U5232 ( .A(n5354), .ZN(n5353) );
  OAI21_X1 U5233 ( .B1(n5356), .B2(n5355), .A(n5930), .ZN(n5354) );
  INV_X1 U5234 ( .A(n5915), .ZN(n5355) );
  INV_X1 U5235 ( .A(SI_18_), .ZN(n10099) );
  OR2_X1 U5236 ( .A1(n7094), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n7095) );
  NAND2_X1 U5237 ( .A1(n5124), .A2(n5122), .ZN(n5786) );
  NAND2_X1 U5238 ( .A1(n5123), .A2(n4883), .ZN(n5122) );
  INV_X1 U5239 ( .A(SI_10_), .ZN(n9993) );
  INV_X1 U5240 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6136) );
  NAND3_X1 U5241 ( .A1(n5089), .A2(n5541), .A3(n5088), .ZN(n5602) );
  NAND2_X1 U5242 ( .A1(n5660), .A2(n5091), .ZN(n5089) );
  INV_X1 U5243 ( .A(n5092), .ZN(n5091) );
  OAI21_X1 U5244 ( .B1(n6718), .B2(n4964), .A(n4963), .ZN(n5533) );
  NAND2_X1 U5245 ( .A1(n6718), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4963) );
  OAI211_X1 U5246 ( .C1(n8865), .C2(n5413), .A(n5408), .B(n5058), .ZN(n6112)
         );
  NAND2_X1 U5247 ( .A1(n5414), .A2(n6063), .ZN(n5413) );
  OAI22_X1 U5248 ( .A1(n5412), .A2(n5411), .B1(n5414), .B2(n5423), .ZN(n5408)
         );
  NAND2_X1 U5249 ( .A1(n8865), .A2(n5410), .ZN(n5058) );
  NOR2_X1 U5250 ( .A1(n10511), .A2(n10512), .ZN(n10509) );
  NAND2_X1 U5251 ( .A1(n4922), .A2(n5441), .ZN(n5437) );
  INV_X1 U5252 ( .A(n5447), .ZN(n5442) );
  OR2_X1 U5253 ( .A1(n5834), .A2(n5833), .ZN(n5836) );
  AOI21_X1 U5254 ( .B1(n8840), .B2(n8839), .A(n5982), .ZN(n6004) );
  OR2_X1 U5255 ( .A1(n5995), .A2(n10081), .ZN(n6006) );
  INV_X1 U5256 ( .A(n7634), .ZN(n5446) );
  NAND2_X1 U5257 ( .A1(n5430), .A2(n5429), .ZN(n5428) );
  INV_X1 U5258 ( .A(n6710), .ZN(n5429) );
  INV_X1 U5259 ( .A(n6709), .ZN(n5430) );
  NAND2_X1 U5260 ( .A1(n8729), .A2(n8592), .ZN(n5263) );
  NAND2_X1 U5261 ( .A1(n8765), .A2(n8592), .ZN(n8586) );
  AND2_X1 U5262 ( .A1(n6050), .A2(n6049), .ZN(n8711) );
  AND3_X1 U5263 ( .A1(n5959), .A2(n5958), .A3(n5957), .ZN(n8859) );
  AND3_X1 U5264 ( .A1(n5947), .A2(n5946), .A3(n5945), .ZN(n8558) );
  AND3_X1 U5265 ( .A1(n5926), .A2(n5925), .A3(n5924), .ZN(n8858) );
  AND4_X1 U5266 ( .A1(n5874), .A2(n5873), .A3(n5872), .A4(n5871), .ZN(n8554)
         );
  NAND2_X1 U5267 ( .A1(n5956), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5613) );
  OR2_X1 U5268 ( .A1(n6237), .A2(n6236), .ZN(n5022) );
  AOI21_X1 U5269 ( .B1(n6401), .B2(P2_REG1_REG_10__SCAN_IN), .A(n6317), .ZN(
        n7165) );
  OR2_X1 U5270 ( .A1(n8955), .A2(n4947), .ZN(n5017) );
  NAND2_X1 U5271 ( .A1(n8583), .A2(n8582), .ZN(n8998) );
  NAND2_X1 U5272 ( .A1(n8551), .A2(n8550), .ZN(n9036) );
  OR2_X1 U5273 ( .A1(n5468), .A2(n5189), .ZN(n5188) );
  AND2_X1 U5274 ( .A1(n5191), .A2(n9030), .ZN(n5189) );
  AND2_X1 U5275 ( .A1(n6056), .A2(n6117), .ZN(n9048) );
  INV_X1 U5276 ( .A(n8697), .ZN(n5250) );
  INV_X1 U5277 ( .A(n8707), .ZN(n5249) );
  NAND2_X1 U5278 ( .A1(n9116), .A2(n5251), .ZN(n5247) );
  NAND2_X1 U5279 ( .A1(n5187), .A2(n5190), .ZN(n9072) );
  NAND2_X1 U5280 ( .A1(n5970), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5995) );
  INV_X1 U5281 ( .A(n5971), .ZN(n5970) );
  NAND2_X1 U5282 ( .A1(n9167), .A2(n4871), .ZN(n9153) );
  OR2_X1 U5283 ( .A1(n9337), .A2(n8554), .ZN(n8662) );
  AND4_X1 U5284 ( .A1(n5894), .A2(n5893), .A3(n5892), .A4(n5891), .ZN(n9215)
         );
  NAND2_X1 U5285 ( .A1(n7975), .A2(n10649), .ZN(n9236) );
  NAND2_X1 U5286 ( .A1(n5195), .A2(n4886), .ZN(n5194) );
  NAND2_X1 U5287 ( .A1(n5199), .A2(n4886), .ZN(n5196) );
  NAND2_X1 U5288 ( .A1(n5200), .A2(n5199), .ZN(n7652) );
  AND2_X1 U5289 ( .A1(n10495), .A2(n8614), .ZN(n7235) );
  NAND2_X1 U5290 ( .A1(n5267), .A2(n4867), .ZN(n7252) );
  NAND2_X1 U5291 ( .A1(n5175), .A2(n7080), .ZN(n5177) );
  NOR2_X1 U5292 ( .A1(n8744), .A2(n5176), .ZN(n5175) );
  INV_X1 U5293 ( .A(n6980), .ZN(n5176) );
  NAND2_X1 U5294 ( .A1(n6989), .A2(n6975), .ZN(n5178) );
  OAI21_X1 U5295 ( .B1(n7238), .B2(n7237), .A(n8611), .ZN(n9248) );
  AND2_X1 U5296 ( .A1(n5157), .A2(n5155), .ZN(n7041) );
  NOR2_X1 U5297 ( .A1(n6568), .A2(n5156), .ZN(n5155) );
  INV_X1 U5298 ( .A(n9214), .ZN(n10587) );
  NAND2_X1 U5299 ( .A1(n7797), .A2(n8763), .ZN(n6877) );
  NAND2_X1 U5300 ( .A1(n5170), .A2(n5169), .ZN(n5487) );
  INV_X1 U5301 ( .A(n5171), .ZN(n5170) );
  NAND2_X1 U5302 ( .A1(n6065), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6095) );
  INV_X1 U5303 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U5304 ( .A1(n5278), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5514) );
  INV_X1 U5305 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5509) );
  INV_X1 U5306 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5513) );
  INV_X1 U5307 ( .A(n5296), .ZN(n5295) );
  AND3_X1 U5308 ( .A1(n5814), .A2(n5818), .A3(n5828), .ZN(n5507) );
  INV_X1 U5309 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5828) );
  NOR2_X1 U5310 ( .A1(n5592), .A2(n5296), .ZN(n5787) );
  AND2_X1 U5311 ( .A1(n7141), .A2(n7068), .ZN(n5051) );
  NOR2_X1 U5312 ( .A1(n7137), .A2(n7140), .ZN(n7141) );
  NAND2_X1 U5313 ( .A1(n9493), .A2(n9494), .ZN(n8046) );
  NOR2_X1 U5314 ( .A1(n8193), .A2(n8192), .ZN(n9393) );
  INV_X1 U5315 ( .A(n8180), .ZN(n5395) );
  AOI21_X1 U5316 ( .B1(n5385), .B2(n5384), .A(n4921), .ZN(n5383) );
  INV_X1 U5317 ( .A(n9411), .ZN(n5384) );
  OR2_X1 U5318 ( .A1(n9403), .A2(n5045), .ZN(n5044) );
  INV_X1 U5319 ( .A(n5042), .ZN(n5041) );
  OAI21_X1 U5320 ( .B1(n9403), .B2(n5043), .A(n9402), .ZN(n5042) );
  OR2_X1 U5321 ( .A1(n9475), .A2(n5045), .ZN(n5043) );
  AND2_X1 U5322 ( .A1(n9403), .A2(n5040), .ZN(n5039) );
  OR2_X1 U5323 ( .A1(n9475), .A2(n5045), .ZN(n5040) );
  OAI21_X1 U5324 ( .B1(n10452), .B2(n6906), .A(n6889), .ZN(n5053) );
  AOI22_X1 U5325 ( .A1(n6883), .A2(n8155), .B1(n7206), .B2(n8191), .ZN(n6896)
         );
  INV_X1 U5326 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7718) );
  INV_X1 U5327 ( .A(n7704), .ZN(n5392) );
  OR2_X1 U5328 ( .A1(n7765), .A2(n7554), .ZN(n5033) );
  INV_X1 U5329 ( .A(n7555), .ZN(n5035) );
  NAND2_X1 U5330 ( .A1(n8045), .A2(n8044), .ZN(n9492) );
  NOR2_X1 U5331 ( .A1(n9503), .A2(n5397), .ZN(n5396) );
  INV_X1 U5332 ( .A(n8159), .ZN(n5397) );
  NAND2_X1 U5333 ( .A1(n4954), .A2(n4952), .ZN(n8362) );
  AND2_X1 U5334 ( .A1(n8130), .A2(n8129), .ZN(n9430) );
  CLKBUF_X1 U5335 ( .A(n6155), .Z(n6780) );
  AND2_X1 U5336 ( .A1(n8172), .A2(n8171), .ZN(n9647) );
  AND2_X1 U5337 ( .A1(n8818), .A2(n8449), .ZN(n9638) );
  OR2_X1 U5338 ( .A1(n8163), .A2(n9506), .ZN(n8165) );
  NAND2_X1 U5339 ( .A1(n5132), .A2(n8796), .ZN(n9655) );
  NAND2_X1 U5340 ( .A1(n4982), .A2(n4981), .ZN(n5132) );
  AOI21_X1 U5341 ( .B1(n4983), .B2(n4986), .A(n9675), .ZN(n4981) );
  NOR2_X1 U5342 ( .A1(n8794), .A2(n4993), .ZN(n4992) );
  INV_X1 U5343 ( .A(n8793), .ZN(n4993) );
  AOI21_X1 U5344 ( .B1(n4991), .B2(n4990), .A(n4989), .ZN(n4988) );
  INV_X1 U5345 ( .A(n8794), .ZN(n4990) );
  NOR2_X1 U5346 ( .A1(n9705), .A2(n9460), .ZN(n4989) );
  AND2_X1 U5347 ( .A1(n8792), .A2(n8793), .ZN(n4991) );
  AND2_X1 U5348 ( .A1(n8815), .A2(n8489), .ZN(n9686) );
  OR2_X1 U5349 ( .A1(n8077), .A2(n8076), .ZN(n8093) );
  NAND2_X1 U5350 ( .A1(n4923), .A2(n8791), .ZN(n5322) );
  OR2_X1 U5351 ( .A1(n9885), .A2(n9780), .ZN(n9738) );
  NAND2_X1 U5352 ( .A1(n7893), .A2(n5120), .ZN(n7926) );
  INV_X1 U5353 ( .A(n4961), .ZN(n7943) );
  OR2_X1 U5354 ( .A1(n7719), .A2(n7718), .ZN(n7773) );
  NAND2_X1 U5355 ( .A1(n7865), .A2(n7864), .ZN(n7866) );
  NAND2_X1 U5356 ( .A1(n7866), .A2(n8510), .ZN(n7893) );
  NAND2_X1 U5357 ( .A1(n5135), .A2(n5133), .ZN(n7903) );
  NAND2_X1 U5358 ( .A1(n5136), .A2(n7805), .ZN(n5135) );
  NAND2_X1 U5359 ( .A1(n5204), .A2(n5201), .ZN(n7806) );
  OR2_X1 U5360 ( .A1(n7753), .A2(n5203), .ZN(n5201) );
  NOR2_X1 U5361 ( .A1(n8507), .A2(n5318), .ZN(n5317) );
  INV_X1 U5362 ( .A(n7747), .ZN(n5318) );
  NAND2_X1 U5363 ( .A1(n5205), .A2(n8389), .ZN(n7804) );
  NAND2_X1 U5364 ( .A1(n7753), .A2(n7752), .ZN(n5205) );
  NAND2_X1 U5365 ( .A1(n7613), .A2(n7612), .ZN(n7614) );
  NAND2_X1 U5366 ( .A1(n7614), .A2(n8290), .ZN(n7748) );
  AND2_X1 U5367 ( .A1(n8388), .A2(n8382), .ZN(n8505) );
  NAND2_X1 U5368 ( .A1(n5131), .A2(n5130), .ZN(n8402) );
  NAND2_X1 U5369 ( .A1(n5321), .A2(n8284), .ZN(n7446) );
  INV_X1 U5370 ( .A(n7296), .ZN(n5321) );
  INV_X1 U5371 ( .A(n7049), .ZN(n8028) );
  NAND2_X1 U5372 ( .A1(n7289), .A2(n5012), .ZN(n7374) );
  AND2_X1 U5373 ( .A1(n8271), .A2(n7288), .ZN(n5012) );
  INV_X1 U5374 ( .A(n10397), .ZN(n9811) );
  AND2_X1 U5375 ( .A1(n8268), .A2(n7319), .ZN(n8494) );
  OR2_X1 U5376 ( .A1(n7210), .A2(n8494), .ZN(n7289) );
  NAND2_X1 U5377 ( .A1(n8496), .A2(n10403), .ZN(n7108) );
  INV_X1 U5378 ( .A(n10393), .ZN(n9779) );
  NAND2_X1 U5379 ( .A1(n10405), .A2(n10389), .ZN(n10391) );
  AOI21_X1 U5380 ( .B1(n5107), .B2(n10393), .A(n5230), .ZN(n5229) );
  AND2_X1 U5381 ( .A1(n9607), .A2(n9532), .ZN(n5230) );
  INV_X1 U5382 ( .A(n7891), .ZN(n10638) );
  AND2_X1 U5383 ( .A1(n7197), .A2(n6677), .ZN(n10501) );
  AOI21_X1 U5384 ( .B1(n5339), .B2(n5341), .A(n5336), .ZN(n5335) );
  INV_X1 U5385 ( .A(n8252), .ZN(n5336) );
  NOR2_X1 U5386 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n5011) );
  INV_X1 U5387 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6406) );
  NAND2_X1 U5388 ( .A1(n6349), .A2(n5224), .ZN(n5008) );
  OR2_X1 U5389 ( .A1(n6161), .A2(n6162), .ZN(n6164) );
  NOR2_X1 U5390 ( .A1(n5402), .A2(n5221), .ZN(n5220) );
  OAI21_X1 U5391 ( .B1(n6374), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6375) );
  NAND2_X1 U5392 ( .A1(n5368), .A2(n5366), .ZN(n5989) );
  NAND2_X1 U5393 ( .A1(n5367), .A2(n4937), .ZN(n5366) );
  NOR2_X1 U5394 ( .A1(n5966), .A2(n5375), .ZN(n5374) );
  INV_X1 U5395 ( .A(n5950), .ZN(n5375) );
  XNOR2_X1 U5396 ( .A(n6166), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8264) );
  NAND2_X1 U5397 ( .A1(n5936), .A2(n5935), .ZN(n5951) );
  AND2_X1 U5398 ( .A1(n6170), .A2(n6169), .ZN(n8483) );
  OR2_X1 U5399 ( .A1(n6168), .A2(n6167), .ZN(n6169) );
  XNOR2_X1 U5400 ( .A(n5931), .B(n5930), .ZN(n8050) );
  NAND2_X1 U5401 ( .A1(n5352), .A2(n5915), .ZN(n5931) );
  OR2_X1 U5402 ( .A1(n6758), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n7094) );
  NAND2_X1 U5403 ( .A1(n5813), .A2(n5567), .ZN(n5826) );
  NAND2_X1 U5404 ( .A1(n5565), .A2(n5363), .ZN(n5813) );
  NOR2_X1 U5405 ( .A1(n5810), .A2(n5364), .ZN(n5363) );
  INV_X1 U5406 ( .A(n5564), .ZN(n5364) );
  XNOR2_X1 U5407 ( .A(n5786), .B(n5785), .ZN(n7767) );
  NAND2_X1 U5408 ( .A1(n5728), .A2(n5727), .ZN(n5324) );
  NAND2_X1 U5409 ( .A1(n5324), .A2(n5323), .ZN(n5752) );
  AND2_X1 U5410 ( .A1(n5559), .A2(n5557), .ZN(n5323) );
  INV_X1 U5411 ( .A(n5749), .ZN(n5559) );
  AOI21_X1 U5412 ( .B1(n8904), .B2(n8900), .A(n8902), .ZN(n8850) );
  NAND2_X1 U5413 ( .A1(n6110), .A2(n6109), .ZN(n9278) );
  OAI21_X1 U5414 ( .B1(n7990), .B2(n5844), .A(n7989), .ZN(n7994) );
  NAND2_X1 U5415 ( .A1(n5581), .A2(n5580), .ZN(n9343) );
  AND4_X1 U5416 ( .A1(n5908), .A2(n5907), .A3(n5906), .A4(n5905), .ZN(n8924)
         );
  NAND2_X1 U5417 ( .A1(n5404), .A2(n5406), .ZN(n5629) );
  INV_X1 U5418 ( .A(n5405), .ZN(n5404) );
  NAND2_X1 U5419 ( .A1(n5887), .A2(n5886), .ZN(n9331) );
  NAND2_X1 U5420 ( .A1(n6971), .A2(n4912), .ZN(n5065) );
  INV_X1 U5421 ( .A(n9216), .ZN(n9230) );
  INV_X1 U5422 ( .A(n8914), .ZN(n9103) );
  INV_X1 U5423 ( .A(n8562), .ZN(n9118) );
  INV_X1 U5424 ( .A(n8894), .ZN(n9139) );
  INV_X1 U5425 ( .A(n8859), .ZN(n9146) );
  INV_X1 U5426 ( .A(n8558), .ZN(n9161) );
  NOR2_X1 U5427 ( .A1(n6247), .A2(n5023), .ZN(n6237) );
  AND2_X1 U5428 ( .A1(n6250), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5023) );
  NOR2_X1 U5429 ( .A1(n6320), .A2(n5024), .ZN(n7161) );
  AND2_X1 U5430 ( .A1(n6401), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5024) );
  NAND2_X1 U5431 ( .A1(n7161), .A2(n7160), .ZN(n7159) );
  NOR2_X1 U5432 ( .A1(n7428), .A2(n7427), .ZN(n7426) );
  NAND2_X1 U5433 ( .A1(n6224), .A2(n6221), .ZN(n10320) );
  AOI21_X1 U5434 ( .B1(n4968), .B2(n9234), .A(n4965), .ZN(n9281) );
  NAND2_X1 U5435 ( .A1(n4967), .A2(n4966), .ZN(n4965) );
  XNOR2_X1 U5436 ( .A(n9045), .B(n9044), .ZN(n4968) );
  NAND2_X1 U5437 ( .A1(n9046), .A2(n10587), .ZN(n4966) );
  NOR2_X1 U5438 ( .A1(n9109), .A2(n4956), .ZN(n9302) );
  AND2_X1 U5439 ( .A1(n9110), .A2(n9111), .ZN(n4956) );
  INV_X1 U5440 ( .A(n10382), .ZN(n9260) );
  AND2_X1 U5441 ( .A1(n10605), .A2(n10596), .ZN(n9263) );
  INV_X1 U5442 ( .A(n9263), .ZN(n9244) );
  AND2_X1 U5443 ( .A1(n5485), .A2(n5174), .ZN(n5173) );
  INV_X1 U5444 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5174) );
  NAND2_X1 U5445 ( .A1(n7877), .A2(n4888), .ZN(n5055) );
  INV_X1 U5446 ( .A(n7876), .ZN(n5057) );
  AND4_X1 U5447 ( .A1(n7861), .A2(n7860), .A3(n7859), .A4(n7858), .ZN(n9441)
         );
  INV_X1 U5448 ( .A(n7225), .ZN(n10426) );
  AND4_X1 U5449 ( .A1(n7942), .A2(n7941), .A3(n7940), .A4(n7939), .ZN(n9497)
         );
  AND2_X1 U5450 ( .A1(n8151), .A2(n8150), .ZN(n9690) );
  INV_X1 U5451 ( .A(n9742), .ZN(n9709) );
  NAND4_X1 U5452 ( .A1(n6444), .A2(n6443), .A3(n6442), .A4(n6441), .ZN(n7322)
         );
  OR2_X1 U5453 ( .A1(n8145), .A2(n7211), .ZN(n6442) );
  AOI21_X1 U5454 ( .B1(n9955), .B2(n8355), .A(n8258), .ZN(n9831) );
  NAND2_X1 U5455 ( .A1(n8121), .A2(n8120), .ZN(n9866) );
  AND2_X1 U5456 ( .A1(n9822), .A2(n7028), .ZN(n9825) );
  NAND2_X1 U5457 ( .A1(n5094), .A2(n5001), .ZN(n9841) );
  NAND2_X1 U5458 ( .A1(n9620), .A2(n5095), .ZN(n5094) );
  INV_X1 U5459 ( .A(n5002), .ZN(n5001) );
  OAI21_X1 U5460 ( .B1(n4873), .B2(n10645), .A(n5104), .ZN(n5100) );
  OR2_X1 U5461 ( .A1(n10491), .A2(n5105), .ZN(n5104) );
  INV_X1 U5462 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5105) );
  AND2_X1 U5463 ( .A1(n10491), .A2(n10397), .ZN(n5098) );
  INV_X1 U5464 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9950) );
  INV_X1 U5465 ( .A(n8483), .ZN(n8525) );
  XNOR2_X1 U5466 ( .A(n6633), .B(n6632), .ZN(n6648) );
  INV_X1 U5467 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6635) );
  NAND2_X1 U5468 ( .A1(n8615), .A2(n8614), .ZN(n5292) );
  AND2_X1 U5469 ( .A1(n5288), .A2(n5287), .ZN(n8623) );
  INV_X1 U5470 ( .A(n8620), .ZN(n5287) );
  NAND2_X1 U5471 ( .A1(n5290), .A2(n5289), .ZN(n5288) );
  NAND2_X1 U5472 ( .A1(n8623), .A2(n5285), .ZN(n8625) );
  NAND2_X1 U5473 ( .A1(n5286), .A2(n8928), .ZN(n5285) );
  NAND2_X1 U5474 ( .A1(n5301), .A2(n8632), .ZN(n5298) );
  AOI21_X1 U5475 ( .B1(n5301), .B2(n5304), .A(n5300), .ZN(n5299) );
  AOI21_X1 U5476 ( .B1(n4915), .B2(n8727), .A(n5305), .ZN(n5304) );
  NOR2_X1 U5477 ( .A1(n8634), .A2(n8727), .ZN(n5305) );
  AOI21_X1 U5478 ( .B1(n5308), .B2(n5306), .A(n8696), .ZN(n8702) );
  NOR2_X1 U5479 ( .A1(n8690), .A2(n5307), .ZN(n5306) );
  NOR2_X1 U5480 ( .A1(n5128), .A2(n10023), .ZN(n5127) );
  INV_X1 U5481 ( .A(n5561), .ZN(n5128) );
  NAND2_X1 U5482 ( .A1(n4893), .A2(n5332), .ZN(n5331) );
  NOR2_X1 U5483 ( .A1(n9843), .A2(n9848), .ZN(n5154) );
  INV_X1 U5484 ( .A(SI_27_), .ZN(n10000) );
  NAND2_X1 U5485 ( .A1(n5372), .A2(n4936), .ZN(n5371) );
  NAND2_X1 U5486 ( .A1(n5984), .A2(n5373), .ZN(n5372) );
  INV_X1 U5487 ( .A(n5965), .ZN(n5373) );
  INV_X1 U5488 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6147) );
  INV_X1 U5489 ( .A(SI_15_), .ZN(n10097) );
  INV_X1 U5490 ( .A(n5825), .ZN(n5365) );
  NOR2_X1 U5491 ( .A1(n5127), .A2(n5126), .ZN(n5125) );
  INV_X1 U5492 ( .A(n5560), .ZN(n5126) );
  INV_X1 U5493 ( .A(n5127), .ZN(n5123) );
  INV_X1 U5494 ( .A(SI_9_), .ZN(n10142) );
  AND2_X1 U5495 ( .A1(n5416), .A2(n5423), .ZN(n5410) );
  NOR2_X1 U5496 ( .A1(n5416), .A2(n5423), .ZN(n5411) );
  AND2_X1 U5497 ( .A1(n5409), .A2(n4931), .ZN(n5414) );
  NAND2_X1 U5498 ( .A1(n5416), .A2(n5420), .ZN(n5409) );
  OR2_X1 U5499 ( .A1(n5949), .A2(n5948), .ZN(n5433) );
  NOR2_X1 U5500 ( .A1(n7607), .A2(n5448), .ZN(n5447) );
  INV_X1 U5501 ( .A(n5450), .ZN(n5448) );
  OAI21_X1 U5502 ( .B1(n7589), .B2(P2_REG1_REG_14__SCAN_IN), .A(n7590), .ZN(
        n6190) );
  NAND2_X1 U5503 ( .A1(n9027), .A2(n8705), .ZN(n5276) );
  INV_X1 U5504 ( .A(n8715), .ZN(n5272) );
  INV_X1 U5505 ( .A(n8705), .ZN(n5273) );
  NOR2_X1 U5506 ( .A1(n9029), .A2(n9028), .ZN(n5468) );
  INV_X1 U5507 ( .A(n9023), .ZN(n5192) );
  INV_X1 U5508 ( .A(n9111), .ZN(n5193) );
  OR2_X1 U5509 ( .A1(n9311), .A2(n8859), .ZN(n8683) );
  INV_X1 U5510 ( .A(n5197), .ZN(n5195) );
  OR2_X1 U5511 ( .A1(n7033), .A2(n8741), .ZN(n8597) );
  NAND2_X1 U5512 ( .A1(n5159), .A2(n5158), .ZN(n7084) );
  INV_X1 U5513 ( .A(n7040), .ZN(n5159) );
  NAND2_X1 U5514 ( .A1(n7035), .A2(n8741), .ZN(n7034) );
  NOR2_X1 U5515 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5474) );
  NOR2_X1 U5516 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5475) );
  INV_X1 U5517 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5454) );
  NOR2_X2 U5518 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5604) );
  OR2_X1 U5519 ( .A1(n5661), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5675) );
  INV_X1 U5520 ( .A(n7543), .ZN(n7544) );
  NAND2_X1 U5521 ( .A1(n5379), .A2(n4908), .ZN(n8042) );
  NAND2_X1 U5522 ( .A1(n4934), .A2(n5381), .ZN(n5380) );
  INV_X1 U5523 ( .A(n8347), .ZN(n8350) );
  OR2_X1 U5524 ( .A1(n9740), .A2(n9760), .ZN(n8516) );
  OR2_X1 U5525 ( .A1(n9901), .A2(n9497), .ZN(n8808) );
  NAND2_X1 U5526 ( .A1(n5110), .A2(n8805), .ZN(n5109) );
  NOR2_X1 U5527 ( .A1(n9908), .A2(n9912), .ZN(n5141) );
  INV_X1 U5528 ( .A(n5203), .ZN(n5202) );
  NAND2_X1 U5529 ( .A1(n5206), .A2(n8392), .ZN(n5204) );
  NAND2_X1 U5530 ( .A1(n8392), .A2(n8389), .ZN(n5203) );
  AND2_X1 U5531 ( .A1(n8393), .A2(n8380), .ZN(n7805) );
  NAND2_X1 U5532 ( .A1(n10562), .A2(n5145), .ZN(n5149) );
  NAND2_X1 U5533 ( .A1(n5219), .A2(n5217), .ZN(n7505) );
  NAND2_X1 U5534 ( .A1(n7450), .A2(n7449), .ZN(n5219) );
  INV_X1 U5535 ( .A(n7378), .ZN(n8499) );
  AND3_X1 U5536 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6426) );
  INV_X1 U5537 ( .A(n8246), .ZN(n5341) );
  INV_X1 U5538 ( .A(n5340), .ZN(n5339) );
  OAI21_X1 U5539 ( .B1(n8244), .B2(n5341), .A(n8353), .ZN(n5340) );
  INV_X1 U5540 ( .A(n5224), .ZN(n5221) );
  OAI21_X1 U5541 ( .B1(n6022), .B2(n5360), .A(n5358), .ZN(n6101) );
  AOI21_X1 U5542 ( .B1(n5361), .B2(n5359), .A(n4945), .ZN(n5358) );
  INV_X1 U5543 ( .A(n5361), .ZN(n5360) );
  NOR2_X1 U5544 ( .A1(n5371), .A2(n5937), .ZN(n5369) );
  INV_X1 U5545 ( .A(n5371), .ZN(n5367) );
  AND2_X1 U5546 ( .A1(n6156), .A2(n6149), .ZN(n6370) );
  NAND2_X1 U5547 ( .A1(n6165), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6168) );
  NOR2_X1 U5548 ( .A1(n5916), .A2(n5357), .ZN(n5356) );
  INV_X1 U5549 ( .A(n5897), .ZN(n5357) );
  INV_X1 U5550 ( .A(SI_13_), .ZN(n10134) );
  AOI21_X1 U5551 ( .B1(n5691), .B2(n5347), .A(n4920), .ZN(n5345) );
  INV_X1 U5552 ( .A(n5347), .ZN(n5346) );
  INV_X1 U5553 ( .A(SI_5_), .ZN(n10034) );
  OAI21_X1 U5554 ( .B1(n6718), .B2(n5525), .A(n5524), .ZN(n5526) );
  INV_X1 U5555 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U5556 ( .A1(n6718), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5524) );
  NOR2_X1 U5557 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6332) );
  INV_X1 U5558 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5049) );
  OR2_X1 U5559 ( .A1(n5689), .A2(n5690), .ZN(n5064) );
  NOR2_X1 U5560 ( .A1(n8911), .A2(n5422), .ZN(n5421) );
  INV_X1 U5561 ( .A(n8866), .ZN(n5422) );
  NAND2_X1 U5562 ( .A1(n5075), .A2(n5072), .ZN(n5979) );
  NOR2_X1 U5563 ( .A1(n5074), .A2(n5073), .ZN(n5072) );
  NOR2_X1 U5564 ( .A1(n5080), .A2(n5076), .ZN(n5074) );
  NAND2_X1 U5565 ( .A1(n5723), .A2(n5451), .ZN(n5450) );
  INV_X1 U5566 ( .A(n5726), .ZN(n5451) );
  INV_X1 U5567 ( .A(n5836), .ZN(n5495) );
  INV_X1 U5568 ( .A(n5943), .ZN(n5942) );
  INV_X1 U5569 ( .A(n8892), .ZN(n5077) );
  NAND2_X1 U5570 ( .A1(n8904), .A2(n5081), .ZN(n5078) );
  NOR2_X1 U5571 ( .A1(n5071), .A2(n5084), .ZN(n5079) );
  INV_X1 U5572 ( .A(n5080), .ZN(n5071) );
  NOR2_X1 U5573 ( .A1(n6849), .A2(n6870), .ZN(n5061) );
  XNOR2_X1 U5574 ( .A(n5863), .B(n6843), .ZN(n5062) );
  OR2_X1 U5575 ( .A1(n5889), .A2(n5888), .ZN(n5903) );
  NAND2_X1 U5576 ( .A1(n5284), .A2(n5283), .ZN(n5282) );
  NOR2_X1 U5577 ( .A1(n5325), .A2(n8761), .ZN(n8762) );
  NAND2_X1 U5578 ( .A1(n8726), .A2(n5326), .ZN(n5325) );
  NOR2_X1 U5579 ( .A1(n9033), .A2(n5327), .ZN(n5326) );
  INV_X1 U5580 ( .A(n6877), .ZN(n8733) );
  NOR2_X1 U5581 ( .A1(n8761), .A2(n8768), .ZN(n5260) );
  AND3_X1 U5582 ( .A1(n8577), .A2(n8576), .A3(n8575), .ZN(n8729) );
  AOI21_X1 U5583 ( .B1(n9048), .B2(n6122), .A(n6060), .ZN(n8923) );
  AND2_X1 U5584 ( .A1(n6002), .A2(n6001), .ZN(n8562) );
  AND4_X1 U5585 ( .A1(n5746), .A2(n5745), .A3(n5744), .A4(n5743), .ZN(n7577)
         );
  AND4_X1 U5586 ( .A1(n5646), .A2(n5645), .A3(n5644), .A4(n5643), .ZN(n6976)
         );
  OR2_X1 U5587 ( .A1(n8572), .A2(n5630), .ZN(n5632) );
  NOR2_X1 U5588 ( .A1(n10309), .A2(n5025), .ZN(n10308) );
  NAND2_X1 U5589 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n5025) );
  OR2_X1 U5590 ( .A1(n6298), .A2(n6297), .ZN(n5028) );
  AOI21_X1 U5591 ( .B1(n6359), .B2(P2_REG1_REG_8__SCAN_IN), .A(n6293), .ZN(
        n6307) );
  NAND2_X1 U5592 ( .A1(n7434), .A2(n7435), .ZN(n7433) );
  NAND2_X1 U5593 ( .A1(n7433), .A2(n4955), .ZN(n7591) );
  NAND2_X1 U5594 ( .A1(n7444), .A2(n6175), .ZN(n4955) );
  NAND2_X1 U5595 ( .A1(n7595), .A2(n5018), .ZN(n6215) );
  NAND2_X1 U5596 ( .A1(n5020), .A2(n5019), .ZN(n5018) );
  OAI21_X1 U5597 ( .B1(n9055), .B2(n5274), .A(n5271), .ZN(n9009) );
  INV_X1 U5598 ( .A(n5275), .ZN(n5274) );
  AOI21_X1 U5599 ( .B1(n5275), .B2(n5273), .A(n5272), .ZN(n5271) );
  AND2_X1 U5600 ( .A1(n9050), .A2(n5276), .ZN(n5275) );
  OAI21_X1 U5601 ( .B1(n9055), .B2(n9027), .A(n8705), .ZN(n9045) );
  NAND2_X1 U5602 ( .A1(n9081), .A2(n9230), .ZN(n4967) );
  OR2_X1 U5603 ( .A1(n9298), .A2(n8562), .ZN(n8697) );
  NAND2_X1 U5604 ( .A1(n9123), .A2(n9107), .ZN(n9089) );
  OAI21_X1 U5605 ( .B1(n9167), .B2(n5181), .A(n5179), .ZN(n9021) );
  INV_X1 U5606 ( .A(n5180), .ZN(n5179) );
  AND2_X1 U5607 ( .A1(n8693), .A2(n9101), .ZN(n9121) );
  NAND2_X1 U5608 ( .A1(n5240), .A2(n5242), .ZN(n9138) );
  AOI21_X1 U5609 ( .B1(n9156), .B2(n8679), .A(n5243), .ZN(n5242) );
  INV_X1 U5610 ( .A(n8559), .ZN(n5243) );
  OR2_X1 U5611 ( .A1(n9148), .A2(n9311), .ZN(n4884) );
  NAND2_X1 U5612 ( .A1(n5164), .A2(n5163), .ZN(n9148) );
  AOI21_X1 U5613 ( .B1(n9204), .B2(n9192), .A(n9016), .ZN(n9179) );
  AOI21_X1 U5614 ( .B1(n5237), .B2(n5239), .A(n4914), .ZN(n5234) );
  AND4_X1 U5615 ( .A1(n5502), .A2(n5501), .A3(n5500), .A4(n5499), .ZN(n9217)
         );
  NOR2_X1 U5616 ( .A1(n8757), .A2(n5186), .ZN(n5185) );
  AND4_X1 U5617 ( .A1(n5840), .A2(n5839), .A3(n5838), .A4(n5837), .ZN(n7983)
         );
  NOR2_X1 U5618 ( .A1(n8737), .A2(n5198), .ZN(n5197) );
  INV_X1 U5619 ( .A(n7651), .ZN(n5198) );
  AND4_X1 U5620 ( .A1(n5779), .A2(n5778), .A3(n5777), .A4(n5776), .ZN(n8224)
         );
  AND4_X1 U5621 ( .A1(n5809), .A2(n5808), .A3(n5807), .A4(n5806), .ZN(n7841)
         );
  NAND2_X1 U5622 ( .A1(n4975), .A2(n4974), .ZN(n10591) );
  AND4_X1 U5623 ( .A1(n5764), .A2(n5763), .A3(n5762), .A4(n5761), .ZN(n7789)
         );
  AND4_X1 U5624 ( .A1(n5798), .A2(n5797), .A3(n5796), .A4(n5795), .ZN(n8210)
         );
  OR2_X1 U5625 ( .A1(n5759), .A2(n10078), .ZN(n5793) );
  AOI21_X1 U5626 ( .B1(n5254), .B2(n5257), .A(n10581), .ZN(n5252) );
  NAND2_X1 U5627 ( .A1(n7469), .A2(n7468), .ZN(n10583) );
  NAND2_X1 U5628 ( .A1(n7334), .A2(n7333), .ZN(n7469) );
  AND4_X1 U5629 ( .A1(n5589), .A2(n5588), .A3(n5587), .A4(n5586), .ZN(n7331)
         );
  AND4_X1 U5630 ( .A1(n5703), .A2(n5702), .A3(n5701), .A4(n5700), .ZN(n7256)
         );
  AND2_X1 U5631 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5679) );
  OR2_X1 U5632 ( .A1(n7076), .A2(n6982), .ZN(n6983) );
  AND2_X1 U5633 ( .A1(n8607), .A2(n8611), .ZN(n8744) );
  NAND2_X1 U5634 ( .A1(n6981), .A2(n8602), .ZN(n7076) );
  INV_X1 U5635 ( .A(n8932), .ZN(n6849) );
  NAND2_X1 U5636 ( .A1(n6125), .A2(n6129), .ZN(n9214) );
  AND2_X1 U5637 ( .A1(n5160), .A2(n5622), .ZN(n5157) );
  OR2_X1 U5638 ( .A1(n5991), .A2(n6719), .ZN(n5160) );
  NAND2_X1 U5639 ( .A1(n6563), .A2(n6562), .ZN(n8590) );
  OR2_X1 U5640 ( .A1(n6173), .A2(n6096), .ZN(n6864) );
  INV_X1 U5641 ( .A(n10648), .ZN(n10628) );
  INV_X1 U5642 ( .A(n10650), .ZN(n10629) );
  NAND2_X1 U5643 ( .A1(n6492), .A2(n8733), .ZN(n10648) );
  AND3_X1 U5644 ( .A1(n6862), .A2(n6865), .A3(n6490), .ZN(n6503) );
  INV_X1 U5645 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10078) );
  MUX2_X1 U5646 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5573), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n5574) );
  NAND2_X1 U5647 ( .A1(n5452), .A2(n5066), .ZN(n5515) );
  XNOR2_X1 U5648 ( .A(n5517), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8592) );
  INV_X1 U5649 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5508) );
  INV_X1 U5650 ( .A(n8155), .ZN(n8196) );
  INV_X1 U5651 ( .A(n6739), .ZN(n6740) );
  OR2_X1 U5652 ( .A1(n8020), .A2(n8019), .ZN(n5382) );
  OR2_X1 U5653 ( .A1(n8049), .A2(n8048), .ZN(n5388) );
  NOR3_X1 U5654 ( .A1(n7555), .A2(n7554), .A3(n7739), .ZN(n7705) );
  XNOR2_X1 U5655 ( .A(n7056), .B(n8188), .ZN(n7060) );
  NAND2_X1 U5656 ( .A1(n7060), .A2(n7059), .ZN(n7139) );
  OR2_X1 U5657 ( .A1(n6631), .A2(n7022), .ZN(n6666) );
  AND4_X1 U5658 ( .A1(n7778), .A2(n7777), .A3(n7776), .A4(n7775), .ZN(n9520)
         );
  OR2_X1 U5659 ( .A1(n7853), .A2(n6789), .ZN(n6790) );
  OR2_X1 U5660 ( .A1(n7853), .A2(n6454), .ZN(n6749) );
  NAND2_X1 U5661 ( .A1(n4916), .A2(n6641), .ZN(n7101) );
  OR2_X1 U5662 ( .A1(n6788), .A2(n6637), .ZN(n6641) );
  NOR2_X1 U5663 ( .A1(n9832), .A2(n5151), .ZN(n5150) );
  INV_X1 U5664 ( .A(n5152), .ZN(n5151) );
  AOI21_X1 U5665 ( .B1(n5115), .B2(n9657), .A(n5114), .ZN(n5113) );
  INV_X1 U5666 ( .A(n8818), .ZN(n5114) );
  AOI21_X1 U5667 ( .B1(n4985), .B2(n4984), .A(n4913), .ZN(n4983) );
  INV_X1 U5668 ( .A(n4992), .ZN(n4984) );
  NOR2_X1 U5669 ( .A1(n9744), .A2(n9874), .ZN(n9726) );
  NAND2_X1 U5670 ( .A1(n9726), .A2(n9705), .ZN(n9699) );
  INV_X1 U5671 ( .A(n8093), .ZN(n6937) );
  AND2_X1 U5672 ( .A1(n8813), .A2(n8375), .ZN(n9718) );
  OR2_X1 U5673 ( .A1(n8055), .A2(n8054), .ZN(n8077) );
  AND2_X1 U5674 ( .A1(n9738), .A2(n8327), .ZN(n9752) );
  AND3_X1 U5675 ( .A1(n8081), .A2(n8080), .A3(n8079), .ZN(n9755) );
  AND4_X1 U5676 ( .A1(n8004), .A2(n8003), .A3(n8002), .A4(n8001), .ZN(n9754)
         );
  INV_X1 U5677 ( .A(n9752), .ZN(n9760) );
  NAND2_X1 U5678 ( .A1(n6935), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8035) );
  AND2_X1 U5679 ( .A1(n8435), .A2(n8436), .ZN(n9777) );
  AND2_X1 U5680 ( .A1(n8432), .A2(n8809), .ZN(n9797) );
  AND2_X1 U5681 ( .A1(n5109), .A2(n8808), .ZN(n5108) );
  INV_X1 U5682 ( .A(n5233), .ZN(n5232) );
  NAND2_X1 U5683 ( .A1(n4863), .A2(n9795), .ZN(n9790) );
  AND2_X1 U5684 ( .A1(n9805), .A2(n8783), .ZN(n9789) );
  INV_X1 U5685 ( .A(n9797), .ZN(n9788) );
  OAI21_X1 U5686 ( .B1(n7865), .B2(n5005), .A(n5003), .ZN(n5457) );
  NAND2_X1 U5687 ( .A1(n4872), .A2(n8510), .ZN(n5005) );
  NAND2_X1 U5688 ( .A1(n5004), .A2(n4872), .ZN(n5003) );
  NAND2_X1 U5689 ( .A1(n5457), .A2(n9812), .ZN(n9805) );
  INV_X1 U5690 ( .A(n5231), .ZN(n9813) );
  OAI21_X1 U5691 ( .B1(n7943), .B2(n5233), .A(n8315), .ZN(n5231) );
  NAND2_X1 U5692 ( .A1(n5111), .A2(n5109), .ZN(n9810) );
  AND4_X1 U5693 ( .A1(n8040), .A2(n8039), .A3(n8038), .A4(n8037), .ZN(n9809)
         );
  NAND2_X1 U5694 ( .A1(n7918), .A2(n7917), .ZN(n7931) );
  NAND2_X1 U5695 ( .A1(n7918), .A2(n5141), .ZN(n9817) );
  AND2_X1 U5696 ( .A1(n7929), .A2(n7928), .ZN(n8009) );
  INV_X1 U5697 ( .A(n7773), .ZN(n6933) );
  NAND2_X1 U5698 ( .A1(n5314), .A2(n7801), .ZN(n5313) );
  INV_X1 U5699 ( .A(n5317), .ZN(n5314) );
  NAND2_X1 U5700 ( .A1(n7803), .A2(n8509), .ZN(n7865) );
  NOR2_X1 U5701 ( .A1(n7800), .A2(n5146), .ZN(n5143) );
  AND4_X1 U5702 ( .A1(n7725), .A2(n7724), .A3(n7723), .A4(n7722), .ZN(n8300)
         );
  INV_X1 U5703 ( .A(n5146), .ZN(n5147) );
  AND4_X1 U5704 ( .A1(n7413), .A2(n7412), .A3(n7411), .A4(n7410), .ZN(n7617)
         );
  NOR2_X1 U5705 ( .A1(n7457), .A2(n5149), .ZN(n7620) );
  NOR2_X1 U5706 ( .A1(n7457), .A2(n10547), .ZN(n7519) );
  OR2_X1 U5707 ( .A1(n7501), .A2(n8505), .ZN(n7613) );
  NAND2_X1 U5708 ( .A1(n7503), .A2(n8505), .ZN(n7753) );
  AND4_X1 U5709 ( .A1(n7515), .A2(n7514), .A3(n7513), .A4(n7512), .ZN(n7754)
         );
  AND2_X1 U5710 ( .A1(n7446), .A2(n7447), .ZN(n5086) );
  NAND2_X1 U5711 ( .A1(n5219), .A2(n8387), .ZN(n7452) );
  INV_X1 U5712 ( .A(n8284), .ZN(n8500) );
  OR2_X1 U5713 ( .A1(n7378), .A2(n7292), .ZN(n7296) );
  NOR2_X1 U5714 ( .A1(n7326), .A2(n7299), .ZN(n7386) );
  NAND2_X1 U5715 ( .A1(n8428), .A2(n8402), .ZN(n7378) );
  NAND2_X1 U5716 ( .A1(n10468), .A2(n5137), .ZN(n7326) );
  INV_X1 U5717 ( .A(n5137), .ZN(n7199) );
  NAND2_X1 U5718 ( .A1(n5208), .A2(n5210), .ZN(n7200) );
  NAND2_X1 U5719 ( .A1(n5209), .A2(n8491), .ZN(n7183) );
  NAND2_X1 U5720 ( .A1(n7217), .A2(n8415), .ZN(n5209) );
  OR2_X1 U5721 ( .A1(n7025), .A2(n7024), .ZN(n7390) );
  AND2_X1 U5722 ( .A1(n6648), .A2(n9781), .ZN(n8531) );
  NAND2_X1 U5723 ( .A1(n8346), .A2(n8345), .ZN(n9837) );
  INV_X1 U5724 ( .A(n5106), .ZN(n5096) );
  AOI21_X1 U5725 ( .B1(n9620), .B2(n5106), .A(n5097), .ZN(n5002) );
  OR2_X1 U5726 ( .A1(n9618), .A2(n9624), .ZN(n9620) );
  OR2_X1 U5727 ( .A1(n9843), .A2(n9648), .ZN(n8819) );
  NAND2_X1 U5728 ( .A1(n7103), .A2(n8263), .ZN(n10397) );
  NAND2_X1 U5729 ( .A1(n8162), .A2(n8161), .ZN(n9854) );
  AND2_X1 U5730 ( .A1(n6888), .A2(n5054), .ZN(n10452) );
  AND2_X1 U5731 ( .A1(n6887), .A2(n6886), .ZN(n5054) );
  INV_X1 U5732 ( .A(n10501), .ZN(n10637) );
  AND2_X1 U5733 ( .A1(n7197), .A2(n6648), .ZN(n10482) );
  AND2_X1 U5734 ( .A1(n8532), .A2(n8525), .ZN(n7197) );
  XNOR2_X1 U5735 ( .A(n8354), .B(n8353), .ZN(n8828) );
  NAND2_X1 U5736 ( .A1(n5338), .A2(n8246), .ZN(n8354) );
  NAND2_X1 U5737 ( .A1(n8239), .A2(n6108), .ZN(n8826) );
  OR2_X1 U5738 ( .A1(n6107), .A2(n6106), .ZN(n6108) );
  XNOR2_X1 U5739 ( .A(n6101), .B(n6100), .ZN(n9382) );
  NAND2_X1 U5740 ( .A1(n6370), .A2(n6369), .ZN(n6374) );
  INV_X1 U5741 ( .A(n6370), .ZN(n6371) );
  XNOR2_X1 U5742 ( .A(n6156), .B(n6159), .ZN(n7823) );
  AOI21_X1 U5743 ( .B1(n5353), .B2(n5355), .A(n4940), .ZN(n5351) );
  NOR2_X1 U5744 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n6145) );
  NOR2_X1 U5745 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n6144) );
  NOR2_X1 U5746 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n6143) );
  AND2_X1 U5747 ( .A1(n6349), .A2(n6141), .ZN(n6361) );
  NAND2_X1 U5748 ( .A1(n5878), .A2(n5877), .ZN(n5883) );
  AND2_X1 U5749 ( .A1(n5897), .A2(n5881), .ZN(n5882) );
  NAND2_X1 U5750 ( .A1(n5883), .A2(n5882), .ZN(n5898) );
  AOI21_X1 U5751 ( .B1(n5850), .B2(n5849), .A(n5848), .ZN(n5855) );
  XNOR2_X1 U5752 ( .A(n5320), .B(n5706), .ZN(n7282) );
  NAND2_X1 U5753 ( .A1(n5349), .A2(n5548), .ZN(n5320) );
  INV_X1 U5754 ( .A(n5537), .ZN(n5093) );
  AND2_X1 U5755 ( .A1(n5537), .A2(n5536), .ZN(n5460) );
  NAND2_X1 U5756 ( .A1(n5415), .A2(n5419), .ZN(n8833) );
  NAND2_X1 U5757 ( .A1(n8865), .A2(n5421), .ZN(n5415) );
  NAND2_X1 U5758 ( .A1(n5822), .A2(n5821), .ZN(n8221) );
  NAND2_X1 U5759 ( .A1(n7495), .A2(n5450), .ZN(n7606) );
  OAI22_X1 U5760 ( .A1(n6577), .A2(n6576), .B1(n5060), .B2(n5059), .ZN(n6703)
         );
  INV_X1 U5761 ( .A(n5062), .ZN(n5060) );
  INV_X1 U5762 ( .A(n5061), .ZN(n5059) );
  AOI21_X1 U5763 ( .B1(n6840), .B2(n8768), .A(n5628), .ZN(n6697) );
  INV_X1 U5764 ( .A(n10510), .ZN(n8873) );
  NAND2_X1 U5765 ( .A1(n5432), .A2(n5437), .ZN(n8857) );
  NAND2_X1 U5766 ( .A1(n8850), .A2(n5438), .ZN(n5432) );
  OAI21_X1 U5767 ( .B1(n7171), .B2(n4868), .A(n5070), .ZN(n8228) );
  NAND2_X1 U5768 ( .A1(n8138), .A2(n8580), .ZN(n4949) );
  NAND2_X1 U5769 ( .A1(n5427), .A2(n6708), .ZN(n6767) );
  NAND2_X1 U5770 ( .A1(n6711), .A2(n6709), .ZN(n5427) );
  AND2_X1 U5771 ( .A1(n5978), .A2(n5977), .ZN(n8894) );
  NAND2_X1 U5772 ( .A1(n7171), .A2(n5725), .ZN(n7495) );
  AND2_X1 U5773 ( .A1(n5440), .A2(n4938), .ZN(n8885) );
  NAND2_X1 U5774 ( .A1(n8850), .A2(n8848), .ZN(n5440) );
  NAND2_X1 U5775 ( .A1(n5789), .A2(n5788), .ZN(n10627) );
  NAND2_X1 U5776 ( .A1(n5078), .A2(n5079), .ZN(n8893) );
  NAND2_X1 U5777 ( .A1(n6116), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10523) );
  NAND2_X1 U5778 ( .A1(n5426), .A2(n4904), .ZN(n6971) );
  INV_X1 U5779 ( .A(n6769), .ZN(n5431) );
  AOI21_X1 U5780 ( .B1(n8865), .B2(n8866), .A(n5462), .ZN(n8912) );
  NAND2_X1 U5781 ( .A1(n6027), .A2(n6026), .ZN(n9289) );
  NAND2_X1 U5782 ( .A1(n5831), .A2(n5830), .ZN(n9347) );
  INV_X1 U5783 ( .A(n7797), .ZN(n8774) );
  INV_X1 U5784 ( .A(n8867), .ZN(n9096) );
  INV_X1 U5785 ( .A(n9215), .ZN(n9174) );
  INV_X1 U5786 ( .A(n7577), .ZN(n10586) );
  INV_X1 U5787 ( .A(n6976), .ZN(n8931) );
  INV_X1 U5788 ( .A(n5168), .ZN(n5167) );
  AND2_X1 U5789 ( .A1(n5633), .A2(n5632), .ZN(n5166) );
  OAI22_X1 U5790 ( .A1(n7042), .A2(n4861), .B1(n8574), .B2(n5631), .ZN(n5168)
         );
  OR2_X1 U5791 ( .A1(n5865), .A2(n5610), .ZN(n5612) );
  OR2_X1 U5792 ( .A1(n4861), .A2(n9983), .ZN(n5614) );
  NAND4_X1 U5793 ( .A1(n5626), .A2(n5625), .A3(n5624), .A4(n5623), .ZN(n8934)
         );
  OR2_X1 U5794 ( .A1(n6030), .A2(n10388), .ZN(n5626) );
  AOI21_X1 U5795 ( .B1(n6287), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6281), .ZN(
        n6259) );
  NOR2_X1 U5796 ( .A1(n6249), .A2(n6248), .ZN(n6247) );
  AOI21_X1 U5797 ( .B1(n6263), .B2(P2_REG1_REG_4__SCAN_IN), .A(n6257), .ZN(
        n6246) );
  INV_X1 U5798 ( .A(n5022), .ZN(n6235) );
  AOI21_X1 U5799 ( .B1(n6238), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6232), .ZN(
        n6271) );
  NAND2_X1 U5800 ( .A1(n6238), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5021) );
  NOR2_X1 U5801 ( .A1(n6272), .A2(n5029), .ZN(n6298) );
  AND2_X1 U5802 ( .A1(n6274), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5029) );
  INV_X1 U5803 ( .A(n5028), .ZN(n6296) );
  NOR2_X1 U5804 ( .A1(n6310), .A2(n6309), .ZN(n6308) );
  AND2_X1 U5805 ( .A1(n5028), .A2(n5027), .ZN(n6310) );
  NAND2_X1 U5806 ( .A1(n6359), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5027) );
  NAND2_X1 U5807 ( .A1(n7159), .A2(n4944), .ZN(n7428) );
  NOR2_X1 U5808 ( .A1(n5592), .A2(n5505), .ZN(n5771) );
  XNOR2_X1 U5809 ( .A(n6215), .B(n8942), .ZN(n8944) );
  NAND2_X1 U5810 ( .A1(n8944), .A2(n5832), .ZN(n8943) );
  NOR2_X1 U5811 ( .A1(n8957), .A2(n8956), .ZN(n8955) );
  AND2_X1 U5812 ( .A1(n5017), .A2(n5016), .ZN(n8973) );
  INV_X1 U5813 ( .A(n6222), .ZN(n5016) );
  INV_X1 U5814 ( .A(n5017), .ZN(n6223) );
  NOR2_X1 U5815 ( .A1(n8973), .A2(n5014), .ZN(n8975) );
  NOR2_X1 U5816 ( .A1(n5015), .A2(n9221), .ZN(n5014) );
  INV_X1 U5817 ( .A(n9047), .ZN(n9035) );
  XNOR2_X1 U5818 ( .A(n9061), .B(n5277), .ZN(n9287) );
  AND2_X1 U5819 ( .A1(n9060), .A2(n9059), .ZN(n9061) );
  NAND2_X1 U5820 ( .A1(n5247), .A2(n5248), .ZN(n9080) );
  NAND2_X1 U5821 ( .A1(n9108), .A2(n9023), .ZN(n9086) );
  OR2_X1 U5822 ( .A1(n9120), .A2(n9121), .ZN(n9304) );
  NAND2_X1 U5823 ( .A1(n9153), .A2(n9019), .ZN(n9131) );
  NAND2_X1 U5824 ( .A1(n9167), .A2(n9018), .ZN(n9155) );
  NAND2_X1 U5825 ( .A1(n5244), .A2(n8675), .ZN(n9144) );
  NAND2_X1 U5826 ( .A1(n9160), .A2(n8557), .ZN(n5244) );
  NAND2_X1 U5827 ( .A1(n5900), .A2(n5899), .ZN(n9327) );
  NAND2_X1 U5828 ( .A1(n9208), .A2(n8756), .ZN(n5236) );
  NAND2_X1 U5829 ( .A1(n7652), .A2(n7651), .ZN(n7653) );
  AND2_X1 U5830 ( .A1(n5267), .A2(n7240), .ZN(n7241) );
  NAND3_X1 U5831 ( .A1(n5177), .A2(n5178), .A3(n7234), .ZN(n10495) );
  NAND2_X1 U5832 ( .A1(n5177), .A2(n5178), .ZN(n9262) );
  NAND2_X1 U5833 ( .A1(n5157), .A2(n5621), .ZN(n7009) );
  INV_X1 U5834 ( .A(n10383), .ZN(n9223) );
  AND2_X2 U5835 ( .A1(n6503), .A2(n6502), .ZN(n10657) );
  NAND2_X1 U5836 ( .A1(n4971), .A2(n4969), .ZN(n9352) );
  INV_X1 U5837 ( .A(n4970), .ZN(n4969) );
  NAND2_X1 U5838 ( .A1(n9267), .A2(n10629), .ZN(n4971) );
  OAI21_X1 U5839 ( .B1(n9268), .B2(n10648), .A(n9270), .ZN(n4970) );
  AND2_X2 U5840 ( .A1(n6503), .A2(n6861), .ZN(n10660) );
  AND2_X1 U5841 ( .A1(n6193), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10300) );
  INV_X1 U5842 ( .A(n5497), .ZN(n9374) );
  MUX2_X1 U5843 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5488), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5489) );
  NAND2_X1 U5844 ( .A1(n6074), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5576) );
  INV_X1 U5845 ( .A(n6080), .ZN(n7958) );
  XNOR2_X1 U5846 ( .A(n6068), .B(n6067), .ZN(n7890) );
  INV_X1 U5847 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6067) );
  XNOR2_X1 U5848 ( .A(n6064), .B(n5063), .ZN(n7797) );
  INV_X1 U5849 ( .A(n8592), .ZN(n8763) );
  INV_X1 U5850 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5511) );
  NOR2_X1 U5851 ( .A1(n5293), .A2(n5592), .ZN(n5578) );
  NAND2_X1 U5852 ( .A1(n5295), .A2(n5507), .ZN(n5293) );
  AND2_X1 U5853 ( .A1(n5735), .A2(n5753), .ZN(n6401) );
  XNOR2_X1 U5854 ( .A(n5639), .B(P2_IR_REG_2__SCAN_IN), .ZN(n10329) );
  NAND2_X1 U5855 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5026) );
  NAND2_X1 U5856 ( .A1(n8046), .A2(n9492), .ZN(n9410) );
  OAI21_X1 U5857 ( .B1(n8160), .B2(n4887), .A(n5393), .ZN(n8203) );
  INV_X1 U5858 ( .A(n5394), .ZN(n5393) );
  OAI21_X1 U5859 ( .B1(n5396), .B2(n4887), .A(n9391), .ZN(n5394) );
  INV_X1 U5860 ( .A(n6721), .ZN(n6722) );
  OAI22_X1 U5861 ( .A1(n6901), .A2(n6720), .B1(n7049), .B2(n10287), .ZN(n6721)
         );
  AND4_X1 U5862 ( .A1(n8061), .A2(n8060), .A3(n8059), .A4(n8058), .ZN(n9780)
         );
  NAND2_X1 U5863 ( .A1(n5030), .A2(n5383), .ZN(n9418) );
  NOR2_X1 U5864 ( .A1(n7705), .A2(n7704), .ZN(n7766) );
  NAND2_X1 U5865 ( .A1(n8141), .A2(n8140), .ZN(n9859) );
  INV_X1 U5866 ( .A(n8009), .ZN(n9908) );
  NAND2_X1 U5867 ( .A1(n9436), .A2(n5382), .ZN(n9448) );
  AND2_X1 U5868 ( .A1(n8118), .A2(n8117), .ZN(n9460) );
  NOR2_X1 U5869 ( .A1(n5041), .A2(n5039), .ZN(n5038) );
  AOI22_X1 U5870 ( .A1(n5041), .A2(n5044), .B1(n5039), .B2(n5045), .ZN(n5037)
         );
  NAND2_X1 U5871 ( .A1(n5387), .A2(n5388), .ZN(n9467) );
  NAND2_X1 U5872 ( .A1(n9410), .A2(n9411), .ZN(n5387) );
  NAND2_X1 U5873 ( .A1(n8053), .A2(n8052), .ZN(n9885) );
  INV_X1 U5874 ( .A(n5391), .ZN(n5390) );
  NAND2_X1 U5875 ( .A1(n5035), .A2(n5032), .ZN(n5389) );
  OAI21_X1 U5876 ( .B1(n7765), .B2(n5392), .A(n7764), .ZN(n5391) );
  AND4_X1 U5877 ( .A1(n7566), .A2(n7565), .A3(n7564), .A4(n7563), .ZN(n7808)
         );
  AND2_X1 U5878 ( .A1(n6745), .A2(n10392), .ZN(n9523) );
  INV_X1 U5879 ( .A(n9530), .ZN(n9485) );
  AOI22_X1 U5880 ( .A1(n9895), .A2(n8185), .B1(n8155), .B2(n9535), .ZN(n9494)
         );
  NAND2_X1 U5881 ( .A1(n7061), .A2(n7139), .ZN(n7137) );
  OR2_X1 U5882 ( .A1(n7060), .A2(n7059), .ZN(n7061) );
  NAND2_X1 U5883 ( .A1(n6745), .A2(n10393), .ZN(n9521) );
  NAND2_X1 U5884 ( .A1(n6661), .A2(n6660), .ZN(n9530) );
  NOR2_X1 U5885 ( .A1(n9781), .A2(n6648), .ZN(n4951) );
  INV_X1 U5886 ( .A(n9690), .ZN(n9533) );
  INV_X1 U5887 ( .A(n9430), .ZN(n9710) );
  INV_X1 U5888 ( .A(n9755), .ZN(n9720) );
  INV_X1 U5889 ( .A(n9754), .ZN(n9798) );
  INV_X1 U5890 ( .A(n9497), .ZN(n9799) );
  OR2_X1 U5891 ( .A1(n6787), .A2(n6688), .ZN(n6646) );
  NAND2_X1 U5892 ( .A1(n5116), .A2(n5115), .ZN(n9650) );
  INV_X1 U5893 ( .A(n9854), .ZN(n9665) );
  AND2_X1 U5894 ( .A1(n8165), .A2(n8164), .ZN(n9662) );
  AOI21_X1 U5895 ( .B1(n9622), .B2(n10392), .A(n4958), .ZN(n4957) );
  NOR2_X1 U5896 ( .A1(n9690), .A2(n9779), .ZN(n4958) );
  NAND2_X1 U5897 ( .A1(n4987), .A2(n4988), .ZN(n9683) );
  NAND2_X1 U5898 ( .A1(n9716), .A2(n4992), .ZN(n4987) );
  OAI21_X1 U5899 ( .B1(n9716), .B2(n8792), .A(n8793), .ZN(n9698) );
  OR2_X1 U5900 ( .A1(n8070), .A2(n6899), .ZN(n8073) );
  NAND2_X1 U5901 ( .A1(n7997), .A2(n7996), .ZN(n9892) );
  NOR2_X1 U5902 ( .A1(n7943), .A2(n8408), .ZN(n8807) );
  NAND2_X1 U5903 ( .A1(n7926), .A2(n7925), .ZN(n8782) );
  NAND2_X1 U5904 ( .A1(n7893), .A2(n7892), .ZN(n7899) );
  NAND2_X1 U5905 ( .A1(n7851), .A2(n7850), .ZN(n7891) );
  NAND2_X1 U5906 ( .A1(n7748), .A2(n5317), .ZN(n7802) );
  NAND2_X1 U5907 ( .A1(n7748), .A2(n7747), .ZN(n7749) );
  NAND2_X1 U5908 ( .A1(n7289), .A2(n7288), .ZN(n7318) );
  INV_X1 U5909 ( .A(n10452), .ZN(n7206) );
  OR2_X1 U5910 ( .A1(n4864), .A2(n6805), .ZN(n6809) );
  OR2_X2 U5911 ( .A1(n6668), .A2(n10504), .ZN(n9819) );
  AND2_X1 U5912 ( .A1(n9822), .A2(n10412), .ZN(n9785) );
  NAND2_X1 U5913 ( .A1(n6377), .A2(n8530), .ZN(n9967) );
  XNOR2_X1 U5914 ( .A(n8257), .B(n8256), .ZN(n9955) );
  NAND2_X1 U5915 ( .A1(n5337), .A2(n5335), .ZN(n8257) );
  NAND2_X1 U5916 ( .A1(n9949), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6404) );
  OR2_X1 U5917 ( .A1(n6405), .A2(n6162), .ZN(n6407) );
  OR2_X1 U5918 ( .A1(n5989), .A2(n5465), .ZN(n5990) );
  NAND2_X1 U5919 ( .A1(n5370), .A2(n5965), .ZN(n5985) );
  NAND2_X1 U5920 ( .A1(n5951), .A2(n5374), .ZN(n5370) );
  INV_X1 U5921 ( .A(n8264), .ZN(n8532) );
  AND2_X1 U5922 ( .A1(n7099), .A2(n7230), .ZN(n9588) );
  AND2_X1 U5923 ( .A1(n6610), .A2(n6689), .ZN(n7707) );
  NAND2_X1 U5924 ( .A1(n5324), .A2(n5557), .ZN(n5750) );
  AND2_X1 U5925 ( .A1(n6351), .A2(n6350), .ZN(n7050) );
  INV_X2 U5926 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5518) );
  NOR2_X1 U5927 ( .A1(n7687), .A2(n7686), .ZN(n10230) );
  NOR2_X1 U5928 ( .A1(n10228), .A2(n10227), .ZN(n7686) );
  NAND2_X1 U5929 ( .A1(n6114), .A2(n6113), .ZN(n6134) );
  AOI211_X1 U5930 ( .C1(n9260), .C2(n9279), .A(n9053), .B(n9052), .ZN(n9054)
         );
  NOR2_X1 U5931 ( .A1(n9302), .A2(n9244), .ZN(n9112) );
  OAI21_X1 U5932 ( .B1(n8543), .B2(n4950), .A(n4962), .ZN(P1_U3240) );
  NAND2_X1 U5933 ( .A1(n8533), .A2(n4951), .ZN(n4950) );
  AOI21_X1 U5934 ( .B1(n8545), .B2(n8546), .A(n8544), .ZN(n4962) );
  INV_X1 U5935 ( .A(n5226), .ZN(n5225) );
  OAI21_X1 U5936 ( .B1(n9841), .B2(n9804), .A(n5227), .ZN(n5226) );
  NAND2_X1 U5937 ( .A1(n4999), .A2(n4998), .ZN(P1_U3552) );
  OR2_X1 U5938 ( .A1(n10644), .A2(n6944), .ZN(n4998) );
  NAND2_X1 U5939 ( .A1(n5000), .A2(n10644), .ZN(n4999) );
  OAI211_X1 U5940 ( .C1(n9841), .C2(n10406), .A(n5103), .B(n4873), .ZN(n5000)
         );
  OAI211_X1 U5941 ( .C1(n9841), .C2(n5102), .A(n5101), .B(n5099), .ZN(P1_U3520) );
  NAND2_X1 U5942 ( .A1(n10491), .A2(n10640), .ZN(n5102) );
  INV_X1 U5943 ( .A(n5100), .ZN(n5099) );
  AND2_X1 U5944 ( .A1(n8639), .A2(n10582), .ZN(n4866) );
  AND2_X1 U5945 ( .A1(n7242), .A2(n7240), .ZN(n4867) );
  OR2_X1 U5946 ( .A1(n5446), .A2(n5442), .ZN(n4868) );
  INV_X1 U5947 ( .A(n9094), .ZN(n5332) );
  AND2_X1 U5948 ( .A1(n8636), .A2(n8633), .ZN(n4869) );
  OR2_X1 U5949 ( .A1(n5172), .A2(n5171), .ZN(n4870) );
  INV_X1 U5950 ( .A(n8624), .ZN(n5286) );
  AND2_X1 U5951 ( .A1(n9145), .A2(n9018), .ZN(n4871) );
  AND2_X1 U5952 ( .A1(n5117), .A2(n4909), .ZN(n4872) );
  AND2_X1 U5953 ( .A1(n9839), .A2(n5229), .ZN(n4873) );
  AND2_X1 U5954 ( .A1(n5067), .A2(n4910), .ZN(n4874) );
  OR2_X1 U5955 ( .A1(n6004), .A2(n6003), .ZN(n4875) );
  INV_X1 U5956 ( .A(n4986), .ZN(n4985) );
  NAND2_X1 U5957 ( .A1(n4988), .A2(n4906), .ZN(n4986) );
  AND2_X1 U5958 ( .A1(n4934), .A2(n5382), .ZN(n4876) );
  INV_X1 U5959 ( .A(n7250), .ZN(n5266) );
  INV_X1 U5960 ( .A(n9812), .ZN(n5110) );
  OR2_X1 U5961 ( .A1(n4868), .A2(n5725), .ZN(n4877) );
  NAND2_X1 U5962 ( .A1(n8548), .A2(n8547), .ZN(n9005) );
  INV_X1 U5963 ( .A(n9005), .ZN(n5333) );
  INV_X1 U5964 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U5965 ( .A1(n8195), .A2(n8194), .ZN(n9843) );
  INV_X1 U5966 ( .A(n7392), .ZN(n5131) );
  AND2_X1 U5967 ( .A1(n5110), .A2(n5232), .ZN(n4878) );
  AND2_X1 U5968 ( .A1(n8726), .A2(n5333), .ZN(n4879) );
  AND2_X1 U5969 ( .A1(n8726), .A2(n5263), .ZN(n4880) );
  AND2_X1 U5970 ( .A1(n7447), .A2(n7734), .ZN(n4881) );
  INV_X1 U5971 ( .A(n9659), .ZN(n9622) );
  AND2_X1 U5972 ( .A1(n7971), .A2(n7970), .ZN(n4882) );
  NOR2_X1 U5973 ( .A1(n5561), .A2(SI_12_), .ZN(n4883) );
  NAND2_X1 U5974 ( .A1(n5756), .A2(n5755), .ZN(n10598) );
  INV_X1 U5975 ( .A(n10598), .ZN(n4974) );
  INV_X1 U5976 ( .A(n8752), .ZN(n5199) );
  INV_X1 U5977 ( .A(n7853), .ZN(n8095) );
  INV_X1 U5978 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9369) );
  OR2_X1 U5979 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4885) );
  OAI211_X1 U5980 ( .C1(n6371), .C2(n6154), .A(n6153), .B(n6152), .ZN(n6155)
         );
  NAND2_X1 U5981 ( .A1(n10627), .A2(n8926), .ZN(n4886) );
  INV_X1 U5982 ( .A(n9027), .ZN(n5277) );
  NAND4_X1 U5983 ( .A1(n5603), .A2(n5604), .A3(n5473), .A4(n5472), .ZN(n5707)
         );
  NAND2_X1 U5984 ( .A1(n4977), .A2(n4976), .ZN(n6788) );
  OR2_X1 U5985 ( .A1(n9393), .A2(n5395), .ZN(n4887) );
  OR2_X1 U5986 ( .A1(n5008), .A2(n5223), .ZN(n6165) );
  NAND2_X1 U5987 ( .A1(n6361), .A2(n6142), .ZN(n6447) );
  NAND2_X1 U5988 ( .A1(n9473), .A2(n8105), .ZN(n9401) );
  XOR2_X1 U5989 ( .A(n7771), .B(n8197), .Z(n4888) );
  OR2_X1 U5990 ( .A1(n8607), .A2(n8727), .ZN(n4889) );
  NAND2_X1 U5991 ( .A1(n5236), .A2(n8662), .ZN(n9191) );
  INV_X1 U5992 ( .A(n8105), .ZN(n5045) );
  AND3_X1 U5993 ( .A1(n5262), .A2(n5261), .A3(n8585), .ZN(n4890) );
  AND2_X1 U5994 ( .A1(n5454), .A2(n5484), .ZN(n4891) );
  NAND4_X1 U5995 ( .A1(n5614), .A2(n5613), .A3(n5612), .A4(n5611), .ZN(n6560)
         );
  OR2_X1 U5996 ( .A1(n6883), .A2(n10452), .ZN(n4892) );
  AND4_X1 U5997 ( .A1(n9111), .A2(n9130), .A3(n9121), .A4(n8759), .ZN(n4893)
         );
  INV_X1 U5998 ( .A(n9901), .ZN(n5140) );
  AND2_X1 U5999 ( .A1(n4891), .A2(n5575), .ZN(n4894) );
  AND4_X1 U6000 ( .A1(n5466), .A2(n5220), .A3(n5398), .A4(n6349), .ZN(n6161)
         );
  OR2_X1 U6001 ( .A1(n6165), .A2(n6148), .ZN(n4895) );
  OR3_X1 U6002 ( .A1(n8673), .A2(n8672), .A3(n9178), .ZN(n4896) );
  NAND2_X1 U6003 ( .A1(n9474), .A2(n9475), .ZN(n9473) );
  INV_X1 U6004 ( .A(n5452), .ZN(n5516) );
  AND2_X1 U6005 ( .A1(n5022), .A2(n5021), .ZN(n4897) );
  OR2_X1 U6006 ( .A1(n6815), .A2(n6814), .ZN(n4898) );
  AND2_X1 U6007 ( .A1(n5210), .A2(n4892), .ZN(n4899) );
  AND2_X1 U6008 ( .A1(n5383), .A2(n5031), .ZN(n4900) );
  AND3_X1 U6009 ( .A1(n5079), .A2(n5077), .A3(n5078), .ZN(n4901) );
  AND2_X1 U6010 ( .A1(n8394), .A2(n8405), .ZN(n7901) );
  NOR2_X1 U6011 ( .A1(n8069), .A2(n5386), .ZN(n5385) );
  NAND2_X1 U6012 ( .A1(n7897), .A2(n7896), .ZN(n9912) );
  NAND2_X1 U6013 ( .A1(n8183), .A2(n8182), .ZN(n9848) );
  AND2_X1 U6014 ( .A1(n5259), .A2(n8767), .ZN(n4902) );
  AND2_X1 U6015 ( .A1(n8277), .A2(n8275), .ZN(n8498) );
  INV_X1 U6016 ( .A(n5165), .ZN(n9074) );
  INV_X1 U6017 ( .A(n5420), .ZN(n5419) );
  OAI21_X1 U6018 ( .B1(n8911), .B2(n5425), .A(n5424), .ZN(n5420) );
  OR2_X1 U6019 ( .A1(n9656), .A2(n8817), .ZN(n4903) );
  INV_X1 U6020 ( .A(n5138), .ZN(n9691) );
  NOR2_X1 U6021 ( .A1(n9699), .A2(n9866), .ZN(n5138) );
  OR2_X1 U6022 ( .A1(n9115), .A2(n8561), .ZN(n9116) );
  INV_X1 U6023 ( .A(n7239), .ZN(n5268) );
  AND2_X1 U6024 ( .A1(n5431), .A2(n6708), .ZN(n4904) );
  AND2_X1 U6025 ( .A1(n8718), .A2(n8717), .ZN(n4905) );
  NAND2_X1 U6026 ( .A1(n9866), .A2(n9710), .ZN(n4906) );
  NAND2_X1 U6027 ( .A1(n9111), .A2(n9101), .ZN(n4907) );
  INV_X1 U6028 ( .A(n9832), .ZN(n9613) );
  NAND2_X1 U6029 ( .A1(n8357), .A2(n8356), .ZN(n9832) );
  AND2_X1 U6030 ( .A1(n5378), .A2(n5380), .ZN(n4908) );
  INV_X1 U6031 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5575) );
  NAND2_X1 U6032 ( .A1(n9908), .A2(n9806), .ZN(n4909) );
  NAND2_X1 U6033 ( .A1(n5782), .A2(n5784), .ZN(n4910) );
  NAND3_X1 U6034 ( .A1(n8722), .A2(n8723), .A3(n8760), .ZN(n4911) );
  OR2_X1 U6035 ( .A1(n5687), .A2(n5686), .ZN(n4912) );
  NOR2_X1 U6036 ( .A1(n9866), .A2(n9710), .ZN(n4913) );
  NOR2_X1 U6037 ( .A1(n9331), .A2(n9215), .ZN(n4914) );
  INV_X1 U6038 ( .A(n5458), .ZN(n5183) );
  OR2_X1 U6039 ( .A1(n9435), .A2(n9438), .ZN(n9436) );
  AND2_X1 U6040 ( .A1(n8751), .A2(n8631), .ZN(n4915) );
  AND3_X1 U6041 ( .A1(n6640), .A2(n6639), .A3(n6642), .ZN(n4916) );
  AND2_X1 U6042 ( .A1(n8644), .A2(n8643), .ZN(n8737) );
  INV_X1 U6043 ( .A(n8737), .ZN(n5300) );
  NAND2_X1 U6044 ( .A1(n5222), .A2(n6361), .ZN(n4917) );
  NAND2_X1 U6045 ( .A1(n5452), .A2(n5270), .ZN(n4918) );
  OR2_X1 U6046 ( .A1(n5077), .A2(n5076), .ZN(n4919) );
  INV_X1 U6047 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6403) );
  AND2_X1 U6048 ( .A1(n8559), .A2(n8677), .ZN(n9156) );
  AND2_X1 U6049 ( .A1(n5550), .A2(n10093), .ZN(n4920) );
  AND2_X1 U6050 ( .A1(n8816), .A2(n8444), .ZN(n9675) );
  INV_X1 U6051 ( .A(n5462), .ZN(n5425) );
  INV_X1 U6052 ( .A(n10468), .ZN(n7287) );
  AND3_X1 U6053 ( .A1(n6905), .A2(n6904), .A3(n6903), .ZN(n10468) );
  NOR2_X1 U6054 ( .A1(n8068), .A2(n8067), .ZN(n4921) );
  NAND2_X1 U6055 ( .A1(n4938), .A2(n8884), .ZN(n4922) );
  NAND2_X1 U6056 ( .A1(n6044), .A2(n6043), .ZN(n9283) );
  OR2_X1 U6057 ( .A1(n8787), .A2(n9760), .ZN(n4923) );
  OR2_X1 U6058 ( .A1(n9321), .A2(n8858), .ZN(n8675) );
  NAND2_X1 U6059 ( .A1(n8715), .A2(n8716), .ZN(n9044) );
  AND2_X1 U6060 ( .A1(n5081), .A2(n5962), .ZN(n4924) );
  AND2_X1 U6061 ( .A1(n8420), .A2(n8422), .ZN(n8491) );
  INV_X1 U6062 ( .A(n8491), .ZN(n5213) );
  AND2_X1 U6063 ( .A1(n9030), .A2(n9023), .ZN(n4925) );
  INV_X1 U6064 ( .A(n6142), .ZN(n5399) );
  NOR2_X1 U6065 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n6142) );
  AND2_X1 U6066 ( .A1(n8731), .A2(n4905), .ZN(n4926) );
  AND2_X1 U6067 ( .A1(n8637), .A2(n8640), .ZN(n8752) );
  AND2_X1 U6068 ( .A1(n5140), .A2(n5141), .ZN(n4927) );
  INV_X1 U6069 ( .A(n5191), .ZN(n5190) );
  OAI21_X1 U6070 ( .B1(n5193), .B2(n5192), .A(n9094), .ZN(n5191) );
  AND2_X1 U6071 ( .A1(n7446), .A2(n4881), .ZN(n4928) );
  AND2_X1 U6072 ( .A1(n5507), .A2(n5508), .ZN(n4929) );
  AND2_X1 U6073 ( .A1(n9624), .A2(n8343), .ZN(n4930) );
  AND2_X1 U6074 ( .A1(n8447), .A2(n9638), .ZN(n5115) );
  NAND2_X1 U6075 ( .A1(n6053), .A2(n6052), .ZN(n4931) );
  INV_X1 U6076 ( .A(n5439), .ZN(n5438) );
  NAND2_X1 U6077 ( .A1(n5441), .A2(n8848), .ZN(n5439) );
  INV_X1 U6078 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5066) );
  NAND2_X1 U6079 ( .A1(n7495), .A2(n5447), .ZN(n5449) );
  AOI21_X1 U6080 ( .B1(n5449), .B2(n5748), .A(n5446), .ZN(n5443) );
  NAND2_X1 U6081 ( .A1(n7652), .A2(n5197), .ZN(n4932) );
  INV_X1 U6082 ( .A(n9648), .ZN(n5107) );
  INV_X1 U6083 ( .A(n9316), .ZN(n5163) );
  OR2_X1 U6084 ( .A1(n9925), .A2(n7754), .ZN(n8389) );
  INV_X1 U6085 ( .A(n8389), .ZN(n5207) );
  OR2_X1 U6086 ( .A1(n5516), .A2(n5455), .ZN(n4933) );
  OR2_X1 U6087 ( .A1(n8026), .A2(n8025), .ZN(n4934) );
  INV_X1 U6088 ( .A(n5937), .ZN(n5935) );
  INV_X1 U6089 ( .A(n7734), .ZN(n9542) );
  AND4_X1 U6090 ( .A1(n7279), .A2(n7278), .A3(n7277), .A4(n7276), .ZN(n7734)
         );
  NAND2_X1 U6091 ( .A1(n4895), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6156) );
  AND2_X1 U6092 ( .A1(n5365), .A2(n5567), .ZN(n4935) );
  INV_X1 U6093 ( .A(n6063), .ZN(n5423) );
  INV_X1 U6094 ( .A(n5164), .ZN(n9163) );
  INV_X1 U6095 ( .A(n5162), .ZN(n9235) );
  OR2_X1 U6096 ( .A1(n5983), .A2(SI_23_), .ZN(n4936) );
  NOR2_X1 U6097 ( .A1(n9774), .A2(n9885), .ZN(n9743) );
  NAND2_X1 U6098 ( .A1(n5374), .A2(n5984), .ZN(n4937) );
  NAND2_X1 U6099 ( .A1(n5912), .A2(n5911), .ZN(n4938) );
  AND2_X1 U6100 ( .A1(n5111), .A2(n5108), .ZN(n4939) );
  INV_X1 U6101 ( .A(n5084), .ZN(n5083) );
  NAND2_X1 U6102 ( .A1(n5434), .A2(n5433), .ZN(n5084) );
  AND2_X1 U6103 ( .A1(n5933), .A2(n10127), .ZN(n4940) );
  AND2_X1 U6104 ( .A1(n5184), .A2(n5183), .ZN(n4941) );
  INV_X1 U6105 ( .A(n9822), .ZN(n10425) );
  INV_X1 U6106 ( .A(n9822), .ZN(n9684) );
  NAND2_X1 U6107 ( .A1(n6669), .A2(n9819), .ZN(n9528) );
  AND2_X1 U6108 ( .A1(n6804), .A2(n6803), .ZN(n6818) );
  OAI21_X1 U6109 ( .B1(n10509), .B2(n5722), .A(n7172), .ZN(n7171) );
  INV_X1 U6110 ( .A(n7171), .ZN(n5069) );
  AND2_X1 U6111 ( .A1(n5148), .A2(n5147), .ZN(n4942) );
  NAND2_X1 U6112 ( .A1(n5052), .A2(n7068), .ZN(n7138) );
  NAND3_X1 U6113 ( .A1(n5452), .A2(n5453), .A3(n5454), .ZN(n4943) );
  OR2_X1 U6114 ( .A1(n6451), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4944) );
  INV_X1 U6115 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4980) );
  NAND2_X1 U6116 ( .A1(n5774), .A2(n5773), .ZN(n10620) );
  INV_X1 U6117 ( .A(n10620), .ZN(n4972) );
  NAND2_X1 U6118 ( .A1(n5065), .A2(n6966), .ZN(n6960) );
  INV_X1 U6119 ( .A(n10590), .ZN(n4975) );
  INV_X1 U6120 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n4979) );
  AND2_X1 U6121 ( .A1(n6042), .A2(n10109), .ZN(n4945) );
  INV_X1 U6122 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5063) );
  OR3_X1 U6123 ( .A1(n6198), .A2(n8999), .A3(n6197), .ZN(n4946) );
  INV_X1 U6124 ( .A(n7367), .ZN(n5130) );
  INV_X1 U6125 ( .A(n10392), .ZN(n9808) );
  AND2_X1 U6126 ( .A1(n6386), .A2(n8540), .ZN(n10392) );
  XNOR2_X1 U6127 ( .A(n6164), .B(n6163), .ZN(n6387) );
  XNOR2_X1 U6128 ( .A(n6728), .B(n8188), .ZN(n6739) );
  INV_X1 U6129 ( .A(n10547), .ZN(n5145) );
  AND2_X1 U6130 ( .A1(n8951), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4947) );
  INV_X1 U6131 ( .A(n8974), .ZN(n5015) );
  XNOR2_X1 U6132 ( .A(n6407), .B(n6406), .ZN(n8243) );
  AND2_X1 U6133 ( .A1(n5820), .A2(n5827), .ZN(n7589) );
  INV_X1 U6134 ( .A(n7589), .ZN(n5020) );
  INV_X1 U6135 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n4964) );
  INV_X1 U6136 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5019) );
  NOR3_X1 U6137 ( .A1(n6198), .A2(n8999), .A3(n6197), .ZN(n4948) );
  NAND2_X1 U6138 ( .A1(n5554), .A2(n5553), .ZN(n5728) );
  AOI21_X1 U6139 ( .B1(n5251), .B2(n5250), .A(n5249), .ZN(n5248) );
  INV_X1 U6140 ( .A(n4953), .ZN(n4952) );
  NAND2_X1 U6141 ( .A1(n8352), .A2(n8351), .ZN(n4954) );
  NAND2_X1 U6142 ( .A1(n8342), .A2(n4930), .ZN(n8347) );
  NOR2_X1 U6143 ( .A1(n8937), .A2(n6191), .ZN(n8950) );
  NAND2_X1 U6144 ( .A1(n7282), .A2(n8355), .ZN(n5319) );
  INV_X1 U6145 ( .A(n5204), .ZN(n5136) );
  AND2_X1 U6146 ( .A1(n9658), .A2(n9657), .ZN(n4960) );
  NAND2_X1 U6147 ( .A1(n9752), .A2(n9756), .ZN(n9757) );
  NAND2_X1 U6148 ( .A1(n9719), .A2(n9718), .ZN(n9717) );
  NAND2_X1 U6149 ( .A1(n5228), .A2(n5225), .ZN(P1_U3355) );
  AND2_X2 U6150 ( .A1(n8392), .A2(n8379), .ZN(n8507) );
  OAI21_X1 U6151 ( .B1(n7752), .B2(n5207), .A(n8507), .ZN(n5206) );
  NAND2_X1 U6152 ( .A1(n9658), .A2(n5115), .ZN(n5112) );
  NAND2_X2 U6153 ( .A1(n4878), .A2(n4961), .ZN(n5111) );
  OR2_X2 U6154 ( .A1(n7904), .A2(n8511), .ZN(n4961) );
  NOR2_X1 U6155 ( .A1(n8014), .A2(n8013), .ZN(n8018) );
  AOI21_X1 U6156 ( .B1(n5051), .B2(n5052), .A(n5461), .ZN(n7355) );
  INV_X1 U6157 ( .A(n7547), .ZN(n5034) );
  NAND2_X1 U6158 ( .A1(n9504), .A2(n8180), .ZN(n9390) );
  OAI21_X2 U6159 ( .B1(n5036), .B2(n5038), .A(n5037), .ZN(n9456) );
  NOR2_X1 U6160 ( .A1(n7739), .A2(n5033), .ZN(n5032) );
  AOI22_X2 U6161 ( .A1(n8370), .A2(n8522), .B1(n8369), .B2(n8480), .ZN(n8541)
         );
  NAND2_X1 U6162 ( .A1(n5091), .A2(n5093), .ZN(n5088) );
  NAND2_X1 U6163 ( .A1(n7965), .A2(n8650), .ZN(n9229) );
  NAND2_X1 U6164 ( .A1(n5235), .A2(n5234), .ZN(n9173) );
  AOI21_X1 U6165 ( .B1(n7468), .B2(n5256), .A(n5255), .ZN(n5254) );
  NAND2_X1 U6166 ( .A1(n5253), .A2(n5252), .ZN(n10585) );
  AND2_X2 U6167 ( .A1(n9196), .A2(n9202), .ZN(n9197) );
  OR2_X2 U6168 ( .A1(n9089), .A2(n9294), .ZN(n9087) );
  NAND2_X2 U6169 ( .A1(n5648), .A2(n5647), .ZN(n5650) );
  OR2_X2 U6170 ( .A1(n9254), .A2(n10525), .ZN(n7262) );
  NOR2_X2 U6171 ( .A1(n9038), .A2(n9005), .ZN(n9004) );
  NAND2_X1 U6172 ( .A1(n5165), .A2(n9067), .ZN(n9063) );
  NOR2_X2 U6173 ( .A1(n9236), .A2(n9347), .ZN(n5162) );
  INV_X1 U6174 ( .A(n5090), .ZN(n5674) );
  NOR2_X1 U6175 ( .A1(n5520), .A2(n10157), .ZN(n5521) );
  NAND2_X1 U6176 ( .A1(n9716), .A2(n4983), .ZN(n4982) );
  OAI21_X1 U6177 ( .B1(n9716), .B2(n4986), .A(n4983), .ZN(n9668) );
  NAND2_X1 U6178 ( .A1(n4994), .A2(n4996), .ZN(n4995) );
  NAND2_X1 U6179 ( .A1(n7501), .A2(n7612), .ZN(n4994) );
  NAND2_X1 U6180 ( .A1(n4995), .A2(n5313), .ZN(n7803) );
  NAND2_X1 U6181 ( .A1(n5119), .A2(n5006), .ZN(n5004) );
  NAND2_X1 U6182 ( .A1(n5466), .A2(n5398), .ZN(n5223) );
  NAND3_X1 U6183 ( .A1(n5401), .A2(n5010), .A3(n6349), .ZN(n5009) );
  NAND2_X1 U6184 ( .A1(n7295), .A2(n7374), .ZN(n7448) );
  MUX2_X1 U6185 ( .A(n6203), .B(P2_REG2_REG_1__SCAN_IN), .S(n10316), .Z(n10309) );
  NOR2_X2 U6186 ( .A1(n7549), .A2(n5034), .ZN(n7739) );
  INV_X1 U6187 ( .A(n9474), .ZN(n5036) );
  AND2_X2 U6188 ( .A1(n5050), .A2(n5046), .ZN(n5577) );
  NAND3_X1 U6189 ( .A1(n5049), .A2(n5048), .A3(n5047), .ZN(n5046) );
  NAND3_X1 U6190 ( .A1(n5518), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5050) );
  NAND2_X1 U6191 ( .A1(n7064), .A2(n7063), .ZN(n5052) );
  XNOR2_X1 U6192 ( .A(n5053), .B(n8197), .ZN(n6895) );
  XNOR2_X1 U6193 ( .A(n5062), .B(n5061), .ZN(n6576) );
  NAND2_X1 U6194 ( .A1(n6960), .A2(n5064), .ZN(n10511) );
  INV_X1 U6195 ( .A(n5068), .ZN(n5070) );
  NAND3_X1 U6196 ( .A1(n4877), .A2(n5444), .A3(n4868), .ZN(n5067) );
  NAND2_X1 U6197 ( .A1(n4877), .A2(n5444), .ZN(n5068) );
  NAND2_X1 U6198 ( .A1(n4924), .A2(n8904), .ZN(n5075) );
  NAND2_X1 U6199 ( .A1(n5085), .A2(n10547), .ZN(n5087) );
  NAND2_X1 U6200 ( .A1(n4928), .A2(n7448), .ZN(n5085) );
  NAND2_X1 U6201 ( .A1(n7448), .A2(n5086), .ZN(n7496) );
  NAND2_X1 U6202 ( .A1(n7497), .A2(n5087), .ZN(n7501) );
  OAI21_X1 U6203 ( .B1(n5460), .B2(n5093), .A(n5467), .ZN(n5092) );
  AOI21_X1 U6204 ( .B1(n5660), .B2(n5460), .A(n5093), .ZN(n5090) );
  NAND2_X1 U6205 ( .A1(n8824), .A2(n10397), .ZN(n5103) );
  NOR2_X1 U6206 ( .A1(n8820), .A2(n5096), .ZN(n5095) );
  INV_X1 U6207 ( .A(n8820), .ZN(n5097) );
  NAND2_X1 U6208 ( .A1(n8824), .A2(n5098), .ZN(n5101) );
  NAND2_X1 U6209 ( .A1(n5112), .A2(n5113), .ZN(n9625) );
  OR2_X2 U6210 ( .A1(n9658), .A2(n9657), .ZN(n5116) );
  NAND2_X1 U6211 ( .A1(n5752), .A2(n5560), .ZN(n5129) );
  NAND2_X1 U6212 ( .A1(n5752), .A2(n5125), .ZN(n5124) );
  NAND3_X1 U6213 ( .A1(n5202), .A2(n5134), .A3(n7805), .ZN(n5133) );
  NAND2_X1 U6214 ( .A1(n7918), .A2(n4927), .ZN(n5142) );
  AND2_X1 U6215 ( .A1(n9660), .A2(n5152), .ZN(n9612) );
  NAND2_X1 U6216 ( .A1(n9660), .A2(n5150), .ZN(n9611) );
  NAND2_X1 U6217 ( .A1(n9660), .A2(n5154), .ZN(n9632) );
  NAND2_X1 U6218 ( .A1(n9660), .A2(n9645), .ZN(n9640) );
  INV_X1 U6219 ( .A(n5621), .ZN(n5156) );
  INV_X2 U6220 ( .A(n6855), .ZN(n5158) );
  NOR2_X2 U6221 ( .A1(n7646), .A2(n10627), .ZN(n7975) );
  NOR2_X2 U6222 ( .A1(n4884), .A2(n9305), .ZN(n9123) );
  NOR2_X2 U6223 ( .A1(n9185), .A2(n9321), .ZN(n5164) );
  NAND3_X1 U6224 ( .A1(n5452), .A2(n4891), .A3(n5453), .ZN(n6074) );
  AND2_X2 U6225 ( .A1(n5482), .A2(n5481), .ZN(n5452) );
  NOR2_X2 U6226 ( .A1(n5480), .A2(n5479), .ZN(n5481) );
  NOR2_X2 U6227 ( .A1(n9063), .A2(n9278), .ZN(n9047) );
  NOR2_X2 U6228 ( .A1(n9087), .A2(n9289), .ZN(n5165) );
  NAND2_X1 U6229 ( .A1(n5482), .A2(n5453), .ZN(n5171) );
  AND3_X1 U6230 ( .A1(n5481), .A2(n4894), .A3(n5485), .ZN(n5169) );
  NAND3_X1 U6231 ( .A1(n5481), .A2(n4894), .A3(n5173), .ZN(n5172) );
  NAND2_X1 U6232 ( .A1(n7080), .A2(n6980), .ZN(n7233) );
  NAND2_X1 U6233 ( .A1(n7971), .A2(n5185), .ZN(n5184) );
  NAND2_X1 U6234 ( .A1(n5184), .A2(n5182), .ZN(n9210) );
  INV_X1 U6235 ( .A(n7970), .ZN(n5186) );
  NAND2_X1 U6236 ( .A1(n9110), .A2(n9023), .ZN(n5187) );
  AOI21_X1 U6237 ( .B1(n9110), .B2(n4925), .A(n5188), .ZN(n9051) );
  OAI21_X1 U6238 ( .B1(n7580), .B2(n5196), .A(n5194), .ZN(n7830) );
  INV_X1 U6239 ( .A(n7580), .ZN(n5200) );
  OR2_X1 U6240 ( .A1(n7217), .A2(n5213), .ZN(n5208) );
  AOI21_X1 U6241 ( .B1(n8491), .B2(n5212), .A(n5211), .ZN(n5210) );
  OAI21_X1 U6242 ( .B1(n7450), .B2(n5216), .A(n5214), .ZN(n7503) );
  INV_X1 U6243 ( .A(n5215), .ZN(n5214) );
  OAI21_X1 U6244 ( .B1(n5216), .B2(n7449), .A(n8381), .ZN(n5215) );
  INV_X1 U6245 ( .A(n5223), .ZN(n5222) );
  AND2_X1 U6246 ( .A1(n6141), .A2(n6632), .ZN(n5224) );
  NAND2_X1 U6247 ( .A1(n6339), .A2(n6136), .ZN(n6346) );
  NAND2_X1 U6248 ( .A1(n9625), .A2(n9624), .ZN(n9623) );
  NAND2_X1 U6249 ( .A1(n9687), .A2(n9686), .ZN(n9685) );
  NAND2_X1 U6250 ( .A1(n9706), .A2(n8814), .ZN(n9687) );
  NAND2_X1 U6251 ( .A1(n7235), .A2(n8747), .ZN(n7258) );
  NAND2_X1 U6252 ( .A1(n9304), .A2(n9022), .ZN(n9110) );
  OAI22_X1 U6253 ( .A1(n7578), .A2(n8751), .B1(n10571), .B2(n7577), .ZN(n10580) );
  NAND2_X1 U6254 ( .A1(n9210), .A2(n9015), .ZN(n9204) );
  NAND2_X1 U6255 ( .A1(n7466), .A2(n7465), .ZN(n7578) );
  NAND2_X1 U6256 ( .A1(n7830), .A2(n8754), .ZN(n7969) );
  NAND2_X1 U6257 ( .A1(n7258), .A2(n7257), .ZN(n7261) );
  NAND2_X1 U6258 ( .A1(n6978), .A2(n6977), .ZN(n7082) );
  NAND2_X1 U6259 ( .A1(n9708), .A2(n9707), .ZN(n9706) );
  NAND2_X1 U6260 ( .A1(n9676), .A2(n9675), .ZN(n9674) );
  NAND2_X1 U6261 ( .A1(n10579), .A2(n7579), .ZN(n7580) );
  NAND2_X1 U6262 ( .A1(n5483), .A2(n5066), .ZN(n5455) );
  INV_X2 U6263 ( .A(n6843), .ZN(n10436) );
  NAND2_X1 U6264 ( .A1(n6979), .A2(n6982), .ZN(n7080) );
  NAND2_X1 U6265 ( .A1(n8266), .A2(n8464), .ZN(n7377) );
  NAND2_X1 U6266 ( .A1(n9674), .A2(n8816), .ZN(n9658) );
  NAND2_X1 U6267 ( .A1(n6138), .A2(n6137), .ZN(n6140) );
  NOR2_X2 U6268 ( .A1(n7084), .A2(n7089), .ZN(n6987) );
  NOR2_X2 U6269 ( .A1(n7262), .A2(n8624), .ZN(n7343) );
  OR2_X1 U6270 ( .A1(n6899), .A2(n6719), .ZN(n6723) );
  NOR2_X2 U6271 ( .A1(n6140), .A2(n6338), .ZN(n6349) );
  NAND2_X1 U6272 ( .A1(n9208), .A2(n5237), .ZN(n5235) );
  NAND2_X1 U6273 ( .A1(n9160), .A2(n5241), .ZN(n5240) );
  OAI21_X1 U6274 ( .B1(n8563), .B2(n4907), .A(n8697), .ZN(n9095) );
  AOI21_X1 U6275 ( .B1(n4907), .B2(n8697), .A(n9094), .ZN(n5251) );
  NAND2_X1 U6276 ( .A1(n7334), .A2(n5254), .ZN(n5253) );
  NAND2_X1 U6277 ( .A1(n8579), .A2(n4879), .ZN(n5261) );
  NAND2_X1 U6278 ( .A1(n5258), .A2(n4880), .ZN(n5262) );
  NAND2_X1 U6279 ( .A1(n8578), .A2(n8760), .ZN(n5258) );
  NAND3_X1 U6280 ( .A1(n5262), .A2(n5261), .A3(n5260), .ZN(n5259) );
  INV_X1 U6281 ( .A(n9248), .ZN(n5269) );
  NAND2_X1 U6282 ( .A1(n5264), .A2(n5265), .ZN(n7251) );
  NAND2_X1 U6283 ( .A1(n9248), .A2(n4867), .ZN(n5264) );
  AND2_X1 U6284 ( .A1(n5453), .A2(n4894), .ZN(n5270) );
  OR2_X1 U6285 ( .A1(n5582), .A2(n8763), .ZN(n8587) );
  XNOR2_X2 U6286 ( .A(n5514), .B(n5513), .ZN(n5582) );
  NAND2_X1 U6287 ( .A1(n5885), .A2(n5509), .ZN(n5278) );
  AOI21_X1 U6288 ( .B1(n5279), .B2(n4926), .A(n5282), .ZN(n8766) );
  NAND3_X1 U6289 ( .A1(n5281), .A2(n5280), .A3(n9050), .ZN(n5279) );
  NAND2_X1 U6290 ( .A1(n8714), .A2(n4860), .ZN(n5280) );
  NAND2_X1 U6291 ( .A1(n8713), .A2(n8727), .ZN(n5281) );
  INV_X1 U6292 ( .A(n5592), .ZN(n5294) );
  NAND3_X1 U6293 ( .A1(n5294), .A2(n5295), .A3(n4929), .ZN(n5859) );
  OAI21_X1 U6294 ( .B1(n8630), .B2(n5298), .A(n5299), .ZN(n8648) );
  NAND2_X1 U6295 ( .A1(n8671), .A2(n8727), .ZN(n5311) );
  NAND2_X1 U6296 ( .A1(n8670), .A2(n4860), .ZN(n5310) );
  NAND4_X1 U6297 ( .A1(n5311), .A2(n5310), .A3(n5309), .A4(n4896), .ZN(n5308)
         );
  NAND2_X2 U6298 ( .A1(n5650), .A2(n5532), .ZN(n5660) );
  NAND2_X1 U6299 ( .A1(n5577), .A2(n5519), .ZN(n5312) );
  OAI21_X1 U6300 ( .B1(n5577), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n5312), .ZN(
        n5520) );
  NAND2_X1 U6301 ( .A1(n8245), .A2(n5339), .ZN(n5337) );
  NAND2_X1 U6302 ( .A1(n8245), .A2(n8244), .ZN(n5338) );
  NAND2_X1 U6303 ( .A1(n5692), .A2(n5547), .ZN(n5349) );
  OAI21_X1 U6304 ( .B1(n5692), .B2(n5346), .A(n5345), .ZN(n5591) );
  NAND2_X1 U6305 ( .A1(n5344), .A2(n5342), .ZN(n5554) );
  NAND2_X1 U6306 ( .A1(n5692), .A2(n5345), .ZN(n5344) );
  NAND2_X1 U6307 ( .A1(n5898), .A2(n5353), .ZN(n5350) );
  NAND2_X1 U6308 ( .A1(n5350), .A2(n5351), .ZN(n5938) );
  NAND2_X1 U6309 ( .A1(n5898), .A2(n5356), .ZN(n5352) );
  NAND2_X1 U6310 ( .A1(n5898), .A2(n5897), .ZN(n5917) );
  OAI21_X1 U6311 ( .B1(n6022), .B2(n6021), .A(n6025), .ZN(n6040) );
  NAND2_X1 U6312 ( .A1(n5565), .A2(n5564), .ZN(n5811) );
  NAND2_X1 U6313 ( .A1(n5936), .A2(n5369), .ZN(n5368) );
  NAND2_X1 U6314 ( .A1(n5951), .A2(n5950), .ZN(n5967) );
  NAND4_X1 U6315 ( .A1(n9484), .A2(n6803), .A3(n6820), .A4(n6804), .ZN(n6894)
         );
  NAND2_X1 U6316 ( .A1(n6951), .A2(n6898), .ZN(n7064) );
  NAND3_X1 U6317 ( .A1(n6894), .A2(n5376), .A3(n6893), .ZN(n6951) );
  AND2_X1 U6318 ( .A1(n6952), .A2(n6949), .ZN(n5376) );
  NAND2_X1 U6319 ( .A1(n6817), .A2(n6820), .ZN(n6893) );
  NAND2_X1 U6320 ( .A1(n5377), .A2(n8137), .ZN(n9427) );
  NAND2_X1 U6321 ( .A1(n9456), .A2(n9457), .ZN(n5377) );
  NAND2_X1 U6322 ( .A1(n9435), .A2(n4876), .ZN(n5379) );
  NAND2_X1 U6323 ( .A1(n8160), .A2(n5396), .ZN(n9504) );
  NAND2_X1 U6324 ( .A1(n8160), .A2(n8159), .ZN(n9502) );
  NAND3_X1 U6325 ( .A1(n5466), .A2(n6361), .A3(n6142), .ZN(n6634) );
  INV_X1 U6326 ( .A(n5863), .ZN(n5407) );
  OR2_X1 U6327 ( .A1(n6038), .A2(n6037), .ZN(n5424) );
  NAND2_X1 U6328 ( .A1(n6711), .A2(n5428), .ZN(n5426) );
  NAND3_X1 U6329 ( .A1(n5436), .A2(n5437), .A3(n5439), .ZN(n5434) );
  NAND2_X1 U6330 ( .A1(n5929), .A2(n5928), .ZN(n5441) );
  INV_X1 U6331 ( .A(n5449), .ZN(n7635) );
  XNOR2_X2 U6332 ( .A(n5456), .B(n5486), .ZN(n5497) );
  OAI211_X1 U6333 ( .C1(n9229), .C2(n8552), .A(n8657), .B(n8653), .ZN(n8553)
         );
  NOR2_X2 U6334 ( .A1(n9337), .A2(n9212), .ZN(n9196) );
  INV_X1 U6335 ( .A(n7082), .ZN(n6979) );
  NAND2_X1 U6336 ( .A1(n7260), .A2(n7259), .ZN(n7341) );
  INV_X1 U6337 ( .A(n7261), .ZN(n7260) );
  NAND2_X1 U6338 ( .A1(n5989), .A2(n5465), .ZN(n6015) );
  NAND2_X1 U6339 ( .A1(n5992), .A2(n8580), .ZN(n5994) );
  INV_X1 U6340 ( .A(n9116), .ZN(n8563) );
  INV_X1 U6341 ( .A(n4861), .ZN(n6122) );
  XNOR2_X1 U6342 ( .A(n8245), .B(n8244), .ZN(n8549) );
  INV_X1 U6343 ( .A(n8998), .ZN(n9268) );
  XNOR2_X1 U6344 ( .A(n6812), .B(n8188), .ZN(n6815) );
  AND2_X1 U6345 ( .A1(n5523), .A2(n5522), .ZN(n5615) );
  INV_X1 U6346 ( .A(n6738), .ZN(n6741) );
  OR2_X1 U6347 ( .A1(n6788), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6791) );
  NAND2_X1 U6348 ( .A1(n6746), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6792) );
  AOI22_X1 U6349 ( .A1(n6813), .A2(n8155), .B1(n10426), .B2(n8191), .ZN(n6814)
         );
  OR2_X2 U6350 ( .A1(n6813), .A2(n7225), .ZN(n8415) );
  INV_X1 U6351 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5818) );
  NAND2_X1 U6352 ( .A1(n8419), .A2(n8490), .ZN(n7217) );
  NOR2_X1 U6353 ( .A1(n5981), .A2(n5980), .ZN(n5982) );
  NAND2_X2 U6354 ( .A1(n7201), .A2(n8423), .ZN(n8266) );
  OR2_X1 U6355 ( .A1(n10650), .A2(n5582), .ZN(n6865) );
  AND2_X2 U6356 ( .A1(n6987), .A2(n6989), .ZN(n9253) );
  NAND2_X1 U6357 ( .A1(n6107), .A2(n6106), .ZN(n8239) );
  NAND2_X1 U6358 ( .A1(n9272), .A2(n10654), .ZN(n9277) );
  AOI21_X1 U6359 ( .B1(n8771), .B2(n8770), .A(n8769), .ZN(n8777) );
  NAND2_X1 U6360 ( .A1(n5470), .A2(n4902), .ZN(n8769) );
  NAND2_X1 U6361 ( .A1(n6815), .A2(n6814), .ZN(n6816) );
  OR2_X1 U6362 ( .A1(n8572), .A2(n10303), .ZN(n5625) );
  OAI21_X1 U6363 ( .B1(n9514), .B2(n9517), .A(n9515), .ZN(n9435) );
  AND2_X2 U6364 ( .A1(n7343), .A2(n10555), .ZN(n7476) );
  INV_X1 U6365 ( .A(n5979), .ZN(n5981) );
  NOR2_X1 U6366 ( .A1(n6112), .A2(n10510), .ZN(n6114) );
  INV_X8 U6367 ( .A(n5577), .ZN(n6718) );
  AND2_X1 U6368 ( .A1(n9343), .A2(n9232), .ZN(n5458) );
  OR2_X1 U6369 ( .A1(n8687), .A2(n8727), .ZN(n5459) );
  NOR2_X1 U6370 ( .A1(n7140), .A2(n7139), .ZN(n5461) );
  AND2_X1 U6371 ( .A1(n6020), .A2(n6019), .ZN(n5462) );
  AND4_X1 U6372 ( .A1(n6160), .A2(n6159), .A3(n6158), .A4(n6157), .ZN(n5463)
         );
  OR2_X1 U6373 ( .A1(n6787), .A2(n6419), .ZN(n5464) );
  AND2_X1 U6374 ( .A1(n6014), .A2(n5988), .ZN(n5465) );
  AND4_X1 U6375 ( .A1(n6146), .A2(n6145), .A3(n6144), .A4(n6143), .ZN(n5466)
         );
  AND2_X1 U6376 ( .A1(n5541), .A2(n5540), .ZN(n5467) );
  AND2_X1 U6377 ( .A1(n9014), .A2(n9013), .ZN(n5469) );
  OR3_X1 U6378 ( .A1(n8734), .A2(n8765), .A3(n8733), .ZN(n5470) );
  INV_X1 U6379 ( .A(n8735), .ZN(n8708) );
  AOI21_X1 U6380 ( .B1(n8710), .B2(n8704), .A(n8564), .ZN(n8706) );
  OAI21_X1 U6381 ( .B1(n7536), .B2(n7539), .A(n7532), .ZN(n7533) );
  INV_X1 U6382 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6157) );
  OAI21_X1 U6383 ( .B1(n7542), .B2(n7541), .A(n7540), .ZN(n7543) );
  OAI21_X1 U6384 ( .B1(P1_IR_REG_24__SCAN_IN), .B2(P1_IR_REG_25__SCAN_IN), .A(
        n6371), .ZN(n6152) );
  INV_X1 U6385 ( .A(n9881), .ZN(n8800) );
  INV_X1 U6386 ( .A(n5804), .ZN(n5494) );
  INV_X1 U6387 ( .A(n5903), .ZN(n5901) );
  INV_X1 U6388 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U6389 ( .A1(n10585), .A2(n8639), .ZN(n7572) );
  INV_X1 U6390 ( .A(n8738), .ZN(n7259) );
  INV_X1 U6391 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5485) );
  INV_X1 U6392 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7407) );
  INV_X1 U6393 ( .A(n6816), .ZN(n6817) );
  NAND2_X1 U6394 ( .A1(n7545), .A2(n7544), .ZN(n7547) );
  INV_X1 U6395 ( .A(n8033), .ZN(n6935) );
  OR2_X1 U6396 ( .A1(n8123), .A2(n8122), .ZN(n8143) );
  INV_X1 U6397 ( .A(n7907), .ZN(n6934) );
  INV_X1 U6398 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7272) );
  NAND2_X1 U6399 ( .A1(n9743), .A2(n8800), .ZN(n9744) );
  OR2_X1 U6400 ( .A1(n4864), .A2(n6885), .ZN(n6887) );
  INV_X1 U6401 ( .A(SI_29_), .ZN(n10102) );
  INV_X1 U6402 ( .A(SI_22_), .ZN(n10122) );
  INV_X1 U6403 ( .A(SI_17_), .ZN(n10021) );
  NAND2_X1 U6404 ( .A1(n5494), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5834) );
  NAND2_X1 U6405 ( .A1(n5901), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5920) );
  NAND2_X1 U6406 ( .A1(n5942), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U6407 ( .A1(n5495), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5868) );
  OR2_X1 U6408 ( .A1(n5954), .A2(n10192), .ZN(n5971) );
  INV_X1 U6409 ( .A(n6773), .ZN(n6130) );
  OR2_X1 U6410 ( .A1(n6055), .A2(n6054), .ZN(n6117) );
  OR2_X1 U6411 ( .A1(n5793), .A2(n5493), .ZN(n5804) );
  NAND2_X1 U6412 ( .A1(n8932), .A2(n10436), .ZN(n8599) );
  OR2_X1 U6413 ( .A1(n6072), .A2(n6080), .ZN(n6077) );
  INV_X1 U6414 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5484) );
  OR2_X1 U6415 ( .A1(n7408), .A2(n7407), .ZN(n7509) );
  INV_X1 U6416 ( .A(n8145), .ZN(n8166) );
  OR2_X1 U6417 ( .A1(n7853), .A2(n6420), .ZN(n6421) );
  OR2_X1 U6418 ( .A1(n7853), .A2(n10291), .ZN(n6645) );
  NAND2_X1 U6419 ( .A1(n6937), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8111) );
  OR2_X1 U6420 ( .A1(n7936), .A2(n9449), .ZN(n8033) );
  NAND2_X1 U6421 ( .A1(n6934), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7936) );
  NAND2_X1 U6422 ( .A1(n6933), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7855) );
  OR2_X1 U6423 ( .A1(n7273), .A2(n7272), .ZN(n7408) );
  INV_X1 U6424 ( .A(n9743), .ZN(n9763) );
  INV_X1 U6425 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6167) );
  NAND2_X1 U6426 ( .A1(n5879), .A2(SI_18_), .ZN(n5897) );
  NAND2_X1 U6427 ( .A1(n5566), .A2(SI_14_), .ZN(n5567) );
  OR2_X1 U6428 ( .A1(n6028), .A2(n8913), .ZN(n6055) );
  INV_X1 U6429 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10081) );
  INV_X1 U6430 ( .A(n9036), .ZN(n9273) );
  AND2_X1 U6431 ( .A1(n8658), .A2(n8657), .ZN(n8757) );
  OR2_X1 U6432 ( .A1(n5741), .A2(n5492), .ZN(n5759) );
  INV_X1 U6433 ( .A(n9261), .ZN(n7234) );
  INV_X1 U6434 ( .A(n6989), .ZN(n10475) );
  INV_X1 U6435 ( .A(n9044), .ZN(n9050) );
  OR2_X1 U6436 ( .A1(n6125), .A2(n6493), .ZN(n9216) );
  NAND2_X1 U6437 ( .A1(n6098), .A2(n8733), .ZN(n10650) );
  AND2_X1 U6438 ( .A1(n6077), .A2(n6076), .ZN(n9969) );
  XNOR2_X1 U6439 ( .A(n6890), .B(n6891), .ZN(n6820) );
  NAND2_X1 U6440 ( .A1(n7355), .A2(n7354), .ZN(n7535) );
  AOI22_X1 U6441 ( .A1(n9917), .A2(n8185), .B1(n8155), .B2(n9538), .ZN(n7876)
         );
  AND2_X1 U6442 ( .A1(n8530), .A2(n6781), .ZN(n6672) );
  OR2_X1 U6443 ( .A1(n6666), .A2(n6665), .ZN(n6669) );
  NAND4_X1 U6444 ( .A1(n6423), .A2(n5464), .A3(n6422), .A4(n6421), .ZN(n6883)
         );
  AOI21_X1 U6445 ( .B1(n6676), .B2(n8155), .A(n6654), .ZN(n6658) );
  INV_X1 U6446 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9449) );
  AND2_X1 U6447 ( .A1(n7019), .A2(n7018), .ZN(n9648) );
  AND2_X1 U6448 ( .A1(n6998), .A2(n6997), .ZN(n9659) );
  INV_X1 U6449 ( .A(n9869), .ZN(n9705) );
  INV_X1 U6450 ( .A(n7805), .ZN(n8509) );
  INV_X1 U6451 ( .A(n9781), .ZN(n10415) );
  AND2_X1 U6452 ( .A1(n10339), .A2(n8540), .ZN(n10393) );
  INV_X1 U6453 ( .A(n7901), .ZN(n8510) );
  AND2_X1 U6454 ( .A1(n6617), .A2(n6616), .ZN(n7023) );
  XNOR2_X1 U6455 ( .A(n5847), .B(n5572), .ZN(n5849) );
  INV_X1 U6456 ( .A(n5634), .ZN(n5636) );
  INV_X1 U6457 ( .A(n7890), .ZN(n6092) );
  XNOR2_X1 U6458 ( .A(n5979), .B(n5980), .ZN(n8840) );
  NOR2_X1 U6459 ( .A1(n8711), .A2(n10514), .ZN(n6131) );
  AOI21_X1 U6460 ( .B1(n7839), .B2(n5841), .A(n7844), .ZN(n7990) );
  AND2_X1 U6461 ( .A1(n6036), .A2(n6035), .ZN(n8867) );
  NAND2_X1 U6462 ( .A1(n6227), .A2(n6226), .ZN(n8968) );
  INV_X1 U6463 ( .A(n10320), .ZN(n8994) );
  NAND2_X1 U6464 ( .A1(n6869), .A2(n10609), .ZN(n10605) );
  INV_X1 U6465 ( .A(n6861), .ZN(n6502) );
  INV_X1 U6466 ( .A(n10654), .ZN(n10530) );
  NAND2_X1 U6467 ( .A1(n7474), .A2(n10435), .ZN(n10654) );
  NAND2_X1 U6468 ( .A1(n6078), .A2(n10297), .ZN(n6861) );
  AND3_X1 U6469 ( .A1(n8098), .A2(n8097), .A3(n8096), .ZN(n9742) );
  INV_X1 U6470 ( .A(n10370), .ZN(n10348) );
  INV_X1 U6471 ( .A(n10364), .ZN(n10288) );
  INV_X1 U6472 ( .A(n10376), .ZN(n10290) );
  AND2_X1 U6473 ( .A1(n8814), .A2(n8469), .ZN(n9707) );
  AND2_X1 U6474 ( .A1(n7926), .A2(n7900), .ZN(n9911) );
  INV_X1 U6475 ( .A(n9836), .ZN(n9816) );
  INV_X1 U6476 ( .A(n9635), .ZN(n9826) );
  NAND2_X1 U6477 ( .A1(n6630), .A2(n9948), .ZN(n7022) );
  INV_X1 U6478 ( .A(n10482), .ZN(n10548) );
  AND2_X1 U6479 ( .A1(n9836), .A2(n10504), .ZN(n10406) );
  OR2_X1 U6480 ( .A1(n8351), .A2(n6667), .ZN(n10504) );
  INV_X1 U6481 ( .A(n10406), .ZN(n10640) );
  AND2_X1 U6482 ( .A1(n6380), .A2(n6780), .ZN(n8530) );
  XNOR2_X1 U6483 ( .A(n6375), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6378) );
  AND2_X1 U6484 ( .A1(n6759), .A2(n7094), .ZN(n10253) );
  AND2_X1 U6485 ( .A1(n6365), .A2(n6397), .ZN(n7283) );
  INV_X1 U6486 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n7657) );
  NOR2_X1 U6487 ( .A1(n10214), .A2(n7665), .ZN(n7666) );
  NOR2_X1 U6488 ( .A1(n10226), .A2(n10225), .ZN(n7683) );
  AND2_X1 U6489 ( .A1(n6093), .A2(n6092), .ZN(n6173) );
  INV_X1 U6490 ( .A(n8711), .ZN(n9081) );
  INV_X1 U6491 ( .A(n8858), .ZN(n9175) );
  INV_X1 U6492 ( .A(n10330), .ZN(n8991) );
  NAND2_X1 U6493 ( .A1(n10605), .A2(n10599), .ZN(n10383) );
  AND2_X1 U6494 ( .A1(n6846), .A2(n6978), .ZN(n6882) );
  OR2_X1 U6495 ( .A1(n6865), .A2(n6864), .ZN(n10609) );
  INV_X1 U6496 ( .A(n10657), .ZN(n10656) );
  AND3_X1 U6497 ( .A1(n10633), .A2(n10632), .A3(n10631), .ZN(n10634) );
  INV_X1 U6498 ( .A(n10660), .ZN(n10658) );
  AND2_X1 U6499 ( .A1(n6786), .A2(n6785), .ZN(n9526) );
  INV_X1 U6500 ( .A(n9528), .ZN(n9513) );
  INV_X1 U6501 ( .A(n9647), .ZN(n9677) );
  INV_X1 U6502 ( .A(n9460), .ZN(n9721) );
  INV_X1 U6503 ( .A(n8300), .ZN(n9538) );
  NAND2_X1 U6504 ( .A1(n6652), .A2(n6380), .ZN(n10340) );
  INV_X1 U6505 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10375) );
  OR2_X1 U6506 ( .A1(P1_U3083), .A2(n6385), .ZN(n10376) );
  INV_X1 U6507 ( .A(n9785), .ZN(n9818) );
  NAND2_X1 U6508 ( .A1(n9822), .A2(n10418), .ZN(n9804) );
  OR2_X1 U6509 ( .A1(n6685), .A2(n7022), .ZN(n10642) );
  AND2_X1 U6510 ( .A1(n10457), .A2(n10456), .ZN(n10459) );
  OR2_X1 U6511 ( .A1(n6685), .A2(n6675), .ZN(n10645) );
  AND2_X1 U6512 ( .A1(n7823), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6380) );
  XNOR2_X1 U6513 ( .A(n6371), .B(P1_IR_REG_24__SCAN_IN), .ZN(n8779) );
  NOR2_X1 U6514 ( .A1(n7684), .A2(n7683), .ZN(n10228) );
  AND2_X1 U6515 ( .A1(n6173), .A2(n10300), .ZN(P2_U3966) );
  INV_X1 U6516 ( .A(n5707), .ZN(n5482) );
  NOR2_X1 U6517 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5477) );
  NAND4_X1 U6518 ( .A1(n5477), .A2(n5476), .A3(n5475), .A4(n5474), .ZN(n5480)
         );
  NAND4_X1 U6519 ( .A1(n5478), .A2(n5729), .A3(n5733), .A4(n5814), .ZN(n5479)
         );
  NAND2_X1 U6520 ( .A1(n5487), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U6521 ( .A1(n8567), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5502) );
  INV_X1 U6522 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n5490) );
  OR2_X1 U6523 ( .A1(n5865), .A2(n5490), .ZN(n5501) );
  NAND2_X1 U6524 ( .A1(n5679), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U6525 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n5491) );
  NOR2_X1 U6526 ( .A1(n5697), .A2(n5491), .ZN(n5711) );
  NAND2_X1 U6527 ( .A1(n5711), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5741) );
  NAND2_X1 U6528 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n5492) );
  NAND2_X1 U6529 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_REG3_REG_13__SCAN_IN), 
        .ZN(n5493) );
  INV_X1 U6530 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10177) );
  NAND2_X1 U6531 ( .A1(n5836), .A2(n10177), .ZN(n5496) );
  NAND2_X1 U6532 ( .A1(n5868), .A2(n5496), .ZN(n7986) );
  OR2_X1 U6533 ( .A1(n4861), .A2(n7986), .ZN(n5500) );
  NAND2_X4 U6534 ( .A1(n5498), .A2(n5497), .ZN(n8572) );
  INV_X1 U6535 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n6192) );
  OR2_X1 U6536 ( .A1(n8572), .A2(n6192), .ZN(n5499) );
  INV_X1 U6537 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5504) );
  NAND3_X1 U6538 ( .A1(n5729), .A2(n5733), .A3(n5504), .ZN(n5505) );
  NAND2_X1 U6539 ( .A1(n5514), .A2(n5513), .ZN(n5510) );
  NAND2_X1 U6540 ( .A1(n5510), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5512) );
  NAND2_X1 U6541 ( .A1(n5515), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U6542 ( .A1(n5516), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5517) );
  OR2_X2 U6543 ( .A1(n6492), .A2(n6877), .ZN(n8768) );
  NOR2_X1 U6544 ( .A1(n9217), .A2(n6870), .ZN(n5846) );
  INV_X1 U6545 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6650) );
  INV_X1 U6546 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U6547 ( .A1(n5521), .A2(SI_1_), .ZN(n5523) );
  MUX2_X1 U6548 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n6718), .Z(n5616) );
  NAND2_X1 U6549 ( .A1(n5615), .A2(n5616), .ZN(n5620) );
  NAND2_X1 U6550 ( .A1(n5620), .A2(n5523), .ZN(n5634) );
  NAND2_X1 U6551 ( .A1(n5526), .A2(SI_2_), .ZN(n5528) );
  OAI21_X1 U6552 ( .B1(n5526), .B2(SI_2_), .A(n5528), .ZN(n5635) );
  INV_X1 U6553 ( .A(n5635), .ZN(n5527) );
  NAND2_X1 U6554 ( .A1(n5634), .A2(n5527), .ZN(n5637) );
  NAND2_X1 U6555 ( .A1(n5637), .A2(n5528), .ZN(n5648) );
  MUX2_X1 U6556 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n6718), .Z(n5529) );
  NAND2_X1 U6557 ( .A1(n5529), .A2(SI_3_), .ZN(n5532) );
  INV_X1 U6558 ( .A(n5529), .ZN(n5530) );
  INV_X1 U6559 ( .A(SI_3_), .ZN(n10151) );
  NAND2_X1 U6560 ( .A1(n5530), .A2(n10151), .ZN(n5531) );
  AND2_X1 U6561 ( .A1(n5532), .A2(n5531), .ZN(n5647) );
  NAND2_X1 U6562 ( .A1(n5533), .A2(SI_4_), .ZN(n5537) );
  INV_X1 U6563 ( .A(n5533), .ZN(n5535) );
  INV_X1 U6564 ( .A(SI_4_), .ZN(n5534) );
  NAND2_X1 U6565 ( .A1(n5535), .A2(n5534), .ZN(n5536) );
  MUX2_X1 U6566 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n6718), .Z(n5538) );
  NAND2_X1 U6567 ( .A1(n5538), .A2(SI_5_), .ZN(n5541) );
  INV_X1 U6568 ( .A(n5538), .ZN(n5539) );
  NAND2_X1 U6569 ( .A1(n5539), .A2(n10034), .ZN(n5540) );
  MUX2_X1 U6570 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6718), .Z(n5542) );
  NAND2_X1 U6571 ( .A1(n5542), .A2(SI_6_), .ZN(n5544) );
  OAI21_X1 U6572 ( .B1(n5542), .B2(SI_6_), .A(n5544), .ZN(n5601) );
  INV_X1 U6573 ( .A(n5601), .ZN(n5543) );
  NAND2_X1 U6574 ( .A1(n5602), .A2(n5543), .ZN(n5545) );
  NAND2_X1 U6575 ( .A1(n5545), .A2(n5544), .ZN(n5692) );
  MUX2_X1 U6576 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6718), .Z(n5546) );
  NAND2_X1 U6577 ( .A1(n5546), .A2(SI_7_), .ZN(n5548) );
  OAI21_X1 U6578 ( .B1(n5546), .B2(SI_7_), .A(n5548), .ZN(n5691) );
  INV_X1 U6579 ( .A(n5691), .ZN(n5547) );
  MUX2_X1 U6580 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n6718), .Z(n5549) );
  XNOR2_X1 U6581 ( .A(n5549), .B(SI_8_), .ZN(n5706) );
  INV_X1 U6582 ( .A(n5549), .ZN(n5550) );
  MUX2_X1 U6583 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n6718), .Z(n5551) );
  XNOR2_X1 U6584 ( .A(n5551), .B(n10142), .ZN(n5590) );
  INV_X1 U6585 ( .A(n5551), .ZN(n5552) );
  NAND2_X1 U6586 ( .A1(n5552), .A2(n10142), .ZN(n5553) );
  MUX2_X1 U6587 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6718), .Z(n5555) );
  XNOR2_X1 U6588 ( .A(n5555), .B(n9993), .ZN(n5727) );
  INV_X1 U6589 ( .A(n5555), .ZN(n5556) );
  NAND2_X1 U6590 ( .A1(n5556), .A2(n9993), .ZN(n5557) );
  MUX2_X1 U6591 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6718), .Z(n5558) );
  NAND2_X1 U6592 ( .A1(n5558), .A2(SI_11_), .ZN(n5560) );
  OAI21_X1 U6593 ( .B1(n5558), .B2(SI_11_), .A(n5560), .ZN(n5749) );
  MUX2_X1 U6594 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6718), .Z(n5561) );
  MUX2_X1 U6595 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6718), .Z(n5562) );
  XNOR2_X1 U6596 ( .A(n5562), .B(n10134), .ZN(n5785) );
  NAND2_X1 U6597 ( .A1(n5786), .A2(n5785), .ZN(n5565) );
  INV_X1 U6598 ( .A(n5562), .ZN(n5563) );
  NAND2_X1 U6599 ( .A1(n5563), .A2(n10134), .ZN(n5564) );
  MUX2_X1 U6600 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6718), .Z(n5566) );
  OAI21_X1 U6601 ( .B1(n5566), .B2(SI_14_), .A(n5567), .ZN(n5810) );
  MUX2_X1 U6602 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6718), .Z(n5568) );
  XNOR2_X1 U6603 ( .A(n5568), .B(SI_15_), .ZN(n5825) );
  INV_X1 U6604 ( .A(n5568), .ZN(n5569) );
  NAND2_X1 U6605 ( .A1(n5569), .A2(n10097), .ZN(n5570) );
  MUX2_X1 U6606 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n6718), .Z(n5847) );
  XNOR2_X1 U6607 ( .A(n5850), .B(n5849), .ZN(n7927) );
  NAND2_X1 U6608 ( .A1(n4918), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U6609 ( .A1(n5574), .A2(n5487), .ZN(n6125) );
  XNOR2_X2 U6610 ( .A(n5576), .B(n5575), .ZN(n9383) );
  NAND2_X2 U6611 ( .A1(n6225), .A2(n8253), .ZN(n5991) );
  NAND2_X1 U6612 ( .A1(n7927), .A2(n8580), .ZN(n5581) );
  OR2_X1 U6613 ( .A1(n5578), .A2(n9369), .ZN(n5579) );
  XNOR2_X1 U6614 ( .A(n5579), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8951) );
  AOI22_X1 U6615 ( .A1(n8581), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6197), .B2(
        n8951), .ZN(n5580) );
  INV_X1 U6616 ( .A(n6098), .ZN(n8765) );
  OR2_X1 U6617 ( .A1(n5582), .A2(n8592), .ZN(n5583) );
  AND2_X4 U6618 ( .A1(n8586), .A2(n5584), .ZN(n5863) );
  XNOR2_X1 U6619 ( .A(n9343), .B(n6061), .ZN(n5843) );
  INV_X1 U6620 ( .A(n5843), .ZN(n5845) );
  NAND2_X1 U6621 ( .A1(n8567), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5589) );
  INV_X1 U6622 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5585) );
  OR2_X1 U6623 ( .A1(n5865), .A2(n5585), .ZN(n5588) );
  INV_X1 U6624 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5740) );
  XNOR2_X1 U6625 ( .A(n5741), .B(n5740), .ZN(n7486) );
  OR2_X1 U6626 ( .A1(n4861), .A2(n7486), .ZN(n5587) );
  INV_X1 U6627 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6187) );
  OR2_X1 U6628 ( .A1(n8572), .A2(n6187), .ZN(n5586) );
  NOR2_X1 U6629 ( .A1(n7331), .A2(n6870), .ZN(n5726) );
  XNOR2_X1 U6630 ( .A(n5591), .B(n5590), .ZN(n7398) );
  NAND2_X1 U6631 ( .A1(n7398), .A2(n8580), .ZN(n5594) );
  NAND2_X1 U6632 ( .A1(n5592), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5730) );
  XNOR2_X1 U6633 ( .A(n5730), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6382) );
  AOI22_X1 U6634 ( .A1(n8581), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6197), .B2(
        n6382), .ZN(n5593) );
  NAND2_X1 U6635 ( .A1(n5594), .A2(n5593), .ZN(n7493) );
  XNOR2_X1 U6636 ( .A(n7493), .B(n6061), .ZN(n5723) );
  NAND2_X1 U6637 ( .A1(n5956), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5600) );
  INV_X1 U6638 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5595) );
  XNOR2_X1 U6639 ( .A(n5697), .B(n5595), .ZN(n9257) );
  OR2_X1 U6640 ( .A1(n4861), .A2(n9257), .ZN(n5599) );
  INV_X1 U6641 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n9252) );
  OR2_X1 U6642 ( .A1(n8574), .A2(n9252), .ZN(n5598) );
  INV_X1 U6643 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5596) );
  OR2_X1 U6644 ( .A1(n5865), .A2(n5596), .ZN(n5597) );
  NAND4_X1 U6645 ( .A1(n5600), .A2(n5599), .A3(n5598), .A4(n5597), .ZN(n8929)
         );
  NAND2_X1 U6646 ( .A1(n8929), .A2(n8768), .ZN(n5688) );
  INV_X1 U6647 ( .A(n5688), .ZN(n5690) );
  XNOR2_X1 U6648 ( .A(n5602), .B(n5601), .ZN(n7051) );
  NAND2_X1 U6649 ( .A1(n7051), .A2(n8580), .ZN(n5609) );
  NAND2_X1 U6650 ( .A1(n5604), .A2(n5603), .ZN(n5661) );
  INV_X1 U6651 ( .A(n5675), .ZN(n5606) );
  INV_X1 U6652 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U6653 ( .A1(n5606), .A2(n5605), .ZN(n5693) );
  NAND2_X1 U6654 ( .A1(n5693), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5607) );
  XNOR2_X1 U6655 ( .A(n5607), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6238) );
  AOI22_X1 U6656 ( .A1(n8581), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6197), .B2(
        n6238), .ZN(n5608) );
  NAND2_X1 U6657 ( .A1(n5609), .A2(n5608), .ZN(n10492) );
  XNOR2_X1 U6658 ( .A(n10492), .B(n5863), .ZN(n5689) );
  INV_X1 U6659 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9983) );
  INV_X1 U6660 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5610) );
  INV_X1 U6661 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6203) );
  OR2_X1 U6662 ( .A1(n8574), .A2(n6203), .ZN(n5611) );
  INV_X1 U6663 ( .A(n5615), .ZN(n5618) );
  INV_X1 U6664 ( .A(n5616), .ZN(n5617) );
  NAND2_X1 U6665 ( .A1(n5618), .A2(n5617), .ZN(n5619) );
  NAND2_X1 U6666 ( .A1(n5620), .A2(n5619), .ZN(n6719) );
  NAND2_X1 U6667 ( .A1(n5651), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5622) );
  NAND2_X1 U6668 ( .A1(n6197), .A2(n10316), .ZN(n5621) );
  INV_X1 U6669 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10388) );
  INV_X1 U6670 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10303) );
  INV_X1 U6671 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10380) );
  OR2_X1 U6672 ( .A1(n8574), .A2(n10380), .ZN(n5624) );
  NAND2_X1 U6673 ( .A1(n5757), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U6674 ( .A1(n8253), .A2(SI_0_), .ZN(n5627) );
  XNOR2_X1 U6675 ( .A(n5627), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9389) );
  MUX2_X1 U6676 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9389), .S(n6225), .Z(n6568) );
  NOR2_X1 U6677 ( .A1(n5863), .A2(n6568), .ZN(n5628) );
  NAND2_X1 U6678 ( .A1(n6695), .A2(n5629), .ZN(n6577) );
  NAND2_X1 U6679 ( .A1(n5757), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5633) );
  INV_X1 U6680 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7042) );
  INV_X1 U6681 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5630) );
  INV_X1 U6682 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5631) );
  NAND2_X1 U6683 ( .A1(n5636), .A2(n5635), .ZN(n5638) );
  NAND2_X1 U6684 ( .A1(n5638), .A2(n5637), .ZN(n6806) );
  NAND2_X1 U6685 ( .A1(n5651), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U6686 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4885), .ZN(n5639) );
  NAND2_X1 U6687 ( .A1(n6197), .A2(n10329), .ZN(n5640) );
  OAI211_X1 U6688 ( .C1(n5991), .C2(n6806), .A(n5641), .B(n5640), .ZN(n6843)
         );
  NAND2_X1 U6689 ( .A1(n5757), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5646) );
  OR2_X1 U6690 ( .A1(n4861), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5645) );
  INV_X1 U6691 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5642) );
  OR2_X1 U6692 ( .A1(n8572), .A2(n5642), .ZN(n5644) );
  INV_X1 U6693 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6873) );
  OR2_X1 U6694 ( .A1(n8574), .A2(n6873), .ZN(n5643) );
  OR2_X1 U6695 ( .A1(n6976), .A2(n6870), .ZN(n5655) );
  OR2_X1 U6696 ( .A1(n5648), .A2(n5647), .ZN(n5649) );
  NAND2_X1 U6697 ( .A1(n5650), .A2(n5649), .ZN(n6795) );
  NAND2_X1 U6698 ( .A1(n5651), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5654) );
  OAI21_X1 U6699 ( .B1(P2_IR_REG_2__SCAN_IN), .B2(n4885), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5652) );
  XNOR2_X1 U6700 ( .A(n5652), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U6701 ( .A1(n6197), .A2(n6287), .ZN(n5653) );
  OAI211_X1 U6702 ( .C1(n5991), .C2(n6795), .A(n5654), .B(n5653), .ZN(n6855)
         );
  XNOR2_X1 U6703 ( .A(n6855), .B(n5863), .ZN(n5656) );
  XNOR2_X1 U6704 ( .A(n5655), .B(n5656), .ZN(n6702) );
  NAND2_X1 U6705 ( .A1(n6703), .A2(n6702), .ZN(n5659) );
  INV_X1 U6706 ( .A(n5655), .ZN(n5657) );
  NAND2_X1 U6707 ( .A1(n5657), .A2(n5656), .ZN(n5658) );
  NAND2_X1 U6708 ( .A1(n5659), .A2(n5658), .ZN(n6711) );
  XNOR2_X1 U6709 ( .A(n5660), .B(n5460), .ZN(n6884) );
  OR2_X1 U6710 ( .A1(n6884), .A2(n5991), .ZN(n5664) );
  NAND2_X1 U6711 ( .A1(n5661), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5662) );
  XNOR2_X1 U6712 ( .A(n5662), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6263) );
  AOI22_X1 U6713 ( .A1(n8581), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n6197), .B2(
        n6263), .ZN(n5663) );
  NAND2_X1 U6714 ( .A1(n5664), .A2(n5663), .ZN(n7089) );
  XNOR2_X1 U6715 ( .A(n7089), .B(n5863), .ZN(n6709) );
  NAND2_X1 U6716 ( .A1(n5956), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5673) );
  INV_X1 U6717 ( .A(n5679), .ZN(n5668) );
  INV_X1 U6718 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5666) );
  INV_X1 U6719 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U6720 ( .A1(n5666), .A2(n5665), .ZN(n5667) );
  NAND2_X1 U6721 ( .A1(n5668), .A2(n5667), .ZN(n7083) );
  OR2_X1 U6722 ( .A1(n4861), .A2(n7083), .ZN(n5672) );
  INV_X1 U6723 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5669) );
  OR2_X1 U6724 ( .A1(n5865), .A2(n5669), .ZN(n5671) );
  INV_X1 U6725 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6206) );
  OR2_X1 U6726 ( .A1(n8574), .A2(n6206), .ZN(n5670) );
  NAND4_X1 U6727 ( .A1(n5673), .A2(n5672), .A3(n5671), .A4(n5670), .ZN(n8930)
         );
  AND2_X1 U6728 ( .A1(n8930), .A2(n8768), .ZN(n6710) );
  NAND2_X1 U6729 ( .A1(n6709), .A2(n6710), .ZN(n6708) );
  OR2_X1 U6730 ( .A1(n6900), .A2(n5991), .ZN(n5678) );
  NAND2_X1 U6731 ( .A1(n5675), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5676) );
  XNOR2_X1 U6732 ( .A(n5676), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6250) );
  AOI22_X1 U6733 ( .A1(n8581), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6197), .B2(
        n6250), .ZN(n5677) );
  AND2_X2 U6734 ( .A1(n5678), .A2(n5677), .ZN(n6989) );
  XNOR2_X1 U6735 ( .A(n6989), .B(n5863), .ZN(n6968) );
  NAND2_X1 U6736 ( .A1(n5956), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5684) );
  OAI21_X1 U6737 ( .B1(n5679), .B2(P2_REG3_REG_5__SCAN_IN), .A(n5697), .ZN(
        n6988) );
  OR2_X1 U6738 ( .A1(n4861), .A2(n6988), .ZN(n5683) );
  INV_X1 U6739 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5680) );
  OR2_X1 U6740 ( .A1(n5865), .A2(n5680), .ZN(n5682) );
  INV_X1 U6741 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6986) );
  OR2_X1 U6742 ( .A1(n8574), .A2(n6986), .ZN(n5681) );
  NAND4_X1 U6743 ( .A1(n5684), .A2(n5683), .A3(n5682), .A4(n5681), .ZN(n9249)
         );
  NAND2_X1 U6744 ( .A1(n9249), .A2(n8768), .ZN(n5685) );
  XNOR2_X1 U6745 ( .A(n6968), .B(n5685), .ZN(n6769) );
  INV_X1 U6746 ( .A(n5685), .ZN(n5687) );
  INV_X1 U6747 ( .A(n6968), .ZN(n5686) );
  XNOR2_X1 U6748 ( .A(n5689), .B(n5688), .ZN(n6966) );
  XNOR2_X1 U6749 ( .A(n5692), .B(n5691), .ZN(n7128) );
  NAND2_X1 U6750 ( .A1(n7128), .A2(n8580), .ZN(n5696) );
  OAI21_X1 U6751 ( .B1(n5693), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5694) );
  XNOR2_X1 U6752 ( .A(n5694), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6274) );
  AOI22_X1 U6753 ( .A1(n8581), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6197), .B2(
        n6274), .ZN(n5695) );
  NAND2_X1 U6754 ( .A1(n5696), .A2(n5695), .ZN(n10525) );
  XNOR2_X1 U6755 ( .A(n10525), .B(n5863), .ZN(n7173) );
  NAND2_X1 U6756 ( .A1(n5738), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5703) );
  INV_X1 U6757 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6185) );
  OR2_X1 U6758 ( .A1(n8572), .A2(n6185), .ZN(n5702) );
  INV_X1 U6759 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7244) );
  OR2_X1 U6760 ( .A1(n8574), .A2(n7244), .ZN(n5701) );
  INV_X1 U6761 ( .A(n5697), .ZN(n5698) );
  AOI21_X1 U6762 ( .B1(n5698), .B2(P2_REG3_REG_6__SCAN_IN), .A(
        P2_REG3_REG_7__SCAN_IN), .ZN(n5699) );
  OR2_X1 U6763 ( .A1(n5699), .A2(n5711), .ZN(n10524) );
  OR2_X1 U6764 ( .A1(n4861), .A2(n10524), .ZN(n5700) );
  NOR2_X1 U6765 ( .A1(n7256), .A2(n6870), .ZN(n5704) );
  NAND2_X1 U6766 ( .A1(n7173), .A2(n5704), .ZN(n5705) );
  OAI21_X1 U6767 ( .B1(n7173), .B2(n5704), .A(n5705), .ZN(n10512) );
  INV_X1 U6768 ( .A(n5705), .ZN(n5722) );
  NAND2_X1 U6769 ( .A1(n7282), .A2(n8580), .ZN(n5710) );
  NAND2_X1 U6770 ( .A1(n5707), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5708) );
  XNOR2_X1 U6771 ( .A(n5708), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6359) );
  AOI22_X1 U6772 ( .A1(n8581), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6197), .B2(
        n6359), .ZN(n5709) );
  NAND2_X1 U6773 ( .A1(n5710), .A2(n5709), .ZN(n8624) );
  XNOR2_X1 U6774 ( .A(n8624), .B(n5863), .ZN(n5718) );
  NAND2_X1 U6775 ( .A1(n5956), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5717) );
  OR2_X1 U6776 ( .A1(n5711), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5712) );
  NAND2_X1 U6777 ( .A1(n5741), .A2(n5712), .ZN(n7265) );
  OR2_X1 U6778 ( .A1(n4861), .A2(n7265), .ZN(n5716) );
  INV_X1 U6779 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7266) );
  OR2_X1 U6780 ( .A1(n8574), .A2(n7266), .ZN(n5715) );
  INV_X1 U6781 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5713) );
  OR2_X1 U6782 ( .A1(n5865), .A2(n5713), .ZN(n5714) );
  NAND4_X1 U6783 ( .A1(n5717), .A2(n5716), .A3(n5715), .A4(n5714), .ZN(n8928)
         );
  AND2_X1 U6784 ( .A1(n8928), .A2(n8768), .ZN(n5719) );
  NAND2_X1 U6785 ( .A1(n5718), .A2(n5719), .ZN(n5724) );
  INV_X1 U6786 ( .A(n5718), .ZN(n7487) );
  INV_X1 U6787 ( .A(n5719), .ZN(n5720) );
  NAND2_X1 U6788 ( .A1(n7487), .A2(n5720), .ZN(n5721) );
  AND2_X1 U6789 ( .A1(n5724), .A2(n5721), .ZN(n7172) );
  XNOR2_X1 U6790 ( .A(n5723), .B(n5726), .ZN(n7489) );
  AND2_X1 U6791 ( .A1(n7489), .A2(n5724), .ZN(n5725) );
  XNOR2_X1 U6792 ( .A(n5728), .B(n5727), .ZN(n7498) );
  NAND2_X1 U6793 ( .A1(n7498), .A2(n8580), .ZN(n5737) );
  NAND2_X1 U6794 ( .A1(n5730), .A2(n5729), .ZN(n5731) );
  NAND2_X1 U6795 ( .A1(n5731), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5734) );
  INV_X1 U6796 ( .A(n5734), .ZN(n5732) );
  NAND2_X1 U6797 ( .A1(n5732), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5735) );
  NAND2_X1 U6798 ( .A1(n5734), .A2(n5733), .ZN(n5753) );
  AOI22_X1 U6799 ( .A1(n8581), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6197), .B2(
        n6401), .ZN(n5736) );
  NAND2_X1 U6800 ( .A1(n5737), .A2(n5736), .ZN(n7610) );
  XNOR2_X1 U6801 ( .A(n7610), .B(n5863), .ZN(n7633) );
  NAND2_X1 U6802 ( .A1(n5738), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5746) );
  INV_X1 U6803 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7475) );
  OR2_X1 U6804 ( .A1(n8574), .A2(n7475), .ZN(n5745) );
  INV_X1 U6805 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5739) );
  OAI21_X1 U6806 ( .B1(n5741), .B2(n5740), .A(n5739), .ZN(n5742) );
  NAND2_X1 U6807 ( .A1(n5742), .A2(n5759), .ZN(n7605) );
  OR2_X1 U6808 ( .A1(n4861), .A2(n7605), .ZN(n5744) );
  INV_X1 U6809 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6188) );
  OR2_X1 U6810 ( .A1(n8572), .A2(n6188), .ZN(n5743) );
  NOR2_X1 U6811 ( .A1(n7577), .A2(n6870), .ZN(n5747) );
  NAND2_X1 U6812 ( .A1(n7633), .A2(n5747), .ZN(n5748) );
  OAI21_X1 U6813 ( .B1(n7633), .B2(n5747), .A(n5748), .ZN(n7607) );
  INV_X1 U6814 ( .A(n5748), .ZN(n5769) );
  NAND2_X1 U6815 ( .A1(n5750), .A2(n5749), .ZN(n5751) );
  NAND2_X1 U6816 ( .A1(n5752), .A2(n5751), .ZN(n7526) );
  OR2_X1 U6817 ( .A1(n7526), .A2(n5991), .ZN(n5756) );
  NAND2_X1 U6818 ( .A1(n5753), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5754) );
  XNOR2_X1 U6819 ( .A(n5754), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6451) );
  AOI22_X1 U6820 ( .A1(n8581), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6197), .B2(
        n6451), .ZN(n5755) );
  XNOR2_X1 U6821 ( .A(n10598), .B(n5863), .ZN(n5765) );
  NAND2_X1 U6822 ( .A1(n5738), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5764) );
  INV_X1 U6823 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5758) );
  OR2_X1 U6824 ( .A1(n8574), .A2(n5758), .ZN(n5763) );
  NAND2_X1 U6825 ( .A1(n5759), .A2(n10078), .ZN(n5760) );
  NAND2_X1 U6826 ( .A1(n5793), .A2(n5760), .ZN(n10610) );
  OR2_X1 U6827 ( .A1(n4861), .A2(n10610), .ZN(n5762) );
  INV_X1 U6828 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6189) );
  OR2_X1 U6829 ( .A1(n8572), .A2(n6189), .ZN(n5761) );
  NOR2_X1 U6830 ( .A1(n7789), .A2(n6870), .ZN(n5766) );
  NAND2_X1 U6831 ( .A1(n5765), .A2(n5766), .ZN(n5780) );
  INV_X1 U6832 ( .A(n5765), .ZN(n7790) );
  INV_X1 U6833 ( .A(n5766), .ZN(n5767) );
  NAND2_X1 U6834 ( .A1(n7790), .A2(n5767), .ZN(n5768) );
  AND2_X1 U6835 ( .A1(n5780), .A2(n5768), .ZN(n7634) );
  NAND2_X1 U6836 ( .A1(n7706), .A2(n8580), .ZN(n5774) );
  OR2_X1 U6837 ( .A1(n5771), .A2(n9369), .ZN(n5772) );
  XNOR2_X1 U6838 ( .A(n5772), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7431) );
  AOI22_X1 U6839 ( .A1(n8581), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6197), .B2(
        n7431), .ZN(n5773) );
  XNOR2_X1 U6840 ( .A(n10620), .B(n6061), .ZN(n5782) );
  NAND2_X1 U6841 ( .A1(n8567), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5779) );
  INV_X1 U6842 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n5775) );
  OR2_X1 U6843 ( .A1(n5865), .A2(n5775), .ZN(n5778) );
  INV_X1 U6844 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5792) );
  XNOR2_X1 U6845 ( .A(n5793), .B(n5792), .ZN(n7788) );
  OR2_X1 U6846 ( .A1(n4861), .A2(n7788), .ZN(n5777) );
  INV_X1 U6847 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6177) );
  OR2_X1 U6848 ( .A1(n8572), .A2(n6177), .ZN(n5776) );
  NOR2_X1 U6849 ( .A1(n8224), .A2(n6870), .ZN(n5783) );
  XNOR2_X1 U6850 ( .A(n5782), .B(n5783), .ZN(n7792) );
  INV_X1 U6851 ( .A(n5782), .ZN(n8229) );
  INV_X1 U6852 ( .A(n5783), .ZN(n5784) );
  NAND2_X1 U6853 ( .A1(n7767), .A2(n8580), .ZN(n5789) );
  OR2_X1 U6854 ( .A1(n5787), .A2(n9369), .ZN(n5815) );
  XNOR2_X1 U6855 ( .A(n5815), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6692) );
  AOI22_X1 U6856 ( .A1(n8581), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6197), .B2(
        n6692), .ZN(n5788) );
  XNOR2_X1 U6857 ( .A(n10627), .B(n6061), .ZN(n5800) );
  NAND2_X1 U6858 ( .A1(n8567), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5798) );
  INV_X1 U6859 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n5790) );
  OR2_X1 U6860 ( .A1(n5865), .A2(n5790), .ZN(n5797) );
  INV_X1 U6861 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5791) );
  OAI21_X1 U6862 ( .B1(n5793), .B2(n5792), .A(n5791), .ZN(n5794) );
  NAND2_X1 U6863 ( .A1(n5804), .A2(n5794), .ZN(n8227) );
  OR2_X1 U6864 ( .A1(n4861), .A2(n8227), .ZN(n5796) );
  INV_X1 U6865 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6175) );
  OR2_X1 U6866 ( .A1(n8572), .A2(n6175), .ZN(n5795) );
  NOR2_X1 U6867 ( .A1(n8210), .A2(n6870), .ZN(n5801) );
  XNOR2_X1 U6868 ( .A(n5800), .B(n5801), .ZN(n8231) );
  NAND2_X1 U6869 ( .A1(n5799), .A2(n8231), .ZN(n8214) );
  INV_X1 U6870 ( .A(n5800), .ZN(n8215) );
  OR2_X1 U6871 ( .A1(n5801), .A2(n8215), .ZN(n5802) );
  NAND2_X1 U6872 ( .A1(n8214), .A2(n5802), .ZN(n5823) );
  NAND2_X1 U6873 ( .A1(n8567), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5809) );
  INV_X1 U6874 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n5803) );
  OR2_X1 U6875 ( .A1(n5865), .A2(n5803), .ZN(n5808) );
  INV_X1 U6876 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10089) );
  NAND2_X1 U6877 ( .A1(n5804), .A2(n10089), .ZN(n5805) );
  NAND2_X1 U6878 ( .A1(n5834), .A2(n5805), .ZN(n8213) );
  OR2_X1 U6879 ( .A1(n4861), .A2(n8213), .ZN(n5807) );
  INV_X1 U6880 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6174) );
  OR2_X1 U6881 ( .A1(n8572), .A2(n6174), .ZN(n5806) );
  INV_X1 U6882 ( .A(n7841), .ZN(n9231) );
  NAND2_X1 U6883 ( .A1(n9231), .A2(n8768), .ZN(n5824) );
  NAND2_X1 U6884 ( .A1(n5811), .A2(n5810), .ZN(n5812) );
  NAND2_X1 U6885 ( .A1(n5813), .A2(n5812), .ZN(n7849) );
  OR2_X1 U6886 ( .A1(n7849), .A2(n5991), .ZN(n5822) );
  NAND2_X1 U6887 ( .A1(n5815), .A2(n5814), .ZN(n5816) );
  NAND2_X1 U6888 ( .A1(n5816), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5819) );
  INV_X1 U6889 ( .A(n5819), .ZN(n5817) );
  NAND2_X1 U6890 ( .A1(n5817), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n5820) );
  NAND2_X1 U6891 ( .A1(n5819), .A2(n5818), .ZN(n5827) );
  AOI22_X1 U6892 ( .A1(n8581), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6197), .B2(
        n7589), .ZN(n5821) );
  XNOR2_X1 U6893 ( .A(n8221), .B(n6061), .ZN(n7842) );
  XOR2_X1 U6894 ( .A(n5824), .B(n7842), .Z(n8217) );
  NAND2_X1 U6895 ( .A1(n5823), .A2(n8217), .ZN(n7839) );
  NAND2_X1 U6896 ( .A1(n7842), .A2(n5824), .ZN(n5841) );
  XNOR2_X1 U6897 ( .A(n5826), .B(n5825), .ZN(n7894) );
  NAND2_X1 U6898 ( .A1(n7894), .A2(n8580), .ZN(n5831) );
  NAND2_X1 U6899 ( .A1(n5827), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5829) );
  XNOR2_X1 U6900 ( .A(n5829), .B(n5828), .ZN(n7003) );
  INV_X1 U6901 ( .A(n7003), .ZN(n8942) );
  AOI22_X1 U6902 ( .A1(n8581), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6197), .B2(
        n8942), .ZN(n5830) );
  XNOR2_X1 U6903 ( .A(n9347), .B(n5863), .ZN(n7987) );
  NAND2_X1 U6904 ( .A1(n5738), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5840) );
  INV_X1 U6905 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n5832) );
  OR2_X1 U6906 ( .A1(n8574), .A2(n5832), .ZN(n5839) );
  NAND2_X1 U6907 ( .A1(n5834), .A2(n5833), .ZN(n5835) );
  NAND2_X1 U6908 ( .A1(n5836), .A2(n5835), .ZN(n9237) );
  OR2_X1 U6909 ( .A1(n4861), .A2(n9237), .ZN(n5838) );
  INV_X1 U6910 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8938) );
  OR2_X1 U6911 ( .A1(n8572), .A2(n8938), .ZN(n5837) );
  NOR2_X1 U6912 ( .A1(n7983), .A2(n6870), .ZN(n5842) );
  XNOR2_X1 U6913 ( .A(n7987), .B(n5842), .ZN(n7844) );
  NOR2_X1 U6914 ( .A1(n7987), .A2(n5842), .ZN(n5844) );
  XNOR2_X1 U6915 ( .A(n5843), .B(n5846), .ZN(n7989) );
  OAI21_X1 U6916 ( .B1(n5846), .B2(n5845), .A(n7994), .ZN(n7951) );
  NOR2_X1 U6917 ( .A1(n5847), .A2(SI_16_), .ZN(n5848) );
  MUX2_X1 U6918 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n6718), .Z(n5851) );
  NAND2_X1 U6919 ( .A1(n5851), .A2(SI_17_), .ZN(n5877) );
  INV_X1 U6920 ( .A(n5851), .ZN(n5852) );
  NAND2_X1 U6921 ( .A1(n5852), .A2(n10021), .ZN(n5853) );
  NAND2_X1 U6922 ( .A1(n5877), .A2(n5853), .ZN(n5856) );
  INV_X1 U6923 ( .A(n5856), .ZN(n5854) );
  NAND2_X1 U6924 ( .A1(n5855), .A2(n5854), .ZN(n5878) );
  INV_X1 U6925 ( .A(n5855), .ZN(n5857) );
  NAND2_X1 U6926 ( .A1(n5857), .A2(n5856), .ZN(n5858) );
  NAND2_X1 U6927 ( .A1(n5878), .A2(n5858), .ZN(n8021) );
  OR2_X1 U6928 ( .A1(n8021), .A2(n5991), .ZN(n5862) );
  NAND2_X1 U6929 ( .A1(n5859), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5860) );
  XNOR2_X1 U6930 ( .A(n5860), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8974) );
  AOI22_X1 U6931 ( .A1(n8581), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6197), .B2(
        n8974), .ZN(n5861) );
  XNOR2_X1 U6932 ( .A(n9337), .B(n5863), .ZN(n5876) );
  NAND2_X1 U6933 ( .A1(n8567), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5874) );
  INV_X1 U6934 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n5864) );
  OR2_X1 U6935 ( .A1(n5865), .A2(n5864), .ZN(n5873) );
  INV_X1 U6936 ( .A(n5868), .ZN(n5866) );
  NAND2_X1 U6937 ( .A1(n5866), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5889) );
  INV_X1 U6938 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U6939 ( .A1(n5868), .A2(n5867), .ZN(n5869) );
  NAND2_X1 U6940 ( .A1(n5889), .A2(n5869), .ZN(n9220) );
  OR2_X1 U6941 ( .A1(n4861), .A2(n9220), .ZN(n5872) );
  INV_X1 U6942 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n5870) );
  OR2_X1 U6943 ( .A1(n8572), .A2(n5870), .ZN(n5871) );
  NOR2_X1 U6944 ( .A1(n8554), .A2(n6870), .ZN(n5875) );
  NOR2_X1 U6945 ( .A1(n5876), .A2(n5875), .ZN(n7947) );
  NAND2_X1 U6946 ( .A1(n5876), .A2(n5875), .ZN(n7948) );
  OAI21_X2 U6947 ( .B1(n7951), .B2(n7947), .A(n7948), .ZN(n8904) );
  MUX2_X1 U6948 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6718), .Z(n5879) );
  INV_X1 U6949 ( .A(n5879), .ZN(n5880) );
  NAND2_X1 U6950 ( .A1(n5880), .A2(n10099), .ZN(n5881) );
  OR2_X1 U6951 ( .A1(n5883), .A2(n5882), .ZN(n5884) );
  NAND2_X1 U6952 ( .A1(n5898), .A2(n5884), .ZN(n8027) );
  OR2_X1 U6953 ( .A1(n8027), .A2(n5991), .ZN(n5887) );
  XNOR2_X1 U6954 ( .A(n5885), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8986) );
  AOI22_X1 U6955 ( .A1(n8581), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6197), .B2(
        n8986), .ZN(n5886) );
  XNOR2_X1 U6956 ( .A(n9331), .B(n6061), .ZN(n5896) );
  NAND2_X1 U6957 ( .A1(n5738), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5894) );
  INV_X1 U6958 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8971) );
  OR2_X1 U6959 ( .A1(n8574), .A2(n8971), .ZN(n5893) );
  INV_X1 U6960 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U6961 ( .A1(n5889), .A2(n5888), .ZN(n5890) );
  NAND2_X1 U6962 ( .A1(n5903), .A2(n5890), .ZN(n9199) );
  OR2_X1 U6963 ( .A1(n4861), .A2(n9199), .ZN(n5892) );
  INV_X1 U6964 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8962) );
  OR2_X1 U6965 ( .A1(n8572), .A2(n8962), .ZN(n5891) );
  OR2_X1 U6966 ( .A1(n9215), .A2(n6870), .ZN(n5895) );
  NAND2_X1 U6967 ( .A1(n5896), .A2(n5895), .ZN(n8900) );
  NOR2_X1 U6968 ( .A1(n5896), .A2(n5895), .ZN(n8902) );
  MUX2_X1 U6969 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n6718), .Z(n5913) );
  XNOR2_X1 U6970 ( .A(n5913), .B(SI_19_), .ZN(n5916) );
  XNOR2_X1 U6971 ( .A(n5917), .B(n5916), .ZN(n7995) );
  NAND2_X1 U6972 ( .A1(n7995), .A2(n8580), .ZN(n5900) );
  INV_X1 U6973 ( .A(n5582), .ZN(n6496) );
  AOI22_X1 U6974 ( .A1(n8581), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6496), .B2(
        n6197), .ZN(n5899) );
  XNOR2_X1 U6975 ( .A(n9327), .B(n6061), .ZN(n5912) );
  INV_X1 U6976 ( .A(n5912), .ZN(n5910) );
  NAND2_X1 U6977 ( .A1(n5738), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5908) );
  INV_X1 U6978 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9181) );
  OR2_X1 U6979 ( .A1(n8574), .A2(n9181), .ZN(n5907) );
  INV_X1 U6980 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5902) );
  NAND2_X1 U6981 ( .A1(n5903), .A2(n5902), .ZN(n5904) );
  NAND2_X1 U6982 ( .A1(n5920), .A2(n5904), .ZN(n9180) );
  OR2_X1 U6983 ( .A1(n4861), .A2(n9180), .ZN(n5906) );
  INV_X1 U6984 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8982) );
  OR2_X1 U6985 ( .A1(n8572), .A2(n8982), .ZN(n5905) );
  OR2_X1 U6986 ( .A1(n8924), .A2(n6870), .ZN(n5911) );
  INV_X1 U6987 ( .A(n5911), .ZN(n5909) );
  NAND2_X1 U6988 ( .A1(n5910), .A2(n5909), .ZN(n8848) );
  INV_X1 U6989 ( .A(n5913), .ZN(n5914) );
  INV_X1 U6990 ( .A(SI_19_), .ZN(n9996) );
  NAND2_X1 U6991 ( .A1(n5914), .A2(n9996), .ZN(n5915) );
  MUX2_X1 U6992 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6718), .Z(n5932) );
  XNOR2_X1 U6993 ( .A(n5932), .B(n10127), .ZN(n5930) );
  NAND2_X1 U6994 ( .A1(n8050), .A2(n8580), .ZN(n5919) );
  NAND2_X1 U6995 ( .A1(n8581), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5918) );
  XNOR2_X1 U6996 ( .A(n9321), .B(n6061), .ZN(n5927) );
  INV_X1 U6997 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10187) );
  NAND2_X1 U6998 ( .A1(n5920), .A2(n10187), .ZN(n5921) );
  AND2_X1 U6999 ( .A1(n5943), .A2(n5921), .ZN(n9164) );
  NAND2_X1 U7000 ( .A1(n9164), .A2(n6122), .ZN(n5926) );
  NAND2_X1 U7001 ( .A1(n5738), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U7002 ( .A1(n8567), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5922) );
  AND2_X1 U7003 ( .A1(n5923), .A2(n5922), .ZN(n5925) );
  NAND2_X1 U7004 ( .A1(n5956), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5924) );
  NOR2_X1 U7005 ( .A1(n8858), .A2(n6870), .ZN(n5928) );
  XNOR2_X1 U7006 ( .A(n5927), .B(n5928), .ZN(n8884) );
  INV_X1 U7007 ( .A(n5927), .ZN(n5929) );
  INV_X1 U7008 ( .A(n5932), .ZN(n5933) );
  MUX2_X1 U7009 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n6718), .Z(n5934) );
  NAND2_X1 U7010 ( .A1(n5934), .A2(SI_21_), .ZN(n5950) );
  OAI21_X1 U7011 ( .B1(n5934), .B2(SI_21_), .A(n5950), .ZN(n5937) );
  NAND2_X1 U7012 ( .A1(n5938), .A2(n5937), .ZN(n5939) );
  NAND2_X1 U7013 ( .A1(n5951), .A2(n5939), .ZN(n8070) );
  OR2_X1 U7014 ( .A1(n8070), .A2(n5991), .ZN(n5941) );
  NAND2_X1 U7015 ( .A1(n8581), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5940) );
  XNOR2_X1 U7016 ( .A(n9316), .B(n6061), .ZN(n5949) );
  INV_X1 U7017 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10172) );
  NAND2_X1 U7018 ( .A1(n5943), .A2(n10172), .ZN(n5944) );
  NAND2_X1 U7019 ( .A1(n5954), .A2(n5944), .ZN(n9150) );
  OR2_X1 U7020 ( .A1(n9150), .A2(n4861), .ZN(n5947) );
  AOI22_X1 U7021 ( .A1(n8567), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n5738), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U7022 ( .A1(n5956), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7023 ( .A1(n9161), .A2(n8768), .ZN(n5948) );
  XNOR2_X1 U7024 ( .A(n5949), .B(n5948), .ZN(n8856) );
  MUX2_X1 U7025 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n6718), .Z(n5963) );
  XNOR2_X1 U7026 ( .A(n5963), .B(SI_22_), .ZN(n5966) );
  XNOR2_X1 U7027 ( .A(n5967), .B(n5966), .ZN(n8088) );
  NAND2_X1 U7028 ( .A1(n8088), .A2(n8580), .ZN(n5953) );
  NAND2_X1 U7029 ( .A1(n8581), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5952) );
  XNOR2_X1 U7030 ( .A(n9311), .B(n6061), .ZN(n5961) );
  INV_X1 U7031 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10192) );
  NAND2_X1 U7032 ( .A1(n5954), .A2(n10192), .ZN(n5955) );
  NAND2_X1 U7033 ( .A1(n5971), .A2(n5955), .ZN(n9133) );
  OR2_X1 U7034 ( .A1(n9133), .A2(n4861), .ZN(n5959) );
  AOI22_X1 U7035 ( .A1(n8567), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n5738), .B2(
        P2_REG0_REG_22__SCAN_IN), .ZN(n5958) );
  NAND2_X1 U7036 ( .A1(n5956), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5957) );
  NAND2_X1 U7037 ( .A1(n9146), .A2(n8768), .ZN(n5960) );
  NAND2_X1 U7038 ( .A1(n5961), .A2(n5960), .ZN(n5962) );
  OAI21_X1 U7039 ( .B1(n5961), .B2(n5960), .A(n5962), .ZN(n8892) );
  INV_X1 U7040 ( .A(n5963), .ZN(n5964) );
  NAND2_X1 U7041 ( .A1(n5964), .A2(n10122), .ZN(n5965) );
  MUX2_X1 U7042 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n6718), .Z(n5983) );
  INV_X1 U7043 ( .A(SI_23_), .ZN(n10118) );
  XNOR2_X1 U7044 ( .A(n5983), .B(n10118), .ZN(n5984) );
  XNOR2_X1 U7045 ( .A(n5985), .B(n5984), .ZN(n8106) );
  NAND2_X1 U7046 ( .A1(n8106), .A2(n8580), .ZN(n5969) );
  NAND2_X1 U7047 ( .A1(n8581), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5968) );
  XNOR2_X1 U7048 ( .A(n9305), .B(n6061), .ZN(n5980) );
  INV_X1 U7049 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10166) );
  NAND2_X1 U7050 ( .A1(n5971), .A2(n10166), .ZN(n5972) );
  NAND2_X1 U7051 ( .A1(n5995), .A2(n5972), .ZN(n9126) );
  OR2_X1 U7052 ( .A1(n9126), .A2(n4861), .ZN(n5978) );
  INV_X1 U7053 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U7054 ( .A1(n8567), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5974) );
  NAND2_X1 U7055 ( .A1(n5738), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5973) );
  OAI211_X1 U7056 ( .C1(n5975), .C2(n8572), .A(n5974), .B(n5973), .ZN(n5976)
         );
  INV_X1 U7057 ( .A(n5976), .ZN(n5977) );
  NOR2_X1 U7058 ( .A1(n8894), .A2(n6870), .ZN(n8839) );
  MUX2_X1 U7059 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n6718), .Z(n5986) );
  NAND2_X1 U7060 ( .A1(n5986), .A2(SI_24_), .ZN(n6014) );
  INV_X1 U7061 ( .A(n5986), .ZN(n5987) );
  INV_X1 U7062 ( .A(SI_24_), .ZN(n10116) );
  NAND2_X1 U7063 ( .A1(n5987), .A2(n10116), .ZN(n5988) );
  NAND2_X1 U7064 ( .A1(n6015), .A2(n5990), .ZN(n8778) );
  INV_X1 U7065 ( .A(n8778), .ZN(n5992) );
  NAND2_X1 U7066 ( .A1(n8581), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5993) );
  XNOR2_X1 U7067 ( .A(n9298), .B(n6061), .ZN(n6003) );
  NAND2_X1 U7068 ( .A1(n5995), .A2(n10081), .ZN(n5996) );
  AND2_X1 U7069 ( .A1(n6006), .A2(n5996), .ZN(n9105) );
  NAND2_X1 U7070 ( .A1(n9105), .A2(n6122), .ZN(n6002) );
  INV_X1 U7071 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n5999) );
  NAND2_X1 U7072 ( .A1(n8567), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U7073 ( .A1(n5738), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5997) );
  OAI211_X1 U7074 ( .C1(n5999), .C2(n8572), .A(n5998), .B(n5997), .ZN(n6000)
         );
  INV_X1 U7075 ( .A(n6000), .ZN(n6001) );
  NAND2_X1 U7076 ( .A1(n9118), .A2(n8768), .ZN(n8874) );
  INV_X1 U7077 ( .A(n6006), .ZN(n6005) );
  NAND2_X1 U7078 ( .A1(n6005), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6028) );
  INV_X1 U7079 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10083) );
  NAND2_X1 U7080 ( .A1(n6006), .A2(n10083), .ZN(n6007) );
  NAND2_X1 U7081 ( .A1(n6028), .A2(n6007), .ZN(n9090) );
  OR2_X1 U7082 ( .A1(n9090), .A2(n4861), .ZN(n6013) );
  INV_X1 U7083 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U7084 ( .A1(n8567), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6009) );
  NAND2_X1 U7085 ( .A1(n5738), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6008) );
  OAI211_X1 U7086 ( .C1(n6010), .C2(n8572), .A(n6009), .B(n6008), .ZN(n6011)
         );
  INV_X1 U7087 ( .A(n6011), .ZN(n6012) );
  NAND2_X1 U7088 ( .A1(n9103), .A2(n8768), .ZN(n6018) );
  MUX2_X1 U7089 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n6718), .Z(n6023) );
  XNOR2_X1 U7090 ( .A(n6023), .B(SI_25_), .ZN(n6021) );
  XNOR2_X1 U7091 ( .A(n6022), .B(n6021), .ZN(n8138) );
  NAND2_X1 U7092 ( .A1(n8581), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6016) );
  XNOR2_X1 U7093 ( .A(n9294), .B(n6061), .ZN(n6017) );
  XOR2_X1 U7094 ( .A(n6018), .B(n6017), .Z(n8866) );
  INV_X1 U7095 ( .A(n6017), .ZN(n6020) );
  INV_X1 U7096 ( .A(n6018), .ZN(n6019) );
  INV_X1 U7097 ( .A(n6023), .ZN(n6024) );
  INV_X1 U7098 ( .A(SI_25_), .ZN(n10113) );
  NAND2_X1 U7099 ( .A1(n6024), .A2(n10113), .ZN(n6025) );
  MUX2_X1 U7100 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .S(n6718), .Z(n6041) );
  XNOR2_X1 U7101 ( .A(n6041), .B(n10109), .ZN(n6039) );
  XNOR2_X1 U7102 ( .A(n6040), .B(n6039), .ZN(n9384) );
  NAND2_X1 U7103 ( .A1(n9384), .A2(n8580), .ZN(n6027) );
  NAND2_X1 U7104 ( .A1(n8581), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6026) );
  XNOR2_X1 U7105 ( .A(n9289), .B(n6061), .ZN(n6038) );
  INV_X1 U7106 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8913) );
  NAND2_X1 U7107 ( .A1(n6028), .A2(n8913), .ZN(n6029) );
  NAND2_X1 U7108 ( .A1(n6055), .A2(n6029), .ZN(n9075) );
  OR2_X1 U7109 ( .A1(n9075), .A2(n4861), .ZN(n6036) );
  INV_X1 U7110 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n6033) );
  NAND2_X1 U7111 ( .A1(n8567), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6032) );
  NAND2_X1 U7112 ( .A1(n5738), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6031) );
  OAI211_X1 U7113 ( .C1(n6033), .C2(n8572), .A(n6032), .B(n6031), .ZN(n6034)
         );
  INV_X1 U7114 ( .A(n6034), .ZN(n6035) );
  NAND2_X1 U7115 ( .A1(n9096), .A2(n8768), .ZN(n6037) );
  XNOR2_X1 U7116 ( .A(n6038), .B(n6037), .ZN(n8911) );
  INV_X1 U7117 ( .A(n6041), .ZN(n6042) );
  MUX2_X1 U7118 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n6718), .Z(n6102) );
  XNOR2_X1 U7119 ( .A(n6102), .B(n10000), .ZN(n6100) );
  NAND2_X1 U7120 ( .A1(n9382), .A2(n8580), .ZN(n6044) );
  NAND2_X1 U7121 ( .A1(n8581), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6043) );
  XNOR2_X1 U7122 ( .A(n9283), .B(n6061), .ZN(n6051) );
  XNOR2_X1 U7123 ( .A(n6055), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n9064) );
  NAND2_X1 U7124 ( .A1(n9064), .A2(n6122), .ZN(n6050) );
  INV_X1 U7125 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6047) );
  NAND2_X1 U7126 ( .A1(n8567), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6046) );
  NAND2_X1 U7127 ( .A1(n5738), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6045) );
  OAI211_X1 U7128 ( .C1(n6047), .C2(n8572), .A(n6046), .B(n6045), .ZN(n6048)
         );
  INV_X1 U7129 ( .A(n6048), .ZN(n6049) );
  NOR2_X1 U7130 ( .A1(n8711), .A2(n6870), .ZN(n6052) );
  XNOR2_X1 U7131 ( .A(n6051), .B(n6052), .ZN(n8832) );
  INV_X1 U7132 ( .A(n6051), .ZN(n6053) );
  INV_X1 U7133 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9986) );
  INV_X1 U7134 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6126) );
  OAI21_X1 U7135 ( .B1(n6055), .B2(n9986), .A(n6126), .ZN(n6056) );
  NAND2_X1 U7136 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n6054) );
  INV_X1 U7137 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U7138 ( .A1(n8567), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7139 ( .A1(n5738), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6057) );
  OAI211_X1 U7140 ( .C1(n6059), .C2(n8572), .A(n6058), .B(n6057), .ZN(n6060)
         );
  NOR2_X1 U7141 ( .A1(n8923), .A2(n6870), .ZN(n6062) );
  MUX2_X1 U7142 ( .A(n8923), .B(n6062), .S(n6061), .Z(n6063) );
  NAND2_X1 U7143 ( .A1(n6064), .A2(n5063), .ZN(n6065) );
  NAND2_X1 U7144 ( .A1(n6095), .A2(n6094), .ZN(n6066) );
  NAND2_X1 U7145 ( .A1(n6066), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6068) );
  INV_X1 U7146 ( .A(P2_B_REG_SCAN_IN), .ZN(n6069) );
  AOI22_X1 U7147 ( .A1(P2_B_REG_SCAN_IN), .A2(n7890), .B1(n6092), .B2(n6069), 
        .ZN(n6072) );
  NAND2_X1 U7148 ( .A1(n4933), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6070) );
  MUX2_X1 U7149 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6070), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6071) );
  AND2_X1 U7150 ( .A1(n6071), .A2(n4943), .ZN(n6080) );
  NAND2_X1 U7151 ( .A1(n4943), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6073) );
  MUX2_X1 U7152 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6073), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6075) );
  NAND2_X1 U7153 ( .A1(n6075), .A2(n6074), .ZN(n9387) );
  INV_X1 U7154 ( .A(n9387), .ZN(n6076) );
  INV_X1 U7155 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10298) );
  NAND2_X1 U7156 ( .A1(n9969), .A2(n10298), .ZN(n6078) );
  NAND2_X1 U7157 ( .A1(n7890), .A2(n9387), .ZN(n10297) );
  INV_X1 U7158 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U7159 ( .A1(n9969), .A2(n6079), .ZN(n6081) );
  NAND2_X1 U7160 ( .A1(n7958), .A2(n9387), .ZN(n9968) );
  NAND2_X1 U7161 ( .A1(n6081), .A2(n9968), .ZN(n6490) );
  INV_X1 U7162 ( .A(n6490), .ZN(n6863) );
  NOR4_X1 U7163 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6085) );
  NOR4_X1 U7164 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6084) );
  NOR4_X1 U7165 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6083) );
  NOR4_X1 U7166 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n6082) );
  NAND4_X1 U7167 ( .A1(n6085), .A2(n6084), .A3(n6083), .A4(n6082), .ZN(n6091)
         );
  NOR2_X1 U7168 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .ZN(
        n6089) );
  NOR4_X1 U7169 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n6088) );
  NOR4_X1 U7170 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6087) );
  NOR4_X1 U7171 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6086) );
  NAND4_X1 U7172 ( .A1(n6089), .A2(n6088), .A3(n6087), .A4(n6086), .ZN(n6090)
         );
  OAI21_X1 U7173 ( .B1(n6091), .B2(n6090), .A(n9969), .ZN(n6489) );
  NAND3_X1 U7174 ( .A1(n6502), .A2(n6863), .A3(n6489), .ZN(n6124) );
  NOR2_X1 U7175 ( .A1(n7958), .A2(n9387), .ZN(n6093) );
  XNOR2_X1 U7176 ( .A(n6095), .B(n6094), .ZN(n6193) );
  INV_X1 U7177 ( .A(n10300), .ZN(n6096) );
  NOR2_X1 U7178 ( .A1(n6864), .A2(n6129), .ZN(n6196) );
  NAND2_X1 U7179 ( .A1(n10648), .A2(n6196), .ZN(n6097) );
  OR2_X2 U7180 ( .A1(n6124), .A2(n6097), .ZN(n10510) );
  NAND2_X1 U7181 ( .A1(n6124), .A2(n6865), .ZN(n6115) );
  INV_X1 U7182 ( .A(n6864), .ZN(n9971) );
  AND2_X1 U7183 ( .A1(n6115), .A2(n9971), .ZN(n6579) );
  AOI21_X1 U7184 ( .B1(n6112), .B2(n8873), .A(n8918), .ZN(n6099) );
  INV_X1 U7185 ( .A(n6099), .ZN(n6111) );
  NAND2_X1 U7186 ( .A1(n6101), .A2(n6100), .ZN(n6105) );
  INV_X1 U7187 ( .A(n6102), .ZN(n6103) );
  NAND2_X1 U7188 ( .A1(n6103), .A2(n10000), .ZN(n6104) );
  NAND2_X1 U7189 ( .A1(n6105), .A2(n6104), .ZN(n6107) );
  MUX2_X1 U7190 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6718), .Z(n8236) );
  INV_X1 U7191 ( .A(SI_28_), .ZN(n10104) );
  XNOR2_X1 U7192 ( .A(n8236), .B(n10104), .ZN(n6106) );
  NAND2_X1 U7193 ( .A1(n8826), .A2(n8580), .ZN(n6110) );
  NAND2_X1 U7194 ( .A1(n8581), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U7195 ( .A1(n6111), .A2(n9278), .ZN(n6135) );
  INV_X1 U7196 ( .A(n9278), .ZN(n6113) );
  INV_X1 U7197 ( .A(n6173), .ZN(n6194) );
  NAND2_X1 U7198 ( .A1(n6492), .A2(n6129), .ZN(n6578) );
  NAND4_X1 U7199 ( .A1(n6115), .A2(n6194), .A3(n6193), .A4(n6578), .ZN(n6116)
         );
  INV_X1 U7200 ( .A(n10523), .ZN(n8886) );
  INV_X1 U7201 ( .A(n6117), .ZN(n9039) );
  INV_X1 U7202 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U7203 ( .A1(n8567), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U7204 ( .A1(n5738), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6118) );
  OAI211_X1 U7205 ( .C1(n6120), .C2(n8572), .A(n6119), .B(n6118), .ZN(n6121)
         );
  AOI21_X1 U7206 ( .B1(n9039), .B2(n6122), .A(n6121), .ZN(n8922) );
  INV_X1 U7207 ( .A(n6492), .ZN(n8772) );
  NAND2_X1 U7208 ( .A1(n8772), .A2(n9971), .ZN(n6123) );
  OR2_X1 U7209 ( .A1(n6124), .A2(n6123), .ZN(n6773) );
  NAND2_X1 U7210 ( .A1(n6130), .A2(n10587), .ZN(n10517) );
  OAI22_X1 U7211 ( .A1(n8922), .A2(n10517), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6126), .ZN(n6127) );
  AOI21_X1 U7212 ( .B1(n9048), .B2(n8886), .A(n6127), .ZN(n6128) );
  INV_X1 U7213 ( .A(n6128), .ZN(n6132) );
  INV_X1 U7214 ( .A(n6129), .ZN(n6493) );
  NAND2_X1 U7215 ( .A1(n6130), .A2(n9230), .ZN(n10514) );
  NOR2_X1 U7216 ( .A1(n6132), .A2(n6131), .ZN(n6133) );
  NAND3_X1 U7217 ( .A1(n6135), .A2(n6134), .A3(n6133), .ZN(P2_U3222) );
  INV_X1 U7218 ( .A(n6346), .ZN(n6138) );
  NAND2_X1 U7219 ( .A1(n6332), .A2(n6139), .ZN(n6338) );
  NAND2_X1 U7220 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n6149) );
  NAND2_X1 U7221 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .ZN(n6369) );
  AOI21_X1 U7222 ( .B1(n6158), .B2(n6369), .A(n6160), .ZN(n6154) );
  INV_X1 U7223 ( .A(n6369), .ZN(n6151) );
  XNOR2_X1 U7224 ( .A(P1_IR_REG_31__SCAN_IN), .B(P1_IR_REG_26__SCAN_IN), .ZN(
        n6150) );
  AOI21_X1 U7225 ( .B1(P1_IR_REG_25__SCAN_IN), .B2(n6151), .A(n6150), .ZN(
        n6153) );
  INV_X1 U7226 ( .A(n6155), .ZN(n6652) );
  INV_X1 U7227 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U7228 ( .A1(n6168), .A2(n6167), .ZN(n6170) );
  NAND2_X1 U7229 ( .A1(n6170), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6166) );
  NAND2_X1 U7230 ( .A1(n8264), .A2(n8483), .ZN(n6678) );
  NAND2_X1 U7231 ( .A1(n6678), .A2(n6780), .ZN(n6171) );
  NAND2_X1 U7232 ( .A1(n6171), .A2(n7823), .ZN(n6465) );
  NAND2_X1 U7233 ( .A1(n7049), .A2(n6465), .ZN(n6172) );
  NAND2_X1 U7234 ( .A1(n6172), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X2 U7235 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  MUX2_X1 U7236 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n6174), .S(n7589), .Z(n7592)
         );
  INV_X1 U7237 ( .A(n6692), .ZN(n7444) );
  NOR2_X1 U7238 ( .A1(n7444), .A2(n6175), .ZN(n6176) );
  AOI21_X1 U7239 ( .B1(n6175), .B2(n7444), .A(n6176), .ZN(n7435) );
  INV_X1 U7240 ( .A(n7431), .ZN(n6612) );
  NOR2_X1 U7241 ( .A1(n6612), .A2(n6177), .ZN(n6178) );
  AOI21_X1 U7242 ( .B1(n6177), .B2(n6612), .A(n6178), .ZN(n7423) );
  INV_X1 U7243 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10301) );
  INV_X1 U7244 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6179) );
  MUX2_X1 U7245 ( .A(n6179), .B(P2_REG1_REG_1__SCAN_IN), .S(n10316), .Z(n10312) );
  NOR3_X1 U7246 ( .A1(n10301), .A2(n10303), .A3(n10312), .ZN(n10311) );
  AOI21_X1 U7247 ( .B1(n10316), .B2(P2_REG1_REG_1__SCAN_IN), .A(n10311), .ZN(
        n10326) );
  NAND2_X1 U7248 ( .A1(n10329), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6180) );
  OAI21_X1 U7249 ( .B1(n10329), .B2(P2_REG1_REG_2__SCAN_IN), .A(n6180), .ZN(
        n10325) );
  NOR2_X1 U7250 ( .A1(n10326), .A2(n10325), .ZN(n10324) );
  AOI21_X1 U7251 ( .B1(n10329), .B2(P2_REG1_REG_2__SCAN_IN), .A(n10324), .ZN(
        n6283) );
  NAND2_X1 U7252 ( .A1(n6287), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6181) );
  OAI21_X1 U7253 ( .B1(n6287), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6181), .ZN(
        n6282) );
  NOR2_X1 U7254 ( .A1(n6283), .A2(n6282), .ZN(n6281) );
  INV_X1 U7255 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6182) );
  MUX2_X1 U7256 ( .A(n6182), .B(P2_REG1_REG_4__SCAN_IN), .S(n6263), .Z(n6258)
         );
  NOR2_X1 U7257 ( .A1(n6259), .A2(n6258), .ZN(n6257) );
  INV_X1 U7258 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6183) );
  MUX2_X1 U7259 ( .A(n6183), .B(P2_REG1_REG_5__SCAN_IN), .S(n6250), .Z(n6245)
         );
  NOR2_X1 U7260 ( .A1(n6246), .A2(n6245), .ZN(n6244) );
  AOI21_X1 U7261 ( .B1(n6250), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6244), .ZN(
        n6234) );
  INV_X1 U7262 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6184) );
  MUX2_X1 U7263 ( .A(n6184), .B(P2_REG1_REG_6__SCAN_IN), .S(n6238), .Z(n6233)
         );
  NOR2_X1 U7264 ( .A1(n6234), .A2(n6233), .ZN(n6232) );
  MUX2_X1 U7265 ( .A(n6185), .B(P2_REG1_REG_7__SCAN_IN), .S(n6274), .Z(n6270)
         );
  NOR2_X1 U7266 ( .A1(n6271), .A2(n6270), .ZN(n6269) );
  AOI21_X1 U7267 ( .B1(n6274), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6269), .ZN(
        n6295) );
  INV_X1 U7268 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6186) );
  MUX2_X1 U7269 ( .A(n6186), .B(P2_REG1_REG_8__SCAN_IN), .S(n6359), .Z(n6294)
         );
  NOR2_X1 U7270 ( .A1(n6295), .A2(n6294), .ZN(n6293) );
  MUX2_X1 U7271 ( .A(n6187), .B(P2_REG1_REG_9__SCAN_IN), .S(n6382), .Z(n6306)
         );
  NOR2_X1 U7272 ( .A1(n6307), .A2(n6306), .ZN(n6305) );
  AOI21_X1 U7273 ( .B1(n6382), .B2(P2_REG1_REG_9__SCAN_IN), .A(n6305), .ZN(
        n6319) );
  MUX2_X1 U7274 ( .A(n6188), .B(P2_REG1_REG_10__SCAN_IN), .S(n6401), .Z(n6318)
         );
  NOR2_X1 U7275 ( .A1(n6319), .A2(n6318), .ZN(n6317) );
  MUX2_X1 U7276 ( .A(n6189), .B(P2_REG1_REG_11__SCAN_IN), .S(n6451), .Z(n7164)
         );
  NOR2_X1 U7277 ( .A1(n7165), .A2(n7164), .ZN(n7163) );
  AOI21_X1 U7278 ( .B1(n6451), .B2(P2_REG1_REG_11__SCAN_IN), .A(n7163), .ZN(
        n7422) );
  NAND2_X1 U7279 ( .A1(n7423), .A2(n7422), .ZN(n7421) );
  OAI21_X1 U7280 ( .B1(n7431), .B2(P2_REG1_REG_12__SCAN_IN), .A(n7421), .ZN(
        n7434) );
  NAND2_X1 U7281 ( .A1(n7592), .A2(n7591), .ZN(n7590) );
  NOR2_X1 U7282 ( .A1(n7003), .A2(n6190), .ZN(n6191) );
  XNOR2_X1 U7283 ( .A(n7003), .B(n6190), .ZN(n8939) );
  NOR2_X1 U7284 ( .A1(n8938), .A2(n8939), .ZN(n8937) );
  XNOR2_X1 U7285 ( .A(n8951), .B(n6192), .ZN(n8949) );
  NAND2_X1 U7286 ( .A1(n8950), .A2(n8949), .ZN(n8948) );
  OAI21_X1 U7287 ( .B1(n8951), .B2(P2_REG1_REG_16__SCAN_IN), .A(n8948), .ZN(
        n6200) );
  XNOR2_X1 U7288 ( .A(n8974), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n6199) );
  NOR2_X1 U7289 ( .A1(n6199), .A2(n6200), .ZN(n8963) );
  OR2_X1 U7290 ( .A1(n6193), .A2(P2_U3152), .ZN(n8776) );
  OAI21_X1 U7291 ( .B1(P2_U3152), .B2(n6194), .A(n8776), .ZN(n6195) );
  OR2_X1 U7292 ( .A1(n6196), .A2(n6195), .ZN(n6219) );
  INV_X1 U7293 ( .A(n6219), .ZN(n6198) );
  INV_X1 U7294 ( .A(n9383), .ZN(n8999) );
  AOI211_X1 U7295 ( .C1(n6200), .C2(n6199), .A(n8963), .B(n4946), .ZN(n6231)
         );
  NOR2_X1 U7296 ( .A1(n7589), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6201) );
  AOI21_X1 U7297 ( .B1(n7589), .B2(P2_REG2_REG_14__SCAN_IN), .A(n6201), .ZN(
        n7597) );
  NAND2_X1 U7298 ( .A1(n7431), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6202) );
  OAI21_X1 U7299 ( .B1(n7431), .B2(P2_REG2_REG_12__SCAN_IN), .A(n6202), .ZN(
        n7427) );
  AOI21_X1 U7300 ( .B1(n10316), .B2(P2_REG2_REG_1__SCAN_IN), .A(n10308), .ZN(
        n10323) );
  NAND2_X1 U7301 ( .A1(n10329), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6204) );
  OAI21_X1 U7302 ( .B1(n10329), .B2(P2_REG2_REG_2__SCAN_IN), .A(n6204), .ZN(
        n10322) );
  NOR2_X1 U7303 ( .A1(n10323), .A2(n10322), .ZN(n10321) );
  AOI21_X1 U7304 ( .B1(n10329), .B2(P2_REG2_REG_2__SCAN_IN), .A(n10321), .ZN(
        n6286) );
  NAND2_X1 U7305 ( .A1(n6287), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6205) );
  OAI21_X1 U7306 ( .B1(n6287), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6205), .ZN(
        n6285) );
  NOR2_X1 U7307 ( .A1(n6286), .A2(n6285), .ZN(n6284) );
  AOI21_X1 U7308 ( .B1(n6287), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6284), .ZN(
        n6262) );
  MUX2_X1 U7309 ( .A(n6206), .B(P2_REG2_REG_4__SCAN_IN), .S(n6263), .Z(n6261)
         );
  NOR2_X1 U7310 ( .A1(n6262), .A2(n6261), .ZN(n6260) );
  AOI21_X1 U7311 ( .B1(n6263), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6260), .ZN(
        n6249) );
  MUX2_X1 U7312 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n6986), .S(n6250), .Z(n6207)
         );
  INV_X1 U7313 ( .A(n6207), .ZN(n6248) );
  MUX2_X1 U7314 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n9252), .S(n6238), .Z(n6208)
         );
  INV_X1 U7315 ( .A(n6208), .ZN(n6236) );
  MUX2_X1 U7316 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7244), .S(n6274), .Z(n6209)
         );
  INV_X1 U7317 ( .A(n6209), .ZN(n6273) );
  NOR2_X1 U7318 ( .A1(n4897), .A2(n6273), .ZN(n6272) );
  MUX2_X1 U7319 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7266), .S(n6359), .Z(n6210)
         );
  INV_X1 U7320 ( .A(n6210), .ZN(n6297) );
  NAND2_X1 U7321 ( .A1(n6382), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6211) );
  OAI21_X1 U7322 ( .B1(n6382), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6211), .ZN(
        n6309) );
  AOI21_X1 U7323 ( .B1(n6382), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6308), .ZN(
        n6322) );
  NAND2_X1 U7324 ( .A1(n6401), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6212) );
  OAI21_X1 U7325 ( .B1(n6401), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6212), .ZN(
        n6321) );
  NOR2_X1 U7326 ( .A1(n6322), .A2(n6321), .ZN(n6320) );
  NOR2_X1 U7327 ( .A1(n6451), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6213) );
  AOI21_X1 U7328 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n6451), .A(n6213), .ZN(
        n7160) );
  AOI21_X1 U7329 ( .B1(n7431), .B2(P2_REG2_REG_12__SCAN_IN), .A(n7426), .ZN(
        n7439) );
  NOR2_X1 U7330 ( .A1(n6692), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6214) );
  AOI21_X1 U7331 ( .B1(n6692), .B2(P2_REG2_REG_13__SCAN_IN), .A(n6214), .ZN(
        n7440) );
  NAND2_X1 U7332 ( .A1(n7439), .A2(n7440), .ZN(n7438) );
  OAI21_X1 U7333 ( .B1(n6692), .B2(P2_REG2_REG_13__SCAN_IN), .A(n7438), .ZN(
        n7596) );
  NAND2_X1 U7334 ( .A1(n7597), .A2(n7596), .ZN(n7595) );
  NAND2_X1 U7335 ( .A1(n7003), .A2(n6215), .ZN(n6216) );
  NAND2_X1 U7336 ( .A1(n6216), .A2(n8943), .ZN(n8957) );
  NAND2_X1 U7337 ( .A1(n8951), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6217) );
  OAI21_X1 U7338 ( .B1(n8951), .B2(P2_REG2_REG_16__SCAN_IN), .A(n6217), .ZN(
        n8956) );
  NAND2_X1 U7339 ( .A1(n8974), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6218) );
  OAI21_X1 U7340 ( .B1(n8974), .B2(P2_REG2_REG_17__SCAN_IN), .A(n6218), .ZN(
        n6222) );
  NAND2_X1 U7341 ( .A1(n6219), .A2(n6225), .ZN(n6220) );
  INV_X2 U7342 ( .A(P2_U3966), .ZN(n8933) );
  NAND2_X1 U7343 ( .A1(n6220), .A2(n8933), .ZN(n6224) );
  NOR2_X1 U7344 ( .A1(n6125), .A2(n9383), .ZN(n6221) );
  AOI211_X1 U7345 ( .C1(n6223), .C2(n6222), .A(n8973), .B(n10320), .ZN(n6230)
         );
  AND2_X1 U7346 ( .A1(n6224), .A2(n6125), .ZN(n10330) );
  NOR2_X1 U7347 ( .A1(n8991), .A2(n5015), .ZN(n6229) );
  OAI21_X1 U7348 ( .B1(n6864), .B2(n6493), .A(n6225), .ZN(n6227) );
  NAND2_X1 U7349 ( .A1(n6864), .A2(n8776), .ZN(n6226) );
  INV_X1 U7350 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7695) );
  NAND2_X1 U7351 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3152), .ZN(n7952) );
  OAI21_X1 U7352 ( .B1(n8968), .B2(n7695), .A(n7952), .ZN(n6228) );
  OR4_X1 U7353 ( .A1(n6231), .A2(n6230), .A3(n6229), .A4(n6228), .ZN(P2_U3262)
         );
  AOI211_X1 U7354 ( .C1(n6234), .C2(n6233), .A(n6232), .B(n4946), .ZN(n6243)
         );
  AOI211_X1 U7355 ( .C1(n6237), .C2(n6236), .A(n6235), .B(n10320), .ZN(n6242)
         );
  INV_X1 U7356 ( .A(n6238), .ZN(n6354) );
  NOR2_X1 U7357 ( .A1(n8991), .A2(n6354), .ZN(n6241) );
  INV_X1 U7358 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6239) );
  NAND2_X1 U7359 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n6961) );
  OAI21_X1 U7360 ( .B1(n8968), .B2(n6239), .A(n6961), .ZN(n6240) );
  OR4_X1 U7361 ( .A1(n6243), .A2(n6242), .A3(n6241), .A4(n6240), .ZN(P2_U3251)
         );
  AOI211_X1 U7362 ( .C1(n6246), .C2(n6245), .A(n6244), .B(n4946), .ZN(n6256)
         );
  AOI211_X1 U7363 ( .C1(n6249), .C2(n6248), .A(n6247), .B(n10320), .ZN(n6255)
         );
  INV_X1 U7364 ( .A(n6250), .ZN(n6345) );
  NOR2_X1 U7365 ( .A1(n8991), .A2(n6345), .ZN(n6254) );
  INV_X1 U7366 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6252) );
  NAND2_X1 U7367 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3152), .ZN(n6251) );
  OAI21_X1 U7368 ( .B1(n8968), .B2(n6252), .A(n6251), .ZN(n6253) );
  OR4_X1 U7369 ( .A1(n6256), .A2(n6255), .A3(n6254), .A4(n6253), .ZN(P2_U3250)
         );
  AOI211_X1 U7370 ( .C1(n6259), .C2(n6258), .A(n6257), .B(n4946), .ZN(n6268)
         );
  AOI211_X1 U7371 ( .C1(n6262), .C2(n6261), .A(n6260), .B(n10320), .ZN(n6267)
         );
  INV_X1 U7372 ( .A(n6263), .ZN(n6342) );
  NOR2_X1 U7373 ( .A1(n8991), .A2(n6342), .ZN(n6266) );
  INV_X1 U7374 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6264) );
  NAND2_X1 U7375 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n6713) );
  OAI21_X1 U7376 ( .B1(n8968), .B2(n6264), .A(n6713), .ZN(n6265) );
  OR4_X1 U7377 ( .A1(n6268), .A2(n6267), .A3(n6266), .A4(n6265), .ZN(P2_U3249)
         );
  AOI211_X1 U7378 ( .C1(n6271), .C2(n6270), .A(n6269), .B(n4946), .ZN(n6280)
         );
  AOI211_X1 U7379 ( .C1(n4897), .C2(n6273), .A(n6272), .B(n10320), .ZN(n6279)
         );
  INV_X1 U7380 ( .A(n6274), .ZN(n6358) );
  NOR2_X1 U7381 ( .A1(n8991), .A2(n6358), .ZN(n6278) );
  INV_X1 U7382 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6276) );
  NAND2_X1 U7383 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3152), .ZN(n6275) );
  OAI21_X1 U7384 ( .B1(n8968), .B2(n6276), .A(n6275), .ZN(n6277) );
  OR4_X1 U7385 ( .A1(n6280), .A2(n6279), .A3(n6278), .A4(n6277), .ZN(P2_U3252)
         );
  AOI211_X1 U7386 ( .C1(n6283), .C2(n6282), .A(n6281), .B(n4946), .ZN(n6292)
         );
  AOI211_X1 U7387 ( .C1(n6286), .C2(n6285), .A(n6284), .B(n10320), .ZN(n6291)
         );
  INV_X1 U7388 ( .A(n6287), .ZN(n6335) );
  NOR2_X1 U7389 ( .A1(n8991), .A2(n6335), .ZN(n6290) );
  NAND2_X1 U7390 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3152), .ZN(n6288) );
  OAI21_X1 U7391 ( .B1(n8968), .B2(n7657), .A(n6288), .ZN(n6289) );
  OR4_X1 U7392 ( .A1(n6292), .A2(n6291), .A3(n6290), .A4(n6289), .ZN(P2_U3248)
         );
  AOI211_X1 U7393 ( .C1(n6295), .C2(n6294), .A(n6293), .B(n4946), .ZN(n6304)
         );
  AOI211_X1 U7394 ( .C1(n6298), .C2(n6297), .A(n6296), .B(n10320), .ZN(n6303)
         );
  INV_X1 U7395 ( .A(n6359), .ZN(n6299) );
  NOR2_X1 U7396 ( .A1(n8991), .A2(n6299), .ZN(n6302) );
  INV_X1 U7397 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n6300) );
  NAND2_X1 U7398 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n7176) );
  OAI21_X1 U7399 ( .B1(n8968), .B2(n6300), .A(n7176), .ZN(n6301) );
  OR4_X1 U7400 ( .A1(n6304), .A2(n6303), .A3(n6302), .A4(n6301), .ZN(P2_U3253)
         );
  AOI211_X1 U7401 ( .C1(n6307), .C2(n6306), .A(n6305), .B(n4946), .ZN(n6316)
         );
  AOI211_X1 U7402 ( .C1(n6310), .C2(n6309), .A(n6308), .B(n10320), .ZN(n6315)
         );
  INV_X1 U7403 ( .A(n6382), .ZN(n6311) );
  NOR2_X1 U7404 ( .A1(n8991), .A2(n6311), .ZN(n6314) );
  INV_X1 U7405 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n6312) );
  NAND2_X1 U7406 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7483) );
  OAI21_X1 U7407 ( .B1(n8968), .B2(n6312), .A(n7483), .ZN(n6313) );
  OR4_X1 U7408 ( .A1(n6316), .A2(n6315), .A3(n6314), .A4(n6313), .ZN(P2_U3254)
         );
  AOI211_X1 U7409 ( .C1(n6319), .C2(n6318), .A(n6317), .B(n4946), .ZN(n6327)
         );
  AOI211_X1 U7410 ( .C1(n6322), .C2(n6321), .A(n6320), .B(n10320), .ZN(n6326)
         );
  INV_X1 U7411 ( .A(n6401), .ZN(n6323) );
  NOR2_X1 U7412 ( .A1(n8991), .A2(n6323), .ZN(n6325) );
  INV_X1 U7413 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7656) );
  NAND2_X1 U7414 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7601) );
  OAI21_X1 U7415 ( .B1(n8968), .B2(n7656), .A(n7601), .ZN(n6324) );
  OR4_X1 U7416 ( .A1(n6327), .A2(n6326), .A3(n6325), .A4(n6324), .ZN(P2_U3255)
         );
  NAND2_X2 U7417 ( .A1(n8253), .A2(P2_U3152), .ZN(n9380) );
  NOR2_X2 U7418 ( .A1(n8253), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9373) );
  AOI22_X1 U7419 ( .A1(n9373), .A2(P1_DATAO_REG_1__SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(n10316), .ZN(n6328) );
  OAI21_X1 U7420 ( .B1(n6719), .B2(n9380), .A(n6328), .ZN(P2_U3357) );
  AOI22_X1 U7421 ( .A1(n9373), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(n10329), .ZN(n6329) );
  OAI21_X1 U7422 ( .B1(n6806), .B2(n9380), .A(n6329), .ZN(P2_U3356) );
  INV_X1 U7423 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n6331) );
  NAND2_X1 U7424 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6330) );
  XNOR2_X1 U7425 ( .A(n6331), .B(n6330), .ZN(n10287) );
  NOR2_X1 U7426 ( .A1(n8253), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9954) );
  INV_X2 U7427 ( .A(n9954), .ZN(n8830) );
  INV_X1 U7428 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6720) );
  NAND2_X2 U7429 ( .A1(n8253), .A2(P1_U3084), .ZN(n9961) );
  OAI222_X1 U7430 ( .A1(P1_U3084), .A2(n10287), .B1(n8830), .B2(n6719), .C1(
        n6720), .C2(n9961), .ZN(P1_U3352) );
  OR2_X1 U7431 ( .A1(n6332), .A2(n6162), .ZN(n6333) );
  XNOR2_X1 U7432 ( .A(n6333), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6471) );
  INV_X1 U7433 ( .A(n6471), .ZN(n10352) );
  INV_X1 U7434 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6805) );
  OAI222_X1 U7435 ( .A1(P1_U3084), .A2(n10352), .B1(n8830), .B2(n6806), .C1(
        n6805), .C2(n9961), .ZN(P1_U3351) );
  INV_X1 U7436 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6334) );
  INV_X1 U7437 ( .A(n9373), .ZN(n9385) );
  OAI222_X1 U7438 ( .A1(n9380), .A2(n6795), .B1(n6335), .B2(P2_U3152), .C1(
        n6334), .C2(n9385), .ZN(P2_U3355) );
  OR3_X1 U7439 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U7440 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n6336), .ZN(n6337) );
  XNOR2_X1 U7441 ( .A(n6337), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6538) );
  INV_X1 U7442 ( .A(n6538), .ZN(n6796) );
  INV_X1 U7443 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6794) );
  OAI222_X1 U7444 ( .A1(P1_U3084), .A2(n6796), .B1(n8830), .B2(n6795), .C1(
        n6794), .C2(n9961), .ZN(P1_U3350) );
  INV_X1 U7445 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6885) );
  NAND2_X1 U7446 ( .A1(n6338), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6340) );
  NAND2_X1 U7447 ( .A1(n6340), .A2(n6339), .ZN(n6343) );
  OR2_X1 U7448 ( .A1(n6340), .A2(n6339), .ZN(n6341) );
  AND2_X1 U7449 ( .A1(n6343), .A2(n6341), .ZN(n6474) );
  INV_X1 U7450 ( .A(n6474), .ZN(n10363) );
  OAI222_X1 U7451 ( .A1(n9961), .A2(n6885), .B1(n8830), .B2(n6884), .C1(
        P1_U3084), .C2(n10363), .ZN(P1_U3349) );
  OAI222_X1 U7452 ( .A1(n6342), .A2(P2_U3152), .B1(n9380), .B2(n6884), .C1(
        n9385), .C2(n4964), .ZN(P2_U3354) );
  INV_X1 U7453 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6902) );
  NAND2_X1 U7454 ( .A1(n6343), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6344) );
  XNOR2_X1 U7455 ( .A(n6344), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6476) );
  INV_X1 U7456 ( .A(n6476), .ZN(n10274) );
  OAI222_X1 U7457 ( .A1(n9961), .A2(n6902), .B1(n8830), .B2(n6900), .C1(
        P1_U3084), .C2(n10274), .ZN(P1_U3348) );
  INV_X1 U7458 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6446) );
  OAI222_X1 U7459 ( .A1(n6345), .A2(P2_U3152), .B1(n9380), .B2(n6900), .C1(
        n9385), .C2(n6446), .ZN(P2_U3353) );
  INV_X1 U7460 ( .A(n8968), .ZN(n10319) );
  NOR2_X1 U7461 ( .A1(n10319), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7462 ( .A(n7051), .ZN(n6353) );
  OR2_X1 U7463 ( .A1(n6338), .A2(n6346), .ZN(n6347) );
  NAND2_X1 U7464 ( .A1(n6347), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6348) );
  MUX2_X1 U7465 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6348), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n6351) );
  INV_X1 U7466 ( .A(n6349), .ZN(n6350) );
  INV_X1 U7467 ( .A(n9961), .ZN(n9958) );
  AOI22_X1 U7468 ( .A1(n7050), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n9958), .ZN(n6352) );
  OAI21_X1 U7469 ( .B1(n6353), .B2(n8830), .A(n6352), .ZN(P1_U3347) );
  INV_X1 U7470 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6435) );
  OAI222_X1 U7471 ( .A1(n6354), .A2(P2_U3152), .B1(n9380), .B2(n6353), .C1(
        n9385), .C2(n6435), .ZN(P2_U3352) );
  INV_X1 U7472 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6356) );
  INV_X1 U7473 ( .A(n7128), .ZN(n6357) );
  OR2_X1 U7474 ( .A1(n6349), .A2(n6162), .ZN(n6355) );
  XNOR2_X1 U7475 ( .A(n6355), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7129) );
  INV_X1 U7476 ( .A(n7129), .ZN(n6482) );
  OAI222_X1 U7477 ( .A1(n9961), .A2(n6356), .B1(n8830), .B2(n6357), .C1(
        P1_U3084), .C2(n6482), .ZN(P1_U3346) );
  INV_X1 U7478 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6418) );
  OAI222_X1 U7479 ( .A1(n6358), .A2(P2_U3152), .B1(n9380), .B2(n6357), .C1(
        n9385), .C2(n6418), .ZN(P2_U3351) );
  INV_X1 U7480 ( .A(n7282), .ZN(n6366) );
  AOI22_X1 U7481 ( .A1(n6359), .A2(P2_STATE_REG_SCAN_IN), .B1(n9373), .B2(
        P1_DATAO_REG_8__SCAN_IN), .ZN(n6360) );
  OAI21_X1 U7482 ( .B1(n6366), .B2(n9380), .A(n6360), .ZN(P2_U3350) );
  INV_X1 U7483 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6367) );
  OR2_X1 U7484 ( .A1(n6361), .A2(n6162), .ZN(n6364) );
  INV_X1 U7485 ( .A(n6364), .ZN(n6362) );
  NAND2_X1 U7486 ( .A1(n6362), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6365) );
  INV_X1 U7487 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6363) );
  NAND2_X1 U7488 ( .A1(n6364), .A2(n6363), .ZN(n6397) );
  INV_X1 U7489 ( .A(n7283), .ZN(n6519) );
  OAI222_X1 U7490 ( .A1(n9961), .A2(n6367), .B1(n8830), .B2(n6366), .C1(
        P1_U3084), .C2(n6519), .ZN(P1_U3345) );
  INV_X1 U7491 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6450) );
  NAND2_X1 U7492 ( .A1(n10586), .A2(P2_U3966), .ZN(n6368) );
  OAI21_X1 U7493 ( .B1(n6450), .B2(P2_U3966), .A(n6368), .ZN(P2_U3562) );
  XNOR2_X1 U7494 ( .A(n6374), .B(P1_IR_REG_25__SCAN_IN), .ZN(n7961) );
  AND2_X1 U7495 ( .A1(n8779), .A2(P1_B_REG_SCAN_IN), .ZN(n6373) );
  INV_X1 U7496 ( .A(P1_B_REG_SCAN_IN), .ZN(n8822) );
  INV_X1 U7497 ( .A(n8779), .ZN(n6372) );
  AOI22_X1 U7498 ( .A1(n7961), .A2(n6373), .B1(n8822), .B2(n6372), .ZN(n6376)
         );
  INV_X1 U7499 ( .A(n6629), .ZN(n6377) );
  INV_X1 U7500 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6615) );
  INV_X1 U7501 ( .A(n6378), .ZN(n9964) );
  NAND2_X1 U7502 ( .A1(n9964), .A2(n7961), .ZN(n6616) );
  INV_X1 U7503 ( .A(n6616), .ZN(n6379) );
  AOI22_X1 U7504 ( .A1(n9967), .A2(n6615), .B1(n6380), .B2(n6379), .ZN(
        P1_U3441) );
  INV_X1 U7505 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6400) );
  INV_X1 U7506 ( .A(n7331), .ZN(n7603) );
  NAND2_X1 U7507 ( .A1(n7603), .A2(P2_U3966), .ZN(n6381) );
  OAI21_X1 U7508 ( .B1(n6400), .B2(P2_U3966), .A(n6381), .ZN(P2_U3561) );
  INV_X1 U7509 ( .A(n7398), .ZN(n6399) );
  AOI22_X1 U7510 ( .A1(n6382), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n9373), .ZN(n6383) );
  OAI21_X1 U7511 ( .B1(n6399), .B2(n9380), .A(n6383), .ZN(P2_U3349) );
  INV_X1 U7512 ( .A(n7823), .ZN(n6384) );
  NOR2_X1 U7513 ( .A1(n6780), .A2(n6384), .ZN(n6385) );
  INV_X1 U7514 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6396) );
  INV_X1 U7515 ( .A(n6386), .ZN(n10339) );
  INV_X1 U7516 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10291) );
  INV_X1 U7517 ( .A(n6387), .ZN(n10338) );
  OR2_X1 U7518 ( .A1(n6386), .A2(n10338), .ZN(n10345) );
  INV_X1 U7519 ( .A(n10345), .ZN(n6388) );
  AOI21_X1 U7520 ( .B1(n10339), .B2(P1_REG2_REG_0__SCAN_IN), .A(n6388), .ZN(
        n10343) );
  INV_X1 U7521 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10342) );
  NOR2_X1 U7522 ( .A1(n10343), .A2(n10342), .ZN(n6391) );
  NAND3_X1 U7523 ( .A1(n7049), .A2(P1_STATE_REG_SCAN_IN), .A3(n6465), .ZN(
        n6390) );
  NOR2_X1 U7524 ( .A1(n10345), .A2(P1_U3084), .ZN(n6389) );
  NAND2_X1 U7525 ( .A1(n6389), .A2(n6465), .ZN(n10333) );
  INV_X1 U7526 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6688) );
  OAI22_X1 U7527 ( .A1(n6391), .A2(n6390), .B1(n10333), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n6394) );
  NOR2_X1 U7528 ( .A1(n10338), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6392) );
  OAI21_X1 U7529 ( .B1(n10343), .B2(n6392), .A(n10342), .ZN(n6393) );
  AOI22_X1 U7530 ( .A1(n6394), .A2(n6393), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3084), .ZN(n6395) );
  OAI21_X1 U7531 ( .B1(n10376), .B2(n6396), .A(n6395), .ZN(P1_U3241) );
  NAND2_X1 U7532 ( .A1(n6397), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6398) );
  XNOR2_X1 U7533 ( .A(n6398), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7399) );
  INV_X1 U7534 ( .A(n7399), .ZN(n6554) );
  OAI222_X1 U7535 ( .A1(P1_U3084), .A2(n6554), .B1(n9961), .B2(n6400), .C1(
        n6399), .C2(n8830), .ZN(P1_U3344) );
  INV_X1 U7536 ( .A(n7498), .ZN(n6449) );
  AOI22_X1 U7537 ( .A1(n6401), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n9373), .ZN(n6402) );
  OAI21_X1 U7538 ( .B1(n6449), .B2(n9380), .A(n6402), .ZN(P2_U3348) );
  INV_X2 U7539 ( .A(n10340), .ZN(P1_U4006) );
  NAND2_X1 U7540 ( .A1(n6405), .A2(n6406), .ZN(n9949) );
  NAND2_X1 U7541 ( .A1(n4862), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6416) );
  INV_X1 U7542 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7385) );
  OR2_X1 U7543 ( .A1(n7853), .A2(n7385), .ZN(n6415) );
  NAND2_X1 U7544 ( .A1(n6426), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6428) );
  INV_X1 U7545 ( .A(n6428), .ZN(n6408) );
  NAND2_X1 U7546 ( .A1(n6408), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7146) );
  INV_X1 U7547 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6409) );
  NAND2_X1 U7548 ( .A1(n6428), .A2(n6409), .ZN(n6410) );
  NAND2_X1 U7549 ( .A1(n7146), .A2(n6410), .ZN(n7391) );
  OR2_X1 U7550 ( .A1(n6788), .A2(n7391), .ZN(n6414) );
  INV_X1 U7551 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6412) );
  OR2_X1 U7552 ( .A1(n6787), .A2(n6412), .ZN(n6413) );
  NAND4_X1 U7553 ( .A1(n6416), .A2(n6415), .A3(n6414), .A4(n6413), .ZN(n7367)
         );
  NAND2_X1 U7554 ( .A1(n7367), .A2(P1_U4006), .ZN(n6417) );
  OAI21_X1 U7555 ( .B1(P1_U4006), .B2(n6418), .A(n6417), .ZN(P1_U3562) );
  NAND2_X1 U7556 ( .A1(n4862), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6423) );
  INV_X1 U7557 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6419) );
  XNOR2_X1 U7558 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7120) );
  OR2_X1 U7559 ( .A1(n6788), .A2(n7120), .ZN(n6422) );
  INV_X1 U7560 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6420) );
  NAND2_X1 U7561 ( .A1(n6883), .A2(P1_U4006), .ZN(n6424) );
  OAI21_X1 U7562 ( .B1(P1_U4006), .B2(n4964), .A(n6424), .ZN(P1_U3559) );
  NAND2_X1 U7563 ( .A1(n4862), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6433) );
  INV_X1 U7564 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6425) );
  OR2_X1 U7565 ( .A1(n7853), .A2(n6425), .ZN(n6432) );
  INV_X1 U7566 ( .A(n6426), .ZN(n6440) );
  INV_X1 U7567 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6523) );
  NAND2_X1 U7568 ( .A1(n6440), .A2(n6523), .ZN(n6427) );
  NAND2_X1 U7569 ( .A1(n6428), .A2(n6427), .ZN(n7327) );
  OR2_X1 U7570 ( .A1(n8145), .A2(n7327), .ZN(n6431) );
  INV_X1 U7571 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6429) );
  OR2_X1 U7572 ( .A1(n6787), .A2(n6429), .ZN(n6430) );
  NAND2_X1 U7573 ( .A1(n7290), .A2(P1_U4006), .ZN(n6434) );
  OAI21_X1 U7574 ( .B1(P1_U4006), .B2(n6435), .A(n6434), .ZN(P1_U3561) );
  NAND2_X1 U7575 ( .A1(n4862), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6444) );
  INV_X1 U7576 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6436) );
  OR2_X1 U7577 ( .A1(n6787), .A2(n6436), .ZN(n6443) );
  INV_X1 U7578 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6438) );
  NAND2_X1 U7579 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6437) );
  NAND2_X1 U7580 ( .A1(n6438), .A2(n6437), .ZN(n6439) );
  NAND2_X1 U7581 ( .A1(n6440), .A2(n6439), .ZN(n7211) );
  INV_X1 U7582 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6459) );
  OR2_X1 U7583 ( .A1(n7853), .A2(n6459), .ZN(n6441) );
  NAND2_X1 U7584 ( .A1(n7322), .A2(P1_U4006), .ZN(n6445) );
  OAI21_X1 U7585 ( .B1(P1_U4006), .B2(n6446), .A(n6445), .ZN(P1_U3560) );
  NAND2_X1 U7586 ( .A1(n6447), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6448) );
  XNOR2_X1 U7587 ( .A(n6448), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10240) );
  INV_X1 U7588 ( .A(n10240), .ZN(n6584) );
  OAI222_X1 U7589 ( .A1(P1_U3084), .A2(n6584), .B1(n9961), .B2(n6450), .C1(
        n6449), .C2(n8830), .ZN(P1_U3343) );
  INV_X1 U7590 ( .A(n6451), .ZN(n7170) );
  INV_X1 U7591 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6452) );
  OAI222_X1 U7592 ( .A1(n9380), .A2(n7526), .B1(n7170), .B2(P2_U3152), .C1(
        n6452), .C2(n9385), .ZN(P2_U3347) );
  NAND2_X1 U7593 ( .A1(n7050), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6461) );
  MUX2_X1 U7594 ( .A(n6425), .B(P1_REG2_REG_6__SCAN_IN), .S(n7050), .Z(n6453)
         );
  INV_X1 U7595 ( .A(n6453), .ZN(n6529) );
  NOR2_X1 U7596 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6476), .ZN(n6460) );
  NOR2_X1 U7597 ( .A1(n6474), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U7598 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(n6538), .ZN(n6457) );
  INV_X1 U7599 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6789) );
  MUX2_X1 U7600 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6789), .S(n6538), .Z(n6540)
         );
  NAND2_X1 U7601 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n6471), .ZN(n6456) );
  INV_X1 U7602 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6454) );
  MUX2_X1 U7603 ( .A(n6454), .B(P1_REG2_REG_2__SCAN_IN), .S(n6471), .Z(n6455)
         );
  INV_X1 U7604 ( .A(n6455), .ZN(n10350) );
  INV_X1 U7605 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10424) );
  MUX2_X1 U7606 ( .A(n10424), .B(P1_REG2_REG_1__SCAN_IN), .S(n10287), .Z(
        n10293) );
  NAND3_X1 U7607 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .A3(n10293), .ZN(n10292) );
  OAI21_X1 U7608 ( .B1(n10287), .B2(n10424), .A(n10292), .ZN(n10349) );
  NAND2_X1 U7609 ( .A1(n10350), .A2(n10349), .ZN(n10347) );
  NAND2_X1 U7610 ( .A1(n6456), .A2(n10347), .ZN(n6541) );
  NAND2_X1 U7611 ( .A1(n6540), .A2(n6541), .ZN(n6539) );
  NAND2_X1 U7612 ( .A1(n6457), .A2(n6539), .ZN(n10359) );
  AOI22_X1 U7613 ( .A1(n6474), .A2(n6420), .B1(P1_REG2_REG_4__SCAN_IN), .B2(
        n10363), .ZN(n10358) );
  NOR2_X1 U7614 ( .A1(n10359), .A2(n10358), .ZN(n10357) );
  NOR2_X1 U7615 ( .A1(n6458), .A2(n10357), .ZN(n10278) );
  MUX2_X1 U7616 ( .A(n6459), .B(P1_REG2_REG_5__SCAN_IN), .S(n6476), .Z(n10277)
         );
  NOR2_X1 U7617 ( .A1(n10278), .A2(n10277), .ZN(n10276) );
  NOR2_X1 U7618 ( .A1(n6460), .A2(n10276), .ZN(n6530) );
  NAND2_X1 U7619 ( .A1(n6529), .A2(n6530), .ZN(n6528) );
  NAND2_X1 U7620 ( .A1(n6461), .A2(n6528), .ZN(n6464) );
  MUX2_X1 U7621 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n7385), .S(n7129), .Z(n6462)
         );
  INV_X1 U7622 ( .A(n6462), .ZN(n6463) );
  NOR2_X1 U7623 ( .A1(n6464), .A2(n6463), .ZN(n6506) );
  AOI21_X1 U7624 ( .B1(n6464), .B2(n6463), .A(n6506), .ZN(n6485) );
  NOR2_X1 U7625 ( .A1(n6387), .A2(P1_U3084), .ZN(n9957) );
  NAND2_X1 U7626 ( .A1(n6465), .A2(n9957), .ZN(n6592) );
  OR2_X1 U7627 ( .A1(n6592), .A2(n6386), .ZN(n10370) );
  OR2_X1 U7628 ( .A1(n6592), .A2(n10339), .ZN(n10364) );
  INV_X1 U7629 ( .A(n10333), .ZN(n10368) );
  NOR2_X1 U7630 ( .A1(n7129), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6466) );
  AOI21_X1 U7631 ( .B1(n7129), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6466), .ZN(
        n6479) );
  OR2_X1 U7632 ( .A1(n6476), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6468) );
  NAND2_X1 U7633 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6476), .ZN(n6467) );
  NAND2_X1 U7634 ( .A1(n6468), .A2(n6467), .ZN(n10265) );
  INV_X1 U7635 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6638) );
  OR2_X1 U7636 ( .A1(n10287), .A2(n6638), .ZN(n6470) );
  MUX2_X1 U7637 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6638), .S(n10287), .Z(n10284) );
  NOR3_X1 U7638 ( .A1(n10342), .A2(n6688), .A3(n10284), .ZN(n10283) );
  INV_X1 U7639 ( .A(n10283), .ZN(n6469) );
  AND2_X1 U7640 ( .A1(n6470), .A2(n6469), .ZN(n10336) );
  XNOR2_X1 U7641 ( .A(n6471), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n10335) );
  NOR2_X1 U7642 ( .A1(n10336), .A2(n10335), .ZN(n10334) );
  AOI21_X1 U7643 ( .B1(n6471), .B2(P1_REG1_REG_2__SCAN_IN), .A(n10334), .ZN(
        n6536) );
  NAND2_X1 U7644 ( .A1(P1_REG1_REG_3__SCAN_IN), .A2(n6538), .ZN(n6472) );
  OAI21_X1 U7645 ( .B1(n6538), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6472), .ZN(
        n6535) );
  NOR2_X1 U7646 ( .A1(n6536), .A2(n6535), .ZN(n6534) );
  AOI21_X1 U7647 ( .B1(n6538), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6534), .ZN(
        n10362) );
  NOR2_X1 U7648 ( .A1(n6474), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6473) );
  AOI21_X1 U7649 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n6474), .A(n6473), .ZN(
        n10361) );
  NAND2_X1 U7650 ( .A1(n10362), .A2(n10361), .ZN(n10360) );
  OR2_X1 U7651 ( .A1(n6474), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6475) );
  NAND2_X1 U7652 ( .A1(n10360), .A2(n6475), .ZN(n10266) );
  NOR2_X1 U7653 ( .A1(n10265), .A2(n10266), .ZN(n10267) );
  AOI21_X1 U7654 ( .B1(n6476), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10267), .ZN(
        n6526) );
  NAND2_X1 U7655 ( .A1(n7050), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6477) );
  OAI21_X1 U7656 ( .B1(n7050), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6477), .ZN(
        n6525) );
  NOR2_X1 U7657 ( .A1(n6526), .A2(n6525), .ZN(n6524) );
  AOI21_X1 U7658 ( .B1(n7050), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6524), .ZN(
        n6478) );
  NAND2_X1 U7659 ( .A1(n6478), .A2(n6479), .ZN(n6513) );
  OAI21_X1 U7660 ( .B1(n6479), .B2(n6478), .A(n6513), .ZN(n6480) );
  AND2_X1 U7661 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7153) );
  AOI21_X1 U7662 ( .B1(n10368), .B2(n6480), .A(n7153), .ZN(n6481) );
  OAI21_X1 U7663 ( .B1(n6482), .B2(n10364), .A(n6481), .ZN(n6483) );
  AOI21_X1 U7664 ( .B1(n10290), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n6483), .ZN(
        n6484) );
  OAI21_X1 U7665 ( .B1(n6485), .B2(n10370), .A(n6484), .ZN(P1_U3248) );
  INV_X1 U7666 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6487) );
  OR2_X1 U7667 ( .A1(n6447), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6606) );
  NAND2_X1 U7668 ( .A1(n6606), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6486) );
  XNOR2_X1 U7669 ( .A(n6486), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7527) );
  INV_X1 U7670 ( .A(n7527), .ZN(n6593) );
  OAI222_X1 U7671 ( .A1(n9961), .A2(n6487), .B1(n8830), .B2(n7526), .C1(n6593), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  AND2_X1 U7672 ( .A1(n6578), .A2(n9971), .ZN(n6488) );
  AND2_X1 U7673 ( .A1(n6489), .A2(n6488), .ZN(n6862) );
  INV_X1 U7674 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6501) );
  INV_X1 U7675 ( .A(n6568), .ZN(n10381) );
  NAND2_X1 U7676 ( .A1(n6496), .A2(n8774), .ZN(n8732) );
  AND2_X1 U7677 ( .A1(n8586), .A2(n8732), .ZN(n7255) );
  NAND2_X1 U7678 ( .A1(n5582), .A2(n8774), .ZN(n6491) );
  NAND2_X1 U7679 ( .A1(n6492), .A2(n6491), .ZN(n6495) );
  AND2_X1 U7680 ( .A1(n6877), .A2(n6493), .ZN(n6494) );
  NAND2_X1 U7681 ( .A1(n6495), .A2(n6494), .ZN(n7474) );
  AND2_X1 U7682 ( .A1(n6496), .A2(n7797), .ZN(n6497) );
  NAND2_X1 U7683 ( .A1(n6098), .A2(n6497), .ZN(n10435) );
  INV_X1 U7684 ( .A(n8934), .ZN(n6498) );
  NAND2_X1 U7685 ( .A1(n6498), .A2(n6568), .ZN(n6563) );
  NAND2_X1 U7686 ( .A1(n8934), .A2(n10381), .ZN(n8591) );
  NAND2_X1 U7687 ( .A1(n6563), .A2(n8591), .ZN(n10377) );
  OAI21_X1 U7688 ( .B1(n9234), .B2(n10654), .A(n10377), .ZN(n6499) );
  NAND2_X1 U7689 ( .A1(n4859), .A2(n10587), .ZN(n10378) );
  OAI211_X1 U7690 ( .C1(n10381), .C2(n6877), .A(n6499), .B(n10378), .ZN(n6504)
         );
  NAND2_X1 U7691 ( .A1(n6504), .A2(n10660), .ZN(n6500) );
  OAI21_X1 U7692 ( .B1(n10660), .B2(n6501), .A(n6500), .ZN(P2_U3451) );
  NAND2_X1 U7693 ( .A1(n6504), .A2(n10657), .ZN(n6505) );
  OAI21_X1 U7694 ( .B1(n10657), .B2(n10303), .A(n6505), .ZN(P2_U3520) );
  NOR2_X1 U7695 ( .A1(n7129), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6507) );
  NOR2_X1 U7696 ( .A1(n6507), .A2(n6506), .ZN(n6511) );
  INV_X1 U7697 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6508) );
  MUX2_X1 U7698 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n6508), .S(n7283), .Z(n6509)
         );
  INV_X1 U7699 ( .A(n6509), .ZN(n6510) );
  NOR2_X1 U7700 ( .A1(n6511), .A2(n6510), .ZN(n6545) );
  AOI21_X1 U7701 ( .B1(n6511), .B2(n6510), .A(n6545), .ZN(n6522) );
  NOR2_X1 U7702 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n7283), .ZN(n6512) );
  AOI21_X1 U7703 ( .B1(n7283), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6512), .ZN(
        n6516) );
  OR2_X1 U7704 ( .A1(n7129), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6514) );
  NAND2_X1 U7705 ( .A1(n6514), .A2(n6513), .ZN(n6515) );
  NAND2_X1 U7706 ( .A1(n6516), .A2(n6515), .ZN(n6551) );
  OAI21_X1 U7707 ( .B1(n6516), .B2(n6515), .A(n6551), .ZN(n6517) );
  INV_X1 U7708 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7145) );
  NOR2_X1 U7709 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7145), .ZN(n7366) );
  AOI21_X1 U7710 ( .B1(n10368), .B2(n6517), .A(n7366), .ZN(n6518) );
  OAI21_X1 U7711 ( .B1(n6519), .B2(n10364), .A(n6518), .ZN(n6520) );
  AOI21_X1 U7712 ( .B1(n10290), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n6520), .ZN(
        n6521) );
  OAI21_X1 U7713 ( .B1(n6522), .B2(n10370), .A(n6521), .ZN(P1_U3249) );
  INV_X1 U7714 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6533) );
  NOR2_X1 U7715 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6523), .ZN(n7071) );
  AOI211_X1 U7716 ( .C1(n6526), .C2(n6525), .A(n6524), .B(n10333), .ZN(n6527)
         );
  AOI211_X1 U7717 ( .C1(n10288), .C2(n7050), .A(n7071), .B(n6527), .ZN(n6532)
         );
  OAI211_X1 U7718 ( .C1(n6530), .C2(n6529), .A(n10348), .B(n6528), .ZN(n6531)
         );
  OAI211_X1 U7719 ( .C1(n6533), .C2(n10376), .A(n6532), .B(n6531), .ZN(
        P1_U3247) );
  INV_X1 U7720 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6544) );
  AND2_X1 U7721 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6822) );
  AOI211_X1 U7722 ( .C1(n6536), .C2(n6535), .A(n6534), .B(n10333), .ZN(n6537)
         );
  AOI211_X1 U7723 ( .C1(n10288), .C2(n6538), .A(n6822), .B(n6537), .ZN(n6543)
         );
  OAI211_X1 U7724 ( .C1(n6541), .C2(n6540), .A(n10348), .B(n6539), .ZN(n6542)
         );
  OAI211_X1 U7725 ( .C1(n6544), .C2(n10376), .A(n6543), .B(n6542), .ZN(
        P1_U3244) );
  INV_X1 U7726 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6559) );
  NOR2_X1 U7727 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n7283), .ZN(n6546) );
  NOR2_X1 U7728 ( .A1(n6546), .A2(n6545), .ZN(n6550) );
  INV_X1 U7729 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6547) );
  MUX2_X1 U7730 ( .A(n6547), .B(P1_REG2_REG_9__SCAN_IN), .S(n7399), .Z(n6548)
         );
  INV_X1 U7731 ( .A(n6548), .ZN(n6549) );
  NAND2_X1 U7732 ( .A1(n6549), .A2(n6550), .ZN(n6589) );
  OAI211_X1 U7733 ( .C1(n6550), .C2(n6549), .A(n10348), .B(n6589), .ZN(n6558)
         );
  INV_X1 U7734 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7275) );
  MUX2_X1 U7735 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n7275), .S(n7399), .Z(n6553)
         );
  OAI21_X1 U7736 ( .B1(n7283), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6551), .ZN(
        n6552) );
  NAND2_X1 U7737 ( .A1(n6553), .A2(n6552), .ZN(n6585) );
  OAI21_X1 U7738 ( .B1(n6553), .B2(n6552), .A(n6585), .ZN(n6556) );
  AND2_X1 U7739 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7415) );
  NOR2_X1 U7740 ( .A1(n10364), .A2(n6554), .ZN(n6555) );
  AOI211_X1 U7741 ( .C1(n10368), .C2(n6556), .A(n7415), .B(n6555), .ZN(n6557)
         );
  OAI211_X1 U7742 ( .C1(n10376), .C2(n6559), .A(n6558), .B(n6557), .ZN(
        P1_U3250) );
  INV_X1 U7743 ( .A(n4859), .ZN(n6561) );
  NAND2_X1 U7744 ( .A1(n6561), .A2(n7009), .ZN(n6562) );
  INV_X1 U7745 ( .A(n7009), .ZN(n6570) );
  NAND2_X1 U7746 ( .A1(n4859), .A2(n6570), .ZN(n6847) );
  NAND2_X1 U7747 ( .A1(n6562), .A2(n6847), .ZN(n8588) );
  XNOR2_X1 U7748 ( .A(n6840), .B(n8588), .ZN(n7012) );
  INV_X1 U7749 ( .A(n6847), .ZN(n8593) );
  INV_X1 U7750 ( .A(n6563), .ZN(n6564) );
  NAND2_X1 U7751 ( .A1(n8588), .A2(n6564), .ZN(n6565) );
  OAI211_X1 U7752 ( .C1(n8590), .C2(n8593), .A(n9234), .B(n6565), .ZN(n6567)
         );
  AOI22_X1 U7753 ( .A1(n8932), .A2(n10587), .B1(n9230), .B2(n8934), .ZN(n6566)
         );
  NAND2_X1 U7754 ( .A1(n6567), .A2(n6566), .ZN(n7008) );
  INV_X1 U7755 ( .A(n7041), .ZN(n6569) );
  OAI21_X1 U7756 ( .B1(n6570), .B2(n10381), .A(n6569), .ZN(n7006) );
  OAI22_X1 U7757 ( .A1(n7006), .A2(n10650), .B1(n6570), .B2(n10648), .ZN(n6571) );
  NOR2_X1 U7758 ( .A1(n7008), .A2(n6571), .ZN(n6572) );
  OAI21_X1 U7759 ( .B1(n10530), .B2(n7012), .A(n6572), .ZN(n6574) );
  NAND2_X1 U7760 ( .A1(n6574), .A2(n10660), .ZN(n6573) );
  OAI21_X1 U7761 ( .B1(n10660), .B2(n5610), .A(n6573), .ZN(P2_U3454) );
  NAND2_X1 U7762 ( .A1(n6574), .A2(n10657), .ZN(n6575) );
  OAI21_X1 U7763 ( .B1(n10657), .B2(n6179), .A(n6575), .ZN(P2_U3521) );
  XNOR2_X1 U7764 ( .A(n6577), .B(n6576), .ZN(n6583) );
  NAND2_X1 U7765 ( .A1(n6579), .A2(n6578), .ZN(n6764) );
  INV_X1 U7766 ( .A(n6764), .ZN(n6701) );
  INV_X1 U7767 ( .A(n10514), .ZN(n8906) );
  INV_X1 U7768 ( .A(n10517), .ZN(n8917) );
  AOI22_X1 U7769 ( .A1(n8906), .A2(n4859), .B1(n8917), .B2(n8931), .ZN(n6580)
         );
  OAI21_X1 U7770 ( .B1(n6701), .B2(n7042), .A(n6580), .ZN(n6581) );
  AOI21_X1 U7771 ( .B1(n8918), .B2(n6843), .A(n6581), .ZN(n6582) );
  OAI21_X1 U7772 ( .B1(n10510), .B2(n6583), .A(n6582), .ZN(P2_U3239) );
  INV_X1 U7773 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10567) );
  AOI22_X1 U7774 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n10240), .B1(n6584), .B2(
        n10567), .ZN(n10242) );
  OAI21_X1 U7775 ( .B1(n7399), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6585), .ZN(
        n10243) );
  NAND2_X1 U7776 ( .A1(n10242), .A2(n10243), .ZN(n10241) );
  OAI21_X1 U7777 ( .B1(n10240), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10241), .ZN(
        n6587) );
  INV_X1 U7778 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7511) );
  MUX2_X1 U7779 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n7511), .S(n7527), .Z(n6586)
         );
  NAND2_X1 U7780 ( .A1(n6586), .A2(n6587), .ZN(n6833) );
  OAI21_X1 U7781 ( .B1(n6587), .B2(n6586), .A(n6833), .ZN(n6588) );
  NAND2_X1 U7782 ( .A1(n6588), .A2(n10368), .ZN(n6605) );
  INV_X1 U7783 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7521) );
  MUX2_X1 U7784 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n7521), .S(n10240), .Z(
        n10246) );
  NAND2_X1 U7785 ( .A1(n7399), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6590) );
  NAND2_X1 U7786 ( .A1(n6590), .A2(n6589), .ZN(n10247) );
  NAND2_X1 U7787 ( .A1(n10246), .A2(n10247), .ZN(n10245) );
  INV_X1 U7788 ( .A(n10245), .ZN(n6591) );
  AOI21_X1 U7789 ( .B1(n10240), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6591), .ZN(
        n6596) );
  INV_X1 U7790 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7507) );
  OR3_X1 U7791 ( .A1(n6592), .A2(n6596), .A3(n7507), .ZN(n6594) );
  AOI21_X1 U7792 ( .B1(n10364), .B2(n6594), .A(n6593), .ZN(n6603) );
  INV_X1 U7793 ( .A(n6596), .ZN(n6599) );
  OR2_X1 U7794 ( .A1(n7527), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6598) );
  NAND2_X1 U7795 ( .A1(n7527), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6595) );
  NAND2_X1 U7796 ( .A1(n6596), .A2(n6595), .ZN(n6597) );
  NAND2_X1 U7797 ( .A1(n6597), .A2(n6598), .ZN(n6926) );
  OAI21_X1 U7798 ( .B1(n6599), .B2(n6598), .A(n6926), .ZN(n6601) );
  AND2_X1 U7799 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7567) );
  INV_X1 U7800 ( .A(n7567), .ZN(n6600) );
  OAI21_X1 U7801 ( .B1(n10370), .B2(n6601), .A(n6600), .ZN(n6602) );
  AOI211_X1 U7802 ( .C1(P1_ADDR_REG_11__SCAN_IN), .C2(n10290), .A(n6603), .B(
        n6602), .ZN(n6604) );
  NAND2_X1 U7803 ( .A1(n6605), .A2(n6604), .ZN(P1_U3252) );
  INV_X1 U7804 ( .A(n7706), .ZN(n6613) );
  NOR2_X1 U7805 ( .A1(n6606), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n6756) );
  OR2_X1 U7806 ( .A1(n6756), .A2(n6162), .ZN(n6609) );
  INV_X1 U7807 ( .A(n6609), .ZN(n6607) );
  NAND2_X1 U7808 ( .A1(n6607), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6610) );
  INV_X1 U7809 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6608) );
  NAND2_X1 U7810 ( .A1(n6609), .A2(n6608), .ZN(n6689) );
  AOI22_X1 U7811 ( .A1(n7707), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9958), .ZN(n6611) );
  OAI21_X1 U7812 ( .B1(n6613), .B2(n8830), .A(n6611), .ZN(P1_U3341) );
  INV_X1 U7813 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6614) );
  OAI222_X1 U7814 ( .A1(n9385), .A2(n6614), .B1(n9380), .B2(n6613), .C1(
        P2_U3152), .C2(n6612), .ZN(P2_U3346) );
  NAND2_X1 U7815 ( .A1(n6629), .A2(n6615), .ZN(n6617) );
  NOR4_X1 U7816 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6626) );
  NOR4_X1 U7817 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6625) );
  OR4_X1 U7818 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6623) );
  NOR4_X1 U7819 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6621) );
  NOR4_X1 U7820 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6620) );
  NOR4_X1 U7821 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6619) );
  NOR4_X1 U7822 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6618) );
  NAND4_X1 U7823 ( .A1(n6621), .A2(n6620), .A3(n6619), .A4(n6618), .ZN(n6622)
         );
  NOR4_X1 U7824 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        n6623), .A4(n6622), .ZN(n6624) );
  NAND3_X1 U7825 ( .A1(n6626), .A2(n6625), .A3(n6624), .ZN(n6627) );
  NAND2_X1 U7826 ( .A1(n6629), .A2(n6627), .ZN(n6673) );
  NAND2_X1 U7827 ( .A1(n7023), .A2(n6673), .ZN(n6631) );
  INV_X1 U7828 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6628) );
  NAND2_X1 U7829 ( .A1(n6629), .A2(n6628), .ZN(n6630) );
  NAND2_X1 U7830 ( .A1(n9964), .A2(n8779), .ZN(n9948) );
  INV_X1 U7831 ( .A(n8530), .ZN(n6662) );
  OR2_X1 U7832 ( .A1(n6666), .A2(n6662), .ZN(n6659) );
  NAND2_X1 U7833 ( .A1(n4917), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6633) );
  NAND2_X1 U7834 ( .A1(n6634), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6636) );
  NOR2_X1 U7835 ( .A1(n6659), .A2(n6677), .ZN(n6745) );
  INV_X1 U7836 ( .A(n6678), .ZN(n8540) );
  NAND2_X1 U7837 ( .A1(n4862), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6642) );
  INV_X1 U7838 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6637) );
  INV_X1 U7839 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7026) );
  OR2_X1 U7840 ( .A1(n6788), .A2(n7026), .ZN(n6644) );
  NAND2_X1 U7841 ( .A1(n4862), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6643) );
  AND2_X1 U7842 ( .A1(n6644), .A2(n6643), .ZN(n6647) );
  OR2_X1 U7843 ( .A1(n8264), .A2(n6677), .ZN(n6649) );
  NAND2_X1 U7844 ( .A1(n6718), .A2(SI_0_), .ZN(n6651) );
  XNOR2_X1 U7845 ( .A(n6651), .B(n6650), .ZN(n9965) );
  MUX2_X1 U7846 ( .A(n10342), .B(n9965), .S(n7049), .Z(n6682) );
  OAI22_X1 U7847 ( .A1(n6682), .A2(n8199), .B1(n10342), .B2(n6780), .ZN(n6654)
         );
  NAND2_X1 U7848 ( .A1(n6676), .A2(n8191), .ZN(n6657) );
  OAI22_X1 U7849 ( .A1(n6682), .A2(n6906), .B1(n6688), .B2(n6780), .ZN(n6655)
         );
  INV_X1 U7850 ( .A(n6655), .ZN(n6656) );
  NAND2_X1 U7851 ( .A1(n6657), .A2(n6656), .ZN(n6729) );
  NAND2_X1 U7852 ( .A1(n6658), .A2(n6729), .ZN(n6731) );
  OAI21_X1 U7853 ( .B1(n6658), .B2(n6729), .A(n6731), .ZN(n10346) );
  INV_X1 U7854 ( .A(n6659), .ZN(n6661) );
  NOR2_X1 U7855 ( .A1(n10501), .A2(n8540), .ZN(n6660) );
  AOI22_X1 U7856 ( .A1(n9523), .A2(n9544), .B1(n10346), .B2(n9485), .ZN(n6671)
         );
  AND2_X1 U7857 ( .A1(n7197), .A2(n6667), .ZN(n10412) );
  INV_X1 U7858 ( .A(n10412), .ZN(n6663) );
  NOR2_X1 U7859 ( .A1(n6663), .A2(n6662), .ZN(n6664) );
  NAND2_X1 U7860 ( .A1(n6666), .A2(n6664), .ZN(n6785) );
  NAND2_X1 U7861 ( .A1(n6666), .A2(n10637), .ZN(n6782) );
  OR2_X1 U7862 ( .A1(n6678), .A2(n8531), .ZN(n6781) );
  NAND3_X1 U7863 ( .A1(n6785), .A2(n6782), .A3(n6672), .ZN(n9487) );
  NAND2_X1 U7864 ( .A1(n10412), .A2(n8530), .ZN(n6665) );
  NAND2_X1 U7865 ( .A1(n8530), .A2(n8525), .ZN(n6668) );
  INV_X1 U7866 ( .A(n6682), .ZN(n10399) );
  AOI22_X1 U7867 ( .A1(n9487), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n9528), .B2(
        n10399), .ZN(n6670) );
  NAND2_X1 U7868 ( .A1(n6671), .A2(n6670), .ZN(P1_U3230) );
  NAND2_X1 U7869 ( .A1(n6673), .A2(n6672), .ZN(n7024) );
  NOR2_X1 U7870 ( .A1(n10504), .A2(n8483), .ZN(n6674) );
  OR3_X1 U7871 ( .A1(n7023), .A2(n7024), .A3(n6674), .ZN(n6685) );
  INV_X1 U7872 ( .A(n7022), .ZN(n6675) );
  INV_X2 U7873 ( .A(n10645), .ZN(n10491) );
  INV_X1 U7874 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6684) );
  INV_X1 U7875 ( .A(n7197), .ZN(n6681) );
  NOR2_X1 U7876 ( .A1(n6676), .A2(n6682), .ZN(n10389) );
  AND2_X1 U7877 ( .A1(n6676), .A2(n6682), .ZN(n8412) );
  NOR2_X1 U7878 ( .A1(n10389), .A2(n8412), .ZN(n8493) );
  OR2_X1 U7879 ( .A1(n6678), .A2(n6677), .ZN(n7115) );
  INV_X1 U7880 ( .A(n7115), .ZN(n6679) );
  NOR3_X1 U7881 ( .A1(n8493), .A2(n6679), .A3(n7197), .ZN(n6680) );
  AOI21_X1 U7882 ( .B1(n10392), .B2(n9544), .A(n6680), .ZN(n7031) );
  OAI21_X1 U7883 ( .B1(n6682), .B2(n6681), .A(n7031), .ZN(n6686) );
  NAND2_X1 U7884 ( .A1(n6686), .A2(n10491), .ZN(n6683) );
  OAI21_X1 U7885 ( .B1(n10491), .B2(n6684), .A(n6683), .ZN(P1_U3454) );
  NAND2_X1 U7886 ( .A1(n6686), .A2(n10644), .ZN(n6687) );
  OAI21_X1 U7887 ( .B1(n10644), .B2(n6688), .A(n6687), .ZN(P1_U3523) );
  INV_X1 U7888 ( .A(n7767), .ZN(n6694) );
  NAND2_X1 U7889 ( .A1(n6689), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6690) );
  XNOR2_X1 U7890 ( .A(n6690), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7768) );
  AOI22_X1 U7891 ( .A1(n7768), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9958), .ZN(n6691) );
  OAI21_X1 U7892 ( .B1(n6694), .B2(n8830), .A(n6691), .ZN(P1_U3340) );
  AOI22_X1 U7893 ( .A1(n6692), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n9373), .ZN(n6693) );
  OAI21_X1 U7894 ( .B1(n6694), .B2(n9380), .A(n6693), .ZN(P2_U3345) );
  AOI22_X1 U7895 ( .A1(n8906), .A2(n8934), .B1(n8917), .B2(n8932), .ZN(n6700)
         );
  OAI21_X1 U7896 ( .B1(n6697), .B2(n6696), .A(n6695), .ZN(n6698) );
  AOI22_X1 U7897 ( .A1(n8918), .A2(n7009), .B1(n8873), .B2(n6698), .ZN(n6699)
         );
  OAI211_X1 U7898 ( .C1(n6701), .C2(n9983), .A(n6700), .B(n6699), .ZN(P2_U3224) );
  XNOR2_X1 U7899 ( .A(n6703), .B(n6702), .ZN(n6707) );
  INV_X1 U7900 ( .A(n8930), .ZN(n6850) );
  OAI22_X1 U7901 ( .A1(n10517), .A2(n6850), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5666), .ZN(n6705) );
  INV_X1 U7902 ( .A(n8918), .ZN(n8883) );
  OAI22_X1 U7903 ( .A1(n8883), .A2(n5158), .B1(n10523), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n6704) );
  AOI211_X1 U7904 ( .C1(n8906), .C2(n8932), .A(n6705), .B(n6704), .ZN(n6706)
         );
  OAI21_X1 U7905 ( .B1(n6707), .B2(n10510), .A(n6706), .ZN(P2_U3220) );
  OAI21_X1 U7906 ( .B1(n6710), .B2(n6709), .A(n6708), .ZN(n6712) );
  XOR2_X1 U7907 ( .A(n6712), .B(n6711), .Z(n6717) );
  INV_X1 U7908 ( .A(n9249), .ZN(n6975) );
  OAI21_X1 U7909 ( .B1(n10517), .B2(n6975), .A(n6713), .ZN(n6715) );
  INV_X1 U7910 ( .A(n7089), .ZN(n10460) );
  OAI22_X1 U7911 ( .A1(n8883), .A2(n10460), .B1(n7083), .B2(n10523), .ZN(n6714) );
  AOI211_X1 U7912 ( .C1(n8906), .C2(n8931), .A(n6715), .B(n6714), .ZN(n6716)
         );
  OAI21_X1 U7913 ( .B1(n6717), .B2(n10510), .A(n6716), .ZN(P2_U3232) );
  NAND2_X1 U7914 ( .A1(n7101), .A2(n8191), .ZN(n6726) );
  NAND2_X1 U7915 ( .A1(n10413), .A2(n8184), .ZN(n6725) );
  NAND2_X1 U7916 ( .A1(n6726), .A2(n6725), .ZN(n6728) );
  NAND2_X1 U7917 ( .A1(n8264), .A2(n9781), .ZN(n6727) );
  INV_X1 U7919 ( .A(n6729), .ZN(n6730) );
  NAND2_X1 U7920 ( .A1(n6730), .A2(n8197), .ZN(n6732) );
  NAND2_X1 U7921 ( .A1(n6732), .A2(n6731), .ZN(n6738) );
  XNOR2_X1 U7922 ( .A(n6739), .B(n6738), .ZN(n6736) );
  NAND2_X1 U7923 ( .A1(n9544), .A2(n8155), .ZN(n6734) );
  NAND2_X1 U7924 ( .A1(n10413), .A2(n8191), .ZN(n6733) );
  NAND2_X1 U7925 ( .A1(n6734), .A2(n6733), .ZN(n6742) );
  INV_X1 U7926 ( .A(n6742), .ZN(n6735) );
  NAND2_X1 U7927 ( .A1(n6736), .A2(n6735), .ZN(n6744) );
  NAND2_X1 U7928 ( .A1(n6738), .A2(n6739), .ZN(n6737) );
  NAND2_X1 U7929 ( .A1(n6737), .A2(n6742), .ZN(n6804) );
  NAND2_X1 U7930 ( .A1(n6741), .A2(n6740), .ZN(n6803) );
  INV_X1 U7931 ( .A(n6803), .ZN(n6743) );
  AOI22_X1 U7932 ( .A1(n6744), .A2(n6804), .B1(n6743), .B2(n6742), .ZN(n6753)
         );
  AOI22_X1 U7933 ( .A1(n9487), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n9528), .B2(
        n10413), .ZN(n6752) );
  INV_X1 U7934 ( .A(n9521), .ZN(n9488) );
  NAND2_X1 U7935 ( .A1(n6746), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6750) );
  INV_X1 U7936 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7224) );
  OR2_X1 U7937 ( .A1(n6788), .A2(n7224), .ZN(n6748) );
  NAND2_X1 U7938 ( .A1(n4862), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6747) );
  AOI22_X1 U7939 ( .A1(n9488), .A2(n6676), .B1(n9523), .B2(n6813), .ZN(n6751)
         );
  OAI211_X1 U7940 ( .C1(n6753), .C2(n9530), .A(n6752), .B(n6751), .ZN(P1_U3220) );
  AOI22_X1 U7941 ( .A1(n7589), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n9373), .ZN(n6754) );
  OAI21_X1 U7942 ( .B1(n7849), .B2(n9380), .A(n6754), .ZN(P2_U3344) );
  INV_X1 U7943 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6760) );
  NOR2_X1 U7944 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n6755) );
  NAND2_X1 U7945 ( .A1(n6756), .A2(n6755), .ZN(n6758) );
  NAND2_X1 U7946 ( .A1(n6758), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6757) );
  MUX2_X1 U7947 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6757), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n6759) );
  INV_X1 U7948 ( .A(n10253), .ZN(n7310) );
  OAI222_X1 U7949 ( .A1(n9961), .A2(n6760), .B1(n8830), .B2(n7849), .C1(n7310), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  AOI21_X1 U7950 ( .B1(n8768), .B2(n8934), .A(n10510), .ZN(n6761) );
  NOR2_X1 U7951 ( .A1(n8918), .A2(n6761), .ZN(n6763) );
  NOR2_X1 U7952 ( .A1(n10510), .A2(n6870), .ZN(n8875) );
  NAND2_X1 U7953 ( .A1(n8875), .A2(n8934), .ZN(n6762) );
  MUX2_X1 U7954 ( .A(n6763), .B(n6762), .S(n10381), .Z(n6766) );
  NAND2_X1 U7955 ( .A1(n6764), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6765) );
  OAI211_X1 U7956 ( .C1(n6773), .C2(n10378), .A(n6766), .B(n6765), .ZN(
        P2_U3234) );
  NAND2_X1 U7957 ( .A1(n6767), .A2(n6769), .ZN(n6768) );
  AOI21_X1 U7958 ( .B1(n6971), .B2(n6768), .A(n10510), .ZN(n6779) );
  NAND4_X1 U7959 ( .A1(n6711), .A2(n8875), .A3(n6769), .A4(n8930), .ZN(n6777)
         );
  INV_X1 U7960 ( .A(n6988), .ZN(n6775) );
  NAND2_X1 U7961 ( .A1(n8929), .A2(n10587), .ZN(n6771) );
  NAND2_X1 U7962 ( .A1(n8930), .A2(n9230), .ZN(n6770) );
  NAND2_X1 U7963 ( .A1(n6771), .A2(n6770), .ZN(n6984) );
  INV_X1 U7964 ( .A(n6984), .ZN(n6772) );
  INV_X1 U7965 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10181) );
  OAI22_X1 U7966 ( .A1(n6773), .A2(n6772), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10181), .ZN(n6774) );
  AOI21_X1 U7967 ( .B1(n8886), .B2(n6775), .A(n6774), .ZN(n6776) );
  OAI211_X1 U7968 ( .C1(n6989), .C2(n8883), .A(n6777), .B(n6776), .ZN(n6778)
         );
  OR2_X1 U7969 ( .A1(n6779), .A2(n6778), .ZN(P2_U3229) );
  AND3_X1 U7970 ( .A1(n6781), .A2(n6780), .A3(n7823), .ZN(n6783) );
  NAND2_X1 U7971 ( .A1(n6783), .A2(n6782), .ZN(n6784) );
  NAND2_X1 U7972 ( .A1(n6784), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6786) );
  NAND2_X1 U7973 ( .A1(n4862), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6793) );
  NAND2_X1 U7974 ( .A1(n6954), .A2(n8191), .ZN(n6801) );
  OR2_X1 U7975 ( .A1(n4864), .A2(n6794), .ZN(n6799) );
  OR2_X1 U7976 ( .A1(n6899), .A2(n6795), .ZN(n6798) );
  OR2_X1 U7977 ( .A1(n7049), .A2(n6796), .ZN(n6797) );
  OR2_X1 U7978 ( .A1(n10443), .A2(n6906), .ZN(n6800) );
  NAND2_X1 U7979 ( .A1(n6801), .A2(n6800), .ZN(n6802) );
  INV_X1 U7980 ( .A(n10443), .ZN(n7193) );
  AOI22_X1 U7981 ( .A1(n6954), .A2(n8155), .B1(n7193), .B2(n8191), .ZN(n6891)
         );
  NAND2_X1 U7982 ( .A1(n6813), .A2(n8191), .ZN(n6811) );
  OR2_X1 U7983 ( .A1(n6899), .A2(n6806), .ZN(n6808) );
  OR2_X1 U7984 ( .A1(n7049), .A2(n10352), .ZN(n6807) );
  NAND2_X1 U7985 ( .A1(n6811), .A2(n6810), .ZN(n6812) );
  AND2_X1 U7986 ( .A1(n4898), .A2(n6816), .ZN(n9484) );
  NAND2_X1 U7987 ( .A1(n6818), .A2(n9484), .ZN(n9483) );
  NAND2_X1 U7988 ( .A1(n9483), .A2(n6816), .ZN(n6819) );
  AND2_X1 U7989 ( .A1(n6893), .A2(n6894), .ZN(n6950) );
  OAI21_X1 U7990 ( .B1(n6820), .B2(n6819), .A(n6950), .ZN(n6821) );
  NAND2_X1 U7991 ( .A1(n6821), .A2(n9485), .ZN(n6827) );
  INV_X1 U7992 ( .A(n6813), .ZN(n6824) );
  AOI21_X1 U7993 ( .B1(n9528), .B2(n7193), .A(n6822), .ZN(n6823) );
  OAI21_X1 U7994 ( .B1(n9521), .B2(n6824), .A(n6823), .ZN(n6825) );
  AOI21_X1 U7995 ( .B1(n9523), .B2(n6883), .A(n6825), .ZN(n6826) );
  OAI211_X1 U7996 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9526), .A(n6827), .B(
        n6826), .ZN(P1_U3216) );
  INV_X1 U7997 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6839) );
  NAND2_X1 U7998 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7707), .ZN(n6828) );
  OAI21_X1 U7999 ( .B1(n7707), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6828), .ZN(
        n6925) );
  NOR2_X1 U8000 ( .A1(n6925), .A2(n6926), .ZN(n6924) );
  AOI21_X1 U8001 ( .B1(n7707), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6924), .ZN(
        n6831) );
  NAND2_X1 U8002 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7768), .ZN(n6829) );
  OAI21_X1 U8003 ( .B1(n7768), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6829), .ZN(
        n6830) );
  NOR2_X1 U8004 ( .A1(n6831), .A2(n6830), .ZN(n7307) );
  AOI211_X1 U8005 ( .C1(n6831), .C2(n6830), .A(n7307), .B(n10370), .ZN(n6832)
         );
  AOI21_X1 U8006 ( .B1(n10288), .B2(n7768), .A(n6832), .ZN(n6838) );
  INV_X1 U8007 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7721) );
  MUX2_X1 U8008 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7721), .S(n7768), .Z(n6835)
         );
  INV_X1 U8009 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7559) );
  MUX2_X1 U8010 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7559), .S(n7707), .Z(n6920)
         );
  OAI21_X1 U8011 ( .B1(n7527), .B2(P1_REG1_REG_11__SCAN_IN), .A(n6833), .ZN(
        n6919) );
  NAND2_X1 U8012 ( .A1(n6920), .A2(n6919), .ZN(n6918) );
  OAI21_X1 U8013 ( .B1(n7707), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6918), .ZN(
        n6834) );
  NAND2_X1 U8014 ( .A1(n6835), .A2(n6834), .ZN(n7311) );
  OAI21_X1 U8015 ( .B1(n6835), .B2(n6834), .A(n7311), .ZN(n6836) );
  AND2_X1 U8016 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7780) );
  AOI21_X1 U8017 ( .B1(n10368), .B2(n6836), .A(n7780), .ZN(n6837) );
  OAI211_X1 U8018 ( .C1(n10376), .C2(n6839), .A(n6838), .B(n6837), .ZN(
        P1_U3254) );
  INV_X1 U8019 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6858) );
  OAI21_X1 U8020 ( .B1(n4859), .B2(n7009), .A(n6840), .ZN(n6842) );
  NAND2_X1 U8021 ( .A1(n4859), .A2(n7009), .ZN(n6841) );
  AND2_X2 U8022 ( .A1(n6842), .A2(n6841), .ZN(n7035) );
  NAND2_X1 U8023 ( .A1(n6849), .A2(n6843), .ZN(n8598) );
  NAND2_X1 U8024 ( .A1(n6849), .A2(n10436), .ZN(n6844) );
  NAND2_X1 U8025 ( .A1(n7034), .A2(n6844), .ZN(n6845) );
  NAND2_X1 U8026 ( .A1(n6976), .A2(n6855), .ZN(n8602) );
  NAND2_X1 U8027 ( .A1(n8931), .A2(n5158), .ZN(n8603) );
  NAND2_X1 U8028 ( .A1(n8602), .A2(n8603), .ZN(n8740) );
  OR2_X1 U8029 ( .A1(n6845), .A2(n8740), .ZN(n6846) );
  NAND2_X1 U8030 ( .A1(n6845), .A2(n8740), .ZN(n6978) );
  INV_X1 U8031 ( .A(n8740), .ZN(n8600) );
  NAND2_X1 U8032 ( .A1(n8590), .A2(n6847), .ZN(n7033) );
  NAND2_X1 U8033 ( .A1(n8597), .A2(n8598), .ZN(n6848) );
  NAND2_X1 U8034 ( .A1(n6848), .A2(n8600), .ZN(n6981) );
  OAI21_X1 U8035 ( .B1(n8600), .B2(n6848), .A(n6981), .ZN(n6853) );
  OAI22_X1 U8036 ( .A1(n6850), .A2(n9214), .B1(n6849), .B2(n9216), .ZN(n6852)
         );
  NOR2_X1 U8037 ( .A1(n6882), .A2(n7474), .ZN(n6851) );
  AOI211_X1 U8038 ( .C1(n9234), .C2(n6853), .A(n6852), .B(n6851), .ZN(n6868)
         );
  NAND2_X1 U8039 ( .A1(n7040), .A2(n6855), .ZN(n6854) );
  AND2_X1 U8040 ( .A1(n7084), .A2(n6854), .ZN(n6872) );
  AOI22_X1 U8041 ( .A1(n6872), .A2(n10629), .B1(n10628), .B2(n6855), .ZN(n6856) );
  OAI211_X1 U8042 ( .C1(n6882), .C2(n10435), .A(n6868), .B(n6856), .ZN(n6859)
         );
  NAND2_X1 U8043 ( .A1(n6859), .A2(n10660), .ZN(n6857) );
  OAI21_X1 U8044 ( .B1(n10660), .B2(n6858), .A(n6857), .ZN(P2_U3460) );
  NAND2_X1 U8045 ( .A1(n6859), .A2(n10657), .ZN(n6860) );
  OAI21_X1 U8046 ( .B1(n10657), .B2(n5642), .A(n6860), .ZN(P2_U3523) );
  NAND3_X1 U8047 ( .A1(n6863), .A2(n6862), .A3(n6861), .ZN(n6869) );
  INV_X1 U8048 ( .A(n8587), .ZN(n6866) );
  NAND2_X1 U8049 ( .A1(n6866), .A2(n6098), .ZN(n6974) );
  INV_X1 U8050 ( .A(n6974), .ZN(n6867) );
  NAND2_X1 U8051 ( .A1(n10605), .A2(n6867), .ZN(n7482) );
  OR2_X1 U8052 ( .A1(n6868), .A2(n10607), .ZN(n6881) );
  INV_X1 U8053 ( .A(n6869), .ZN(n6871) );
  NAND2_X1 U8054 ( .A1(n6871), .A2(n6870), .ZN(n10382) );
  INV_X1 U8055 ( .A(n6872), .ZN(n6876) );
  OR2_X1 U8056 ( .A1(n10605), .A2(n6873), .ZN(n6875) );
  INV_X1 U8057 ( .A(n10609), .ZN(n9238) );
  NAND2_X1 U8058 ( .A1(n9238), .A2(n5666), .ZN(n6874) );
  OAI211_X1 U8059 ( .C1(n10382), .C2(n6876), .A(n6875), .B(n6874), .ZN(n6879)
         );
  NOR2_X1 U8060 ( .A1(n6098), .A2(n6877), .ZN(n10599) );
  NOR2_X1 U8061 ( .A1(n10383), .A2(n5158), .ZN(n6878) );
  NOR2_X1 U8062 ( .A1(n6879), .A2(n6878), .ZN(n6880) );
  OAI211_X1 U8063 ( .C1(n6882), .C2(n7482), .A(n6881), .B(n6880), .ZN(P2_U3293) );
  NAND2_X1 U8064 ( .A1(n6883), .A2(n8191), .ZN(n6889) );
  OR2_X1 U8065 ( .A1(n6899), .A2(n6884), .ZN(n6888) );
  OR2_X1 U8066 ( .A1(n7049), .A2(n10363), .ZN(n6886) );
  XNOR2_X1 U8067 ( .A(n6895), .B(n6896), .ZN(n6952) );
  INV_X1 U8068 ( .A(n6890), .ZN(n6892) );
  NAND2_X1 U8069 ( .A1(n6892), .A2(n6891), .ZN(n6949) );
  INV_X1 U8070 ( .A(n6895), .ZN(n6897) );
  OR2_X1 U8071 ( .A1(n6897), .A2(n6896), .ZN(n6898) );
  NAND2_X1 U8072 ( .A1(n7322), .A2(n8191), .ZN(n6908) );
  OR2_X1 U8073 ( .A1(n6899), .A2(n6900), .ZN(n6905) );
  OR2_X1 U8074 ( .A1(n4864), .A2(n6902), .ZN(n6904) );
  OR2_X1 U8075 ( .A1(n7049), .A2(n10274), .ZN(n6903) );
  OR2_X1 U8076 ( .A1(n10468), .A2(n6906), .ZN(n6907) );
  NAND2_X1 U8077 ( .A1(n6908), .A2(n6907), .ZN(n6909) );
  XNOR2_X1 U8078 ( .A(n6909), .B(n8188), .ZN(n7065) );
  NAND2_X1 U8079 ( .A1(n7322), .A2(n8155), .ZN(n6911) );
  OR2_X1 U8080 ( .A1(n10468), .A2(n8199), .ZN(n6910) );
  AND2_X1 U8081 ( .A1(n6911), .A2(n6910), .ZN(n7062) );
  INV_X1 U8082 ( .A(n7062), .ZN(n7066) );
  XNOR2_X1 U8083 ( .A(n7065), .B(n7066), .ZN(n6912) );
  XNOR2_X1 U8084 ( .A(n7064), .B(n6912), .ZN(n6917) );
  NOR2_X1 U8085 ( .A1(n9526), .A2(n7211), .ZN(n6915) );
  INV_X1 U8086 ( .A(n9523), .ZN(n9507) );
  INV_X1 U8087 ( .A(n7290), .ZN(n7376) );
  AND2_X1 U8088 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10271) );
  AOI21_X1 U8089 ( .B1(n9528), .B2(n7287), .A(n10271), .ZN(n6913) );
  OAI21_X1 U8090 ( .B1(n9507), .B2(n7376), .A(n6913), .ZN(n6914) );
  AOI211_X1 U8091 ( .C1(n9488), .C2(n6883), .A(n6915), .B(n6914), .ZN(n6916)
         );
  OAI21_X1 U8092 ( .B1(n6917), .B2(n9530), .A(n6916), .ZN(P1_U3225) );
  INV_X1 U8093 ( .A(n7707), .ZN(n6923) );
  OAI21_X1 U8094 ( .B1(n6920), .B2(n6919), .A(n6918), .ZN(n6921) );
  NAND2_X1 U8095 ( .A1(n10368), .A2(n6921), .ZN(n6922) );
  NAND2_X1 U8096 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7726) );
  OAI211_X1 U8097 ( .C1(n10364), .C2(n6923), .A(n6922), .B(n7726), .ZN(n6928)
         );
  AOI211_X1 U8098 ( .C1(n6926), .C2(n6925), .A(n6924), .B(n10370), .ZN(n6927)
         );
  AOI211_X1 U8099 ( .C1(P1_ADDR_REG_12__SCAN_IN), .C2(n10290), .A(n6928), .B(
        n6927), .ZN(n6929) );
  INV_X1 U8100 ( .A(n6929), .ZN(P1_U3253) );
  INV_X1 U8101 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9378) );
  INV_X1 U8102 ( .A(n7146), .ZN(n6930) );
  NAND2_X1 U8103 ( .A1(n6930), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7273) );
  INV_X1 U8104 ( .A(n7509), .ZN(n6931) );
  NAND2_X1 U8105 ( .A1(n6931), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7561) );
  INV_X1 U8106 ( .A(n7561), .ZN(n6932) );
  NAND2_X1 U8107 ( .A1(n6932), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7719) );
  INV_X1 U8108 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7854) );
  INV_X1 U8109 ( .A(n8035), .ZN(n6936) );
  NAND2_X1 U8110 ( .A1(n6936), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8055) );
  INV_X1 U8111 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8054) );
  INV_X1 U8112 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8076) );
  INV_X1 U8113 ( .A(n8111), .ZN(n6938) );
  NAND2_X1 U8114 ( .A1(n6938), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8123) );
  INV_X1 U8115 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8122) );
  INV_X1 U8116 ( .A(n8143), .ZN(n6939) );
  NAND2_X1 U8117 ( .A1(n6939), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8163) );
  INV_X1 U8118 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9506) );
  INV_X1 U8119 ( .A(n8165), .ZN(n6941) );
  AND2_X1 U8120 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .ZN(n6940) );
  NAND2_X1 U8121 ( .A1(n6941), .A2(n6940), .ZN(n8801) );
  OR2_X1 U8122 ( .A1(n8801), .A2(n8145), .ZN(n6947) );
  INV_X1 U8123 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6944) );
  NAND2_X1 U8124 ( .A1(n4862), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6943) );
  NAND2_X1 U8125 ( .A1(n8095), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6942) );
  OAI211_X1 U8126 ( .C1(n6944), .C2(n6787), .A(n6943), .B(n6942), .ZN(n6945)
         );
  INV_X1 U8127 ( .A(n6945), .ZN(n6946) );
  NAND2_X1 U8128 ( .A1(n6947), .A2(n6946), .ZN(n9621) );
  NAND2_X1 U8129 ( .A1(n9621), .A2(P1_U4006), .ZN(n6948) );
  OAI21_X1 U8130 ( .B1(n9378), .B2(P1_U4006), .A(n6948), .ZN(P1_U3584) );
  AND2_X1 U8131 ( .A1(n6950), .A2(n6949), .ZN(n6953) );
  OAI211_X1 U8132 ( .C1(n6953), .C2(n6952), .A(n9485), .B(n6951), .ZN(n6959)
         );
  INV_X1 U8133 ( .A(n7322), .ZN(n6956) );
  AND2_X1 U8134 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10366) );
  AOI21_X1 U8135 ( .B1(n9528), .B2(n7206), .A(n10366), .ZN(n6955) );
  OAI21_X1 U8136 ( .B1(n9507), .B2(n6956), .A(n6955), .ZN(n6957) );
  AOI21_X1 U8137 ( .B1(n9488), .B2(n6954), .A(n6957), .ZN(n6958) );
  OAI211_X1 U8138 ( .C1(n9526), .C2(n7120), .A(n6959), .B(n6958), .ZN(P1_U3228) );
  NAND2_X1 U8139 ( .A1(n8906), .A2(n9249), .ZN(n6962) );
  OAI211_X1 U8140 ( .C1(n7256), .C2(n10517), .A(n6962), .B(n6961), .ZN(n6965)
         );
  NAND2_X1 U8141 ( .A1(n8918), .A2(n10492), .ZN(n6963) );
  OAI21_X1 U8142 ( .B1(n10523), .B2(n9257), .A(n6963), .ZN(n6964) );
  NOR2_X1 U8143 ( .A1(n6965), .A2(n6964), .ZN(n6973) );
  INV_X1 U8144 ( .A(n6966), .ZN(n6970) );
  NAND2_X1 U8145 ( .A1(n8875), .A2(n9249), .ZN(n6967) );
  OAI21_X1 U8146 ( .B1(n10510), .B2(n6968), .A(n6967), .ZN(n6969) );
  NAND3_X1 U8147 ( .A1(n6971), .A2(n6970), .A3(n6969), .ZN(n6972) );
  OAI211_X1 U8148 ( .C1(n6960), .C2(n10510), .A(n6973), .B(n6972), .ZN(
        P2_U3241) );
  NAND2_X1 U8149 ( .A1(n7474), .A2(n6974), .ZN(n10596) );
  NAND2_X1 U8150 ( .A1(n6989), .A2(n9249), .ZN(n8607) );
  NAND2_X1 U8151 ( .A1(n6975), .A2(n10475), .ZN(n8611) );
  NAND2_X1 U8152 ( .A1(n6976), .A2(n5158), .ZN(n6977) );
  XNOR2_X1 U8153 ( .A(n8930), .B(n7089), .ZN(n8743) );
  NAND2_X1 U8154 ( .A1(n8930), .A2(n7089), .ZN(n6980) );
  XOR2_X1 U8155 ( .A(n8744), .B(n7233), .Z(n10478) );
  INV_X1 U8156 ( .A(n8743), .ZN(n6982) );
  NAND2_X1 U8157 ( .A1(n8930), .A2(n10460), .ZN(n8609) );
  NAND2_X1 U8158 ( .A1(n6983), .A2(n8609), .ZN(n7238) );
  XOR2_X1 U8159 ( .A(n8744), .B(n7238), .Z(n6985) );
  AOI21_X1 U8160 ( .B1(n6985), .B2(n9234), .A(n6984), .ZN(n10477) );
  MUX2_X1 U8161 ( .A(n10477), .B(n6986), .S(n10607), .Z(n6992) );
  INV_X1 U8162 ( .A(n6987), .ZN(n7085) );
  AOI211_X1 U8163 ( .C1(n10475), .C2(n7085), .A(n10650), .B(n9253), .ZN(n10474) );
  AND2_X1 U8164 ( .A1(n10605), .A2(n5582), .ZN(n9186) );
  OAI22_X1 U8165 ( .A1(n10383), .A2(n6989), .B1(n6988), .B2(n10609), .ZN(n6990) );
  AOI21_X1 U8166 ( .B1(n10474), .B2(n9186), .A(n6990), .ZN(n6991) );
  OAI211_X1 U8167 ( .C1(n9244), .C2(n10478), .A(n6992), .B(n6991), .ZN(
        P2_U3291) );
  INV_X1 U8168 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7000) );
  XNOR2_X1 U8169 ( .A(n8165), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9643) );
  NAND2_X1 U8170 ( .A1(n9643), .A2(n8166), .ZN(n6998) );
  INV_X1 U8171 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6995) );
  NAND2_X1 U8172 ( .A1(n4862), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6994) );
  NAND2_X1 U8173 ( .A1(n6746), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6993) );
  OAI211_X1 U8174 ( .C1(n6995), .C2(n7853), .A(n6994), .B(n6993), .ZN(n6996)
         );
  INV_X1 U8175 ( .A(n6996), .ZN(n6997) );
  NAND2_X1 U8176 ( .A1(n9622), .A2(P1_U4006), .ZN(n6999) );
  OAI21_X1 U8177 ( .B1(P1_U4006), .B2(n7000), .A(n6999), .ZN(P1_U3582) );
  INV_X1 U8178 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7002) );
  INV_X1 U8179 ( .A(n7894), .ZN(n7004) );
  NAND2_X1 U8180 ( .A1(n7094), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7001) );
  XNOR2_X1 U8181 ( .A(n7001), .B(n4980), .ZN(n9553) );
  OAI222_X1 U8182 ( .A1(n9961), .A2(n7002), .B1(n8830), .B2(n7004), .C1(
        P1_U3084), .C2(n9553), .ZN(P1_U3338) );
  INV_X1 U8183 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7005) );
  OAI222_X1 U8184 ( .A1(n9385), .A2(n7005), .B1(n9380), .B2(n7004), .C1(
        P2_U3152), .C2(n7003), .ZN(P2_U3343) );
  OAI22_X1 U8185 ( .A1(n10382), .A2(n7006), .B1(n9983), .B2(n10609), .ZN(n7007) );
  AOI21_X1 U8186 ( .B1(n10607), .B2(P2_REG2_REG_1__SCAN_IN), .A(n7007), .ZN(
        n7011) );
  AOI22_X1 U8187 ( .A1(n9223), .A2(n7009), .B1(n7008), .B2(n10605), .ZN(n7010)
         );
  OAI211_X1 U8188 ( .C1(n7012), .C2(n9244), .A(n7011), .B(n7010), .ZN(P2_U3295) );
  INV_X1 U8189 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7021) );
  INV_X1 U8190 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9395) );
  INV_X1 U8191 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7013) );
  OAI21_X1 U8192 ( .B1(n8165), .B2(n9395), .A(n7013), .ZN(n7014) );
  NAND2_X1 U8193 ( .A1(n7014), .A2(n8801), .ZN(n9629) );
  OR2_X1 U8194 ( .A1(n9629), .A2(n8145), .ZN(n7019) );
  INV_X1 U8195 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9628) );
  NAND2_X1 U8196 ( .A1(n4862), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n7016) );
  NAND2_X1 U8197 ( .A1(n6746), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n7015) );
  OAI211_X1 U8198 ( .C1(n9628), .C2(n7853), .A(n7016), .B(n7015), .ZN(n7017)
         );
  INV_X1 U8199 ( .A(n7017), .ZN(n7018) );
  NAND2_X1 U8200 ( .A1(n5107), .A2(P1_U4006), .ZN(n7020) );
  OAI21_X1 U8201 ( .B1(P1_U4006), .B2(n7021), .A(n7020), .ZN(P1_U3583) );
  NAND2_X1 U8202 ( .A1(n7023), .A2(n7022), .ZN(n7025) );
  OAI22_X1 U8203 ( .A1(n9822), .A2(n10291), .B1(n7026), .B2(n9819), .ZN(n7027)
         );
  INV_X1 U8204 ( .A(n7027), .ZN(n7030) );
  AND2_X1 U8205 ( .A1(n7197), .A2(n8531), .ZN(n7028) );
  OAI21_X1 U8206 ( .B1(n9825), .B2(n9785), .A(n10399), .ZN(n7029) );
  OAI211_X1 U8207 ( .C1(n7031), .C2(n10425), .A(n7030), .B(n7029), .ZN(
        P1_U3291) );
  INV_X1 U8208 ( .A(n8597), .ZN(n7032) );
  AOI21_X1 U8209 ( .B1(n8741), .B2(n7033), .A(n7032), .ZN(n7039) );
  AOI22_X1 U8210 ( .A1(n8931), .A2(n10587), .B1(n9230), .B2(n4859), .ZN(n7038)
         );
  OAI21_X1 U8211 ( .B1(n7035), .B2(n8741), .A(n7034), .ZN(n10440) );
  INV_X1 U8212 ( .A(n7474), .ZN(n7036) );
  NAND2_X1 U8213 ( .A1(n10440), .A2(n7036), .ZN(n7037) );
  OAI211_X1 U8214 ( .C1(n7039), .C2(n7255), .A(n7038), .B(n7037), .ZN(n10438)
         );
  INV_X1 U8215 ( .A(n10438), .ZN(n7047) );
  OAI21_X1 U8216 ( .B1(n7041), .B2(n10436), .A(n7040), .ZN(n10437) );
  OAI22_X1 U8217 ( .A1(n10382), .A2(n10437), .B1(n7042), .B2(n10609), .ZN(
        n7045) );
  INV_X1 U8218 ( .A(n10440), .ZN(n7043) );
  OAI22_X1 U8219 ( .A1(n7043), .A2(n7482), .B1(n10436), .B2(n10383), .ZN(n7044) );
  AOI211_X1 U8220 ( .C1(P2_REG2_REG_2__SCAN_IN), .C2(n10607), .A(n7045), .B(
        n7044), .ZN(n7046) );
  OAI21_X1 U8221 ( .B1(n10607), .B2(n7047), .A(n7046), .ZN(P2_U3294) );
  INV_X1 U8222 ( .A(n7927), .ZN(n7126) );
  AOI22_X1 U8223 ( .A1(n8951), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n9373), .ZN(n7048) );
  OAI21_X1 U8224 ( .B1(n7126), .B2(n9380), .A(n7048), .ZN(P2_U3342) );
  NAND2_X1 U8225 ( .A1(n7290), .A2(n8191), .ZN(n7055) );
  AOI22_X1 U8226 ( .A1(n8029), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8028), .B2(
        n7050), .ZN(n7053) );
  NAND2_X1 U8227 ( .A1(n7051), .A2(n8355), .ZN(n7052) );
  OR2_X1 U8228 ( .A1(n10485), .A2(n6906), .ZN(n7054) );
  NAND2_X1 U8229 ( .A1(n7055), .A2(n7054), .ZN(n7056) );
  NAND2_X1 U8230 ( .A1(n7290), .A2(n8155), .ZN(n7058) );
  OR2_X1 U8231 ( .A1(n10485), .A2(n8199), .ZN(n7057) );
  AND2_X1 U8232 ( .A1(n7058), .A2(n7057), .ZN(n7059) );
  NAND2_X1 U8233 ( .A1(n7065), .A2(n7062), .ZN(n7063) );
  INV_X1 U8234 ( .A(n7065), .ZN(n7067) );
  NAND2_X1 U8235 ( .A1(n7067), .A2(n7066), .ZN(n7068) );
  OR2_X1 U8236 ( .A1(n7138), .A2(n7137), .ZN(n7136) );
  INV_X1 U8237 ( .A(n7136), .ZN(n7069) );
  AOI21_X1 U8238 ( .B1(n7137), .B2(n7138), .A(n7069), .ZN(n7075) );
  OAI22_X1 U8239 ( .A1(n9507), .A2(n5130), .B1(n10485), .B2(n9513), .ZN(n7070)
         );
  AOI211_X1 U8240 ( .C1(n9488), .C2(n7322), .A(n7071), .B(n7070), .ZN(n7074)
         );
  INV_X1 U8241 ( .A(n9526), .ZN(n9510) );
  INV_X1 U8242 ( .A(n7327), .ZN(n7072) );
  NAND2_X1 U8243 ( .A1(n9510), .A2(n7072), .ZN(n7073) );
  OAI211_X1 U8244 ( .C1(n7075), .C2(n9530), .A(n7074), .B(n7073), .ZN(P1_U3237) );
  XNOR2_X1 U8245 ( .A(n7076), .B(n8743), .ZN(n7077) );
  INV_X2 U8246 ( .A(n7255), .ZN(n9234) );
  NAND2_X1 U8247 ( .A1(n7077), .A2(n9234), .ZN(n7079) );
  AOI22_X1 U8248 ( .A1(n8931), .A2(n9230), .B1(n10587), .B2(n9249), .ZN(n7078)
         );
  NAND2_X1 U8249 ( .A1(n7079), .A2(n7078), .ZN(n10462) );
  INV_X1 U8250 ( .A(n10462), .ZN(n7092) );
  INV_X1 U8251 ( .A(n7080), .ZN(n7081) );
  AOI21_X1 U8252 ( .B1(n8743), .B2(n7082), .A(n7081), .ZN(n10464) );
  NAND2_X1 U8253 ( .A1(n10464), .A2(n9263), .ZN(n7091) );
  OAI22_X1 U8254 ( .A1(n7083), .A2(n10609), .B1(n6206), .B2(n10605), .ZN(n7088) );
  INV_X1 U8255 ( .A(n7084), .ZN(n7086) );
  OAI21_X1 U8256 ( .B1(n10460), .B2(n7086), .A(n7085), .ZN(n10461) );
  NOR2_X1 U8257 ( .A1(n10461), .A2(n10382), .ZN(n7087) );
  AOI211_X1 U8258 ( .C1(n9223), .C2(n7089), .A(n7088), .B(n7087), .ZN(n7090)
         );
  OAI211_X1 U8259 ( .C1(n7092), .C2(n10607), .A(n7091), .B(n7090), .ZN(
        P2_U3292) );
  AOI22_X1 U8260 ( .A1(n8974), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n9373), .ZN(n7093) );
  OAI21_X1 U8261 ( .B1(n8021), .B2(n9380), .A(n7093), .ZN(P2_U3341) );
  NAND2_X1 U8262 ( .A1(n7095), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7125) );
  INV_X1 U8263 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n7096) );
  AOI21_X1 U8264 ( .B1(n7125), .B2(n7096), .A(n6162), .ZN(n7097) );
  NAND2_X1 U8265 ( .A1(n7097), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n7099) );
  INV_X1 U8266 ( .A(n7097), .ZN(n7098) );
  NAND2_X1 U8267 ( .A1(n7098), .A2(n4979), .ZN(n7230) );
  AOI22_X1 U8268 ( .A1(n9588), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9958), .ZN(n7100) );
  OAI21_X1 U8269 ( .B1(n8021), .B2(n8830), .A(n7100), .ZN(P1_U3336) );
  OR2_X1 U8270 ( .A1(n9544), .A2(n5013), .ZN(n7102) );
  NAND2_X1 U8271 ( .A1(n6813), .A2(n7225), .ZN(n8417) );
  NAND2_X1 U8272 ( .A1(n8415), .A2(n8417), .ZN(n7109) );
  OR2_X1 U8273 ( .A1(n6954), .A2(n10443), .ZN(n8420) );
  NAND2_X1 U8274 ( .A1(n6954), .A2(n10443), .ZN(n8422) );
  NAND2_X1 U8275 ( .A1(n6883), .A2(n10452), .ZN(n8423) );
  NAND2_X1 U8276 ( .A1(n4892), .A2(n8423), .ZN(n7204) );
  INV_X1 U8277 ( .A(n7204), .ZN(n8492) );
  XNOR2_X1 U8278 ( .A(n7200), .B(n8492), .ZN(n7104) );
  NAND2_X1 U8279 ( .A1(n8264), .A2(n10415), .ZN(n7103) );
  OR2_X1 U8280 ( .A1(n6648), .A2(n8525), .ZN(n8263) );
  NAND2_X1 U8281 ( .A1(n7104), .A2(n10397), .ZN(n7106) );
  AOI22_X1 U8282 ( .A1(n10393), .A2(n6954), .B1(n7322), .B2(n10392), .ZN(n7105) );
  AND2_X1 U8283 ( .A1(n7106), .A2(n7105), .ZN(n10457) );
  NAND2_X1 U8284 ( .A1(n6676), .A2(n10399), .ZN(n10403) );
  OR2_X1 U8285 ( .A1(n9544), .A2(n10413), .ZN(n7107) );
  NAND2_X1 U8286 ( .A1(n7108), .A2(n7107), .ZN(n7216) );
  NAND2_X1 U8287 ( .A1(n7216), .A2(n7109), .ZN(n7111) );
  OR2_X1 U8288 ( .A1(n6813), .A2(n10426), .ZN(n7110) );
  NAND2_X1 U8289 ( .A1(n7111), .A2(n7110), .ZN(n7188) );
  NAND2_X1 U8290 ( .A1(n7188), .A2(n5213), .ZN(n7113) );
  OR2_X1 U8291 ( .A1(n6954), .A2(n7193), .ZN(n7112) );
  NAND2_X1 U8292 ( .A1(n7113), .A2(n7112), .ZN(n7205) );
  XNOR2_X1 U8293 ( .A(n7205), .B(n7204), .ZN(n10455) );
  AOI21_X1 U8294 ( .B1(n8532), .B2(n7116), .A(n10415), .ZN(n7114) );
  NAND2_X1 U8295 ( .A1(n7115), .A2(n7114), .ZN(n9836) );
  NOR2_X1 U8296 ( .A1(n7116), .A2(n9781), .ZN(n7191) );
  INV_X1 U8297 ( .A(n7191), .ZN(n7117) );
  NAND2_X1 U8298 ( .A1(n9836), .A2(n7117), .ZN(n10418) );
  INV_X1 U8299 ( .A(n9804), .ZN(n7867) );
  INV_X1 U8300 ( .A(n9825), .ZN(n9728) );
  OR2_X1 U8301 ( .A1(n10413), .A2(n10399), .ZN(n10400) );
  NAND2_X1 U8302 ( .A1(n7223), .A2(n10443), .ZN(n7118) );
  NAND2_X1 U8303 ( .A1(n7118), .A2(n7206), .ZN(n7119) );
  NAND2_X1 U8304 ( .A1(n7199), .A2(n7119), .ZN(n10453) );
  OAI22_X1 U8305 ( .A1(n9822), .A2(n6420), .B1(n7120), .B2(n9819), .ZN(n7121)
         );
  AOI21_X1 U8306 ( .B1(n9785), .B2(n7206), .A(n7121), .ZN(n7122) );
  OAI21_X1 U8307 ( .B1(n9728), .B2(n10453), .A(n7122), .ZN(n7123) );
  AOI21_X1 U8308 ( .B1(n10455), .B2(n7867), .A(n7123), .ZN(n7124) );
  OAI21_X1 U8309 ( .B1(n10457), .B2(n9684), .A(n7124), .ZN(P1_U3287) );
  INV_X1 U8310 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7127) );
  XNOR2_X1 U8311 ( .A(n7125), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9570) );
  INV_X1 U8312 ( .A(n9570), .ZN(n9560) );
  OAI222_X1 U8313 ( .A1(n9961), .A2(n7127), .B1(n8830), .B2(n7126), .C1(n9560), 
        .C2(P1_U3084), .ZN(P1_U3337) );
  NAND2_X1 U8314 ( .A1(n7128), .A2(n8355), .ZN(n7131) );
  AOI22_X1 U8315 ( .A1(n8029), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8028), .B2(
        n7129), .ZN(n7130) );
  NAND2_X1 U8316 ( .A1(n7367), .A2(n8191), .ZN(n7132) );
  OAI21_X1 U8317 ( .B1(n7392), .B2(n6906), .A(n7132), .ZN(n7133) );
  XNOR2_X1 U8318 ( .A(n7133), .B(n8188), .ZN(n7353) );
  OR2_X1 U8319 ( .A1(n7392), .A2(n8199), .ZN(n7135) );
  NAND2_X1 U8320 ( .A1(n7367), .A2(n8155), .ZN(n7134) );
  NAND2_X1 U8321 ( .A1(n7135), .A2(n7134), .ZN(n7351) );
  XNOR2_X1 U8322 ( .A(n7353), .B(n7351), .ZN(n7143) );
  NAND2_X1 U8323 ( .A1(n7136), .A2(n7139), .ZN(n7142) );
  INV_X1 U8324 ( .A(n7143), .ZN(n7140) );
  OAI21_X1 U8325 ( .B1(n7143), .B2(n7142), .A(n7355), .ZN(n7144) );
  NAND2_X1 U8326 ( .A1(n7144), .A2(n9485), .ZN(n7158) );
  INV_X1 U8327 ( .A(n7391), .ZN(n7156) );
  NAND2_X1 U8328 ( .A1(n4862), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7152) );
  OR2_X1 U8329 ( .A1(n7853), .A2(n6508), .ZN(n7151) );
  NAND2_X1 U8330 ( .A1(n7146), .A2(n7145), .ZN(n7147) );
  NAND2_X1 U8331 ( .A1(n7273), .A2(n7147), .ZN(n7369) );
  OR2_X1 U8332 ( .A1(n8145), .A2(n7369), .ZN(n7150) );
  INV_X1 U8333 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7148) );
  OR2_X1 U8334 ( .A1(n6787), .A2(n7148), .ZN(n7149) );
  AOI21_X1 U8335 ( .B1(n9488), .B2(n7290), .A(n7153), .ZN(n7154) );
  OAI21_X1 U8336 ( .B1(n7445), .B2(n9507), .A(n7154), .ZN(n7155) );
  AOI21_X1 U8337 ( .B1(n7156), .B2(n9510), .A(n7155), .ZN(n7157) );
  OAI211_X1 U8338 ( .C1(n7392), .C2(n9513), .A(n7158), .B(n7157), .ZN(P1_U3211) );
  OAI21_X1 U8339 ( .B1(n7161), .B2(n7160), .A(n7159), .ZN(n7162) );
  NAND2_X1 U8340 ( .A1(n7162), .A2(n8994), .ZN(n7169) );
  NAND2_X1 U8341 ( .A1(P2_U3152), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7630) );
  INV_X1 U8342 ( .A(n7630), .ZN(n7167) );
  AOI211_X1 U8343 ( .C1(n7165), .C2(n7164), .A(n7163), .B(n4946), .ZN(n7166)
         );
  AOI211_X1 U8344 ( .C1(n10319), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n7167), .B(
        n7166), .ZN(n7168) );
  OAI211_X1 U8345 ( .C1(n8991), .C2(n7170), .A(n7169), .B(n7168), .ZN(P2_U3256) );
  OAI21_X1 U8346 ( .B1(n10509), .B2(n7172), .A(n8873), .ZN(n7175) );
  INV_X1 U8347 ( .A(n7256), .ZN(n9250) );
  NAND3_X1 U8348 ( .A1(n7173), .A2(n8875), .A3(n9250), .ZN(n7174) );
  AND2_X1 U8349 ( .A1(n7175), .A2(n7174), .ZN(n7181) );
  NOR2_X1 U8350 ( .A1(n10523), .A2(n7265), .ZN(n7179) );
  NAND2_X1 U8351 ( .A1(n8906), .A2(n9250), .ZN(n7177) );
  OAI211_X1 U8352 ( .C1(n7331), .C2(n10517), .A(n7177), .B(n7176), .ZN(n7178)
         );
  AOI211_X1 U8353 ( .C1(n8918), .C2(n8624), .A(n7179), .B(n7178), .ZN(n7180)
         );
  OAI21_X1 U8354 ( .B1(n5069), .B2(n7181), .A(n7180), .ZN(P2_U3223) );
  NAND3_X1 U8355 ( .A1(n7217), .A2(n5213), .A3(n8415), .ZN(n7182) );
  NAND2_X1 U8356 ( .A1(n7183), .A2(n7182), .ZN(n7187) );
  NAND2_X1 U8357 ( .A1(n6813), .A2(n10393), .ZN(n7185) );
  NAND2_X1 U8358 ( .A1(n6883), .A2(n10392), .ZN(n7184) );
  NAND2_X1 U8359 ( .A1(n7185), .A2(n7184), .ZN(n7186) );
  AOI21_X1 U8360 ( .B1(n7187), .B2(n10397), .A(n7186), .ZN(n7190) );
  XNOR2_X1 U8361 ( .A(n7188), .B(n5213), .ZN(n10446) );
  NAND2_X1 U8362 ( .A1(n10446), .A2(n9816), .ZN(n7189) );
  AND2_X1 U8363 ( .A1(n7190), .A2(n7189), .ZN(n10448) );
  NAND2_X1 U8364 ( .A1(n9822), .A2(n7191), .ZN(n9635) );
  XNOR2_X1 U8365 ( .A(n7223), .B(n10443), .ZN(n10444) );
  OAI22_X1 U8366 ( .A1(n9822), .A2(n6789), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9819), .ZN(n7192) );
  AOI21_X1 U8367 ( .B1(n9785), .B2(n7193), .A(n7192), .ZN(n7194) );
  OAI21_X1 U8368 ( .B1(n9728), .B2(n10444), .A(n7194), .ZN(n7195) );
  AOI21_X1 U8369 ( .B1(n10446), .B2(n9826), .A(n7195), .ZN(n7196) );
  OAI21_X1 U8370 ( .B1(n10448), .B2(n9684), .A(n7196), .ZN(P1_U3288) );
  INV_X1 U8371 ( .A(n7326), .ZN(n7198) );
  AOI211_X1 U8372 ( .C1(n7287), .C2(n7199), .A(n10548), .B(n7198), .ZN(n10466)
         );
  INV_X1 U8373 ( .A(n6883), .ZN(n7203) );
  OR2_X1 U8374 ( .A1(n7322), .A2(n10468), .ZN(n8268) );
  NAND2_X1 U8375 ( .A1(n7322), .A2(n10468), .ZN(n7319) );
  XNOR2_X1 U8376 ( .A(n8266), .B(n8494), .ZN(n7202) );
  OAI222_X1 U8377 ( .A1(n9808), .A2(n7376), .B1(n9779), .B2(n7203), .C1(n9811), 
        .C2(n7202), .ZN(n10469) );
  AOI21_X1 U8378 ( .B1(n10466), .B2(n9781), .A(n10469), .ZN(n7215) );
  NAND2_X1 U8379 ( .A1(n7205), .A2(n7204), .ZN(n7208) );
  OR2_X1 U8380 ( .A1(n6883), .A2(n7206), .ZN(n7207) );
  NAND2_X1 U8381 ( .A1(n7208), .A2(n7207), .ZN(n7210) );
  INV_X1 U8382 ( .A(n7289), .ZN(n7209) );
  AOI21_X1 U8383 ( .B1(n8494), .B2(n7210), .A(n7209), .ZN(n10471) );
  NOR2_X1 U8384 ( .A1(n9818), .A2(n10468), .ZN(n7213) );
  OAI22_X1 U8385 ( .A1(n9822), .A2(n6459), .B1(n7211), .B2(n9819), .ZN(n7212)
         );
  AOI211_X1 U8386 ( .C1(n10471), .C2(n7867), .A(n7213), .B(n7212), .ZN(n7214)
         );
  OAI21_X1 U8387 ( .B1(n7215), .B2(n9684), .A(n7214), .ZN(P1_U3286) );
  XNOR2_X1 U8388 ( .A(n7216), .B(n8490), .ZN(n10430) );
  OAI21_X1 U8389 ( .B1(n8490), .B2(n8419), .A(n7217), .ZN(n7222) );
  INV_X1 U8390 ( .A(n9544), .ZN(n7219) );
  INV_X1 U8391 ( .A(n6954), .ZN(n7218) );
  OAI22_X1 U8392 ( .A1(n7219), .A2(n9779), .B1(n7218), .B2(n9808), .ZN(n7221)
         );
  NOR2_X1 U8393 ( .A1(n10430), .A2(n9836), .ZN(n7220) );
  AOI211_X1 U8394 ( .C1(n10397), .C2(n7222), .A(n7221), .B(n7220), .ZN(n10429)
         );
  MUX2_X1 U8395 ( .A(n6454), .B(n10429), .S(n9822), .Z(n7228) );
  AOI21_X1 U8396 ( .B1(n10426), .B2(n10400), .A(n7223), .ZN(n10427) );
  OAI22_X1 U8397 ( .A1(n9818), .A2(n7225), .B1(n9819), .B2(n7224), .ZN(n7226)
         );
  AOI21_X1 U8398 ( .B1(n9825), .B2(n10427), .A(n7226), .ZN(n7227) );
  OAI211_X1 U8399 ( .C1(n10430), .C2(n9635), .A(n7228), .B(n7227), .ZN(
        P1_U3289) );
  AOI22_X1 U8400 ( .A1(n8986), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n9373), .ZN(n7229) );
  OAI21_X1 U8401 ( .B1(n8027), .B2(n9380), .A(n7229), .ZN(P2_U3340) );
  NAND2_X1 U8402 ( .A1(n7230), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7231) );
  XNOR2_X1 U8403 ( .A(n7231), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9598) );
  AOI22_X1 U8404 ( .A1(n9598), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9958), .ZN(n7232) );
  OAI21_X1 U8405 ( .B1(n8027), .B2(n8830), .A(n7232), .ZN(P1_U3335) );
  OR2_X1 U8406 ( .A1(n10492), .A2(n8929), .ZN(n8616) );
  NAND2_X1 U8407 ( .A1(n10492), .A2(n8929), .ZN(n8614) );
  NAND2_X1 U8408 ( .A1(n8616), .A2(n8614), .ZN(n9261) );
  OR2_X1 U8409 ( .A1(n10525), .A2(n7256), .ZN(n8618) );
  NAND2_X1 U8410 ( .A1(n10525), .A2(n7256), .ZN(n7250) );
  NAND2_X1 U8411 ( .A1(n8618), .A2(n7250), .ZN(n8747) );
  OAI21_X1 U8412 ( .B1(n7235), .B2(n8747), .A(n7258), .ZN(n7236) );
  INV_X1 U8413 ( .A(n7236), .ZN(n10529) );
  INV_X1 U8414 ( .A(n8747), .ZN(n7242) );
  INV_X1 U8415 ( .A(n8607), .ZN(n7237) );
  INV_X1 U8416 ( .A(n8929), .ZN(n10513) );
  AND2_X1 U8417 ( .A1(n10492), .A2(n10513), .ZN(n7239) );
  OR2_X1 U8418 ( .A1(n10492), .A2(n10513), .ZN(n7240) );
  OAI21_X1 U8419 ( .B1(n7242), .B2(n7241), .A(n7252), .ZN(n7243) );
  AOI222_X1 U8420 ( .A1(n9234), .A2(n7243), .B1(n8928), .B2(n10587), .C1(n8929), .C2(n9230), .ZN(n10528) );
  MUX2_X1 U8421 ( .A(n7244), .B(n10528), .S(n10605), .Z(n7248) );
  INV_X1 U8422 ( .A(n10492), .ZN(n9258) );
  NAND2_X1 U8423 ( .A1(n9253), .A2(n9258), .ZN(n9254) );
  INV_X1 U8424 ( .A(n7262), .ZN(n7264) );
  AOI21_X1 U8425 ( .B1(n10525), .B2(n9254), .A(n7264), .ZN(n10526) );
  INV_X1 U8426 ( .A(n10525), .ZN(n7245) );
  OAI22_X1 U8427 ( .A1(n10383), .A2(n7245), .B1(n10609), .B2(n10524), .ZN(
        n7246) );
  AOI21_X1 U8428 ( .B1(n10526), .B2(n9260), .A(n7246), .ZN(n7247) );
  OAI211_X1 U8429 ( .C1(n10529), .C2(n9244), .A(n7248), .B(n7247), .ZN(
        P2_U3289) );
  NAND2_X1 U8430 ( .A1(n8624), .A2(n8928), .ZN(n7339) );
  OR2_X1 U8431 ( .A1(n8624), .A2(n8928), .ZN(n7249) );
  NAND2_X1 U8432 ( .A1(n7339), .A2(n7249), .ZN(n8738) );
  NOR2_X1 U8433 ( .A1(n8738), .A2(n5266), .ZN(n7253) );
  NAND2_X1 U8434 ( .A1(n7251), .A2(n8738), .ZN(n7334) );
  INV_X1 U8435 ( .A(n7334), .ZN(n7332) );
  AOI21_X1 U8436 ( .B1(n7253), .B2(n7252), .A(n7332), .ZN(n7254) );
  OAI222_X1 U8437 ( .A1(n9214), .A2(n7331), .B1(n9216), .B2(n7256), .C1(n7255), 
        .C2(n7254), .ZN(n10543) );
  INV_X1 U8438 ( .A(n10543), .ZN(n7271) );
  OR2_X1 U8439 ( .A1(n10525), .A2(n9250), .ZN(n7257) );
  INV_X1 U8440 ( .A(n7341), .ZN(n7338) );
  AOI21_X1 U8441 ( .B1(n8738), .B2(n7261), .A(n7338), .ZN(n10545) );
  INV_X1 U8442 ( .A(n7343), .ZN(n7263) );
  OAI211_X1 U8443 ( .C1(n5286), .C2(n7264), .A(n7263), .B(n10629), .ZN(n10542)
         );
  INV_X1 U8444 ( .A(n9186), .ZN(n9225) );
  OAI22_X1 U8445 ( .A1(n10605), .A2(n7266), .B1(n7265), .B2(n10609), .ZN(n7267) );
  AOI21_X1 U8446 ( .B1(n9223), .B2(n8624), .A(n7267), .ZN(n7268) );
  OAI21_X1 U8447 ( .B1(n10542), .B2(n9225), .A(n7268), .ZN(n7269) );
  AOI21_X1 U8448 ( .B1(n10545), .B2(n9263), .A(n7269), .ZN(n7270) );
  OAI21_X1 U8449 ( .B1(n7271), .B2(n10607), .A(n7270), .ZN(P2_U3288) );
  NAND2_X1 U8450 ( .A1(n4862), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7279) );
  OR2_X1 U8451 ( .A1(n7853), .A2(n6547), .ZN(n7278) );
  NAND2_X1 U8452 ( .A1(n7273), .A2(n7272), .ZN(n7274) );
  NAND2_X1 U8453 ( .A1(n7408), .A2(n7274), .ZN(n7456) );
  OR2_X1 U8454 ( .A1(n8145), .A2(n7456), .ZN(n7277) );
  OR2_X1 U8455 ( .A1(n6787), .A2(n7275), .ZN(n7276) );
  OR2_X1 U8456 ( .A1(n7290), .A2(n10485), .ZN(n8277) );
  AND2_X1 U8457 ( .A1(n8277), .A2(n8268), .ZN(n8464) );
  NAND2_X1 U8458 ( .A1(n7392), .A2(n7367), .ZN(n8428) );
  NAND2_X1 U8459 ( .A1(n7290), .A2(n10485), .ZN(n8275) );
  NAND2_X1 U8460 ( .A1(n7319), .A2(n8275), .ZN(n7280) );
  NAND2_X1 U8461 ( .A1(n7280), .A2(n8277), .ZN(n8427) );
  AND2_X1 U8462 ( .A1(n8499), .A2(n8427), .ZN(n7281) );
  NAND2_X1 U8463 ( .A1(n7450), .A2(n8402), .ZN(n7285) );
  AOI22_X1 U8464 ( .A1(n8029), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8028), .B2(
        n7283), .ZN(n7284) );
  OR2_X1 U8465 ( .A1(n10534), .A2(n7445), .ZN(n8387) );
  NAND2_X1 U8466 ( .A1(n10534), .A2(n7445), .ZN(n8403) );
  NAND2_X1 U8467 ( .A1(n8387), .A2(n8403), .ZN(n8284) );
  XNOR2_X1 U8468 ( .A(n7285), .B(n8284), .ZN(n7286) );
  OAI222_X1 U8469 ( .A1(n9808), .A2(n7734), .B1(n9779), .B2(n5130), .C1(n7286), 
        .C2(n9811), .ZN(n10537) );
  INV_X1 U8470 ( .A(n10537), .ZN(n7305) );
  NAND2_X1 U8471 ( .A1(n7322), .A2(n7287), .ZN(n7288) );
  INV_X1 U8472 ( .A(n10485), .ZN(n7299) );
  OR2_X1 U8473 ( .A1(n7290), .A2(n7299), .ZN(n7373) );
  OR2_X1 U8474 ( .A1(n7367), .A2(n5131), .ZN(n7291) );
  AND2_X1 U8475 ( .A1(n7373), .A2(n7291), .ZN(n7294) );
  NAND2_X1 U8476 ( .A1(n7374), .A2(n7294), .ZN(n7293) );
  INV_X1 U8477 ( .A(n7291), .ZN(n7292) );
  AND2_X1 U8478 ( .A1(n7293), .A2(n7296), .ZN(n7298) );
  AND2_X1 U8479 ( .A1(n7294), .A2(n8284), .ZN(n7295) );
  NAND2_X1 U8480 ( .A1(n7448), .A2(n7446), .ZN(n7297) );
  AOI21_X1 U8481 ( .B1(n8500), .B2(n7298), .A(n7297), .ZN(n10539) );
  NAND2_X1 U8482 ( .A1(n7386), .A2(n7392), .ZN(n7387) );
  OR2_X2 U8483 ( .A1(n7387), .A2(n10534), .ZN(n7457) );
  NAND2_X1 U8484 ( .A1(n7387), .A2(n10534), .ZN(n7300) );
  NAND2_X1 U8485 ( .A1(n7457), .A2(n7300), .ZN(n10536) );
  OAI22_X1 U8486 ( .A1(n9822), .A2(n6508), .B1(n7369), .B2(n9819), .ZN(n7301)
         );
  AOI21_X1 U8487 ( .B1(n9785), .B2(n10534), .A(n7301), .ZN(n7302) );
  OAI21_X1 U8488 ( .B1(n10536), .B2(n9728), .A(n7302), .ZN(n7303) );
  AOI21_X1 U8489 ( .B1(n10539), .B2(n7867), .A(n7303), .ZN(n7304) );
  OAI21_X1 U8490 ( .B1(n10425), .B2(n7305), .A(n7304), .ZN(P1_U3283) );
  NOR2_X1 U8491 ( .A1(n10253), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7306) );
  AOI21_X1 U8492 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n10253), .A(n7306), .ZN(
        n10256) );
  AOI21_X1 U8493 ( .B1(n7768), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7307), .ZN(
        n10255) );
  NAND2_X1 U8494 ( .A1(n10256), .A2(n10255), .ZN(n10254) );
  OAI21_X1 U8495 ( .B1(n10253), .B2(P1_REG2_REG_14__SCAN_IN), .A(n10254), .ZN(
        n9546) );
  XNOR2_X1 U8496 ( .A(n9546), .B(n9553), .ZN(n7309) );
  INV_X1 U8497 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7308) );
  NOR2_X1 U8498 ( .A1(n7308), .A2(n7309), .ZN(n9547) );
  AOI211_X1 U8499 ( .C1(n7309), .C2(n7308), .A(n9547), .B(n10370), .ZN(n7316)
         );
  INV_X1 U8500 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10643) );
  AOI22_X1 U8501 ( .A1(n10253), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n10643), 
        .B2(n7310), .ZN(n10259) );
  OAI21_X1 U8502 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n7768), .A(n7311), .ZN(
        n10258) );
  NAND2_X1 U8503 ( .A1(n10259), .A2(n10258), .ZN(n10257) );
  OAI21_X1 U8504 ( .B1(n10253), .B2(P1_REG1_REG_14__SCAN_IN), .A(n10257), .ZN(
        n9552) );
  XNOR2_X1 U8505 ( .A(n9552), .B(n9553), .ZN(n7312) );
  INV_X1 U8506 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7857) );
  NOR2_X1 U8507 ( .A1(n7857), .A2(n7312), .ZN(n9554) );
  AOI211_X1 U8508 ( .C1(n7312), .C2(n7857), .A(n9554), .B(n10333), .ZN(n7315)
         );
  NAND2_X1 U8509 ( .A1(n10290), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n7313) );
  NAND2_X1 U8510 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9519) );
  OAI211_X1 U8511 ( .C1(n9553), .C2(n10364), .A(n7313), .B(n9519), .ZN(n7314)
         );
  OR3_X1 U8512 ( .A1(n7316), .A2(n7315), .A3(n7314), .ZN(P1_U3256) );
  INV_X1 U8513 ( .A(n7374), .ZN(n7317) );
  AOI21_X1 U8514 ( .B1(n8498), .B2(n7318), .A(n7317), .ZN(n10481) );
  INV_X1 U8515 ( .A(n7319), .ZN(n8269) );
  OR2_X1 U8516 ( .A1(n8266), .A2(n8269), .ZN(n8465) );
  NAND2_X1 U8517 ( .A1(n8465), .A2(n8268), .ZN(n7320) );
  XNOR2_X1 U8518 ( .A(n7320), .B(n8498), .ZN(n7321) );
  NAND2_X1 U8519 ( .A1(n7321), .A2(n10397), .ZN(n7324) );
  AOI22_X1 U8520 ( .A1(n10393), .A2(n7322), .B1(n7367), .B2(n10392), .ZN(n7323) );
  NAND2_X1 U8521 ( .A1(n7324), .A2(n7323), .ZN(n10486) );
  MUX2_X1 U8522 ( .A(n10486), .B(P1_REG2_REG_6__SCAN_IN), .S(n10425), .Z(n7325) );
  INV_X1 U8523 ( .A(n7325), .ZN(n7330) );
  XNOR2_X1 U8524 ( .A(n7326), .B(n10485), .ZN(n10483) );
  OAI22_X1 U8525 ( .A1(n9818), .A2(n10485), .B1(n9819), .B2(n7327), .ZN(n7328)
         );
  AOI21_X1 U8526 ( .B1(n10483), .B2(n9825), .A(n7328), .ZN(n7329) );
  OAI211_X1 U8527 ( .C1(n10481), .C2(n9804), .A(n7330), .B(n7329), .ZN(
        P1_U3285) );
  INV_X1 U8528 ( .A(n8928), .ZN(n10516) );
  AND2_X1 U8529 ( .A1(n8624), .A2(n10516), .ZN(n8621) );
  OR2_X1 U8530 ( .A1(n7493), .A2(n7331), .ZN(n8632) );
  NAND2_X1 U8531 ( .A1(n7493), .A2(n7331), .ZN(n8631) );
  NAND2_X1 U8532 ( .A1(n8632), .A2(n8631), .ZN(n8748) );
  OAI21_X1 U8533 ( .B1(n7332), .B2(n8621), .A(n8748), .ZN(n7335) );
  NOR2_X1 U8534 ( .A1(n8748), .A2(n8621), .ZN(n7333) );
  NAND3_X1 U8535 ( .A1(n7335), .A2(n7469), .A3(n9234), .ZN(n7337) );
  AOI22_X1 U8536 ( .A1(n10586), .A2(n10587), .B1(n9230), .B2(n8928), .ZN(n7336) );
  NAND2_X1 U8537 ( .A1(n7337), .A2(n7336), .ZN(n10557) );
  INV_X1 U8538 ( .A(n10557), .ZN(n7350) );
  INV_X1 U8539 ( .A(n7339), .ZN(n8626) );
  NOR2_X1 U8540 ( .A1(n7338), .A2(n8626), .ZN(n7342) );
  AND2_X1 U8541 ( .A1(n8748), .A2(n7339), .ZN(n7340) );
  NAND2_X1 U8542 ( .A1(n7341), .A2(n7340), .ZN(n7466) );
  OAI21_X1 U8543 ( .B1(n7342), .B2(n8748), .A(n7466), .ZN(n10559) );
  INV_X1 U8544 ( .A(n7493), .ZN(n10555) );
  NOR2_X1 U8545 ( .A1(n7343), .A2(n10555), .ZN(n7344) );
  OR2_X1 U8546 ( .A1(n7476), .A2(n7344), .ZN(n10556) );
  INV_X1 U8547 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7345) );
  OAI22_X1 U8548 ( .A1(n10605), .A2(n7345), .B1(n7486), .B2(n10609), .ZN(n7346) );
  AOI21_X1 U8549 ( .B1(n7493), .B2(n9223), .A(n7346), .ZN(n7347) );
  OAI21_X1 U8550 ( .B1(n10556), .B2(n10382), .A(n7347), .ZN(n7348) );
  AOI21_X1 U8551 ( .B1(n10559), .B2(n9263), .A(n7348), .ZN(n7349) );
  OAI21_X1 U8552 ( .B1(n10607), .B2(n7350), .A(n7349), .ZN(P2_U3287) );
  INV_X1 U8553 ( .A(n7351), .ZN(n7352) );
  NAND2_X1 U8554 ( .A1(n7353), .A2(n7352), .ZN(n7354) );
  INV_X1 U8555 ( .A(n7535), .ZN(n7358) );
  NAND2_X1 U8556 ( .A1(n10534), .A2(n8185), .ZN(n7357) );
  OR2_X1 U8557 ( .A1(n7445), .A2(n8196), .ZN(n7356) );
  NAND2_X1 U8558 ( .A1(n7357), .A2(n7356), .ZN(n7530) );
  NAND2_X1 U8559 ( .A1(n7358), .A2(n7530), .ZN(n7362) );
  NAND2_X1 U8560 ( .A1(n10534), .A2(n8184), .ZN(n7360) );
  OR2_X1 U8561 ( .A1(n7445), .A2(n8199), .ZN(n7359) );
  NAND2_X1 U8562 ( .A1(n7360), .A2(n7359), .ZN(n7361) );
  XNOR2_X1 U8563 ( .A(n7361), .B(n8197), .ZN(n7531) );
  INV_X1 U8564 ( .A(n7531), .ZN(n7537) );
  NAND2_X1 U8565 ( .A1(n7362), .A2(n7537), .ZN(n7397) );
  INV_X1 U8566 ( .A(n7397), .ZN(n7364) );
  INV_X1 U8567 ( .A(n7530), .ZN(n7538) );
  NAND2_X1 U8568 ( .A1(n7535), .A2(n7538), .ZN(n7396) );
  AOI21_X1 U8569 ( .B1(n7362), .B2(n7396), .A(n7537), .ZN(n7363) );
  AOI21_X1 U8570 ( .B1(n7364), .B2(n7396), .A(n7363), .ZN(n7372) );
  NOR2_X1 U8571 ( .A1(n9507), .A2(n7734), .ZN(n7365) );
  AOI211_X1 U8572 ( .C1(n9488), .C2(n7367), .A(n7366), .B(n7365), .ZN(n7368)
         );
  OAI21_X1 U8573 ( .B1(n9526), .B2(n7369), .A(n7368), .ZN(n7370) );
  AOI21_X1 U8574 ( .B1(n10534), .B2(n9528), .A(n7370), .ZN(n7371) );
  OAI21_X1 U8575 ( .B1(n7372), .B2(n9530), .A(n7371), .ZN(P1_U3219) );
  NAND2_X1 U8576 ( .A1(n7374), .A2(n7373), .ZN(n7375) );
  XNOR2_X1 U8577 ( .A(n7375), .B(n7378), .ZN(n7384) );
  INV_X1 U8578 ( .A(n7384), .ZN(n10505) );
  OAI22_X1 U8579 ( .A1(n7376), .A2(n9779), .B1(n7445), .B2(n9808), .ZN(n7383)
         );
  INV_X1 U8580 ( .A(n7377), .ZN(n7380) );
  INV_X1 U8581 ( .A(n8427), .ZN(n7379) );
  OAI21_X1 U8582 ( .B1(n7380), .B2(n7379), .A(n7378), .ZN(n7381) );
  AOI21_X1 U8583 ( .B1(n7381), .B2(n7450), .A(n9811), .ZN(n7382) );
  AOI211_X1 U8584 ( .C1(n9816), .C2(n7384), .A(n7383), .B(n7382), .ZN(n10503)
         );
  MUX2_X1 U8585 ( .A(n7385), .B(n10503), .S(n9822), .Z(n7395) );
  INV_X1 U8586 ( .A(n7386), .ZN(n7389) );
  INV_X1 U8587 ( .A(n7387), .ZN(n7388) );
  AOI211_X1 U8588 ( .C1(n5131), .C2(n7389), .A(n10548), .B(n7388), .ZN(n10500)
         );
  NOR2_X1 U8589 ( .A1(n7390), .A2(n10415), .ZN(n7935) );
  OAI22_X1 U8590 ( .A1(n9818), .A2(n7392), .B1(n9819), .B2(n7391), .ZN(n7393)
         );
  AOI21_X1 U8591 ( .B1(n10500), .B2(n7935), .A(n7393), .ZN(n7394) );
  OAI211_X1 U8592 ( .C1(n10505), .C2(n9635), .A(n7395), .B(n7394), .ZN(
        P1_U3284) );
  NAND2_X1 U8593 ( .A1(n7397), .A2(n7396), .ZN(n7406) );
  NAND2_X1 U8594 ( .A1(n7398), .A2(n8355), .ZN(n7401) );
  AOI22_X1 U8595 ( .A1(n8029), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8028), .B2(
        n7399), .ZN(n7400) );
  NAND2_X1 U8596 ( .A1(n10547), .A2(n8184), .ZN(n7403) );
  OR2_X1 U8597 ( .A1(n7734), .A2(n8199), .ZN(n7402) );
  NAND2_X1 U8598 ( .A1(n7403), .A2(n7402), .ZN(n7404) );
  XNOR2_X1 U8599 ( .A(n7404), .B(n8188), .ZN(n7536) );
  AOI22_X1 U8600 ( .A1(n10547), .A2(n8185), .B1(n8155), .B2(n9542), .ZN(n7539)
         );
  XNOR2_X1 U8601 ( .A(n7536), .B(n7539), .ZN(n7405) );
  XNOR2_X1 U8602 ( .A(n7406), .B(n7405), .ZN(n7419) );
  NAND2_X1 U8603 ( .A1(n4862), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7413) );
  OR2_X1 U8604 ( .A1(n7853), .A2(n7521), .ZN(n7412) );
  NAND2_X1 U8605 ( .A1(n7408), .A2(n7407), .ZN(n7409) );
  NAND2_X1 U8606 ( .A1(n7509), .A2(n7409), .ZN(n7737) );
  OR2_X1 U8607 ( .A1(n8145), .A2(n7737), .ZN(n7411) );
  OR2_X1 U8608 ( .A1(n6787), .A2(n10567), .ZN(n7410) );
  INV_X1 U8609 ( .A(n7617), .ZN(n9541) );
  NOR2_X1 U8610 ( .A1(n9521), .A2(n7445), .ZN(n7414) );
  AOI211_X1 U8611 ( .C1(n9523), .C2(n9541), .A(n7415), .B(n7414), .ZN(n7416)
         );
  OAI21_X1 U8612 ( .B1(n9526), .B2(n7456), .A(n7416), .ZN(n7417) );
  AOI21_X1 U8613 ( .B1(n10547), .B2(n9528), .A(n7417), .ZN(n7418) );
  OAI21_X1 U8614 ( .B1(n7419), .B2(n9530), .A(n7418), .ZN(P1_U3229) );
  INV_X1 U8615 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7420) );
  INV_X1 U8616 ( .A(n7995), .ZN(n7981) );
  OAI222_X1 U8617 ( .A1(n9961), .A2(n7420), .B1(n8830), .B2(n7981), .C1(
        P1_U3084), .C2(n9781), .ZN(P1_U3334) );
  INV_X1 U8618 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7682) );
  OAI21_X1 U8619 ( .B1(n7423), .B2(n7422), .A(n7421), .ZN(n7424) );
  NAND2_X1 U8620 ( .A1(n4948), .A2(n7424), .ZN(n7425) );
  NAND2_X1 U8621 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7785) );
  OAI211_X1 U8622 ( .C1(n7682), .C2(n8968), .A(n7425), .B(n7785), .ZN(n7430)
         );
  AOI211_X1 U8623 ( .C1(n7428), .C2(n7427), .A(n7426), .B(n10320), .ZN(n7429)
         );
  AOI211_X1 U8624 ( .C1(n10330), .C2(n7431), .A(n7430), .B(n7429), .ZN(n7432)
         );
  INV_X1 U8625 ( .A(n7432), .ZN(P2_U3257) );
  OAI21_X1 U8626 ( .B1(n7435), .B2(n7434), .A(n7433), .ZN(n7437) );
  INV_X1 U8627 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7685) );
  NAND2_X1 U8628 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3152), .ZN(n8223) );
  OAI21_X1 U8629 ( .B1(n8968), .B2(n7685), .A(n8223), .ZN(n7436) );
  AOI21_X1 U8630 ( .B1(n4948), .B2(n7437), .A(n7436), .ZN(n7443) );
  OAI21_X1 U8631 ( .B1(n7440), .B2(n7439), .A(n7438), .ZN(n7441) );
  NAND2_X1 U8632 ( .A1(n8994), .A2(n7441), .ZN(n7442) );
  OAI211_X1 U8633 ( .C1(n8991), .C2(n7444), .A(n7443), .B(n7442), .ZN(P2_U3258) );
  INV_X1 U8634 ( .A(n7445), .ZN(n9543) );
  NAND2_X1 U8635 ( .A1(n10534), .A2(n9543), .ZN(n7447) );
  OR2_X1 U8636 ( .A1(n10547), .A2(n7734), .ZN(n8386) );
  NAND2_X1 U8637 ( .A1(n10547), .A2(n7734), .ZN(n8381) );
  NAND2_X1 U8638 ( .A1(n8386), .A2(n8381), .ZN(n8502) );
  INV_X1 U8639 ( .A(n8502), .ZN(n8286) );
  XNOR2_X1 U8640 ( .A(n7496), .B(n8286), .ZN(n10552) );
  INV_X1 U8641 ( .A(n10552), .ZN(n7464) );
  INV_X1 U8642 ( .A(n8402), .ZN(n8276) );
  INV_X1 U8643 ( .A(n7505), .ZN(n7451) );
  AOI21_X1 U8644 ( .B1(n7452), .B2(n8502), .A(n7451), .ZN(n7455) );
  NAND2_X1 U8645 ( .A1(n10552), .A2(n9816), .ZN(n7454) );
  AOI22_X1 U8646 ( .A1(n10393), .A2(n9543), .B1(n9541), .B2(n10392), .ZN(n7453) );
  OAI211_X1 U8647 ( .C1(n9811), .C2(n7455), .A(n7454), .B(n7453), .ZN(n10550)
         );
  NAND2_X1 U8648 ( .A1(n10550), .A2(n9822), .ZN(n7463) );
  OAI22_X1 U8649 ( .A1(n9822), .A2(n6547), .B1(n7456), .B2(n9819), .ZN(n7461)
         );
  INV_X1 U8650 ( .A(n7519), .ZN(n7459) );
  NAND2_X1 U8651 ( .A1(n7457), .A2(n10547), .ZN(n7458) );
  NAND2_X1 U8652 ( .A1(n7459), .A2(n7458), .ZN(n10549) );
  NOR2_X1 U8653 ( .A1(n10549), .A2(n9728), .ZN(n7460) );
  AOI211_X1 U8654 ( .C1(n9785), .C2(n10547), .A(n7461), .B(n7460), .ZN(n7462)
         );
  OAI211_X1 U8655 ( .C1(n7464), .C2(n9635), .A(n7463), .B(n7462), .ZN(P1_U3282) );
  OR2_X1 U8656 ( .A1(n7493), .A2(n7603), .ZN(n7465) );
  OR2_X1 U8657 ( .A1(n7610), .A2(n7577), .ZN(n8633) );
  NAND2_X1 U8658 ( .A1(n7610), .A2(n7577), .ZN(n10582) );
  XNOR2_X1 U8659 ( .A(n7578), .B(n8751), .ZN(n10570) );
  INV_X1 U8660 ( .A(n7789), .ZN(n8927) );
  AOI22_X1 U8661 ( .A1(n9230), .A2(n7603), .B1(n8927), .B2(n10587), .ZN(n7473)
         );
  INV_X1 U8662 ( .A(n8751), .ZN(n7467) );
  INV_X1 U8663 ( .A(n8632), .ZN(n8629) );
  NOR2_X1 U8664 ( .A1(n7467), .A2(n8629), .ZN(n7468) );
  INV_X1 U8665 ( .A(n10583), .ZN(n7471) );
  AOI21_X1 U8666 ( .B1(n7469), .B2(n8632), .A(n8751), .ZN(n7470) );
  OAI21_X1 U8667 ( .B1(n7471), .B2(n7470), .A(n9234), .ZN(n7472) );
  OAI211_X1 U8668 ( .C1(n10570), .C2(n7474), .A(n7473), .B(n7472), .ZN(n10573)
         );
  NAND2_X1 U8669 ( .A1(n10573), .A2(n10605), .ZN(n7481) );
  OAI22_X1 U8670 ( .A1(n10605), .A2(n7475), .B1(n7605), .B2(n10609), .ZN(n7479) );
  INV_X1 U8671 ( .A(n7610), .ZN(n10571) );
  NAND2_X1 U8672 ( .A1(n7476), .A2(n10571), .ZN(n10590) );
  OR2_X1 U8673 ( .A1(n7476), .A2(n10571), .ZN(n7477) );
  NAND2_X1 U8674 ( .A1(n10590), .A2(n7477), .ZN(n10572) );
  NOR2_X1 U8675 ( .A1(n10572), .A2(n10382), .ZN(n7478) );
  AOI211_X1 U8676 ( .C1(n9223), .C2(n7610), .A(n7479), .B(n7478), .ZN(n7480)
         );
  OAI211_X1 U8677 ( .C1(n10570), .C2(n7482), .A(n7481), .B(n7480), .ZN(
        P2_U3286) );
  OAI21_X1 U8678 ( .B1(n10514), .B2(n10516), .A(n7483), .ZN(n7484) );
  AOI21_X1 U8679 ( .B1(n8917), .B2(n10586), .A(n7484), .ZN(n7485) );
  OAI21_X1 U8680 ( .B1(n7486), .B2(n10523), .A(n7485), .ZN(n7492) );
  INV_X1 U8681 ( .A(n8875), .ZN(n7840) );
  NOR3_X1 U8682 ( .A1(n7487), .A2(n10516), .A3(n7840), .ZN(n7488) );
  AOI21_X1 U8683 ( .B1(n5069), .B2(n8873), .A(n7488), .ZN(n7490) );
  NOR2_X1 U8684 ( .A1(n7490), .A2(n7489), .ZN(n7491) );
  AOI211_X1 U8685 ( .C1(n8918), .C2(n7493), .A(n7492), .B(n7491), .ZN(n7494)
         );
  OAI21_X1 U8686 ( .B1(n7495), .B2(n10510), .A(n7494), .ZN(P2_U3233) );
  NAND2_X1 U8687 ( .A1(n7496), .A2(n9542), .ZN(n7497) );
  NAND2_X1 U8688 ( .A1(n7498), .A2(n8355), .ZN(n7500) );
  AOI22_X1 U8689 ( .A1(n8029), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n8028), .B2(
        n10240), .ZN(n7499) );
  NAND2_X1 U8690 ( .A1(n7500), .A2(n7499), .ZN(n7745) );
  OR2_X1 U8691 ( .A1(n7745), .A2(n7617), .ZN(n8388) );
  NAND2_X1 U8692 ( .A1(n7745), .A2(n7617), .ZN(n8382) );
  NAND2_X1 U8693 ( .A1(n7501), .A2(n8505), .ZN(n7502) );
  NAND2_X1 U8694 ( .A1(n7613), .A2(n7502), .ZN(n10564) );
  INV_X1 U8695 ( .A(n8505), .ZN(n7504) );
  NAND3_X1 U8696 ( .A1(n7505), .A2(n7504), .A3(n8381), .ZN(n7506) );
  AOI21_X1 U8697 ( .B1(n7753), .B2(n7506), .A(n9811), .ZN(n7517) );
  NAND2_X1 U8698 ( .A1(n4862), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7515) );
  OR2_X1 U8699 ( .A1(n7853), .A2(n7507), .ZN(n7514) );
  INV_X1 U8700 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7508) );
  NAND2_X1 U8701 ( .A1(n7509), .A2(n7508), .ZN(n7510) );
  NAND2_X1 U8702 ( .A1(n7561), .A2(n7510), .ZN(n7558) );
  OR2_X1 U8703 ( .A1(n8145), .A2(n7558), .ZN(n7513) );
  OR2_X1 U8704 ( .A1(n6787), .A2(n7511), .ZN(n7512) );
  OAI22_X1 U8705 ( .A1(n7734), .A2(n9779), .B1(n7754), .B2(n9808), .ZN(n7516)
         );
  OR2_X1 U8706 ( .A1(n7517), .A2(n7516), .ZN(n7518) );
  AOI21_X1 U8707 ( .B1(n10564), .B2(n9816), .A(n7518), .ZN(n10566) );
  INV_X1 U8708 ( .A(n7745), .ZN(n10562) );
  OAI21_X1 U8709 ( .B1(n7519), .B2(n10562), .A(n10482), .ZN(n7520) );
  OR2_X1 U8710 ( .A1(n7520), .A2(n7620), .ZN(n10561) );
  INV_X1 U8711 ( .A(n7935), .ZN(n7871) );
  OAI22_X1 U8712 ( .A1(n9822), .A2(n7521), .B1(n7737), .B2(n9819), .ZN(n7522)
         );
  AOI21_X1 U8713 ( .B1(n7745), .B2(n9785), .A(n7522), .ZN(n7523) );
  OAI21_X1 U8714 ( .B1(n10561), .B2(n7871), .A(n7523), .ZN(n7524) );
  AOI21_X1 U8715 ( .B1(n10564), .B2(n9826), .A(n7524), .ZN(n7525) );
  OAI21_X1 U8716 ( .B1(n10566), .B2(n10425), .A(n7525), .ZN(P1_U3281) );
  OR2_X1 U8717 ( .A1(n7526), .A2(n6899), .ZN(n7529) );
  AOI22_X1 U8718 ( .A1(n8029), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8028), .B2(
        n7527), .ZN(n7528) );
  INV_X1 U8719 ( .A(n9925), .ZN(n7625) );
  NAND2_X1 U8720 ( .A1(n7531), .A2(n7530), .ZN(n7532) );
  NAND2_X1 U8721 ( .A1(n7535), .A2(n7534), .ZN(n7545) );
  AOI21_X1 U8722 ( .B1(n7537), .B2(n7538), .A(n7539), .ZN(n7542) );
  INV_X1 U8723 ( .A(n7536), .ZN(n7541) );
  NAND3_X1 U8724 ( .A1(n7539), .A2(n7538), .A3(n7537), .ZN(n7540) );
  OAI22_X1 U8725 ( .A1(n10562), .A2(n6906), .B1(n7617), .B2(n8199), .ZN(n7546)
         );
  XOR2_X1 U8726 ( .A(n8197), .B(n7546), .Z(n7548) );
  OAI22_X1 U8727 ( .A1(n10562), .A2(n8199), .B1(n7617), .B2(n8196), .ZN(n7740)
         );
  INV_X1 U8728 ( .A(n7548), .ZN(n7549) );
  NAND2_X1 U8729 ( .A1(n9925), .A2(n8184), .ZN(n7551) );
  OR2_X1 U8730 ( .A1(n7754), .A2(n8199), .ZN(n7550) );
  NAND2_X1 U8731 ( .A1(n7551), .A2(n7550), .ZN(n7552) );
  XNOR2_X1 U8732 ( .A(n7552), .B(n8188), .ZN(n7703) );
  NOR2_X1 U8733 ( .A1(n7754), .A2(n8196), .ZN(n7553) );
  AOI21_X1 U8734 ( .B1(n9925), .B2(n8185), .A(n7553), .ZN(n7702) );
  XNOR2_X1 U8735 ( .A(n7703), .B(n7702), .ZN(n7554) );
  INV_X1 U8736 ( .A(n7705), .ZN(n7557) );
  OAI21_X1 U8737 ( .B1(n7555), .B2(n7739), .A(n7554), .ZN(n7556) );
  NAND3_X1 U8738 ( .A1(n7557), .A2(n9485), .A3(n7556), .ZN(n7571) );
  INV_X1 U8739 ( .A(n7558), .ZN(n7622) );
  NAND2_X1 U8740 ( .A1(n4862), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7566) );
  OR2_X1 U8741 ( .A1(n6787), .A2(n7559), .ZN(n7565) );
  INV_X1 U8742 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7560) );
  NAND2_X1 U8743 ( .A1(n7561), .A2(n7560), .ZN(n7562) );
  NAND2_X1 U8744 ( .A1(n7719), .A2(n7562), .ZN(n7758) );
  OR2_X1 U8745 ( .A1(n8145), .A2(n7758), .ZN(n7564) );
  INV_X1 U8746 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7759) );
  OR2_X1 U8747 ( .A1(n7853), .A2(n7759), .ZN(n7563) );
  AOI21_X1 U8748 ( .B1(n9488), .B2(n9541), .A(n7567), .ZN(n7568) );
  OAI21_X1 U8749 ( .B1(n7808), .B2(n9507), .A(n7568), .ZN(n7569) );
  AOI21_X1 U8750 ( .B1(n7622), .B2(n9510), .A(n7569), .ZN(n7570) );
  OAI211_X1 U8751 ( .C1(n7625), .C2(n9513), .A(n7571), .B(n7570), .ZN(P1_U3234) );
  INV_X1 U8752 ( .A(n8050), .ZN(n7629) );
  INV_X1 U8753 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8051) );
  OAI222_X1 U8754 ( .A1(P1_U3084), .A2(n6648), .B1(n8830), .B2(n7629), .C1(
        n8051), .C2(n9961), .ZN(P1_U3333) );
  OR2_X1 U8755 ( .A1(n10620), .A2(n8224), .ZN(n8637) );
  NAND2_X1 U8756 ( .A1(n10620), .A2(n8224), .ZN(n8640) );
  OR2_X1 U8757 ( .A1(n10598), .A2(n7789), .ZN(n8636) );
  NAND2_X1 U8758 ( .A1(n10598), .A2(n7789), .ZN(n8639) );
  NAND2_X1 U8759 ( .A1(n8636), .A2(n8639), .ZN(n10581) );
  INV_X1 U8760 ( .A(n10581), .ZN(n8750) );
  NAND2_X1 U8761 ( .A1(n7572), .A2(n8752), .ZN(n7641) );
  OAI21_X1 U8762 ( .B1(n8752), .B2(n7572), .A(n7641), .ZN(n7573) );
  NAND2_X1 U8763 ( .A1(n7573), .A2(n9234), .ZN(n7576) );
  OAI22_X1 U8764 ( .A1(n8210), .A2(n9214), .B1(n7789), .B2(n9216), .ZN(n7574)
         );
  INV_X1 U8765 ( .A(n7574), .ZN(n7575) );
  NAND2_X1 U8766 ( .A1(n7576), .A2(n7575), .ZN(n10622) );
  INV_X1 U8767 ( .A(n10622), .ZN(n7587) );
  NAND2_X1 U8768 ( .A1(n10580), .A2(n10581), .ZN(n10579) );
  NAND2_X1 U8769 ( .A1(n10598), .A2(n8927), .ZN(n7579) );
  OAI21_X1 U8770 ( .B1(n5200), .B2(n5199), .A(n7652), .ZN(n10624) );
  NAND2_X1 U8771 ( .A1(n10620), .A2(n10591), .ZN(n7581) );
  NAND2_X1 U8772 ( .A1(n7646), .A2(n7581), .ZN(n10621) );
  INV_X1 U8773 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7582) );
  OAI22_X1 U8774 ( .A1(n10605), .A2(n7582), .B1(n7788), .B2(n10609), .ZN(n7583) );
  AOI21_X1 U8775 ( .B1(n10620), .B2(n9223), .A(n7583), .ZN(n7584) );
  OAI21_X1 U8776 ( .B1(n10621), .B2(n10382), .A(n7584), .ZN(n7585) );
  AOI21_X1 U8777 ( .B1(n10624), .B2(n9263), .A(n7585), .ZN(n7586) );
  OAI21_X1 U8778 ( .B1(n10607), .B2(n7587), .A(n7586), .ZN(P2_U3284) );
  INV_X1 U8779 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7588) );
  OAI222_X1 U8780 ( .A1(n9380), .A2(n8070), .B1(P2_U3152), .B2(n8763), .C1(
        n7588), .C2(n9385), .ZN(P2_U3337) );
  OAI21_X1 U8781 ( .B1(n7592), .B2(n7591), .A(n7590), .ZN(n7594) );
  INV_X1 U8782 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7688) );
  NAND2_X1 U8783 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n8209) );
  OAI21_X1 U8784 ( .B1(n8968), .B2(n7688), .A(n8209), .ZN(n7593) );
  AOI21_X1 U8785 ( .B1(n4948), .B2(n7594), .A(n7593), .ZN(n7600) );
  OAI21_X1 U8786 ( .B1(n7597), .B2(n7596), .A(n7595), .ZN(n7598) );
  NAND2_X1 U8787 ( .A1(n8994), .A2(n7598), .ZN(n7599) );
  OAI211_X1 U8788 ( .C1(n8991), .C2(n5020), .A(n7600), .B(n7599), .ZN(P2_U3259) );
  INV_X1 U8789 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8071) );
  OAI222_X1 U8790 ( .A1(P1_U3084), .A2(n8525), .B1(n8830), .B2(n8070), .C1(
        n8071), .C2(n9961), .ZN(P1_U3332) );
  OAI21_X1 U8791 ( .B1(n10517), .B2(n7789), .A(n7601), .ZN(n7602) );
  AOI21_X1 U8792 ( .B1(n8906), .B2(n7603), .A(n7602), .ZN(n7604) );
  OAI21_X1 U8793 ( .B1(n7605), .B2(n10523), .A(n7604), .ZN(n7609) );
  AOI211_X1 U8794 ( .C1(n7607), .C2(n7606), .A(n10510), .B(n7635), .ZN(n7608)
         );
  AOI211_X1 U8795 ( .C1(n8918), .C2(n7610), .A(n7609), .B(n7608), .ZN(n7611)
         );
  INV_X1 U8796 ( .A(n7611), .ZN(P2_U3219) );
  OR2_X1 U8797 ( .A1(n7745), .A2(n9541), .ZN(n7612) );
  NAND2_X1 U8798 ( .A1(n9925), .A2(n7754), .ZN(n8385) );
  NAND2_X1 U8799 ( .A1(n8389), .A2(n8385), .ZN(n8290) );
  OAI21_X1 U8800 ( .B1(n7614), .B2(n8290), .A(n7748), .ZN(n9924) );
  NAND2_X1 U8801 ( .A1(n7753), .A2(n8382), .ZN(n7615) );
  XNOR2_X1 U8802 ( .A(n7615), .B(n8290), .ZN(n7616) );
  NOR2_X1 U8803 ( .A1(n7616), .A2(n9811), .ZN(n7619) );
  OAI22_X1 U8804 ( .A1(n7617), .A2(n9779), .B1(n7808), .B2(n9808), .ZN(n7618)
         );
  AOI211_X1 U8805 ( .C1(n9924), .C2(n9816), .A(n7619), .B(n7618), .ZN(n9928)
         );
  INV_X1 U8806 ( .A(n7620), .ZN(n7621) );
  AOI21_X1 U8807 ( .B1(n9925), .B2(n7621), .A(n4942), .ZN(n9926) );
  NAND2_X1 U8808 ( .A1(n9926), .A2(n9825), .ZN(n7624) );
  INV_X1 U8809 ( .A(n9819), .ZN(n10411) );
  AOI22_X1 U8810 ( .A1(n10425), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7622), .B2(
        n10411), .ZN(n7623) );
  OAI211_X1 U8811 ( .C1(n7625), .C2(n9818), .A(n7624), .B(n7623), .ZN(n7626)
         );
  AOI21_X1 U8812 ( .B1(n9924), .B2(n9826), .A(n7626), .ZN(n7627) );
  OAI21_X1 U8813 ( .B1(n9928), .B2(n9684), .A(n7627), .ZN(P1_U3280) );
  INV_X1 U8814 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7628) );
  OAI222_X1 U8815 ( .A1(n9380), .A2(n7629), .B1(P2_U3152), .B2(n6098), .C1(
        n7628), .C2(n9385), .ZN(P2_U3338) );
  OAI21_X1 U8816 ( .B1(n10517), .B2(n8224), .A(n7630), .ZN(n7631) );
  AOI21_X1 U8817 ( .B1(n8906), .B2(n10586), .A(n7631), .ZN(n7632) );
  OAI21_X1 U8818 ( .B1(n10610), .B2(n10523), .A(n7632), .ZN(n7639) );
  NAND3_X1 U8819 ( .A1(n7633), .A2(n8875), .A3(n10586), .ZN(n7637) );
  OAI21_X1 U8820 ( .B1(n7635), .B2(n7634), .A(n8873), .ZN(n7636) );
  AOI21_X1 U8821 ( .B1(n7637), .B2(n7636), .A(n5443), .ZN(n7638) );
  AOI211_X1 U8822 ( .C1(n8918), .C2(n10598), .A(n7639), .B(n7638), .ZN(n7640)
         );
  INV_X1 U8823 ( .A(n7640), .ZN(P2_U3238) );
  NAND2_X1 U8824 ( .A1(n7641), .A2(n8640), .ZN(n7642) );
  OR2_X1 U8825 ( .A1(n10627), .A2(n8210), .ZN(n8644) );
  NAND2_X1 U8826 ( .A1(n10627), .A2(n8210), .ZN(n8643) );
  NAND2_X1 U8827 ( .A1(n7642), .A2(n8737), .ZN(n7964) );
  OR2_X1 U8828 ( .A1(n7642), .A2(n8737), .ZN(n7643) );
  NAND2_X1 U8829 ( .A1(n7964), .A2(n7643), .ZN(n7645) );
  OAI22_X1 U8830 ( .A1(n7841), .A2(n9214), .B1(n8224), .B2(n9216), .ZN(n7644)
         );
  AOI21_X1 U8831 ( .B1(n7645), .B2(n9234), .A(n7644), .ZN(n10632) );
  AOI21_X1 U8832 ( .B1(n10627), .B2(n7646), .A(n7975), .ZN(n10630) );
  INV_X1 U8833 ( .A(n10627), .ZN(n7647) );
  NOR2_X1 U8834 ( .A1(n7647), .A2(n10383), .ZN(n7650) );
  INV_X1 U8835 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7648) );
  OAI22_X1 U8836 ( .A1(n10605), .A2(n7648), .B1(n8227), .B2(n10609), .ZN(n7649) );
  AOI211_X1 U8837 ( .C1(n10630), .C2(n9260), .A(n7650), .B(n7649), .ZN(n7655)
         );
  INV_X1 U8838 ( .A(n8224), .ZN(n10588) );
  OR2_X1 U8839 ( .A1(n10620), .A2(n10588), .ZN(n7651) );
  NAND2_X1 U8840 ( .A1(n7653), .A2(n8737), .ZN(n10626) );
  NAND3_X1 U8841 ( .A1(n4932), .A2(n10626), .A3(n9263), .ZN(n7654) );
  OAI211_X1 U8842 ( .C1(n10632), .C2(n10607), .A(n7655), .B(n7654), .ZN(
        P2_U3283) );
  NOR2_X1 U8843 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7697) );
  NOR2_X1 U8844 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7694) );
  NOR2_X1 U8845 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7692) );
  NOR2_X1 U8846 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7690) );
  NOR2_X1 U8847 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7687) );
  NOR2_X1 U8848 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7684) );
  NAND2_X1 U8849 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7681) );
  XOR2_X1 U8850 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n10224) );
  NAND2_X1 U8851 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7679) );
  XNOR2_X1 U8852 ( .A(n7656), .B(P1_ADDR_REG_10__SCAN_IN), .ZN(n10222) );
  NOR2_X1 U8853 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7663) );
  XOR2_X1 U8854 ( .A(n10375), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10213) );
  NAND2_X1 U8855 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7661) );
  XNOR2_X1 U8856 ( .A(n7657), .B(P1_ADDR_REG_3__SCAN_IN), .ZN(n10211) );
  NAND2_X1 U8857 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7659) );
  INV_X1 U8858 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10356) );
  XNOR2_X1 U8859 ( .A(n10356), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(n10209) );
  AOI21_X1 U8860 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10203) );
  INV_X1 U8861 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10207) );
  NAND3_X1 U8862 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10205) );
  OAI21_X1 U8863 ( .B1(n10203), .B2(n10207), .A(n10205), .ZN(n10208) );
  NAND2_X1 U8864 ( .A1(n10209), .A2(n10208), .ZN(n7658) );
  NAND2_X1 U8865 ( .A1(n7659), .A2(n7658), .ZN(n10210) );
  NAND2_X1 U8866 ( .A1(n10211), .A2(n10210), .ZN(n7660) );
  NAND2_X1 U8867 ( .A1(n7661), .A2(n7660), .ZN(n10212) );
  NOR2_X1 U8868 ( .A1(n10213), .A2(n10212), .ZN(n7662) );
  NOR2_X1 U8869 ( .A1(n7663), .A2(n7662), .ZN(n7664) );
  NOR2_X1 U8870 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7664), .ZN(n10214) );
  AND2_X1 U8871 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7664), .ZN(n10215) );
  NOR2_X1 U8872 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10215), .ZN(n7665) );
  NAND2_X1 U8873 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n7666), .ZN(n7668) );
  XOR2_X1 U8874 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n7666), .Z(n10217) );
  NAND2_X1 U8875 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10217), .ZN(n7667) );
  NAND2_X1 U8876 ( .A1(n7668), .A2(n7667), .ZN(n7669) );
  NAND2_X1 U8877 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7669), .ZN(n7671) );
  XOR2_X1 U8878 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7669), .Z(n10218) );
  NAND2_X1 U8879 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10218), .ZN(n7670) );
  NAND2_X1 U8880 ( .A1(n7671), .A2(n7670), .ZN(n7672) );
  NAND2_X1 U8881 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7672), .ZN(n7674) );
  XOR2_X1 U8882 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7672), .Z(n10219) );
  NAND2_X1 U8883 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10219), .ZN(n7673) );
  NAND2_X1 U8884 ( .A1(n7674), .A2(n7673), .ZN(n7675) );
  NAND2_X1 U8885 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n7675), .ZN(n7677) );
  XOR2_X1 U8886 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n7675), .Z(n10220) );
  NAND2_X1 U8887 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10220), .ZN(n7676) );
  NAND2_X1 U8888 ( .A1(n7677), .A2(n7676), .ZN(n10221) );
  NAND2_X1 U8889 ( .A1(n10222), .A2(n10221), .ZN(n7678) );
  NAND2_X1 U8890 ( .A1(n7679), .A2(n7678), .ZN(n10223) );
  NAND2_X1 U8891 ( .A1(n10224), .A2(n10223), .ZN(n7680) );
  NAND2_X1 U8892 ( .A1(n7681), .A2(n7680), .ZN(n10226) );
  XOR2_X1 U8893 ( .A(n7682), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n10225) );
  XOR2_X1 U8894 ( .A(n7685), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n10227) );
  XOR2_X1 U8895 ( .A(n7688), .B(P1_ADDR_REG_14__SCAN_IN), .Z(n10229) );
  NOR2_X1 U8896 ( .A1(n10230), .A2(n10229), .ZN(n7689) );
  NOR2_X1 U8897 ( .A1(n7690), .A2(n7689), .ZN(n10232) );
  INV_X1 U8898 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8936) );
  XOR2_X1 U8899 ( .A(n8936), .B(P1_ADDR_REG_15__SCAN_IN), .Z(n10231) );
  NOR2_X1 U8900 ( .A1(n10232), .A2(n10231), .ZN(n7691) );
  NOR2_X1 U8901 ( .A1(n7692), .A2(n7691), .ZN(n10234) );
  INV_X1 U8902 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8954) );
  XOR2_X1 U8903 ( .A(n8954), .B(P1_ADDR_REG_16__SCAN_IN), .Z(n10233) );
  NOR2_X1 U8904 ( .A1(n10234), .A2(n10233), .ZN(n7693) );
  NOR2_X1 U8905 ( .A1(n7694), .A2(n7693), .ZN(n10236) );
  XOR2_X1 U8906 ( .A(n7695), .B(P1_ADDR_REG_17__SCAN_IN), .Z(n10235) );
  NOR2_X1 U8907 ( .A1(n10236), .A2(n10235), .ZN(n7696) );
  NOR2_X1 U8908 ( .A1(n7697), .A2(n7696), .ZN(n7698) );
  AND2_X1 U8909 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n7698), .ZN(n10237) );
  NOR2_X1 U8910 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10237), .ZN(n7699) );
  NOR2_X1 U8911 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n7698), .ZN(n10238) );
  NOR2_X1 U8912 ( .A1(n7699), .A2(n10238), .ZN(n7701) );
  XNOR2_X1 U8913 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7700) );
  XNOR2_X1 U8914 ( .A(n7701), .B(n7700), .ZN(ADD_1071_U4) );
  NOR2_X1 U8915 ( .A1(n7703), .A2(n7702), .ZN(n7704) );
  NAND2_X1 U8916 ( .A1(n7706), .A2(n8355), .ZN(n7709) );
  AOI22_X1 U8917 ( .A1(n8029), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n8028), .B2(
        n7707), .ZN(n7708) );
  NAND2_X2 U8918 ( .A1(n7709), .A2(n7708), .ZN(n7800) );
  NAND2_X1 U8919 ( .A1(n7800), .A2(n8184), .ZN(n7711) );
  OR2_X1 U8920 ( .A1(n7808), .A2(n8199), .ZN(n7710) );
  NAND2_X1 U8921 ( .A1(n7711), .A2(n7710), .ZN(n7712) );
  XNOR2_X1 U8922 ( .A(n7712), .B(n8188), .ZN(n7715) );
  NOR2_X1 U8923 ( .A1(n7808), .A2(n8196), .ZN(n7713) );
  AOI21_X1 U8924 ( .B1(n7800), .B2(n8185), .A(n7713), .ZN(n7714) );
  AND2_X1 U8925 ( .A1(n7715), .A2(n7714), .ZN(n7765) );
  INV_X1 U8926 ( .A(n7765), .ZN(n7716) );
  OR2_X1 U8927 ( .A1(n7715), .A2(n7714), .ZN(n7764) );
  NAND2_X1 U8928 ( .A1(n7716), .A2(n7764), .ZN(n7717) );
  XNOR2_X1 U8929 ( .A(n7766), .B(n7717), .ZN(n7732) );
  NAND2_X1 U8930 ( .A1(n4862), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7725) );
  INV_X1 U8931 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7816) );
  OR2_X1 U8932 ( .A1(n7853), .A2(n7816), .ZN(n7724) );
  NAND2_X1 U8933 ( .A1(n7719), .A2(n7718), .ZN(n7720) );
  NAND2_X1 U8934 ( .A1(n7773), .A2(n7720), .ZN(n7815) );
  OR2_X1 U8935 ( .A1(n8145), .A2(n7815), .ZN(n7723) );
  OR2_X1 U8936 ( .A1(n6787), .A2(n7721), .ZN(n7722) );
  INV_X1 U8937 ( .A(n7726), .ZN(n7728) );
  NOR2_X1 U8938 ( .A1(n9521), .A2(n7754), .ZN(n7727) );
  AOI211_X1 U8939 ( .C1(n9523), .C2(n9538), .A(n7728), .B(n7727), .ZN(n7729)
         );
  OAI21_X1 U8940 ( .B1(n9526), .B2(n7758), .A(n7729), .ZN(n7730) );
  AOI21_X1 U8941 ( .B1(n7800), .B2(n9528), .A(n7730), .ZN(n7731) );
  OAI21_X1 U8942 ( .B1(n7732), .B2(n9530), .A(n7731), .ZN(P1_U3222) );
  INV_X1 U8943 ( .A(n7754), .ZN(n9540) );
  NAND2_X1 U8944 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10250) );
  INV_X1 U8945 ( .A(n10250), .ZN(n7733) );
  AOI21_X1 U8946 ( .B1(n9523), .B2(n9540), .A(n7733), .ZN(n7736) );
  OR2_X1 U8947 ( .A1(n9521), .A2(n7734), .ZN(n7735) );
  OAI211_X1 U8948 ( .C1(n9526), .C2(n7737), .A(n7736), .B(n7735), .ZN(n7744)
         );
  NOR2_X1 U8949 ( .A1(n7739), .A2(n7738), .ZN(n7741) );
  XNOR2_X1 U8950 ( .A(n7741), .B(n7740), .ZN(n7742) );
  NOR2_X1 U8951 ( .A1(n7742), .A2(n9530), .ZN(n7743) );
  AOI211_X1 U8952 ( .C1(n7745), .C2(n9528), .A(n7744), .B(n7743), .ZN(n7746)
         );
  INV_X1 U8953 ( .A(n7746), .ZN(P1_U3215) );
  OR2_X1 U8954 ( .A1(n9925), .A2(n9540), .ZN(n7747) );
  NAND2_X1 U8955 ( .A1(n7800), .A2(n7808), .ZN(n8379) );
  NAND2_X1 U8956 ( .A1(n7749), .A2(n8507), .ZN(n7750) );
  NAND2_X1 U8957 ( .A1(n7802), .A2(n7750), .ZN(n10611) );
  INV_X1 U8958 ( .A(n8382), .ZN(n7751) );
  NOR2_X1 U8959 ( .A1(n8290), .A2(n7751), .ZN(n7752) );
  XOR2_X1 U8960 ( .A(n8507), .B(n7804), .Z(n7756) );
  OAI22_X1 U8961 ( .A1(n7754), .A2(n9779), .B1(n8300), .B2(n9808), .ZN(n7755)
         );
  AOI21_X1 U8962 ( .B1(n7756), .B2(n10397), .A(n7755), .ZN(n7757) );
  OAI21_X1 U8963 ( .B1(n10611), .B2(n9836), .A(n7757), .ZN(n10614) );
  NAND2_X1 U8964 ( .A1(n10614), .A2(n9822), .ZN(n7763) );
  OAI22_X1 U8965 ( .A1(n9822), .A2(n7759), .B1(n7758), .B2(n9819), .ZN(n7761)
         );
  INV_X1 U8966 ( .A(n7800), .ZN(n10613) );
  OAI211_X1 U8967 ( .C1(n4942), .C2(n10613), .A(n10482), .B(n7813), .ZN(n10612) );
  NOR2_X1 U8968 ( .A1(n10612), .A2(n7871), .ZN(n7760) );
  AOI211_X1 U8969 ( .C1(n9785), .C2(n7800), .A(n7761), .B(n7760), .ZN(n7762)
         );
  OAI211_X1 U8970 ( .C1(n10611), .C2(n9635), .A(n7763), .B(n7762), .ZN(
        P1_U3279) );
  NAND2_X1 U8971 ( .A1(n7767), .A2(n8355), .ZN(n7770) );
  AOI22_X1 U8972 ( .A1(n8029), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n8028), .B2(
        n7768), .ZN(n7769) );
  AOI22_X1 U8973 ( .A1(n9917), .A2(n8184), .B1(n8185), .B2(n9538), .ZN(n7771)
         );
  XNOR2_X1 U8974 ( .A(n4888), .B(n7876), .ZN(n7772) );
  XNOR2_X1 U8975 ( .A(n7877), .B(n7772), .ZN(n7784) );
  NAND2_X1 U8976 ( .A1(n4862), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7778) );
  INV_X1 U8977 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7868) );
  OR2_X1 U8978 ( .A1(n7853), .A2(n7868), .ZN(n7777) );
  INV_X1 U8979 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7882) );
  NAND2_X1 U8980 ( .A1(n7773), .A2(n7882), .ZN(n7774) );
  NAND2_X1 U8981 ( .A1(n7855), .A2(n7774), .ZN(n7885) );
  OR2_X1 U8982 ( .A1(n8145), .A2(n7885), .ZN(n7776) );
  OR2_X1 U8983 ( .A1(n6787), .A2(n10643), .ZN(n7775) );
  INV_X1 U8984 ( .A(n9520), .ZN(n9537) );
  NOR2_X1 U8985 ( .A1(n9521), .A2(n7808), .ZN(n7779) );
  AOI211_X1 U8986 ( .C1(n9523), .C2(n9537), .A(n7780), .B(n7779), .ZN(n7781)
         );
  OAI21_X1 U8987 ( .B1(n9526), .B2(n7815), .A(n7781), .ZN(n7782) );
  AOI21_X1 U8988 ( .B1(n9917), .B2(n9528), .A(n7782), .ZN(n7783) );
  OAI21_X1 U8989 ( .B1(n7784), .B2(n9530), .A(n7783), .ZN(P1_U3232) );
  INV_X1 U8990 ( .A(n8210), .ZN(n8926) );
  OAI21_X1 U8991 ( .B1(n10514), .B2(n7789), .A(n7785), .ZN(n7786) );
  AOI21_X1 U8992 ( .B1(n8917), .B2(n8926), .A(n7786), .ZN(n7787) );
  OAI21_X1 U8993 ( .B1(n7788), .B2(n10523), .A(n7787), .ZN(n7795) );
  NOR3_X1 U8994 ( .A1(n7790), .A2(n7789), .A3(n7840), .ZN(n7791) );
  AOI21_X1 U8995 ( .B1(n5443), .B2(n8873), .A(n7791), .ZN(n7793) );
  NOR2_X1 U8996 ( .A1(n7793), .A2(n7792), .ZN(n7794) );
  AOI211_X1 U8997 ( .C1(n8918), .C2(n10620), .A(n7795), .B(n7794), .ZN(n7796)
         );
  OAI21_X1 U8998 ( .B1(n8228), .B2(n10510), .A(n7796), .ZN(P2_U3226) );
  INV_X1 U8999 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8089) );
  INV_X1 U9000 ( .A(n8088), .ZN(n7798) );
  OAI222_X1 U9001 ( .A1(n9961), .A2(n8089), .B1(n8830), .B2(n7798), .C1(
        P1_U3084), .C2(n8532), .ZN(P1_U3331) );
  INV_X1 U9002 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7799) );
  OAI222_X1 U9003 ( .A1(n9385), .A2(n7799), .B1(n9380), .B2(n7798), .C1(n7797), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  INV_X1 U9004 ( .A(n7808), .ZN(n9539) );
  NAND2_X1 U9005 ( .A1(n7800), .A2(n9539), .ZN(n7801) );
  OR2_X1 U9006 ( .A1(n9917), .A2(n8300), .ZN(n8393) );
  NAND2_X1 U9007 ( .A1(n9917), .A2(n8300), .ZN(n8380) );
  OAI21_X1 U9008 ( .B1(n7803), .B2(n8509), .A(n7865), .ZN(n9921) );
  NOR2_X1 U9009 ( .A1(n7806), .A2(n7805), .ZN(n7807) );
  OAI21_X1 U9010 ( .B1(n7807), .B2(n7903), .A(n10397), .ZN(n7811) );
  OAI22_X1 U9011 ( .A1(n7808), .A2(n9779), .B1(n9520), .B2(n9808), .ZN(n7809)
         );
  INV_X1 U9012 ( .A(n7809), .ZN(n7810) );
  NAND2_X1 U9013 ( .A1(n7811), .A2(n7810), .ZN(n7812) );
  AOI21_X1 U9014 ( .B1(n9921), .B2(n9816), .A(n7812), .ZN(n9923) );
  AND2_X1 U9015 ( .A1(n7813), .A2(n9917), .ZN(n7814) );
  NOR2_X2 U9016 ( .A1(n7813), .A2(n9917), .ZN(n7870) );
  OR2_X1 U9017 ( .A1(n7814), .A2(n7870), .ZN(n9919) );
  OAI22_X1 U9018 ( .A1(n9822), .A2(n7816), .B1(n7815), .B2(n9819), .ZN(n7817)
         );
  AOI21_X1 U9019 ( .B1(n9917), .B2(n9785), .A(n7817), .ZN(n7818) );
  OAI21_X1 U9020 ( .B1(n9919), .B2(n9728), .A(n7818), .ZN(n7819) );
  AOI21_X1 U9021 ( .B1(n9921), .B2(n9826), .A(n7819), .ZN(n7820) );
  OAI21_X1 U9022 ( .B1(n9923), .B2(n9684), .A(n7820), .ZN(P1_U3278) );
  INV_X1 U9023 ( .A(n8106), .ZN(n7822) );
  NAND2_X1 U9024 ( .A1(n9373), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7821) );
  OAI211_X1 U9025 ( .C1(n7822), .C2(n9380), .A(n8776), .B(n7821), .ZN(P2_U3335) );
  INV_X1 U9026 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8107) );
  NAND2_X1 U9027 ( .A1(n8106), .A2(n9954), .ZN(n7824) );
  OR2_X1 U9028 ( .A1(n7823), .A2(P1_U3084), .ZN(n8542) );
  OAI211_X1 U9029 ( .C1(n8107), .C2(n9961), .A(n7824), .B(n8542), .ZN(P1_U3330) );
  NAND2_X1 U9030 ( .A1(n7964), .A2(n8643), .ZN(n7825) );
  NAND2_X1 U9031 ( .A1(n8221), .A2(n7841), .ZN(n8649) );
  NAND2_X1 U9032 ( .A1(n8650), .A2(n8649), .ZN(n8754) );
  INV_X1 U9033 ( .A(n8754), .ZN(n8646) );
  XNOR2_X1 U9034 ( .A(n7825), .B(n8646), .ZN(n7826) );
  NAND2_X1 U9035 ( .A1(n7826), .A2(n9234), .ZN(n7829) );
  OAI22_X1 U9036 ( .A1(n7983), .A2(n9214), .B1(n8210), .B2(n9216), .ZN(n7827)
         );
  INV_X1 U9037 ( .A(n7827), .ZN(n7828) );
  NAND2_X1 U9038 ( .A1(n7829), .A2(n7828), .ZN(n10653) );
  INV_X1 U9039 ( .A(n10653), .ZN(n7835) );
  OAI21_X1 U9040 ( .B1(n7830), .B2(n8754), .A(n7969), .ZN(n10655) );
  INV_X1 U9041 ( .A(n8221), .ZN(n10649) );
  XNOR2_X1 U9042 ( .A(n10649), .B(n7975), .ZN(n10651) );
  OAI22_X1 U9043 ( .A1(n10605), .A2(n5019), .B1(n8213), .B2(n10609), .ZN(n7831) );
  AOI21_X1 U9044 ( .B1(n8221), .B2(n9223), .A(n7831), .ZN(n7832) );
  OAI21_X1 U9045 ( .B1(n10651), .B2(n10382), .A(n7832), .ZN(n7833) );
  AOI21_X1 U9046 ( .B1(n10655), .B2(n9263), .A(n7833), .ZN(n7834) );
  OAI21_X1 U9047 ( .B1(n10607), .B2(n7835), .A(n7834), .ZN(P2_U3282) );
  INV_X1 U9048 ( .A(n7990), .ZN(n7847) );
  INV_X1 U9049 ( .A(n9217), .ZN(n9232) );
  NAND2_X1 U9050 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n8935) );
  OAI21_X1 U9051 ( .B1(n10514), .B2(n7841), .A(n8935), .ZN(n7836) );
  AOI21_X1 U9052 ( .B1(n8917), .B2(n9232), .A(n7836), .ZN(n7837) );
  OAI21_X1 U9053 ( .B1(n9237), .B2(n10523), .A(n7837), .ZN(n7838) );
  AOI21_X1 U9054 ( .B1(n9347), .B2(n8918), .A(n7838), .ZN(n7846) );
  OAI22_X1 U9055 ( .A1(n7842), .A2(n10510), .B1(n7841), .B2(n7840), .ZN(n7843)
         );
  NAND3_X1 U9056 ( .A1(n7839), .A2(n7844), .A3(n7843), .ZN(n7845) );
  OAI211_X1 U9057 ( .C1(n7847), .C2(n10510), .A(n7846), .B(n7845), .ZN(
        P2_U3243) );
  INV_X1 U9058 ( .A(n8380), .ZN(n7848) );
  OR2_X1 U9059 ( .A1(n7903), .A2(n7848), .ZN(n7852) );
  OR2_X1 U9060 ( .A1(n7849), .A2(n6899), .ZN(n7851) );
  AOI22_X1 U9061 ( .A1(n8029), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n8028), .B2(
        n10253), .ZN(n7850) );
  NAND2_X1 U9062 ( .A1(n7891), .A2(n9520), .ZN(n8405) );
  XNOR2_X1 U9063 ( .A(n7852), .B(n7901), .ZN(n7863) );
  NAND2_X1 U9064 ( .A1(n4862), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7861) );
  OR2_X1 U9065 ( .A1(n7853), .A2(n7308), .ZN(n7860) );
  NAND2_X1 U9066 ( .A1(n7855), .A2(n7854), .ZN(n7856) );
  NAND2_X1 U9067 ( .A1(n7907), .A2(n7856), .ZN(n9525) );
  OR2_X1 U9068 ( .A1(n8145), .A2(n9525), .ZN(n7859) );
  OR2_X1 U9069 ( .A1(n6787), .A2(n7857), .ZN(n7858) );
  OAI22_X1 U9070 ( .A1(n8300), .A2(n9779), .B1(n9441), .B2(n9808), .ZN(n7862)
         );
  AOI21_X1 U9071 ( .B1(n7863), .B2(n10397), .A(n7862), .ZN(n10636) );
  OR2_X1 U9072 ( .A1(n9917), .A2(n9538), .ZN(n7864) );
  OAI21_X1 U9073 ( .B1(n7866), .B2(n8510), .A(n7893), .ZN(n10641) );
  NAND2_X1 U9074 ( .A1(n10641), .A2(n7867), .ZN(n7875) );
  OAI22_X1 U9075 ( .A1(n9822), .A2(n7868), .B1(n7885), .B2(n9819), .ZN(n7873)
         );
  AND2_X2 U9076 ( .A1(n7870), .A2(n10638), .ZN(n7918) );
  INV_X1 U9077 ( .A(n7918), .ZN(n7869) );
  OAI211_X1 U9078 ( .C1(n10638), .C2(n7870), .A(n7869), .B(n10482), .ZN(n10635) );
  NOR2_X1 U9079 ( .A1(n10635), .A2(n7871), .ZN(n7872) );
  AOI211_X1 U9080 ( .C1(n9785), .C2(n7891), .A(n7873), .B(n7872), .ZN(n7874)
         );
  OAI211_X1 U9081 ( .C1(n10425), .C2(n10636), .A(n7875), .B(n7874), .ZN(
        P1_U3277) );
  NAND2_X1 U9082 ( .A1(n7891), .A2(n8185), .ZN(n7879) );
  OR2_X1 U9083 ( .A1(n9520), .A2(n8196), .ZN(n7878) );
  NAND2_X1 U9084 ( .A1(n7879), .A2(n7878), .ZN(n8017) );
  OAI22_X1 U9085 ( .A1(n10638), .A2(n6906), .B1(n9520), .B2(n8199), .ZN(n7880)
         );
  XOR2_X1 U9086 ( .A(n8197), .B(n7880), .Z(n8013) );
  XOR2_X1 U9087 ( .A(n8017), .B(n8013), .Z(n7881) );
  XNOR2_X1 U9088 ( .A(n8014), .B(n7881), .ZN(n7888) );
  INV_X1 U9089 ( .A(n9441), .ZN(n9536) );
  NOR2_X1 U9090 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7882), .ZN(n10252) );
  NOR2_X1 U9091 ( .A1(n9521), .A2(n8300), .ZN(n7883) );
  AOI211_X1 U9092 ( .C1(n9523), .C2(n9536), .A(n10252), .B(n7883), .ZN(n7884)
         );
  OAI21_X1 U9093 ( .B1(n9526), .B2(n7885), .A(n7884), .ZN(n7886) );
  AOI21_X1 U9094 ( .B1(n7891), .B2(n9528), .A(n7886), .ZN(n7887) );
  OAI21_X1 U9095 ( .B1(n7888), .B2(n9530), .A(n7887), .ZN(P1_U3213) );
  INV_X1 U9096 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7889) );
  OAI222_X1 U9097 ( .A1(n9380), .A2(n8778), .B1(P2_U3152), .B2(n7890), .C1(
        n7889), .C2(n9385), .ZN(P2_U3334) );
  OR2_X1 U9098 ( .A1(n7891), .A2(n9537), .ZN(n7892) );
  NAND2_X1 U9099 ( .A1(n7894), .A2(n8355), .ZN(n7897) );
  INV_X1 U9100 ( .A(n9553), .ZN(n7895) );
  AOI22_X1 U9101 ( .A1(n8029), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8028), .B2(
        n7895), .ZN(n7896) );
  OR2_X1 U9102 ( .A1(n9912), .A2(n9441), .ZN(n8398) );
  NAND2_X1 U9103 ( .A1(n9912), .A2(n9441), .ZN(n8397) );
  NAND2_X1 U9104 ( .A1(n8398), .A2(n8397), .ZN(n8511) );
  INV_X1 U9105 ( .A(n8511), .ZN(n7898) );
  NAND2_X1 U9106 ( .A1(n7899), .A2(n7898), .ZN(n7900) );
  NAND2_X1 U9107 ( .A1(n7901), .A2(n8380), .ZN(n7902) );
  AOI21_X1 U9108 ( .B1(n8511), .B2(n7904), .A(n7943), .ZN(n7915) );
  NAND2_X1 U9109 ( .A1(n8095), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7913) );
  INV_X1 U9110 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n7905) );
  OR2_X1 U9111 ( .A1(n4858), .A2(n7905), .ZN(n7912) );
  INV_X1 U9112 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7906) );
  NAND2_X1 U9113 ( .A1(n7907), .A2(n7906), .ZN(n7908) );
  NAND2_X1 U9114 ( .A1(n7936), .A2(n7908), .ZN(n9439) );
  OR2_X1 U9115 ( .A1(n8145), .A2(n9439), .ZN(n7911) );
  INV_X1 U9116 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7909) );
  OR2_X1 U9117 ( .A1(n6787), .A2(n7909), .ZN(n7910) );
  NAND4_X1 U9118 ( .A1(n7913), .A2(n7912), .A3(n7911), .A4(n7910), .ZN(n9806)
         );
  AOI22_X1 U9119 ( .A1(n9537), .A2(n10393), .B1(n10392), .B2(n9806), .ZN(n7914) );
  OAI21_X1 U9120 ( .B1(n7915), .B2(n9811), .A(n7914), .ZN(n7916) );
  AOI21_X1 U9121 ( .B1(n9911), .B2(n9816), .A(n7916), .ZN(n9915) );
  INV_X1 U9122 ( .A(n9912), .ZN(n7917) );
  OR2_X1 U9123 ( .A1(n7917), .A2(n7918), .ZN(n7919) );
  AND2_X1 U9124 ( .A1(n7919), .A2(n7931), .ZN(n9913) );
  NAND2_X1 U9125 ( .A1(n9913), .A2(n9825), .ZN(n7922) );
  OAI22_X1 U9126 ( .A1(n9822), .A2(n7308), .B1(n9525), .B2(n9819), .ZN(n7920)
         );
  AOI21_X1 U9127 ( .B1(n9912), .B2(n9785), .A(n7920), .ZN(n7921) );
  NAND2_X1 U9128 ( .A1(n7922), .A2(n7921), .ZN(n7923) );
  AOI21_X1 U9129 ( .B1(n9911), .B2(n9826), .A(n7923), .ZN(n7924) );
  OAI21_X1 U9130 ( .B1(n9915), .B2(n10425), .A(n7924), .ZN(P1_U3276) );
  NAND2_X1 U9131 ( .A1(n9912), .A2(n9536), .ZN(n7925) );
  NAND2_X1 U9132 ( .A1(n7927), .A2(n8355), .ZN(n7929) );
  AOI22_X1 U9133 ( .A1(n8029), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8028), .B2(
        n9570), .ZN(n7928) );
  AND2_X1 U9134 ( .A1(n8009), .A2(n9806), .ZN(n8805) );
  INV_X1 U9135 ( .A(n8805), .ZN(n8315) );
  INV_X1 U9136 ( .A(n9806), .ZN(n9450) );
  NAND2_X1 U9137 ( .A1(n9908), .A2(n9450), .ZN(n8806) );
  NAND2_X1 U9138 ( .A1(n8315), .A2(n8806), .ZN(n8781) );
  XNOR2_X1 U9139 ( .A(n8782), .B(n8781), .ZN(n9910) );
  INV_X1 U9140 ( .A(n9817), .ZN(n7930) );
  AOI211_X1 U9141 ( .C1(n9908), .C2(n7931), .A(n10548), .B(n7930), .ZN(n9907)
         );
  NOR2_X1 U9142 ( .A1(n8009), .A2(n9818), .ZN(n7934) );
  INV_X1 U9143 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7932) );
  OAI22_X1 U9144 ( .A1(n9822), .A2(n7932), .B1(n9439), .B2(n9819), .ZN(n7933)
         );
  AOI211_X1 U9145 ( .C1(n9907), .C2(n7935), .A(n7934), .B(n7933), .ZN(n7946)
         );
  NAND2_X1 U9146 ( .A1(n4862), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n7942) );
  INV_X1 U9147 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9821) );
  OR2_X1 U9148 ( .A1(n7853), .A2(n9821), .ZN(n7941) );
  NAND2_X1 U9149 ( .A1(n7936), .A2(n9449), .ZN(n7937) );
  NAND2_X1 U9150 ( .A1(n8033), .A2(n7937), .ZN(n9820) );
  OR2_X1 U9151 ( .A1(n8145), .A2(n9820), .ZN(n7940) );
  INV_X1 U9152 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n7938) );
  OR2_X1 U9153 ( .A1(n6787), .A2(n7938), .ZN(n7939) );
  INV_X1 U9154 ( .A(n8397), .ZN(n8408) );
  INV_X1 U9155 ( .A(n8781), .ZN(n8514) );
  XNOR2_X1 U9156 ( .A(n8807), .B(n8514), .ZN(n7944) );
  OAI222_X1 U9157 ( .A1(n9808), .A2(n9497), .B1(n9779), .B2(n9441), .C1(n7944), 
        .C2(n9811), .ZN(n9906) );
  NAND2_X1 U9158 ( .A1(n9906), .A2(n9822), .ZN(n7945) );
  OAI211_X1 U9159 ( .C1(n9910), .C2(n9804), .A(n7946), .B(n7945), .ZN(P1_U3275) );
  INV_X1 U9160 ( .A(n7947), .ZN(n7949) );
  NAND2_X1 U9161 ( .A1(n7949), .A2(n7948), .ZN(n7950) );
  XNOR2_X1 U9162 ( .A(n7951), .B(n7950), .ZN(n7957) );
  OAI21_X1 U9163 ( .B1(n10517), .B2(n9215), .A(n7952), .ZN(n7953) );
  AOI21_X1 U9164 ( .B1(n8906), .B2(n9232), .A(n7953), .ZN(n7954) );
  OAI21_X1 U9165 ( .B1(n9220), .B2(n10523), .A(n7954), .ZN(n7955) );
  AOI21_X1 U9166 ( .B1(n9337), .B2(n8918), .A(n7955), .ZN(n7956) );
  OAI21_X1 U9167 ( .B1(n7957), .B2(n10510), .A(n7956), .ZN(P2_U3230) );
  INV_X1 U9168 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7959) );
  INV_X1 U9169 ( .A(n8138), .ZN(n7960) );
  OAI222_X1 U9170 ( .A1(n9385), .A2(n7959), .B1(n9380), .B2(n7960), .C1(n7958), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  INV_X1 U9171 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8139) );
  OAI222_X1 U9172 ( .A1(n8139), .A2(n9961), .B1(P1_U3084), .B2(n7961), .C1(
        n8830), .C2(n7960), .ZN(P1_U3328) );
  INV_X1 U9173 ( .A(n8643), .ZN(n7962) );
  NOR2_X1 U9174 ( .A1(n8754), .A2(n7962), .ZN(n7963) );
  NAND2_X1 U9175 ( .A1(n7964), .A2(n7963), .ZN(n7965) );
  NAND2_X1 U9176 ( .A1(n9347), .A2(n7983), .ZN(n8653) );
  OR2_X1 U9177 ( .A1(n9347), .A2(n7983), .ZN(n8654) );
  INV_X1 U9178 ( .A(n8654), .ZN(n8552) );
  AOI21_X1 U9179 ( .B1(n9229), .B2(n8653), .A(n8552), .ZN(n7966) );
  OR2_X1 U9180 ( .A1(n9343), .A2(n9217), .ZN(n8658) );
  NAND2_X1 U9181 ( .A1(n9343), .A2(n9217), .ZN(n8657) );
  XNOR2_X1 U9182 ( .A(n7966), .B(n8757), .ZN(n7967) );
  INV_X1 U9183 ( .A(n8554), .ZN(n9193) );
  INV_X1 U9184 ( .A(n7983), .ZN(n8925) );
  AOI222_X1 U9185 ( .A1(n9234), .A2(n7967), .B1(n9193), .B2(n10587), .C1(n8925), .C2(n9230), .ZN(n9345) );
  OR2_X1 U9186 ( .A1(n8221), .A2(n9231), .ZN(n7968) );
  NAND2_X1 U9187 ( .A1(n7969), .A2(n7968), .ZN(n9243) );
  NAND2_X1 U9188 ( .A1(n8654), .A2(n8653), .ZN(n9228) );
  NAND2_X1 U9189 ( .A1(n9243), .A2(n9228), .ZN(n7971) );
  OR2_X1 U9190 ( .A1(n9347), .A2(n8925), .ZN(n7970) );
  INV_X1 U9191 ( .A(n8757), .ZN(n7972) );
  OAI21_X1 U9192 ( .B1(n4882), .B2(n7972), .A(n5184), .ZN(n9346) );
  INV_X1 U9193 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7973) );
  OAI22_X1 U9194 ( .A1(n10605), .A2(n7973), .B1(n7986), .B2(n10609), .ZN(n7974) );
  AOI21_X1 U9195 ( .B1(n9343), .B2(n9223), .A(n7974), .ZN(n7978) );
  AOI21_X1 U9196 ( .B1(n9343), .B2(n9235), .A(n10650), .ZN(n7976) );
  AND2_X1 U9197 ( .A1(n7976), .A2(n9212), .ZN(n9342) );
  NAND2_X1 U9198 ( .A1(n9342), .A2(n9186), .ZN(n7977) );
  OAI211_X1 U9199 ( .C1(n9346), .C2(n9244), .A(n7978), .B(n7977), .ZN(n7979)
         );
  INV_X1 U9200 ( .A(n7979), .ZN(n7980) );
  OAI21_X1 U9201 ( .B1(n10607), .B2(n9345), .A(n7980), .ZN(P2_U3280) );
  INV_X1 U9202 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7982) );
  OAI222_X1 U9203 ( .A1(n9385), .A2(n7982), .B1(n9380), .B2(n7981), .C1(n5582), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  NAND2_X1 U9204 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8952) );
  OAI21_X1 U9205 ( .B1(n10514), .B2(n7983), .A(n8952), .ZN(n7984) );
  AOI21_X1 U9206 ( .B1(n8917), .B2(n9193), .A(n7984), .ZN(n7985) );
  OAI21_X1 U9207 ( .B1(n7986), .B2(n10523), .A(n7985), .ZN(n7992) );
  AOI22_X1 U9208 ( .A1(n7987), .A2(n8873), .B1(n8875), .B2(n8925), .ZN(n7988)
         );
  NOR3_X1 U9209 ( .A1(n7990), .A2(n7989), .A3(n7988), .ZN(n7991) );
  AOI211_X1 U9210 ( .C1(n8918), .C2(n9343), .A(n7992), .B(n7991), .ZN(n7993)
         );
  OAI21_X1 U9211 ( .B1(n7994), .B2(n10510), .A(n7993), .ZN(P2_U3228) );
  NAND2_X1 U9212 ( .A1(n7995), .A2(n8355), .ZN(n7997) );
  AOI22_X1 U9213 ( .A1(n8029), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n8028), .B2(
        n10415), .ZN(n7996) );
  NAND2_X1 U9214 ( .A1(n9892), .A2(n8184), .ZN(n8006) );
  NAND2_X1 U9215 ( .A1(n4862), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8004) );
  INV_X1 U9216 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n7998) );
  OR2_X1 U9217 ( .A1(n6787), .A2(n7998), .ZN(n8003) );
  INV_X1 U9218 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7999) );
  NAND2_X1 U9219 ( .A1(n8035), .A2(n7999), .ZN(n8000) );
  NAND2_X1 U9220 ( .A1(n8055), .A2(n8000), .ZN(n9772) );
  OR2_X1 U9221 ( .A1(n8145), .A2(n9772), .ZN(n8002) );
  INV_X1 U9222 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9773) );
  OR2_X1 U9223 ( .A1(n7853), .A2(n9773), .ZN(n8001) );
  OR2_X1 U9224 ( .A1(n9754), .A2(n8199), .ZN(n8005) );
  NAND2_X1 U9225 ( .A1(n8006), .A2(n8005), .ZN(n8007) );
  XNOR2_X1 U9226 ( .A(n8007), .B(n8197), .ZN(n8049) );
  AOI22_X1 U9227 ( .A1(n9892), .A2(n8185), .B1(n8155), .B2(n9798), .ZN(n8047)
         );
  INV_X1 U9228 ( .A(n8047), .ZN(n8048) );
  OAI22_X1 U9229 ( .A1(n8009), .A2(n6906), .B1(n9450), .B2(n8199), .ZN(n8008)
         );
  XNOR2_X1 U9230 ( .A(n8008), .B(n8197), .ZN(n8020) );
  OAI22_X1 U9231 ( .A1(n8009), .A2(n8199), .B1(n9450), .B2(n8196), .ZN(n8019)
         );
  NAND2_X1 U9232 ( .A1(n8014), .A2(n8013), .ZN(n8016) );
  NAND2_X1 U9233 ( .A1(n9912), .A2(n8184), .ZN(n8011) );
  OR2_X1 U9234 ( .A1(n9441), .A2(n8199), .ZN(n8010) );
  NAND2_X1 U9235 ( .A1(n8011), .A2(n8010), .ZN(n8012) );
  XNOR2_X1 U9236 ( .A(n8012), .B(n8197), .ZN(n8015) );
  AOI211_X2 U9237 ( .C1(n8017), .C2(n8016), .A(n8015), .B(n8018), .ZN(n9514)
         );
  AOI22_X1 U9238 ( .A1(n9912), .A2(n8185), .B1(n8155), .B2(n9536), .ZN(n9517)
         );
  OAI211_X1 U9239 ( .C1(n8018), .C2(n8017), .A(n8016), .B(n8015), .ZN(n9515)
         );
  XNOR2_X1 U9240 ( .A(n8020), .B(n8019), .ZN(n9438) );
  OR2_X1 U9241 ( .A1(n8021), .A2(n6899), .ZN(n8023) );
  AOI22_X1 U9242 ( .A1(n8029), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8028), .B2(
        n9588), .ZN(n8022) );
  AOI22_X1 U9243 ( .A1(n9901), .A2(n8184), .B1(n8185), .B2(n9799), .ZN(n8024)
         );
  XOR2_X1 U9244 ( .A(n8197), .B(n8024), .Z(n8026) );
  OAI22_X1 U9245 ( .A1(n5140), .A2(n8199), .B1(n9497), .B2(n8196), .ZN(n8025)
         );
  NAND2_X1 U9246 ( .A1(n8026), .A2(n8025), .ZN(n9446) );
  OR2_X1 U9247 ( .A1(n8027), .A2(n6899), .ZN(n8031) );
  AOI22_X1 U9248 ( .A1(n8029), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n8028), .B2(
        n9598), .ZN(n8030) );
  INV_X1 U9249 ( .A(n9895), .ZN(n9795) );
  NAND2_X1 U9250 ( .A1(n4862), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8040) );
  INV_X1 U9251 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9586) );
  OR2_X1 U9252 ( .A1(n6787), .A2(n9586), .ZN(n8039) );
  INV_X1 U9253 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8032) );
  NAND2_X1 U9254 ( .A1(n8033), .A2(n8032), .ZN(n8034) );
  NAND2_X1 U9255 ( .A1(n8035), .A2(n8034), .ZN(n9792) );
  OR2_X1 U9256 ( .A1(n8145), .A2(n9792), .ZN(n8038) );
  INV_X1 U9257 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8036) );
  OR2_X1 U9258 ( .A1(n7853), .A2(n8036), .ZN(n8037) );
  OAI22_X1 U9259 ( .A1(n9795), .A2(n6906), .B1(n9809), .B2(n8199), .ZN(n8041)
         );
  XNOR2_X1 U9260 ( .A(n8041), .B(n8197), .ZN(n8043) );
  INV_X1 U9261 ( .A(n9809), .ZN(n9535) );
  INV_X1 U9262 ( .A(n8042), .ZN(n8045) );
  INV_X1 U9263 ( .A(n8043), .ZN(n8044) );
  XNOR2_X1 U9264 ( .A(n8049), .B(n8047), .ZN(n9411) );
  NAND2_X1 U9265 ( .A1(n8050), .A2(n8355), .ZN(n8053) );
  OR2_X1 U9266 ( .A1(n4865), .A2(n8051), .ZN(n8052) );
  NAND2_X1 U9267 ( .A1(n9885), .A2(n8184), .ZN(n8063) );
  NAND2_X1 U9268 ( .A1(n4862), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8061) );
  NAND2_X1 U9269 ( .A1(n8055), .A2(n8054), .ZN(n8056) );
  NAND2_X1 U9270 ( .A1(n8077), .A2(n8056), .ZN(n9765) );
  OR2_X1 U9271 ( .A1(n9765), .A2(n8145), .ZN(n8060) );
  INV_X1 U9272 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n8057) );
  OR2_X1 U9273 ( .A1(n6787), .A2(n8057), .ZN(n8059) );
  INV_X1 U9274 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9766) );
  OR2_X1 U9275 ( .A1(n7853), .A2(n9766), .ZN(n8058) );
  OR2_X1 U9276 ( .A1(n9780), .A2(n8199), .ZN(n8062) );
  NAND2_X1 U9277 ( .A1(n8063), .A2(n8062), .ZN(n8064) );
  XNOR2_X1 U9278 ( .A(n8064), .B(n8197), .ZN(n9465) );
  NAND2_X1 U9279 ( .A1(n9885), .A2(n8185), .ZN(n8066) );
  OR2_X1 U9280 ( .A1(n9780), .A2(n8196), .ZN(n8065) );
  NAND2_X1 U9281 ( .A1(n8066), .A2(n8065), .ZN(n9464) );
  NOR2_X1 U9282 ( .A1(n9465), .A2(n9464), .ZN(n8069) );
  INV_X1 U9283 ( .A(n9465), .ZN(n8068) );
  INV_X1 U9284 ( .A(n9464), .ZN(n8067) );
  OR2_X1 U9285 ( .A1(n4864), .A2(n8071), .ZN(n8072) );
  NAND2_X1 U9286 ( .A1(n9881), .A2(n8184), .ZN(n8083) );
  NAND2_X1 U9287 ( .A1(n8095), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8075) );
  NAND2_X1 U9288 ( .A1(n4862), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8074) );
  AND2_X1 U9289 ( .A1(n8075), .A2(n8074), .ZN(n8081) );
  NAND2_X1 U9290 ( .A1(n8077), .A2(n8076), .ZN(n8078) );
  AND2_X1 U9291 ( .A1(n8093), .A2(n8078), .ZN(n9746) );
  NAND2_X1 U9292 ( .A1(n9746), .A2(n8166), .ZN(n8080) );
  NAND2_X1 U9293 ( .A1(n6746), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n8079) );
  NAND2_X1 U9294 ( .A1(n9720), .A2(n8185), .ZN(n8082) );
  NAND2_X1 U9295 ( .A1(n8083), .A2(n8082), .ZN(n8084) );
  XNOR2_X1 U9296 ( .A(n8084), .B(n8188), .ZN(n8087) );
  NOR2_X1 U9297 ( .A1(n9755), .A2(n8196), .ZN(n8085) );
  AOI21_X1 U9298 ( .B1(n9881), .B2(n8185), .A(n8085), .ZN(n8086) );
  NOR2_X1 U9299 ( .A1(n8087), .A2(n8086), .ZN(n9419) );
  NAND2_X1 U9300 ( .A1(n8087), .A2(n8086), .ZN(n9417) );
  NAND2_X1 U9301 ( .A1(n8088), .A2(n8355), .ZN(n8091) );
  OR2_X1 U9302 ( .A1(n4865), .A2(n8089), .ZN(n8090) );
  NAND2_X1 U9303 ( .A1(n9874), .A2(n8184), .ZN(n8100) );
  INV_X1 U9304 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8092) );
  NAND2_X1 U9305 ( .A1(n8093), .A2(n8092), .ZN(n8094) );
  NAND2_X1 U9306 ( .A1(n8111), .A2(n8094), .ZN(n9724) );
  OR2_X1 U9307 ( .A1(n9724), .A2(n8145), .ZN(n8098) );
  AOI22_X1 U9308 ( .A1(n4862), .A2(P1_REG0_REG_22__SCAN_IN), .B1(n6746), .B2(
        P1_REG1_REG_22__SCAN_IN), .ZN(n8097) );
  NAND2_X1 U9309 ( .A1(n8095), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8096) );
  NAND2_X1 U9310 ( .A1(n9709), .A2(n8185), .ZN(n8099) );
  NAND2_X1 U9311 ( .A1(n8100), .A2(n8099), .ZN(n8101) );
  XNOR2_X1 U9312 ( .A(n8101), .B(n8197), .ZN(n8102) );
  AOI22_X1 U9313 ( .A1(n9874), .A2(n8185), .B1(n8155), .B2(n9709), .ZN(n8103)
         );
  XNOR2_X1 U9314 ( .A(n8102), .B(n8103), .ZN(n9475) );
  INV_X1 U9315 ( .A(n8102), .ZN(n8104) );
  NAND2_X1 U9316 ( .A1(n8104), .A2(n8103), .ZN(n8105) );
  NAND2_X1 U9317 ( .A1(n8106), .A2(n8355), .ZN(n8109) );
  OR2_X1 U9318 ( .A1(n4864), .A2(n8107), .ZN(n8108) );
  INV_X1 U9319 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8110) );
  NAND2_X1 U9320 ( .A1(n8111), .A2(n8110), .ZN(n8112) );
  NAND2_X1 U9321 ( .A1(n8123), .A2(n8112), .ZN(n9702) );
  OR2_X1 U9322 ( .A1(n9702), .A2(n8145), .ZN(n8118) );
  INV_X1 U9323 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n8115) );
  NAND2_X1 U9324 ( .A1(n6746), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8114) );
  NAND2_X1 U9325 ( .A1(n4862), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8113) );
  OAI211_X1 U9326 ( .C1(n7853), .C2(n8115), .A(n8114), .B(n8113), .ZN(n8116)
         );
  INV_X1 U9327 ( .A(n8116), .ZN(n8117) );
  OAI22_X1 U9328 ( .A1(n9705), .A2(n6906), .B1(n9460), .B2(n8199), .ZN(n8119)
         );
  XOR2_X1 U9329 ( .A(n8197), .B(n8119), .Z(n9403) );
  AOI22_X1 U9330 ( .A1(n9869), .A2(n8185), .B1(n8155), .B2(n9721), .ZN(n9402)
         );
  OR2_X1 U9331 ( .A1(n8778), .A2(n6899), .ZN(n8121) );
  INV_X1 U9332 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8780) );
  OR2_X1 U9333 ( .A1(n4865), .A2(n8780), .ZN(n8120) );
  NAND2_X1 U9334 ( .A1(n9866), .A2(n8184), .ZN(n8132) );
  NAND2_X1 U9335 ( .A1(n8123), .A2(n8122), .ZN(n8124) );
  AND2_X1 U9336 ( .A1(n8143), .A2(n8124), .ZN(n9692) );
  NAND2_X1 U9337 ( .A1(n9692), .A2(n8166), .ZN(n8130) );
  INV_X1 U9338 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n8127) );
  NAND2_X1 U9339 ( .A1(n4862), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8126) );
  NAND2_X1 U9340 ( .A1(n6746), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8125) );
  OAI211_X1 U9341 ( .C1(n8127), .C2(n7853), .A(n8126), .B(n8125), .ZN(n8128)
         );
  INV_X1 U9342 ( .A(n8128), .ZN(n8129) );
  NAND2_X1 U9343 ( .A1(n9710), .A2(n8185), .ZN(n8131) );
  NAND2_X1 U9344 ( .A1(n8132), .A2(n8131), .ZN(n8133) );
  XNOR2_X1 U9345 ( .A(n8133), .B(n8197), .ZN(n8134) );
  AOI22_X1 U9346 ( .A1(n9866), .A2(n8185), .B1(n8155), .B2(n9710), .ZN(n8135)
         );
  XNOR2_X1 U9347 ( .A(n8134), .B(n8135), .ZN(n9457) );
  INV_X1 U9348 ( .A(n8134), .ZN(n8136) );
  NAND2_X1 U9349 ( .A1(n8136), .A2(n8135), .ZN(n8137) );
  NAND2_X1 U9350 ( .A1(n8138), .A2(n8355), .ZN(n8141) );
  OR2_X1 U9351 ( .A1(n4864), .A2(n8139), .ZN(n8140) );
  NAND2_X1 U9352 ( .A1(n9859), .A2(n8184), .ZN(n8153) );
  INV_X1 U9353 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8142) );
  NAND2_X1 U9354 ( .A1(n8143), .A2(n8142), .ZN(n8144) );
  NAND2_X1 U9355 ( .A1(n8163), .A2(n8144), .ZN(n9670) );
  OR2_X1 U9356 ( .A1(n9670), .A2(n8145), .ZN(n8151) );
  INV_X1 U9357 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n8148) );
  NAND2_X1 U9358 ( .A1(n6746), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8147) );
  NAND2_X1 U9359 ( .A1(n4862), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8146) );
  OAI211_X1 U9360 ( .C1(n7853), .C2(n8148), .A(n8147), .B(n8146), .ZN(n8149)
         );
  INV_X1 U9361 ( .A(n8149), .ZN(n8150) );
  NAND2_X1 U9362 ( .A1(n9533), .A2(n8185), .ZN(n8152) );
  NAND2_X1 U9363 ( .A1(n8153), .A2(n8152), .ZN(n8154) );
  XNOR2_X1 U9364 ( .A(n8154), .B(n8197), .ZN(n8156) );
  AOI22_X1 U9365 ( .A1(n9859), .A2(n8185), .B1(n8155), .B2(n9533), .ZN(n8157)
         );
  XNOR2_X1 U9366 ( .A(n8156), .B(n8157), .ZN(n9428) );
  NAND2_X1 U9367 ( .A1(n9427), .A2(n9428), .ZN(n8160) );
  INV_X1 U9368 ( .A(n8156), .ZN(n8158) );
  NAND2_X1 U9369 ( .A1(n8158), .A2(n8157), .ZN(n8159) );
  NAND2_X1 U9370 ( .A1(n9384), .A2(n8355), .ZN(n8162) );
  INV_X1 U9371 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9962) );
  OR2_X1 U9372 ( .A1(n4865), .A2(n9962), .ZN(n8161) );
  NAND2_X1 U9373 ( .A1(n8163), .A2(n9506), .ZN(n8164) );
  NAND2_X1 U9374 ( .A1(n9662), .A2(n8166), .ZN(n8172) );
  INV_X1 U9375 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n8169) );
  NAND2_X1 U9376 ( .A1(n6746), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8168) );
  NAND2_X1 U9377 ( .A1(n4862), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8167) );
  OAI211_X1 U9378 ( .C1(n7853), .C2(n8169), .A(n8168), .B(n8167), .ZN(n8170)
         );
  INV_X1 U9379 ( .A(n8170), .ZN(n8171) );
  NOR2_X1 U9380 ( .A1(n9647), .A2(n8196), .ZN(n8173) );
  AOI21_X1 U9381 ( .B1(n9854), .B2(n8185), .A(n8173), .ZN(n8178) );
  NAND2_X1 U9382 ( .A1(n9854), .A2(n8184), .ZN(n8175) );
  NAND2_X1 U9383 ( .A1(n9677), .A2(n8185), .ZN(n8174) );
  NAND2_X1 U9384 ( .A1(n8175), .A2(n8174), .ZN(n8176) );
  XNOR2_X1 U9385 ( .A(n8176), .B(n8197), .ZN(n8177) );
  XOR2_X1 U9386 ( .A(n8178), .B(n8177), .Z(n9503) );
  INV_X1 U9387 ( .A(n8177), .ZN(n8179) );
  OR2_X1 U9388 ( .A1(n8179), .A2(n8178), .ZN(n8180) );
  NAND2_X1 U9389 ( .A1(n9382), .A2(n8355), .ZN(n8183) );
  INV_X1 U9390 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8181) );
  OR2_X1 U9391 ( .A1(n4864), .A2(n8181), .ZN(n8182) );
  NAND2_X1 U9392 ( .A1(n9848), .A2(n8184), .ZN(n8187) );
  NAND2_X1 U9393 ( .A1(n9622), .A2(n8185), .ZN(n8186) );
  NAND2_X1 U9394 ( .A1(n8187), .A2(n8186), .ZN(n8189) );
  XNOR2_X1 U9395 ( .A(n8189), .B(n8188), .ZN(n8193) );
  NOR2_X1 U9396 ( .A1(n9659), .A2(n8196), .ZN(n8190) );
  AOI21_X1 U9397 ( .B1(n9848), .B2(n8185), .A(n8190), .ZN(n8192) );
  NAND2_X1 U9398 ( .A1(n8193), .A2(n8192), .ZN(n9391) );
  NAND2_X1 U9399 ( .A1(n8826), .A2(n8355), .ZN(n8195) );
  INV_X1 U9400 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8827) );
  OR2_X1 U9401 ( .A1(n4865), .A2(n8827), .ZN(n8194) );
  INV_X1 U9402 ( .A(n9843), .ZN(n8799) );
  OAI22_X1 U9403 ( .A1(n8799), .A2(n8199), .B1(n9648), .B2(n8196), .ZN(n8198)
         );
  XNOR2_X1 U9404 ( .A(n8198), .B(n8197), .ZN(n8201) );
  OAI22_X1 U9405 ( .A1(n8799), .A2(n6906), .B1(n9648), .B2(n8199), .ZN(n8200)
         );
  XNOR2_X1 U9406 ( .A(n8201), .B(n8200), .ZN(n8202) );
  XNOR2_X1 U9407 ( .A(n8203), .B(n8202), .ZN(n8208) );
  NOR2_X1 U9408 ( .A1(n9659), .A2(n9521), .ZN(n8206) );
  AOI22_X1 U9409 ( .A1(n9621), .A2(n9523), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8204) );
  OAI21_X1 U9410 ( .B1(n9526), .B2(n9629), .A(n8204), .ZN(n8205) );
  AOI211_X1 U9411 ( .C1(n9843), .C2(n9528), .A(n8206), .B(n8205), .ZN(n8207)
         );
  OAI21_X1 U9412 ( .B1(n8208), .B2(n9530), .A(n8207), .ZN(P1_U3218) );
  OAI21_X1 U9413 ( .B1(n10514), .B2(n8210), .A(n8209), .ZN(n8211) );
  AOI21_X1 U9414 ( .B1(n8917), .B2(n8925), .A(n8211), .ZN(n8212) );
  OAI21_X1 U9415 ( .B1(n8213), .B2(n10523), .A(n8212), .ZN(n8220) );
  INV_X1 U9416 ( .A(n8214), .ZN(n8218) );
  AOI22_X1 U9417 ( .A1(n8215), .A2(n8873), .B1(n8875), .B2(n8926), .ZN(n8216)
         );
  NOR3_X1 U9418 ( .A1(n8218), .A2(n8217), .A3(n8216), .ZN(n8219) );
  AOI211_X1 U9419 ( .C1(n8918), .C2(n8221), .A(n8220), .B(n8219), .ZN(n8222)
         );
  OAI21_X1 U9420 ( .B1(n7839), .B2(n10510), .A(n8222), .ZN(P2_U3217) );
  OAI21_X1 U9421 ( .B1(n10514), .B2(n8224), .A(n8223), .ZN(n8225) );
  AOI21_X1 U9422 ( .B1(n8917), .B2(n9231), .A(n8225), .ZN(n8226) );
  OAI21_X1 U9423 ( .B1(n8227), .B2(n10523), .A(n8226), .ZN(n8234) );
  INV_X1 U9424 ( .A(n8228), .ZN(n8232) );
  AOI22_X1 U9425 ( .A1(n8229), .A2(n8873), .B1(n8875), .B2(n10588), .ZN(n8230)
         );
  NOR3_X1 U9426 ( .A1(n8232), .A2(n8231), .A3(n8230), .ZN(n8233) );
  AOI211_X1 U9427 ( .C1(n8918), .C2(n10627), .A(n8234), .B(n8233), .ZN(n8235)
         );
  OAI21_X1 U9428 ( .B1(n8214), .B2(n10510), .A(n8235), .ZN(P2_U3236) );
  INV_X1 U9429 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8344) );
  INV_X1 U9430 ( .A(n8236), .ZN(n8237) );
  NAND2_X1 U9431 ( .A1(n8237), .A2(n10104), .ZN(n8238) );
  MUX2_X1 U9432 ( .A(n8344), .B(n9378), .S(n8253), .Z(n8240) );
  NAND2_X1 U9433 ( .A1(n8240), .A2(n10102), .ZN(n8246) );
  INV_X1 U9434 ( .A(n8240), .ZN(n8241) );
  NAND2_X1 U9435 ( .A1(n8241), .A2(SI_29_), .ZN(n8242) );
  INV_X1 U9436 ( .A(n8549), .ZN(n9379) );
  OAI222_X1 U9437 ( .A1(n9961), .A2(n8344), .B1(n8830), .B2(n9379), .C1(n8243), 
        .C2(P1_U3084), .ZN(P1_U3324) );
  INV_X1 U9438 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8829) );
  INV_X1 U9439 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8247) );
  MUX2_X1 U9440 ( .A(n8829), .B(n8247), .S(n8253), .Z(n8249) );
  INV_X1 U9441 ( .A(SI_30_), .ZN(n8248) );
  NAND2_X1 U9442 ( .A1(n8249), .A2(n8248), .ZN(n8252) );
  INV_X1 U9443 ( .A(n8249), .ZN(n8250) );
  NAND2_X1 U9444 ( .A1(n8250), .A2(SI_30_), .ZN(n8251) );
  MUX2_X1 U9445 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8253), .Z(n8255) );
  INV_X1 U9446 ( .A(SI_31_), .ZN(n8254) );
  XNOR2_X1 U9447 ( .A(n8255), .B(n8254), .ZN(n8256) );
  INV_X1 U9448 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9951) );
  NOR2_X1 U9449 ( .A1(n4865), .A2(n9951), .ZN(n8258) );
  INV_X1 U9450 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n8262) );
  NAND2_X1 U9451 ( .A1(n4862), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8261) );
  INV_X1 U9452 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n8259) );
  OR2_X1 U9453 ( .A1(n6787), .A2(n8259), .ZN(n8260) );
  OAI211_X1 U9454 ( .C1(n7853), .C2(n8262), .A(n8261), .B(n8260), .ZN(n9608)
         );
  AND2_X1 U9455 ( .A1(n9831), .A2(n9608), .ZN(n8456) );
  NOR4_X1 U9456 ( .A1(n8456), .A2(n8264), .A3(n8263), .A4(n8542), .ZN(n8546)
         );
  NAND2_X1 U9457 ( .A1(n9843), .A2(n9648), .ZN(n8450) );
  NAND2_X1 U9458 ( .A1(n9848), .A2(n9659), .ZN(n8449) );
  INV_X1 U9459 ( .A(n8351), .ZN(n8369) );
  MUX2_X1 U9460 ( .A(n8449), .B(n8818), .S(n8369), .Z(n8343) );
  NAND2_X1 U9461 ( .A1(n9854), .A2(n9647), .ZN(n8447) );
  OR2_X1 U9462 ( .A1(n9854), .A2(n9647), .ZN(n8371) );
  MUX2_X1 U9463 ( .A(n8447), .B(n8371), .S(n8351), .Z(n8341) );
  NAND2_X1 U9464 ( .A1(n8371), .A2(n8447), .ZN(n9657) );
  INV_X1 U9465 ( .A(n9657), .ZN(n8339) );
  NAND2_X1 U9466 ( .A1(n9859), .A2(n9690), .ZN(n8444) );
  MUX2_X1 U9467 ( .A(n8444), .B(n8816), .S(n8369), .Z(n8338) );
  NAND2_X1 U9468 ( .A1(n9866), .A2(n9430), .ZN(n8489) );
  NAND2_X1 U9469 ( .A1(n9869), .A2(n9460), .ZN(n8469) );
  NAND2_X1 U9470 ( .A1(n8489), .A2(n8469), .ZN(n8265) );
  OR2_X1 U9471 ( .A1(n9866), .A2(n9430), .ZN(n8815) );
  OR2_X1 U9472 ( .A1(n9869), .A2(n9460), .ZN(n8814) );
  NAND2_X1 U9473 ( .A1(n8815), .A2(n8814), .ZN(n8443) );
  MUX2_X1 U9474 ( .A(n8265), .B(n8443), .S(n8369), .Z(n8336) );
  XNOR2_X1 U9475 ( .A(n8266), .B(n8351), .ZN(n8267) );
  NAND2_X1 U9476 ( .A1(n8267), .A2(n8494), .ZN(n8274) );
  INV_X1 U9477 ( .A(n8268), .ZN(n8270) );
  MUX2_X1 U9478 ( .A(n8270), .B(n8269), .S(n8351), .Z(n8272) );
  INV_X1 U9479 ( .A(n8498), .ZN(n8271) );
  NOR2_X1 U9480 ( .A1(n8272), .A2(n8271), .ZN(n8273) );
  NAND2_X1 U9481 ( .A1(n8274), .A2(n8273), .ZN(n8280) );
  AND2_X1 U9482 ( .A1(n8428), .A2(n8275), .ZN(n8462) );
  AOI21_X1 U9483 ( .B1(n8280), .B2(n8462), .A(n8276), .ZN(n8282) );
  AND2_X1 U9484 ( .A1(n8402), .A2(n8277), .ZN(n8279) );
  INV_X1 U9485 ( .A(n8428), .ZN(n8278) );
  AOI21_X1 U9486 ( .B1(n8280), .B2(n8279), .A(n8278), .ZN(n8281) );
  MUX2_X1 U9487 ( .A(n8282), .B(n8281), .S(n8351), .Z(n8285) );
  MUX2_X1 U9488 ( .A(n8403), .B(n8387), .S(n8351), .Z(n8283) );
  OAI21_X1 U9489 ( .B1(n8285), .B2(n8284), .A(n8283), .ZN(n8287) );
  NAND2_X1 U9490 ( .A1(n8287), .A2(n8286), .ZN(n8289) );
  MUX2_X1 U9491 ( .A(n8381), .B(n8386), .S(n8351), .Z(n8288) );
  NAND3_X1 U9492 ( .A1(n8289), .A2(n8505), .A3(n8288), .ZN(n8292) );
  INV_X1 U9493 ( .A(n8290), .ZN(n8506) );
  MUX2_X1 U9494 ( .A(n8382), .B(n8388), .S(n8369), .Z(n8291) );
  NAND3_X1 U9495 ( .A1(n8292), .A2(n8506), .A3(n8291), .ZN(n8295) );
  MUX2_X1 U9496 ( .A(n8385), .B(n8389), .S(n8351), .Z(n8293) );
  AND2_X1 U9497 ( .A1(n8507), .A2(n8293), .ZN(n8294) );
  NAND2_X1 U9498 ( .A1(n8295), .A2(n8294), .ZN(n8297) );
  NAND2_X1 U9499 ( .A1(n8297), .A2(n8379), .ZN(n8296) );
  NAND4_X1 U9500 ( .A1(n8296), .A2(n8394), .A3(n8393), .A4(n8351), .ZN(n8312)
         );
  NAND2_X1 U9501 ( .A1(n8297), .A2(n8392), .ZN(n8298) );
  NAND4_X1 U9502 ( .A1(n8298), .A2(n8369), .A3(n8405), .A4(n8380), .ZN(n8311)
         );
  NAND2_X1 U9503 ( .A1(n8300), .A2(n8351), .ZN(n8303) );
  INV_X1 U9504 ( .A(n8303), .ZN(n8299) );
  AOI22_X1 U9505 ( .A1(n9917), .A2(n8299), .B1(n9520), .B2(n8351), .ZN(n8308)
         );
  OR2_X1 U9506 ( .A1(n8300), .A2(n8351), .ZN(n8302) );
  OAI22_X1 U9507 ( .A1(n9917), .A2(n8302), .B1(n9520), .B2(n8351), .ZN(n8301)
         );
  NAND2_X1 U9508 ( .A1(n10638), .A2(n8301), .ZN(n8307) );
  NOR2_X1 U9509 ( .A1(n8302), .A2(n9520), .ZN(n8305) );
  OAI21_X1 U9510 ( .B1(n9537), .B2(n8303), .A(n9917), .ZN(n8304) );
  OAI21_X1 U9511 ( .B1(n8305), .B2(n9917), .A(n8304), .ZN(n8306) );
  OAI211_X1 U9512 ( .C1(n10638), .C2(n8308), .A(n8307), .B(n8306), .ZN(n8309)
         );
  NOR2_X1 U9513 ( .A1(n8511), .A2(n8309), .ZN(n8310) );
  NAND3_X1 U9514 ( .A1(n8312), .A2(n8311), .A3(n8310), .ZN(n8314) );
  MUX2_X1 U9515 ( .A(n8397), .B(n8398), .S(n8351), .Z(n8313) );
  NAND3_X1 U9516 ( .A1(n8314), .A2(n8514), .A3(n8313), .ZN(n8317) );
  MUX2_X1 U9517 ( .A(n8806), .B(n8315), .S(n8369), .Z(n8316) );
  NAND2_X1 U9518 ( .A1(n9901), .A2(n9497), .ZN(n8377) );
  AOI21_X1 U9519 ( .B1(n8317), .B2(n8316), .A(n9812), .ZN(n8321) );
  OR2_X1 U9520 ( .A1(n9895), .A2(n9809), .ZN(n8432) );
  NAND2_X1 U9521 ( .A1(n9895), .A2(n9809), .ZN(n8809) );
  MUX2_X1 U9522 ( .A(n8377), .B(n8808), .S(n8369), .Z(n8318) );
  NAND2_X1 U9523 ( .A1(n9797), .A2(n8318), .ZN(n8320) );
  OR2_X1 U9524 ( .A1(n9892), .A2(n9754), .ZN(n8435) );
  NAND2_X1 U9525 ( .A1(n9892), .A2(n9754), .ZN(n8436) );
  MUX2_X1 U9526 ( .A(n8809), .B(n8432), .S(n8351), .Z(n8319) );
  OAI211_X1 U9527 ( .C1(n8321), .C2(n8320), .A(n9777), .B(n8319), .ZN(n8323)
         );
  MUX2_X1 U9528 ( .A(n8436), .B(n8435), .S(n8369), .Z(n8322) );
  AND2_X1 U9529 ( .A1(n8323), .A2(n8322), .ZN(n8329) );
  AND2_X1 U9530 ( .A1(n9881), .A2(n9755), .ZN(n8811) );
  INV_X1 U9531 ( .A(n8811), .ZN(n8326) );
  OR2_X1 U9532 ( .A1(n9881), .A2(n9755), .ZN(n8431) );
  NAND2_X1 U9533 ( .A1(n9885), .A2(n9780), .ZN(n8327) );
  INV_X1 U9534 ( .A(n8327), .ZN(n8324) );
  NAND2_X1 U9535 ( .A1(n8431), .A2(n8324), .ZN(n8325) );
  NAND2_X1 U9536 ( .A1(n8326), .A2(n8325), .ZN(n8374) );
  OR2_X1 U9537 ( .A1(n8374), .A2(n8351), .ZN(n8328) );
  NAND2_X1 U9538 ( .A1(n8431), .A2(n8326), .ZN(n9740) );
  MUX2_X1 U9539 ( .A(n8329), .B(n8328), .S(n8516), .Z(n8331) );
  OR2_X1 U9540 ( .A1(n9874), .A2(n9742), .ZN(n8813) );
  NAND2_X1 U9541 ( .A1(n9874), .A2(n9742), .ZN(n8375) );
  NAND2_X1 U9542 ( .A1(n8374), .A2(n8351), .ZN(n8330) );
  NAND3_X1 U9543 ( .A1(n8331), .A2(n9718), .A3(n8330), .ZN(n8333) );
  MUX2_X1 U9544 ( .A(n8375), .B(n8813), .S(n8351), .Z(n8332) );
  AND3_X1 U9545 ( .A1(n9707), .A2(n8333), .A3(n8332), .ZN(n8335) );
  MUX2_X1 U9546 ( .A(n8489), .B(n8815), .S(n8351), .Z(n8334) );
  OAI211_X1 U9547 ( .C1(n8336), .C2(n8335), .A(n9675), .B(n8334), .ZN(n8337)
         );
  NAND3_X1 U9548 ( .A1(n8339), .A2(n8338), .A3(n8337), .ZN(n8340) );
  NAND3_X1 U9549 ( .A1(n9638), .A2(n8341), .A3(n8340), .ZN(n8342) );
  NAND2_X1 U9550 ( .A1(n8549), .A2(n8355), .ZN(n8346) );
  OR2_X1 U9551 ( .A1(n4864), .A2(n8344), .ZN(n8345) );
  INV_X1 U9552 ( .A(n9621), .ZN(n8348) );
  NAND2_X1 U9553 ( .A1(n9837), .A2(n8348), .ZN(n8487) );
  NAND3_X1 U9554 ( .A1(n8347), .A2(n8487), .A3(n8450), .ZN(n8349) );
  NAND2_X1 U9555 ( .A1(n8488), .A2(n8819), .ZN(n8452) );
  OAI21_X1 U9556 ( .B1(n8350), .B2(n8452), .A(n8487), .ZN(n8352) );
  NAND2_X1 U9557 ( .A1(n8828), .A2(n8355), .ZN(n8357) );
  OR2_X1 U9558 ( .A1(n4864), .A2(n8829), .ZN(n8356) );
  INV_X1 U9559 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9614) );
  INV_X1 U9560 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8358) );
  OR2_X1 U9561 ( .A1(n6787), .A2(n8358), .ZN(n8360) );
  NAND2_X1 U9562 ( .A1(n4862), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8359) );
  OAI211_X1 U9563 ( .C1(n7853), .C2(n9614), .A(n8360), .B(n8359), .ZN(n9532)
         );
  INV_X1 U9564 ( .A(n9532), .ZN(n8363) );
  NAND2_X1 U9565 ( .A1(n9832), .A2(n8363), .ZN(n8485) );
  INV_X1 U9566 ( .A(n9608), .ZN(n8367) );
  NAND2_X1 U9567 ( .A1(n9832), .A2(n8367), .ZN(n8361) );
  AND2_X1 U9568 ( .A1(n8485), .A2(n8361), .ZN(n8476) );
  OR2_X1 U9569 ( .A1(n9832), .A2(n8363), .ZN(n8486) );
  NOR2_X1 U9570 ( .A1(n9831), .A2(n8486), .ZN(n8364) );
  OAI22_X1 U9571 ( .A1(n8365), .A2(n8364), .B1(n8369), .B2(n8476), .ZN(n8370)
         );
  INV_X1 U9572 ( .A(n9831), .ZN(n8366) );
  NAND2_X1 U9573 ( .A1(n8366), .A2(n8367), .ZN(n8522) );
  OR2_X1 U9574 ( .A1(n8486), .A2(n8367), .ZN(n8368) );
  NAND2_X1 U9575 ( .A1(n8522), .A2(n8368), .ZN(n8480) );
  INV_X1 U9576 ( .A(n8541), .ZN(n8545) );
  INV_X1 U9577 ( .A(n8542), .ZN(n8533) );
  NAND2_X1 U9578 ( .A1(n8533), .A2(n8531), .ZN(n8461) );
  NAND3_X1 U9579 ( .A1(n8533), .A2(n10415), .A3(n6648), .ZN(n8460) );
  INV_X1 U9580 ( .A(n8816), .ZN(n8373) );
  INV_X1 U9581 ( .A(n8371), .ZN(n8372) );
  OR3_X1 U9582 ( .A1(n8452), .A2(n8373), .A3(n8372), .ZN(n8478) );
  INV_X1 U9583 ( .A(n8374), .ZN(n8376) );
  NAND2_X1 U9584 ( .A1(n8376), .A2(n8375), .ZN(n8440) );
  INV_X1 U9585 ( .A(n8436), .ZN(n8810) );
  AND2_X1 U9586 ( .A1(n8377), .A2(n8806), .ZN(n8378) );
  NAND2_X1 U9587 ( .A1(n8809), .A2(n8378), .ZN(n8409) );
  NAND2_X1 U9588 ( .A1(n8380), .A2(n8379), .ZN(n8407) );
  NAND2_X1 U9589 ( .A1(n8382), .A2(n8381), .ZN(n8383) );
  NAND2_X1 U9590 ( .A1(n8383), .A2(n8388), .ZN(n8384) );
  AND2_X1 U9591 ( .A1(n8385), .A2(n8384), .ZN(n8404) );
  NAND3_X1 U9592 ( .A1(n8388), .A2(n8387), .A3(n8386), .ZN(n8390) );
  AOI21_X1 U9593 ( .B1(n8404), .B2(n8390), .A(n5207), .ZN(n8391) );
  AND2_X1 U9594 ( .A1(n8392), .A2(n8391), .ZN(n8395) );
  OAI211_X1 U9595 ( .C1(n8407), .C2(n8395), .A(n8394), .B(n8393), .ZN(n8396)
         );
  NAND3_X1 U9596 ( .A1(n8397), .A2(n8405), .A3(n8396), .ZN(n8399) );
  NAND2_X1 U9597 ( .A1(n8399), .A2(n8398), .ZN(n8400) );
  NOR2_X1 U9598 ( .A1(n8805), .A2(n8400), .ZN(n8401) );
  OR2_X1 U9599 ( .A1(n8409), .A2(n8401), .ZN(n8467) );
  NAND4_X1 U9600 ( .A1(n8405), .A2(n8404), .A3(n8403), .A4(n8402), .ZN(n8406)
         );
  OR4_X1 U9601 ( .A1(n8409), .A2(n8408), .A3(n8407), .A4(n8406), .ZN(n8410) );
  AND2_X1 U9602 ( .A1(n8467), .A2(n8410), .ZN(n8411) );
  OR3_X1 U9603 ( .A1(n8440), .A2(n8810), .A3(n8411), .ZN(n8471) );
  INV_X1 U9604 ( .A(n8412), .ZN(n8414) );
  NAND2_X1 U9605 ( .A1(n9544), .A2(n5013), .ZN(n8413) );
  NAND3_X1 U9606 ( .A1(n8414), .A2(n8483), .A3(n8413), .ZN(n8416) );
  NAND2_X1 U9607 ( .A1(n8416), .A2(n8415), .ZN(n8418) );
  OAI21_X1 U9608 ( .B1(n8419), .B2(n8418), .A(n8417), .ZN(n8421) );
  NAND2_X1 U9609 ( .A1(n8421), .A2(n8420), .ZN(n8424) );
  NAND3_X1 U9610 ( .A1(n8424), .A2(n8423), .A3(n8422), .ZN(n8425) );
  NAND3_X1 U9611 ( .A1(n8425), .A2(n8464), .A3(n4892), .ZN(n8426) );
  NAND4_X1 U9612 ( .A1(n8467), .A2(n8428), .A3(n8427), .A4(n8426), .ZN(n8429)
         );
  NAND2_X1 U9613 ( .A1(n8469), .A2(n8429), .ZN(n8430) );
  NOR2_X1 U9614 ( .A1(n8471), .A2(n8430), .ZN(n8445) );
  AND2_X1 U9615 ( .A1(n8431), .A2(n9738), .ZN(n8812) );
  NAND2_X1 U9616 ( .A1(n8432), .A2(n8808), .ZN(n8433) );
  NAND2_X1 U9617 ( .A1(n8433), .A2(n8809), .ZN(n8434) );
  NAND2_X1 U9618 ( .A1(n8435), .A2(n8434), .ZN(n8437) );
  NAND2_X1 U9619 ( .A1(n8437), .A2(n8436), .ZN(n8438) );
  AND2_X1 U9620 ( .A1(n8812), .A2(n8438), .ZN(n8439) );
  OAI21_X1 U9621 ( .B1(n8440), .B2(n8439), .A(n8813), .ZN(n8441) );
  AND2_X1 U9622 ( .A1(n8441), .A2(n8469), .ZN(n8442) );
  OR2_X1 U9623 ( .A1(n8443), .A2(n8442), .ZN(n8473) );
  AND2_X1 U9624 ( .A1(n8444), .A2(n8489), .ZN(n8472) );
  OAI21_X1 U9625 ( .B1(n8445), .B2(n8473), .A(n8472), .ZN(n8446) );
  NAND2_X1 U9626 ( .A1(n9638), .A2(n8446), .ZN(n8454) );
  INV_X1 U9627 ( .A(n8447), .ZN(n8817) );
  NAND2_X1 U9628 ( .A1(n8818), .A2(n8817), .ZN(n8448) );
  AND3_X1 U9629 ( .A1(n8450), .A2(n8449), .A3(n8448), .ZN(n8451) );
  OR2_X1 U9630 ( .A1(n8452), .A2(n8451), .ZN(n8453) );
  AND2_X1 U9631 ( .A1(n8453), .A2(n8487), .ZN(n8477) );
  OAI211_X1 U9632 ( .C1(n8478), .C2(n8454), .A(n8477), .B(n8485), .ZN(n8455)
         );
  NAND2_X1 U9633 ( .A1(n8455), .A2(n8486), .ZN(n8457) );
  INV_X1 U9634 ( .A(n8456), .ZN(n8524) );
  NAND2_X1 U9635 ( .A1(n8457), .A2(n8524), .ZN(n8458) );
  NAND2_X1 U9636 ( .A1(n8458), .A2(n8522), .ZN(n8459) );
  MUX2_X1 U9637 ( .A(n8461), .B(n8460), .S(n8459), .Z(n8538) );
  INV_X1 U9638 ( .A(n8462), .ZN(n8463) );
  AOI21_X1 U9639 ( .B1(n8465), .B2(n8464), .A(n8463), .ZN(n8466) );
  NAND2_X1 U9640 ( .A1(n8467), .A2(n8466), .ZN(n8468) );
  NAND2_X1 U9641 ( .A1(n8469), .A2(n8468), .ZN(n8470) );
  NOR2_X1 U9642 ( .A1(n8471), .A2(n8470), .ZN(n8474) );
  OAI21_X1 U9643 ( .B1(n8474), .B2(n8473), .A(n8472), .ZN(n8475) );
  NAND2_X1 U9644 ( .A1(n8818), .A2(n8475), .ZN(n8479) );
  OAI211_X1 U9645 ( .C1(n8479), .C2(n8478), .A(n8477), .B(n8476), .ZN(n8482)
         );
  INV_X1 U9646 ( .A(n8480), .ZN(n8481) );
  NAND2_X1 U9647 ( .A1(n8482), .A2(n8481), .ZN(n8484) );
  NAND3_X1 U9648 ( .A1(n8484), .A2(n8483), .A3(n8524), .ZN(n8529) );
  NOR2_X1 U9649 ( .A1(n6648), .A2(n10415), .ZN(n8528) );
  AND2_X1 U9650 ( .A1(n8486), .A2(n8485), .ZN(n8523) );
  NAND2_X1 U9651 ( .A1(n8488), .A2(n8487), .ZN(n8820) );
  INV_X1 U9652 ( .A(n9624), .ZN(n8520) );
  INV_X1 U9653 ( .A(n9638), .ZN(n9646) );
  INV_X1 U9654 ( .A(n9675), .ZN(n8795) );
  NAND4_X1 U9655 ( .A1(n8493), .A2(n8492), .A3(n8491), .A4(n8490), .ZN(n8497)
         );
  INV_X1 U9656 ( .A(n8494), .ZN(n8495) );
  NOR3_X1 U9657 ( .A1(n8497), .A2(n8496), .A3(n8495), .ZN(n8501) );
  NAND4_X1 U9658 ( .A1(n8501), .A2(n8500), .A3(n8499), .A4(n8498), .ZN(n8503)
         );
  NOR2_X1 U9659 ( .A1(n8503), .A2(n8502), .ZN(n8504) );
  NAND4_X1 U9660 ( .A1(n8507), .A2(n8506), .A3(n8505), .A4(n8504), .ZN(n8508)
         );
  OR4_X1 U9661 ( .A1(n8511), .A2(n8510), .A3(n8509), .A4(n8508), .ZN(n8512) );
  NOR2_X1 U9662 ( .A1(n9812), .A2(n8512), .ZN(n8513) );
  NAND4_X1 U9663 ( .A1(n9777), .A2(n9797), .A3(n8514), .A4(n8513), .ZN(n8515)
         );
  NOR2_X1 U9664 ( .A1(n8516), .A2(n8515), .ZN(n8517) );
  NAND4_X1 U9665 ( .A1(n9686), .A2(n9718), .A3(n9707), .A4(n8517), .ZN(n8518)
         );
  OR3_X1 U9666 ( .A1(n9657), .A2(n8795), .A3(n8518), .ZN(n8519) );
  NOR4_X1 U9667 ( .A1(n8820), .A2(n8520), .A3(n9646), .A4(n8519), .ZN(n8521)
         );
  NAND4_X1 U9668 ( .A1(n8524), .A2(n8523), .A3(n8522), .A4(n8521), .ZN(n8526)
         );
  AND2_X1 U9669 ( .A1(n8526), .A2(n8525), .ZN(n8539) );
  INV_X1 U9670 ( .A(n8539), .ZN(n8527) );
  NAND4_X1 U9671 ( .A1(n8529), .A2(n8533), .A3(n8528), .A4(n8527), .ZN(n8537)
         );
  NAND4_X1 U9672 ( .A1(n10393), .A2(n10338), .A3(n8531), .A4(n8530), .ZN(n8535) );
  AOI21_X1 U9673 ( .B1(n8533), .B2(n8532), .A(n8822), .ZN(n8534) );
  NAND2_X1 U9674 ( .A1(n8535), .A2(n8534), .ZN(n8536) );
  NAND3_X1 U9675 ( .A1(n8538), .A2(n8537), .A3(n8536), .ZN(n8544) );
  AOI21_X1 U9676 ( .B1(n8541), .B2(n8540), .A(n8539), .ZN(n8543) );
  NAND2_X1 U9677 ( .A1(n8828), .A2(n8580), .ZN(n8548) );
  NAND2_X1 U9678 ( .A1(n8581), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8547) );
  NAND2_X1 U9679 ( .A1(n8549), .A2(n8580), .ZN(n8551) );
  NAND2_X1 U9680 ( .A1(n8581), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8550) );
  XNOR2_X1 U9681 ( .A(n9036), .B(n8922), .ZN(n9033) );
  INV_X1 U9682 ( .A(n9033), .ZN(n8718) );
  NAND2_X1 U9683 ( .A1(n8553), .A2(n8658), .ZN(n9208) );
  NAND2_X1 U9684 ( .A1(n9337), .A2(n8554), .ZN(n8661) );
  NAND2_X1 U9685 ( .A1(n8662), .A2(n8661), .ZN(n9211) );
  INV_X1 U9686 ( .A(n9211), .ZN(n8756) );
  XNOR2_X1 U9687 ( .A(n9331), .B(n9215), .ZN(n9192) );
  INV_X1 U9688 ( .A(n9192), .ZN(n9203) );
  NAND2_X1 U9689 ( .A1(n9327), .A2(n8924), .ZN(n8666) );
  NAND2_X1 U9690 ( .A1(n8668), .A2(n8666), .ZN(n9178) );
  INV_X1 U9691 ( .A(n9178), .ZN(n8555) );
  NAND2_X1 U9692 ( .A1(n9173), .A2(n8555), .ZN(n8556) );
  NAND2_X1 U9693 ( .A1(n8556), .A2(n8668), .ZN(n9160) );
  NAND2_X1 U9694 ( .A1(n9321), .A2(n8858), .ZN(n8676) );
  NAND2_X1 U9695 ( .A1(n8675), .A2(n8676), .ZN(n9168) );
  INV_X1 U9696 ( .A(n9168), .ZN(n8557) );
  OR2_X1 U9697 ( .A1(n9316), .A2(n8558), .ZN(n8559) );
  NAND2_X1 U9698 ( .A1(n9316), .A2(n8558), .ZN(n8677) );
  NAND2_X1 U9699 ( .A1(n9311), .A2(n8859), .ZN(n8687) );
  NAND2_X1 U9700 ( .A1(n8683), .A2(n8687), .ZN(n9137) );
  INV_X1 U9701 ( .A(n9137), .ZN(n9130) );
  NAND2_X1 U9702 ( .A1(n9138), .A2(n9130), .ZN(n8560) );
  NAND2_X1 U9703 ( .A1(n8560), .A2(n8683), .ZN(n9115) );
  NAND2_X1 U9704 ( .A1(n9305), .A2(n8894), .ZN(n9101) );
  INV_X1 U9705 ( .A(n9121), .ZN(n8561) );
  NAND2_X1 U9706 ( .A1(n9298), .A2(n8562), .ZN(n8692) );
  NAND2_X1 U9707 ( .A1(n9294), .A2(n8914), .ZN(n8703) );
  NAND2_X1 U9708 ( .A1(n8707), .A2(n8703), .ZN(n9094) );
  INV_X1 U9709 ( .A(n8736), .ZN(n8564) );
  NAND2_X1 U9710 ( .A1(n9289), .A2(n8867), .ZN(n8735) );
  XNOR2_X1 U9711 ( .A(n9283), .B(n8711), .ZN(n9027) );
  OR2_X1 U9712 ( .A1(n9283), .A2(n8711), .ZN(n8705) );
  NAND2_X1 U9713 ( .A1(n9278), .A2(n8923), .ZN(n8716) );
  OR2_X1 U9714 ( .A1(n9036), .A2(n8922), .ZN(n8720) );
  INV_X1 U9715 ( .A(n8720), .ZN(n8566) );
  AOI21_X1 U9716 ( .B1(n8718), .B2(n9009), .A(n8566), .ZN(n8578) );
  INV_X1 U9717 ( .A(n8578), .ZN(n8579) );
  INV_X1 U9718 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8570) );
  NAND2_X1 U9719 ( .A1(n8567), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U9720 ( .A1(n5738), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8568) );
  OAI211_X1 U9721 ( .C1(n8572), .C2(n8570), .A(n8569), .B(n8568), .ZN(n9011)
         );
  INV_X1 U9722 ( .A(n9011), .ZN(n8584) );
  NAND2_X1 U9723 ( .A1(n5738), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8577) );
  INV_X1 U9724 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8571) );
  OR2_X1 U9725 ( .A1(n8572), .A2(n8571), .ZN(n8576) );
  INV_X1 U9726 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8573) );
  OR2_X1 U9727 ( .A1(n8574), .A2(n8573), .ZN(n8575) );
  NAND2_X1 U9728 ( .A1(n9955), .A2(n8580), .ZN(n8583) );
  NAND2_X1 U9729 ( .A1(n8581), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8582) );
  NAND2_X1 U9730 ( .A1(n9005), .A2(n8584), .ZN(n8723) );
  INV_X1 U9731 ( .A(n8761), .ZN(n8585) );
  XNOR2_X1 U9732 ( .A(n4890), .B(n5582), .ZN(n8771) );
  INV_X1 U9733 ( .A(n8586), .ZN(n8770) );
  MUX2_X1 U9734 ( .A(n8929), .B(n10492), .S(n8727), .Z(n8615) );
  INV_X1 U9735 ( .A(n8615), .ZN(n8617) );
  NOR2_X1 U9736 ( .A1(n10377), .A2(n8588), .ZN(n8739) );
  INV_X1 U9737 ( .A(n8741), .ZN(n8589) );
  OAI21_X1 U9738 ( .B1(n8739), .B2(n8727), .A(n8589), .ZN(n8596) );
  AOI21_X1 U9739 ( .B1(n8592), .B2(n8591), .A(n8590), .ZN(n8594) );
  NOR3_X1 U9740 ( .A1(n8594), .A2(n4860), .A3(n8593), .ZN(n8595) );
  AOI21_X1 U9741 ( .B1(n8597), .B2(n8596), .A(n8595), .ZN(n8606) );
  MUX2_X1 U9742 ( .A(n8599), .B(n8598), .S(n4860), .Z(n8601) );
  NAND2_X1 U9743 ( .A1(n8601), .A2(n8600), .ZN(n8605) );
  MUX2_X1 U9744 ( .A(n8603), .B(n8602), .S(n8727), .Z(n8604) );
  OAI211_X1 U9745 ( .C1(n8606), .C2(n8605), .A(n8743), .B(n8604), .ZN(n8608)
         );
  OAI211_X1 U9746 ( .C1(n4860), .C2(n8609), .A(n8608), .B(n8607), .ZN(n8612)
         );
  OAI21_X1 U9747 ( .B1(n10460), .B2(n8930), .A(n8611), .ZN(n8610) );
  AOI22_X1 U9748 ( .A1(n8612), .A2(n8611), .B1(n4860), .B2(n8610), .ZN(n8613)
         );
  INV_X1 U9749 ( .A(n8618), .ZN(n8619) );
  MUX2_X1 U9750 ( .A(n8619), .B(n5266), .S(n8727), .Z(n8620) );
  INV_X1 U9751 ( .A(n8623), .ZN(n8622) );
  OAI22_X1 U9752 ( .A1(n8622), .A2(n8621), .B1(n10516), .B2(n8626), .ZN(n8628)
         );
  OAI211_X1 U9753 ( .C1(n5286), .C2(n8626), .A(n8625), .B(n8631), .ZN(n8627)
         );
  MUX2_X1 U9754 ( .A(n8628), .B(n8627), .S(n4860), .Z(n8630) );
  NAND2_X1 U9755 ( .A1(n8633), .A2(n8632), .ZN(n8634) );
  INV_X1 U9756 ( .A(n8640), .ZN(n8635) );
  AOI21_X1 U9757 ( .B1(n8637), .B2(n8636), .A(n8635), .ZN(n8642) );
  INV_X1 U9758 ( .A(n8637), .ZN(n8638) );
  AOI21_X1 U9759 ( .B1(n8640), .B2(n8639), .A(n8638), .ZN(n8641) );
  MUX2_X1 U9760 ( .A(n8642), .B(n8641), .S(n8727), .Z(n8647) );
  MUX2_X1 U9761 ( .A(n8644), .B(n8643), .S(n4860), .Z(n8645) );
  OAI211_X1 U9762 ( .C1(n8648), .C2(n8647), .A(n8646), .B(n8645), .ZN(n8652)
         );
  INV_X1 U9763 ( .A(n9228), .ZN(n9242) );
  MUX2_X1 U9764 ( .A(n8650), .B(n8649), .S(n8727), .Z(n8651) );
  NAND3_X1 U9765 ( .A1(n8652), .A2(n9242), .A3(n8651), .ZN(n8656) );
  MUX2_X1 U9766 ( .A(n8654), .B(n8653), .S(n4860), .Z(n8655) );
  NAND3_X1 U9767 ( .A1(n8656), .A2(n8757), .A3(n8655), .ZN(n8660) );
  MUX2_X1 U9768 ( .A(n8658), .B(n8657), .S(n8727), .Z(n8659) );
  NAND3_X1 U9769 ( .A1(n8660), .A2(n8756), .A3(n8659), .ZN(n8664) );
  MUX2_X1 U9770 ( .A(n8662), .B(n8661), .S(n4860), .Z(n8663) );
  NAND2_X1 U9771 ( .A1(n8664), .A2(n8663), .ZN(n8673) );
  MUX2_X1 U9772 ( .A(n9331), .B(n9174), .S(n8727), .Z(n8672) );
  NAND2_X1 U9773 ( .A1(n8673), .A2(n8672), .ZN(n8667) );
  NAND3_X1 U9774 ( .A1(n8667), .A2(n9331), .A3(n8668), .ZN(n8665) );
  NAND3_X1 U9775 ( .A1(n8665), .A2(n8676), .A3(n8666), .ZN(n8671) );
  NAND3_X1 U9776 ( .A1(n8667), .A2(n9174), .A3(n8666), .ZN(n8669) );
  NAND3_X1 U9777 ( .A1(n8669), .A2(n8675), .A3(n8668), .ZN(n8670) );
  OR2_X1 U9778 ( .A1(n9316), .A2(n9161), .ZN(n9019) );
  OAI21_X1 U9779 ( .B1(n4860), .B2(n9161), .A(n9316), .ZN(n8674) );
  AND2_X1 U9780 ( .A1(n9019), .A2(n8674), .ZN(n8680) );
  INV_X1 U9781 ( .A(n9101), .ZN(n8691) );
  INV_X1 U9782 ( .A(n8675), .ZN(n8679) );
  NAND2_X1 U9783 ( .A1(n8677), .A2(n8676), .ZN(n8678) );
  MUX2_X1 U9784 ( .A(n8679), .B(n8678), .S(n4860), .Z(n8682) );
  INV_X1 U9785 ( .A(n8680), .ZN(n8681) );
  AND4_X1 U9786 ( .A1(n8683), .A2(n8687), .A3(n8682), .A4(n8681), .ZN(n8690)
         );
  INV_X1 U9787 ( .A(n9311), .ZN(n9136) );
  NAND2_X1 U9788 ( .A1(n9161), .A2(n8727), .ZN(n8684) );
  OAI22_X1 U9789 ( .A1(n9316), .A2(n8684), .B1(n8859), .B2(n4860), .ZN(n8686)
         );
  NOR3_X1 U9790 ( .A1(n9316), .A2(n8859), .A3(n8684), .ZN(n8685) );
  AOI21_X1 U9791 ( .B1(n9136), .B2(n8686), .A(n8685), .ZN(n8688) );
  NAND3_X1 U9792 ( .A1(n8688), .A2(n8693), .A3(n5459), .ZN(n8689) );
  NAND2_X1 U9793 ( .A1(n8692), .A2(n9101), .ZN(n8695) );
  NAND2_X1 U9794 ( .A1(n8697), .A2(n8693), .ZN(n8694) );
  MUX2_X1 U9795 ( .A(n8695), .B(n8694), .S(n4860), .Z(n8696) );
  OAI21_X1 U9796 ( .B1(n8727), .B2(n9118), .A(n8697), .ZN(n8701) );
  INV_X1 U9797 ( .A(n8703), .ZN(n8699) );
  OAI21_X1 U9798 ( .B1(n8702), .B2(n9298), .A(n5332), .ZN(n8698) );
  OAI21_X1 U9799 ( .B1(n4860), .B2(n8699), .A(n8698), .ZN(n8700) );
  OAI21_X1 U9800 ( .B1(n8702), .B2(n8701), .A(n8700), .ZN(n8710) );
  OAI21_X1 U9801 ( .B1(n8706), .B2(n9027), .A(n8705), .ZN(n8714) );
  AOI21_X1 U9802 ( .B1(n8710), .B2(n8709), .A(n8708), .ZN(n8712) );
  INV_X1 U9803 ( .A(n9283), .ZN(n9067) );
  OAI22_X1 U9804 ( .A1(n8712), .A2(n9027), .B1(n9067), .B2(n9081), .ZN(n8713)
         );
  MUX2_X1 U9805 ( .A(n8716), .B(n8715), .S(n8727), .Z(n8717) );
  NAND2_X1 U9806 ( .A1(n9036), .A2(n8922), .ZN(n8721) );
  MUX2_X1 U9807 ( .A(n8721), .B(n8720), .S(n4860), .Z(n8722) );
  INV_X1 U9808 ( .A(n8760), .ZN(n8724) );
  NOR2_X1 U9809 ( .A1(n8761), .A2(n8724), .ZN(n8725) );
  MUX2_X1 U9810 ( .A(n8726), .B(n8725), .S(n8727), .Z(n8731) );
  INV_X1 U9811 ( .A(n8729), .ZN(n9001) );
  MUX2_X1 U9812 ( .A(n9001), .B(n8998), .S(n8727), .Z(n8728) );
  AOI21_X1 U9813 ( .B1(n8729), .B2(n9268), .A(n8728), .ZN(n8730) );
  XNOR2_X1 U9814 ( .A(n8766), .B(n8732), .ZN(n8734) );
  NAND2_X1 U9815 ( .A1(n8736), .A2(n8735), .ZN(n9079) );
  INV_X1 U9816 ( .A(n9156), .ZN(n9145) );
  INV_X1 U9817 ( .A(n8739), .ZN(n8742) );
  NOR4_X1 U9818 ( .A1(n8742), .A2(n6098), .A3(n8741), .A4(n8740), .ZN(n8745)
         );
  NAND4_X1 U9819 ( .A1(n9261), .A2(n8745), .A3(n8744), .A4(n8743), .ZN(n8746)
         );
  NOR4_X1 U9820 ( .A1(n8748), .A2(n7259), .A3(n8747), .A4(n8746), .ZN(n8749)
         );
  NAND4_X1 U9821 ( .A1(n8752), .A2(n8751), .A3(n8750), .A4(n8749), .ZN(n8753)
         );
  NOR4_X1 U9822 ( .A1(n8754), .A2(n5300), .A3(n9228), .A4(n8753), .ZN(n8755)
         );
  NAND4_X1 U9823 ( .A1(n9203), .A2(n8757), .A3(n8756), .A4(n8755), .ZN(n8758)
         );
  NOR4_X1 U9824 ( .A1(n9145), .A2(n9178), .A3(n9168), .A4(n8758), .ZN(n8759)
         );
  XNOR2_X1 U9825 ( .A(n8762), .B(n5582), .ZN(n8764) );
  OAI211_X1 U9826 ( .C1(n8766), .C2(n8765), .A(n8764), .B(n8763), .ZN(n8767)
         );
  NAND4_X1 U9827 ( .A1(n8772), .A2(n9971), .A3(n8999), .A4(n9230), .ZN(n8773)
         );
  OAI211_X1 U9828 ( .C1(n8774), .C2(n8776), .A(n8773), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8775) );
  OAI21_X1 U9829 ( .B1(n8777), .B2(n8776), .A(n8775), .ZN(P2_U3244) );
  OAI222_X1 U9830 ( .A1(n9961), .A2(n8780), .B1(P1_U3084), .B2(n8779), .C1(
        n8778), .C2(n8830), .ZN(P1_U3329) );
  OR2_X1 U9831 ( .A1(n9901), .A2(n9799), .ZN(n8783) );
  NAND2_X1 U9832 ( .A1(n9789), .A2(n9788), .ZN(n9787) );
  NAND2_X1 U9833 ( .A1(n9895), .A2(n9535), .ZN(n8784) );
  NAND2_X1 U9834 ( .A1(n9787), .A2(n8784), .ZN(n9771) );
  OR2_X1 U9835 ( .A1(n9892), .A2(n9798), .ZN(n8785) );
  NAND2_X1 U9836 ( .A1(n9771), .A2(n8785), .ZN(n9734) );
  NAND2_X1 U9837 ( .A1(n9892), .A2(n9798), .ZN(n9733) );
  INV_X1 U9838 ( .A(n9780), .ZN(n9534) );
  NAND2_X1 U9839 ( .A1(n9885), .A2(n9534), .ZN(n9735) );
  NAND2_X1 U9840 ( .A1(n9881), .A2(n9720), .ZN(n8789) );
  AND2_X1 U9841 ( .A1(n9735), .A2(n8789), .ZN(n8786) );
  AND2_X1 U9842 ( .A1(n9733), .A2(n8786), .ZN(n8788) );
  INV_X1 U9843 ( .A(n8786), .ZN(n8787) );
  INV_X1 U9844 ( .A(n8789), .ZN(n8790) );
  OR2_X1 U9845 ( .A1(n8790), .A2(n9740), .ZN(n8791) );
  AND2_X1 U9846 ( .A1(n9874), .A2(n9709), .ZN(n8792) );
  OR2_X1 U9847 ( .A1(n9874), .A2(n9709), .ZN(n8793) );
  NOR2_X1 U9848 ( .A1(n9869), .A2(n9721), .ZN(n8794) );
  OR2_X1 U9849 ( .A1(n9859), .A2(n9533), .ZN(n8796) );
  NOR2_X1 U9850 ( .A1(n9854), .A2(n9677), .ZN(n8797) );
  NAND2_X1 U9851 ( .A1(n9854), .A2(n9677), .ZN(n8798) );
  OAI22_X1 U9852 ( .A1(n9639), .A2(n9638), .B1(n9622), .B2(n9848), .ZN(n9618)
         );
  INV_X1 U9853 ( .A(n9848), .ZN(n9645) );
  AND2_X2 U9854 ( .A1(n9665), .A2(n9669), .ZN(n9660) );
  AOI21_X1 U9855 ( .B1(n9837), .B2(n9632), .A(n9612), .ZN(n9838) );
  INV_X1 U9856 ( .A(n9837), .ZN(n8804) );
  INV_X1 U9857 ( .A(n8801), .ZN(n8802) );
  AOI22_X1 U9858 ( .A1(n8802), .A2(n10411), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9684), .ZN(n8803) );
  OAI21_X1 U9859 ( .B1(n8804), .B2(n9818), .A(n8803), .ZN(n8825) );
  NAND2_X1 U9860 ( .A1(n9717), .A2(n8813), .ZN(n9708) );
  NAND2_X1 U9861 ( .A1(n9685), .A2(n8815), .ZN(n9676) );
  NAND2_X1 U9862 ( .A1(n9623), .A2(n8819), .ZN(n8821) );
  XNOR2_X1 U9863 ( .A(n8821), .B(n8820), .ZN(n8824) );
  OR2_X1 U9864 ( .A1(n6387), .A2(n8822), .ZN(n8823) );
  AND2_X1 U9865 ( .A1(n10392), .A2(n8823), .ZN(n9607) );
  INV_X1 U9866 ( .A(n8826), .ZN(n9381) );
  OAI222_X1 U9867 ( .A1(n9961), .A2(n8827), .B1(n8830), .B2(n9381), .C1(
        P1_U3084), .C2(n6386), .ZN(P1_U3325) );
  INV_X1 U9868 ( .A(n8828), .ZN(n9376) );
  XNOR2_X1 U9869 ( .A(n8833), .B(n8832), .ZN(n8838) );
  NOR2_X1 U9870 ( .A1(n8867), .A2(n10514), .ZN(n8835) );
  OAI22_X1 U9871 ( .A1(n8923), .A2(n10517), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9986), .ZN(n8834) );
  AOI211_X1 U9872 ( .C1(n8886), .C2(n9064), .A(n8835), .B(n8834), .ZN(n8837)
         );
  NAND2_X1 U9873 ( .A1(n9283), .A2(n8918), .ZN(n8836) );
  OAI211_X1 U9874 ( .C1(n8838), .C2(n10510), .A(n8837), .B(n8836), .ZN(
        P2_U3216) );
  INV_X1 U9875 ( .A(n9305), .ZN(n8847) );
  NAND2_X1 U9876 ( .A1(n8875), .A2(n9139), .ZN(n8842) );
  OR2_X1 U9877 ( .A1(n10510), .A2(n8839), .ZN(n8841) );
  MUX2_X1 U9878 ( .A(n8842), .B(n8841), .S(n8840), .Z(n8846) );
  NOR2_X1 U9879 ( .A1(n10523), .A2(n9126), .ZN(n8844) );
  OAI22_X1 U9880 ( .A1(n10514), .A2(n8859), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10166), .ZN(n8843) );
  AOI211_X1 U9881 ( .C1(n8917), .C2(n9118), .A(n8844), .B(n8843), .ZN(n8845)
         );
  OAI211_X1 U9882 ( .C1(n8847), .C2(n8883), .A(n8846), .B(n8845), .ZN(P2_U3218) );
  NAND2_X1 U9883 ( .A1(n4938), .A2(n8848), .ZN(n8849) );
  XNOR2_X1 U9884 ( .A(n8850), .B(n8849), .ZN(n8855) );
  NAND2_X1 U9885 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8990) );
  OAI21_X1 U9886 ( .B1(n10517), .B2(n8858), .A(n8990), .ZN(n8851) );
  AOI21_X1 U9887 ( .B1(n8906), .B2(n9174), .A(n8851), .ZN(n8852) );
  OAI21_X1 U9888 ( .B1(n9180), .B2(n10523), .A(n8852), .ZN(n8853) );
  AOI21_X1 U9889 ( .B1(n9327), .B2(n8918), .A(n8853), .ZN(n8854) );
  OAI21_X1 U9890 ( .B1(n8855), .B2(n10510), .A(n8854), .ZN(P2_U3221) );
  XNOR2_X1 U9891 ( .A(n8857), .B(n8856), .ZN(n8864) );
  OAI22_X1 U9892 ( .A1(n10517), .A2(n8859), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10172), .ZN(n8860) );
  AOI21_X1 U9893 ( .B1(n8906), .B2(n9175), .A(n8860), .ZN(n8861) );
  OAI21_X1 U9894 ( .B1(n9150), .B2(n10523), .A(n8861), .ZN(n8862) );
  AOI21_X1 U9895 ( .B1(n9316), .B2(n8918), .A(n8862), .ZN(n8863) );
  OAI21_X1 U9896 ( .B1(n8864), .B2(n10510), .A(n8863), .ZN(P2_U3225) );
  XNOR2_X1 U9897 ( .A(n8865), .B(n8866), .ZN(n8872) );
  OAI22_X1 U9898 ( .A1(n8867), .A2(n10517), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10083), .ZN(n8868) );
  AOI21_X1 U9899 ( .B1(n8906), .B2(n9118), .A(n8868), .ZN(n8869) );
  OAI21_X1 U9900 ( .B1(n9090), .B2(n10523), .A(n8869), .ZN(n8870) );
  AOI21_X1 U9901 ( .B1(n9294), .B2(n8918), .A(n8870), .ZN(n8871) );
  OAI21_X1 U9902 ( .B1(n8872), .B2(n10510), .A(n8871), .ZN(P2_U3227) );
  INV_X1 U9903 ( .A(n9298), .ZN(n9107) );
  NAND2_X1 U9904 ( .A1(n8874), .A2(n8873), .ZN(n8878) );
  NAND2_X1 U9905 ( .A1(n9118), .A2(n8875), .ZN(n8877) );
  MUX2_X1 U9906 ( .A(n8878), .B(n8877), .S(n8876), .Z(n8882) );
  OAI22_X1 U9907 ( .A1(n10514), .A2(n8894), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10081), .ZN(n8880) );
  NOR2_X1 U9908 ( .A1(n8914), .A2(n10517), .ZN(n8879) );
  AOI211_X1 U9909 ( .C1(n8886), .C2(n9105), .A(n8880), .B(n8879), .ZN(n8881)
         );
  OAI211_X1 U9910 ( .C1(n9107), .C2(n8883), .A(n8882), .B(n8881), .ZN(P2_U3231) );
  XNOR2_X1 U9911 ( .A(n8885), .B(n8884), .ZN(n8891) );
  AOI22_X1 U9912 ( .A1(n8917), .A2(n9161), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8888) );
  NAND2_X1 U9913 ( .A1(n8886), .A2(n9164), .ZN(n8887) );
  OAI211_X1 U9914 ( .C1(n8924), .C2(n10514), .A(n8888), .B(n8887), .ZN(n8889)
         );
  AOI21_X1 U9915 ( .B1(n9321), .B2(n8918), .A(n8889), .ZN(n8890) );
  OAI21_X1 U9916 ( .B1(n8891), .B2(n10510), .A(n8890), .ZN(P2_U3235) );
  AOI21_X1 U9917 ( .B1(n8893), .B2(n8892), .A(n4901), .ZN(n8899) );
  OAI22_X1 U9918 ( .A1(n10517), .A2(n8894), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10192), .ZN(n8895) );
  AOI21_X1 U9919 ( .B1(n8906), .B2(n9161), .A(n8895), .ZN(n8896) );
  OAI21_X1 U9920 ( .B1(n9133), .B2(n10523), .A(n8896), .ZN(n8897) );
  AOI21_X1 U9921 ( .B1(n9311), .B2(n8918), .A(n8897), .ZN(n8898) );
  OAI21_X1 U9922 ( .B1(n8899), .B2(n10510), .A(n8898), .ZN(P2_U3237) );
  INV_X1 U9923 ( .A(n8900), .ZN(n8901) );
  NOR2_X1 U9924 ( .A1(n8902), .A2(n8901), .ZN(n8903) );
  XNOR2_X1 U9925 ( .A(n8904), .B(n8903), .ZN(n8910) );
  NAND2_X1 U9926 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8966) );
  OAI21_X1 U9927 ( .B1(n10517), .B2(n8924), .A(n8966), .ZN(n8905) );
  AOI21_X1 U9928 ( .B1(n8906), .B2(n9193), .A(n8905), .ZN(n8907) );
  OAI21_X1 U9929 ( .B1(n9199), .B2(n10523), .A(n8907), .ZN(n8908) );
  AOI21_X1 U9930 ( .B1(n9331), .B2(n8918), .A(n8908), .ZN(n8909) );
  OAI21_X1 U9931 ( .B1(n8910), .B2(n10510), .A(n8909), .ZN(P2_U3240) );
  XNOR2_X1 U9932 ( .A(n8912), .B(n8911), .ZN(n8921) );
  NOR2_X1 U9933 ( .A1(n9075), .A2(n10523), .ZN(n8916) );
  OAI22_X1 U9934 ( .A1(n8914), .A2(n10514), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8913), .ZN(n8915) );
  AOI211_X1 U9935 ( .C1(n9081), .C2(n8917), .A(n8916), .B(n8915), .ZN(n8920)
         );
  NAND2_X1 U9936 ( .A1(n9289), .A2(n8918), .ZN(n8919) );
  OAI211_X1 U9937 ( .C1(n8921), .C2(n10510), .A(n8920), .B(n8919), .ZN(
        P2_U3242) );
  MUX2_X1 U9938 ( .A(n9001), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8933), .Z(
        P2_U3583) );
  MUX2_X1 U9939 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n9011), .S(P2_U3966), .Z(
        P2_U3582) );
  INV_X1 U9940 ( .A(n8922), .ZN(n9046) );
  MUX2_X1 U9941 ( .A(n9046), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8933), .Z(
        P2_U3581) );
  INV_X1 U9942 ( .A(n8923), .ZN(n9056) );
  MUX2_X1 U9943 ( .A(n9056), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8933), .Z(
        P2_U3580) );
  MUX2_X1 U9944 ( .A(n9081), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8933), .Z(
        P2_U3579) );
  MUX2_X1 U9945 ( .A(n9096), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8933), .Z(
        P2_U3578) );
  MUX2_X1 U9946 ( .A(n9103), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8933), .Z(
        P2_U3577) );
  MUX2_X1 U9947 ( .A(n9118), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8933), .Z(
        P2_U3576) );
  MUX2_X1 U9948 ( .A(n9139), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8933), .Z(
        P2_U3575) );
  MUX2_X1 U9949 ( .A(n9146), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8933), .Z(
        P2_U3574) );
  MUX2_X1 U9950 ( .A(n9161), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8933), .Z(
        P2_U3573) );
  MUX2_X1 U9951 ( .A(n9175), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8933), .Z(
        P2_U3572) );
  INV_X1 U9952 ( .A(n8924), .ZN(n9194) );
  MUX2_X1 U9953 ( .A(n9194), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8933), .Z(
        P2_U3571) );
  MUX2_X1 U9954 ( .A(n9174), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8933), .Z(
        P2_U3570) );
  MUX2_X1 U9955 ( .A(n9193), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8933), .Z(
        P2_U3569) );
  MUX2_X1 U9956 ( .A(n9232), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8933), .Z(
        P2_U3568) );
  MUX2_X1 U9957 ( .A(n8925), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8933), .Z(
        P2_U3567) );
  MUX2_X1 U9958 ( .A(n9231), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8933), .Z(
        P2_U3566) );
  MUX2_X1 U9959 ( .A(n8926), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8933), .Z(
        P2_U3565) );
  MUX2_X1 U9960 ( .A(n10588), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8933), .Z(
        P2_U3564) );
  MUX2_X1 U9961 ( .A(n8927), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8933), .Z(
        P2_U3563) );
  MUX2_X1 U9962 ( .A(n8928), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8933), .Z(
        P2_U3560) );
  MUX2_X1 U9963 ( .A(n9250), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8933), .Z(
        P2_U3559) );
  MUX2_X1 U9964 ( .A(n8929), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8933), .Z(
        P2_U3558) );
  MUX2_X1 U9965 ( .A(n9249), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8933), .Z(
        P2_U3557) );
  MUX2_X1 U9966 ( .A(n8930), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8933), .Z(
        P2_U3556) );
  MUX2_X1 U9967 ( .A(n8931), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8933), .Z(
        P2_U3555) );
  MUX2_X1 U9968 ( .A(n8932), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8933), .Z(
        P2_U3554) );
  MUX2_X1 U9969 ( .A(n4859), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8933), .Z(
        P2_U3553) );
  MUX2_X1 U9970 ( .A(n8934), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8933), .Z(
        P2_U3552) );
  OAI21_X1 U9971 ( .B1(n8968), .B2(n8936), .A(n8935), .ZN(n8941) );
  AOI211_X1 U9972 ( .C1(n8939), .C2(n8938), .A(n8937), .B(n4946), .ZN(n8940)
         );
  AOI211_X1 U9973 ( .C1(n10330), .C2(n8942), .A(n8941), .B(n8940), .ZN(n8947)
         );
  OAI21_X1 U9974 ( .B1(n8944), .B2(n5832), .A(n8943), .ZN(n8945) );
  NAND2_X1 U9975 ( .A1(n8994), .A2(n8945), .ZN(n8946) );
  NAND2_X1 U9976 ( .A1(n8947), .A2(n8946), .ZN(P2_U3260) );
  OAI21_X1 U9977 ( .B1(n8950), .B2(n8949), .A(n8948), .ZN(n8960) );
  NAND2_X1 U9978 ( .A1(n10330), .A2(n8951), .ZN(n8953) );
  OAI211_X1 U9979 ( .C1(n8954), .C2(n8968), .A(n8953), .B(n8952), .ZN(n8959)
         );
  AOI211_X1 U9980 ( .C1(n8957), .C2(n8956), .A(n8955), .B(n10320), .ZN(n8958)
         );
  AOI211_X1 U9981 ( .C1(n4948), .C2(n8960), .A(n8959), .B(n8958), .ZN(n8961)
         );
  INV_X1 U9982 ( .A(n8961), .ZN(P2_U3261) );
  INV_X1 U9983 ( .A(n8986), .ZN(n8980) );
  XNOR2_X1 U9984 ( .A(n8986), .B(n8962), .ZN(n8965) );
  AOI21_X1 U9985 ( .B1(n8974), .B2(P2_REG1_REG_17__SCAN_IN), .A(n8963), .ZN(
        n8964) );
  NAND2_X1 U9986 ( .A1(n8965), .A2(n8964), .ZN(n8981) );
  OAI21_X1 U9987 ( .B1(n8965), .B2(n8964), .A(n8981), .ZN(n8970) );
  INV_X1 U9988 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8967) );
  OAI21_X1 U9989 ( .B1(n8968), .B2(n8967), .A(n8966), .ZN(n8969) );
  AOI21_X1 U9990 ( .B1(n4948), .B2(n8970), .A(n8969), .ZN(n8979) );
  NOR2_X1 U9991 ( .A1(n8980), .A2(n8971), .ZN(n8972) );
  AOI21_X1 U9992 ( .B1(n8971), .B2(n8980), .A(n8972), .ZN(n8976) );
  NAND2_X1 U9993 ( .A1(n8976), .A2(n8975), .ZN(n8985) );
  OAI21_X1 U9994 ( .B1(n8976), .B2(n8975), .A(n8985), .ZN(n8977) );
  NAND2_X1 U9995 ( .A1(n8994), .A2(n8977), .ZN(n8978) );
  OAI211_X1 U9996 ( .C1(n8991), .C2(n8980), .A(n8979), .B(n8978), .ZN(P2_U3263) );
  OAI21_X1 U9997 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n8986), .A(n8981), .ZN(
        n8984) );
  XNOR2_X1 U9998 ( .A(n5582), .B(n8982), .ZN(n8983) );
  XNOR2_X1 U9999 ( .A(n8984), .B(n8983), .ZN(n8996) );
  OAI21_X1 U10000 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8986), .A(n8985), .ZN(
        n8988) );
  XNOR2_X1 U10001 ( .A(n5582), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8987) );
  XNOR2_X1 U10002 ( .A(n8988), .B(n8987), .ZN(n8993) );
  NAND2_X1 U10003 ( .A1(n10319), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8989) );
  OAI211_X1 U10004 ( .C1(n8991), .C2(n5582), .A(n8990), .B(n8989), .ZN(n8992)
         );
  AOI21_X1 U10005 ( .B1(n8994), .B2(n8993), .A(n8992), .ZN(n8995) );
  OAI21_X1 U10006 ( .B1(n4946), .B2(n8996), .A(n8995), .ZN(P2_U3264) );
  INV_X1 U10007 ( .A(n9327), .ZN(n8997) );
  INV_X1 U10008 ( .A(n9331), .ZN(n9202) );
  NAND2_X1 U10009 ( .A1(n8997), .A2(n9197), .ZN(n9185) );
  XNOR2_X1 U10010 ( .A(n9004), .B(n8998), .ZN(n9267) );
  NAND2_X1 U10011 ( .A1(n9267), .A2(n9260), .ZN(n9003) );
  AND2_X1 U10012 ( .A1(n8999), .A2(P2_B_REG_SCAN_IN), .ZN(n9000) );
  NOR2_X1 U10013 ( .A1(n9214), .A2(n9000), .ZN(n9012) );
  NAND2_X1 U10014 ( .A1(n9001), .A2(n9012), .ZN(n9270) );
  NOR2_X1 U10015 ( .A1(n10607), .A2(n9270), .ZN(n9006) );
  AOI21_X1 U10016 ( .B1(n10607), .B2(P2_REG2_REG_31__SCAN_IN), .A(n9006), .ZN(
        n9002) );
  OAI211_X1 U10017 ( .C1(n9268), .C2(n10383), .A(n9003), .B(n9002), .ZN(
        P2_U3265) );
  AOI21_X1 U10018 ( .B1(n9005), .B2(n9038), .A(n9004), .ZN(n9269) );
  NAND2_X1 U10019 ( .A1(n9269), .A2(n9260), .ZN(n9008) );
  AOI21_X1 U10020 ( .B1(n10607), .B2(P2_REG2_REG_30__SCAN_IN), .A(n9006), .ZN(
        n9007) );
  OAI211_X1 U10021 ( .C1(n5333), .C2(n10383), .A(n9008), .B(n9007), .ZN(
        P2_U3266) );
  XNOR2_X1 U10022 ( .A(n9033), .B(n9009), .ZN(n9010) );
  NAND2_X1 U10023 ( .A1(n9010), .A2(n9234), .ZN(n9014) );
  AOI22_X1 U10024 ( .A1(n9056), .A2(n9230), .B1(n9012), .B2(n9011), .ZN(n9013)
         );
  OR2_X1 U10025 ( .A1(n9337), .A2(n9193), .ZN(n9015) );
  NOR2_X1 U10026 ( .A1(n9331), .A2(n9174), .ZN(n9016) );
  NAND2_X1 U10027 ( .A1(n9179), .A2(n9178), .ZN(n9177) );
  NAND2_X1 U10028 ( .A1(n9327), .A2(n9194), .ZN(n9017) );
  NAND2_X1 U10029 ( .A1(n9177), .A2(n9017), .ZN(n9169) );
  NAND2_X1 U10030 ( .A1(n9321), .A2(n9175), .ZN(n9018) );
  OR2_X1 U10031 ( .A1(n9311), .A2(n9146), .ZN(n9020) );
  NAND2_X1 U10032 ( .A1(n9021), .A2(n9020), .ZN(n9120) );
  NAND2_X1 U10033 ( .A1(n9305), .A2(n9139), .ZN(n9022) );
  OR2_X1 U10034 ( .A1(n9298), .A2(n9118), .ZN(n9023) );
  OR2_X1 U10035 ( .A1(n9294), .A2(n9103), .ZN(n9071) );
  OR2_X1 U10036 ( .A1(n9289), .A2(n9096), .ZN(n9025) );
  AND2_X1 U10037 ( .A1(n9071), .A2(n9025), .ZN(n9058) );
  OR2_X1 U10038 ( .A1(n9283), .A2(n9081), .ZN(n9024) );
  AND2_X1 U10039 ( .A1(n9058), .A2(n9024), .ZN(n9030) );
  INV_X1 U10040 ( .A(n9024), .ZN(n9029) );
  INV_X1 U10041 ( .A(n9025), .ZN(n9026) );
  OR2_X1 U10042 ( .A1(n9026), .A2(n9079), .ZN(n9059) );
  AND2_X1 U10043 ( .A1(n9027), .A2(n9059), .ZN(n9028) );
  NAND2_X1 U10044 ( .A1(n9051), .A2(n9044), .ZN(n9032) );
  OR2_X1 U10045 ( .A1(n9278), .A2(n9056), .ZN(n9031) );
  NAND2_X1 U10046 ( .A1(n9032), .A2(n9031), .ZN(n9034) );
  XNOR2_X1 U10047 ( .A(n9034), .B(n9033), .ZN(n9272) );
  NAND2_X1 U10048 ( .A1(n9036), .A2(n9035), .ZN(n9037) );
  NAND2_X1 U10049 ( .A1(n9038), .A2(n9037), .ZN(n9274) );
  NOR2_X1 U10050 ( .A1(n9274), .A2(n10382), .ZN(n9042) );
  AOI22_X1 U10051 ( .A1(n9039), .A2(n9238), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n10607), .ZN(n9040) );
  OAI21_X1 U10052 ( .B1(n9273), .B2(n10383), .A(n9040), .ZN(n9041) );
  AOI211_X1 U10053 ( .C1(n9272), .C2(n9263), .A(n9042), .B(n9041), .ZN(n9043)
         );
  OAI21_X1 U10054 ( .B1(n5469), .B2(n10607), .A(n9043), .ZN(P2_U3267) );
  AOI21_X1 U10055 ( .B1(n9278), .B2(n9063), .A(n9047), .ZN(n9279) );
  AOI22_X1 U10056 ( .A1(n9048), .A2(n9238), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n10607), .ZN(n9049) );
  OAI21_X1 U10057 ( .B1(n6113), .B2(n10383), .A(n9049), .ZN(n9053) );
  XNOR2_X1 U10058 ( .A(n9051), .B(n9050), .ZN(n9282) );
  NOR2_X1 U10059 ( .A1(n9282), .A2(n9244), .ZN(n9052) );
  OAI21_X1 U10060 ( .B1(n9281), .B2(n10607), .A(n9054), .ZN(P2_U3268) );
  XNOR2_X1 U10061 ( .A(n5277), .B(n9055), .ZN(n9057) );
  AOI222_X1 U10062 ( .A1(n9234), .A2(n9057), .B1(n9056), .B2(n10587), .C1(
        n9096), .C2(n9230), .ZN(n9286) );
  NAND2_X1 U10063 ( .A1(n9072), .A2(n9058), .ZN(n9060) );
  INV_X1 U10064 ( .A(n9287), .ZN(n9069) );
  NAND2_X1 U10065 ( .A1(n9283), .A2(n9074), .ZN(n9062) );
  AND2_X1 U10066 ( .A1(n9063), .A2(n9062), .ZN(n9284) );
  NAND2_X1 U10067 ( .A1(n9284), .A2(n9260), .ZN(n9066) );
  AOI22_X1 U10068 ( .A1(n9064), .A2(n9238), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n10607), .ZN(n9065) );
  OAI211_X1 U10069 ( .C1(n9067), .C2(n10383), .A(n9066), .B(n9065), .ZN(n9068)
         );
  AOI21_X1 U10070 ( .B1(n9069), .B2(n9263), .A(n9068), .ZN(n9070) );
  OAI21_X1 U10071 ( .B1(n10607), .B2(n9286), .A(n9070), .ZN(P2_U3269) );
  NAND2_X1 U10072 ( .A1(n9072), .A2(n9071), .ZN(n9073) );
  XOR2_X1 U10073 ( .A(n9079), .B(n9073), .Z(n9292) );
  AOI211_X1 U10074 ( .C1(n9289), .C2(n9087), .A(n10650), .B(n5165), .ZN(n9288)
         );
  INV_X1 U10075 ( .A(n9289), .ZN(n9078) );
  INV_X1 U10076 ( .A(n9075), .ZN(n9076) );
  AOI22_X1 U10077 ( .A1(n9076), .A2(n9238), .B1(P2_REG2_REG_26__SCAN_IN), .B2(
        n10607), .ZN(n9077) );
  OAI21_X1 U10078 ( .B1(n9078), .B2(n10383), .A(n9077), .ZN(n9084) );
  XNOR2_X1 U10079 ( .A(n9080), .B(n9079), .ZN(n9082) );
  AOI222_X1 U10080 ( .A1(n9234), .A2(n9082), .B1(n9081), .B2(n10587), .C1(
        n9103), .C2(n9230), .ZN(n9291) );
  NOR2_X1 U10081 ( .A1(n9291), .A2(n10607), .ZN(n9083) );
  AOI211_X1 U10082 ( .C1(n9288), .C2(n9186), .A(n9084), .B(n9083), .ZN(n9085)
         );
  OAI21_X1 U10083 ( .B1(n9292), .B2(n9244), .A(n9085), .ZN(P2_U3270) );
  XNOR2_X1 U10084 ( .A(n9086), .B(n5332), .ZN(n9297) );
  INV_X1 U10085 ( .A(n9087), .ZN(n9088) );
  AOI211_X1 U10086 ( .C1(n9294), .C2(n9089), .A(n10650), .B(n9088), .ZN(n9293)
         );
  INV_X1 U10087 ( .A(n9294), .ZN(n9093) );
  INV_X1 U10088 ( .A(n9090), .ZN(n9091) );
  AOI22_X1 U10089 ( .A1(n9091), .A2(n9238), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n10607), .ZN(n9092) );
  OAI21_X1 U10090 ( .B1(n9093), .B2(n10383), .A(n9092), .ZN(n9099) );
  XNOR2_X1 U10091 ( .A(n9095), .B(n9094), .ZN(n9097) );
  AOI222_X1 U10092 ( .A1(n9234), .A2(n9097), .B1(n9096), .B2(n10587), .C1(
        n9118), .C2(n9230), .ZN(n9296) );
  NOR2_X1 U10093 ( .A1(n9296), .A2(n10607), .ZN(n9098) );
  AOI211_X1 U10094 ( .C1(n9186), .C2(n9293), .A(n9099), .B(n9098), .ZN(n9100)
         );
  OAI21_X1 U10095 ( .B1(n9297), .B2(n9244), .A(n9100), .ZN(P2_U3271) );
  NAND2_X1 U10096 ( .A1(n9116), .A2(n9101), .ZN(n9102) );
  XNOR2_X1 U10097 ( .A(n9111), .B(n9102), .ZN(n9104) );
  AOI222_X1 U10098 ( .A1(n9234), .A2(n9104), .B1(n9103), .B2(n10587), .C1(
        n9139), .C2(n9230), .ZN(n9301) );
  XNOR2_X1 U10099 ( .A(n9123), .B(n9298), .ZN(n9299) );
  AOI22_X1 U10100 ( .A1(n10607), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n9105), 
        .B2(n9238), .ZN(n9106) );
  OAI21_X1 U10101 ( .B1(n9107), .B2(n10383), .A(n9106), .ZN(n9113) );
  INV_X1 U10102 ( .A(n9108), .ZN(n9109) );
  AOI211_X1 U10103 ( .C1(n9299), .C2(n9260), .A(n9113), .B(n9112), .ZN(n9114)
         );
  OAI21_X1 U10104 ( .B1(n10607), .B2(n9301), .A(n9114), .ZN(P2_U3272) );
  INV_X1 U10105 ( .A(n9115), .ZN(n9117) );
  OAI21_X1 U10106 ( .B1(n9117), .B2(n9121), .A(n9116), .ZN(n9119) );
  AOI222_X1 U10107 ( .A1(n9234), .A2(n9119), .B1(n9146), .B2(n9230), .C1(n9118), .C2(n10587), .ZN(n9309) );
  NAND2_X1 U10108 ( .A1(n9120), .A2(n9121), .ZN(n9303) );
  NAND3_X1 U10109 ( .A1(n9304), .A2(n9303), .A3(n9263), .ZN(n9129) );
  AND2_X1 U10110 ( .A1(n9305), .A2(n4884), .ZN(n9122) );
  NOR2_X1 U10111 ( .A1(n9123), .A2(n9122), .ZN(n9306) );
  NAND2_X1 U10112 ( .A1(n9305), .A2(n9223), .ZN(n9125) );
  NAND2_X1 U10113 ( .A1(n10607), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n9124) );
  OAI211_X1 U10114 ( .C1(n10609), .C2(n9126), .A(n9125), .B(n9124), .ZN(n9127)
         );
  AOI21_X1 U10115 ( .B1(n9306), .B2(n9260), .A(n9127), .ZN(n9128) );
  OAI211_X1 U10116 ( .C1(n10607), .C2(n9309), .A(n9129), .B(n9128), .ZN(
        P2_U3273) );
  XNOR2_X1 U10117 ( .A(n9131), .B(n9130), .ZN(n9315) );
  INV_X1 U10118 ( .A(n4884), .ZN(n9132) );
  AOI21_X1 U10119 ( .B1(n9311), .B2(n9148), .A(n9132), .ZN(n9312) );
  INV_X1 U10120 ( .A(n9133), .ZN(n9134) );
  AOI22_X1 U10121 ( .A1(n10607), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9134), 
        .B2(n9238), .ZN(n9135) );
  OAI21_X1 U10122 ( .B1(n9136), .B2(n10383), .A(n9135), .ZN(n9142) );
  XNOR2_X1 U10123 ( .A(n9138), .B(n9137), .ZN(n9140) );
  AOI222_X1 U10124 ( .A1(n9234), .A2(n9140), .B1(n9161), .B2(n9230), .C1(n9139), .C2(n10587), .ZN(n9314) );
  NOR2_X1 U10125 ( .A1(n9314), .A2(n10607), .ZN(n9141) );
  AOI211_X1 U10126 ( .C1(n9312), .C2(n9260), .A(n9142), .B(n9141), .ZN(n9143)
         );
  OAI21_X1 U10127 ( .B1(n9315), .B2(n9244), .A(n9143), .ZN(P2_U3274) );
  XNOR2_X1 U10128 ( .A(n9145), .B(n9144), .ZN(n9147) );
  AOI222_X1 U10129 ( .A1(n9234), .A2(n9147), .B1(n9146), .B2(n10587), .C1(
        n9175), .C2(n9230), .ZN(n9319) );
  INV_X1 U10130 ( .A(n9148), .ZN(n9149) );
  AOI21_X1 U10131 ( .B1(n9316), .B2(n9163), .A(n9149), .ZN(n9317) );
  INV_X1 U10132 ( .A(n9150), .ZN(n9151) );
  AOI22_X1 U10133 ( .A1(n10607), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9151), 
        .B2(n9238), .ZN(n9152) );
  OAI21_X1 U10134 ( .B1(n5163), .B2(n10383), .A(n9152), .ZN(n9158) );
  INV_X1 U10135 ( .A(n9153), .ZN(n9154) );
  AOI21_X1 U10136 ( .B1(n9156), .B2(n9155), .A(n9154), .ZN(n9320) );
  NOR2_X1 U10137 ( .A1(n9320), .A2(n9244), .ZN(n9157) );
  AOI211_X1 U10138 ( .C1(n9317), .C2(n9260), .A(n9158), .B(n9157), .ZN(n9159)
         );
  OAI21_X1 U10139 ( .B1(n10607), .B2(n9319), .A(n9159), .ZN(P2_U3275) );
  XNOR2_X1 U10140 ( .A(n9160), .B(n9168), .ZN(n9162) );
  AOI222_X1 U10141 ( .A1(n9234), .A2(n9162), .B1(n9161), .B2(n10587), .C1(
        n9194), .C2(n9230), .ZN(n9324) );
  AOI21_X1 U10142 ( .B1(n9321), .B2(n9185), .A(n5164), .ZN(n9322) );
  INV_X1 U10143 ( .A(n9321), .ZN(n9166) );
  AOI22_X1 U10144 ( .A1(n10607), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9164), 
        .B2(n9238), .ZN(n9165) );
  OAI21_X1 U10145 ( .B1(n9166), .B2(n10383), .A(n9165), .ZN(n9171) );
  OAI21_X1 U10146 ( .B1(n9169), .B2(n9168), .A(n9167), .ZN(n9325) );
  NOR2_X1 U10147 ( .A1(n9325), .A2(n9244), .ZN(n9170) );
  AOI211_X1 U10148 ( .C1(n9322), .C2(n9260), .A(n9171), .B(n9170), .ZN(n9172)
         );
  OAI21_X1 U10149 ( .B1(n10607), .B2(n9324), .A(n9172), .ZN(P2_U3276) );
  XNOR2_X1 U10150 ( .A(n9173), .B(n9178), .ZN(n9176) );
  AOI222_X1 U10151 ( .A1(n9234), .A2(n9176), .B1(n9175), .B2(n10587), .C1(
        n9174), .C2(n9230), .ZN(n9329) );
  OAI21_X1 U10152 ( .B1(n9179), .B2(n9178), .A(n9177), .ZN(n9330) );
  OAI22_X1 U10153 ( .A1(n10605), .A2(n9181), .B1(n9180), .B2(n10609), .ZN(
        n9182) );
  AOI21_X1 U10154 ( .B1(n9327), .B2(n9223), .A(n9182), .ZN(n9188) );
  INV_X1 U10155 ( .A(n9197), .ZN(n9183) );
  NAND2_X1 U10156 ( .A1(n9183), .A2(n9327), .ZN(n9184) );
  AND3_X1 U10157 ( .A1(n9185), .A2(n10629), .A3(n9184), .ZN(n9326) );
  NAND2_X1 U10158 ( .A1(n9326), .A2(n9186), .ZN(n9187) );
  OAI211_X1 U10159 ( .C1(n9330), .C2(n9244), .A(n9188), .B(n9187), .ZN(n9189)
         );
  INV_X1 U10160 ( .A(n9189), .ZN(n9190) );
  OAI21_X1 U10161 ( .B1(n10607), .B2(n9329), .A(n9190), .ZN(P2_U3277) );
  XNOR2_X1 U10162 ( .A(n9191), .B(n9192), .ZN(n9195) );
  AOI222_X1 U10163 ( .A1(n9234), .A2(n9195), .B1(n9194), .B2(n10587), .C1(
        n9193), .C2(n9230), .ZN(n9334) );
  NOR2_X1 U10164 ( .A1(n9202), .A2(n9196), .ZN(n9198) );
  NOR2_X1 U10165 ( .A1(n9198), .A2(n9197), .ZN(n9332) );
  INV_X1 U10166 ( .A(n9199), .ZN(n9200) );
  AOI22_X1 U10167 ( .A1(n10607), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9200), 
        .B2(n9238), .ZN(n9201) );
  OAI21_X1 U10168 ( .B1(n9202), .B2(n10383), .A(n9201), .ZN(n9206) );
  XNOR2_X1 U10169 ( .A(n9204), .B(n9203), .ZN(n9335) );
  NOR2_X1 U10170 ( .A1(n9335), .A2(n9244), .ZN(n9205) );
  AOI211_X1 U10171 ( .C1(n9332), .C2(n9260), .A(n9206), .B(n9205), .ZN(n9207)
         );
  OAI21_X1 U10172 ( .B1(n10607), .B2(n9334), .A(n9207), .ZN(P2_U3278) );
  XNOR2_X1 U10173 ( .A(n9208), .B(n9211), .ZN(n9209) );
  NAND2_X1 U10174 ( .A1(n9209), .A2(n9234), .ZN(n9339) );
  OAI21_X1 U10175 ( .B1(n4941), .B2(n9211), .A(n9210), .ZN(n9336) );
  INV_X1 U10176 ( .A(n9212), .ZN(n9213) );
  XNOR2_X1 U10177 ( .A(n9213), .B(n9337), .ZN(n9219) );
  OAI22_X1 U10178 ( .A1(n9217), .A2(n9216), .B1(n9215), .B2(n9214), .ZN(n9218)
         );
  AOI21_X1 U10179 ( .B1(n9219), .B2(n10629), .A(n9218), .ZN(n9340) );
  INV_X1 U10180 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9221) );
  OAI22_X1 U10181 ( .A1(n10605), .A2(n9221), .B1(n9220), .B2(n10609), .ZN(
        n9222) );
  AOI21_X1 U10182 ( .B1(n9337), .B2(n9223), .A(n9222), .ZN(n9224) );
  OAI21_X1 U10183 ( .B1(n9340), .B2(n9225), .A(n9224), .ZN(n9226) );
  AOI21_X1 U10184 ( .B1(n9336), .B2(n9263), .A(n9226), .ZN(n9227) );
  OAI21_X1 U10185 ( .B1(n10607), .B2(n9339), .A(n9227), .ZN(P2_U3279) );
  XNOR2_X1 U10186 ( .A(n9229), .B(n9228), .ZN(n9233) );
  AOI222_X1 U10187 ( .A1(n9234), .A2(n9233), .B1(n9232), .B2(n10587), .C1(
        n9231), .C2(n9230), .ZN(n9350) );
  AOI21_X1 U10188 ( .B1(n9347), .B2(n9236), .A(n5162), .ZN(n9348) );
  INV_X1 U10189 ( .A(n9347), .ZN(n9241) );
  INV_X1 U10190 ( .A(n9237), .ZN(n9239) );
  AOI22_X1 U10191 ( .A1(n10607), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n9239), 
        .B2(n9238), .ZN(n9240) );
  OAI21_X1 U10192 ( .B1(n9241), .B2(n10383), .A(n9240), .ZN(n9246) );
  XNOR2_X1 U10193 ( .A(n9243), .B(n9242), .ZN(n9351) );
  NOR2_X1 U10194 ( .A1(n9351), .A2(n9244), .ZN(n9245) );
  AOI211_X1 U10195 ( .C1(n9348), .C2(n9260), .A(n9246), .B(n9245), .ZN(n9247)
         );
  OAI21_X1 U10196 ( .B1(n10607), .B2(n9350), .A(n9247), .ZN(P2_U3281) );
  XNOR2_X1 U10197 ( .A(n9248), .B(n9261), .ZN(n9251) );
  AOI222_X1 U10198 ( .A1(n9234), .A2(n9251), .B1(n9250), .B2(n10587), .C1(
        n9249), .C2(n9230), .ZN(n10498) );
  MUX2_X1 U10199 ( .A(n9252), .B(n10498), .S(n10605), .Z(n9266) );
  INV_X1 U10200 ( .A(n9253), .ZN(n9256) );
  INV_X1 U10201 ( .A(n9254), .ZN(n9255) );
  AOI21_X1 U10202 ( .B1(n10492), .B2(n9256), .A(n9255), .ZN(n10493) );
  OAI22_X1 U10203 ( .A1(n10383), .A2(n9258), .B1(n9257), .B2(n10609), .ZN(
        n9259) );
  AOI21_X1 U10204 ( .B1(n10493), .B2(n9260), .A(n9259), .ZN(n9265) );
  NAND2_X1 U10205 ( .A1(n9262), .A2(n9261), .ZN(n10494) );
  NAND3_X1 U10206 ( .A1(n10495), .A2(n10494), .A3(n9263), .ZN(n9264) );
  NAND3_X1 U10207 ( .A1(n9266), .A2(n9265), .A3(n9264), .ZN(P2_U3290) );
  MUX2_X1 U10208 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9352), .S(n10657), .Z(
        P2_U3551) );
  NAND2_X1 U10209 ( .A1(n9269), .A2(n10629), .ZN(n9271) );
  OAI211_X1 U10210 ( .C1(n5333), .C2(n10648), .A(n9271), .B(n9270), .ZN(n9353)
         );
  MUX2_X1 U10211 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9353), .S(n10657), .Z(
        P2_U3550) );
  OAI22_X1 U10212 ( .A1(n9274), .A2(n10650), .B1(n9273), .B2(n10648), .ZN(
        n9275) );
  INV_X1 U10213 ( .A(n9275), .ZN(n9276) );
  NAND3_X1 U10214 ( .A1(n9277), .A2(n5469), .A3(n9276), .ZN(n9354) );
  MUX2_X1 U10215 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9354), .S(n10657), .Z(
        P2_U3549) );
  AOI22_X1 U10216 ( .A1(n9279), .A2(n10629), .B1(n10628), .B2(n9278), .ZN(
        n9280) );
  OAI211_X1 U10217 ( .C1(n9282), .C2(n10530), .A(n9281), .B(n9280), .ZN(n9355)
         );
  MUX2_X1 U10218 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9355), .S(n10657), .Z(
        P2_U3548) );
  AOI22_X1 U10219 ( .A1(n9284), .A2(n10629), .B1(n10628), .B2(n9283), .ZN(
        n9285) );
  OAI211_X1 U10220 ( .C1(n9287), .C2(n10530), .A(n9286), .B(n9285), .ZN(n9356)
         );
  MUX2_X1 U10221 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9356), .S(n10657), .Z(
        P2_U3547) );
  AOI21_X1 U10222 ( .B1(n10628), .B2(n9289), .A(n9288), .ZN(n9290) );
  OAI211_X1 U10223 ( .C1(n9292), .C2(n10530), .A(n9291), .B(n9290), .ZN(n9357)
         );
  MUX2_X1 U10224 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9357), .S(n10657), .Z(
        P2_U3546) );
  AOI21_X1 U10225 ( .B1(n10628), .B2(n9294), .A(n9293), .ZN(n9295) );
  OAI211_X1 U10226 ( .C1(n9297), .C2(n10530), .A(n9296), .B(n9295), .ZN(n9358)
         );
  MUX2_X1 U10227 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9358), .S(n10657), .Z(
        P2_U3545) );
  AOI22_X1 U10228 ( .A1(n9299), .A2(n10629), .B1(n10628), .B2(n9298), .ZN(
        n9300) );
  OAI211_X1 U10229 ( .C1(n9302), .C2(n10530), .A(n9301), .B(n9300), .ZN(n9359)
         );
  MUX2_X1 U10230 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9359), .S(n10657), .Z(
        P2_U3544) );
  NAND3_X1 U10231 ( .A1(n9304), .A2(n10654), .A3(n9303), .ZN(n9310) );
  NAND2_X1 U10232 ( .A1(n9305), .A2(n10628), .ZN(n9308) );
  NAND2_X1 U10233 ( .A1(n9306), .A2(n10629), .ZN(n9307) );
  NAND4_X1 U10234 ( .A1(n9310), .A2(n9309), .A3(n9308), .A4(n9307), .ZN(n9360)
         );
  MUX2_X1 U10235 ( .A(n9360), .B(P2_REG1_REG_23__SCAN_IN), .S(n10656), .Z(
        P2_U3543) );
  AOI22_X1 U10236 ( .A1(n9312), .A2(n10629), .B1(n10628), .B2(n9311), .ZN(
        n9313) );
  OAI211_X1 U10237 ( .C1(n9315), .C2(n10530), .A(n9314), .B(n9313), .ZN(n9361)
         );
  MUX2_X1 U10238 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9361), .S(n10657), .Z(
        P2_U3542) );
  AOI22_X1 U10239 ( .A1(n9317), .A2(n10629), .B1(n10628), .B2(n9316), .ZN(
        n9318) );
  OAI211_X1 U10240 ( .C1(n9320), .C2(n10530), .A(n9319), .B(n9318), .ZN(n9362)
         );
  MUX2_X1 U10241 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9362), .S(n10657), .Z(
        P2_U3541) );
  AOI22_X1 U10242 ( .A1(n9322), .A2(n10629), .B1(n10628), .B2(n9321), .ZN(
        n9323) );
  OAI211_X1 U10243 ( .C1(n9325), .C2(n10530), .A(n9324), .B(n9323), .ZN(n9363)
         );
  MUX2_X1 U10244 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9363), .S(n10657), .Z(
        P2_U3540) );
  AOI21_X1 U10245 ( .B1(n10628), .B2(n9327), .A(n9326), .ZN(n9328) );
  OAI211_X1 U10246 ( .C1(n9330), .C2(n10530), .A(n9329), .B(n9328), .ZN(n9364)
         );
  MUX2_X1 U10247 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9364), .S(n10657), .Z(
        P2_U3539) );
  AOI22_X1 U10248 ( .A1(n9332), .A2(n10629), .B1(n10628), .B2(n9331), .ZN(
        n9333) );
  OAI211_X1 U10249 ( .C1(n9335), .C2(n10530), .A(n9334), .B(n9333), .ZN(n9365)
         );
  MUX2_X1 U10250 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9365), .S(n10657), .Z(
        P2_U3538) );
  NAND2_X1 U10251 ( .A1(n9336), .A2(n10654), .ZN(n9341) );
  NAND2_X1 U10252 ( .A1(n9337), .A2(n10628), .ZN(n9338) );
  NAND4_X1 U10253 ( .A1(n9341), .A2(n9340), .A3(n9339), .A4(n9338), .ZN(n9366)
         );
  MUX2_X1 U10254 ( .A(n9366), .B(P2_REG1_REG_17__SCAN_IN), .S(n10656), .Z(
        P2_U3537) );
  AOI21_X1 U10255 ( .B1(n10628), .B2(n9343), .A(n9342), .ZN(n9344) );
  OAI211_X1 U10256 ( .C1(n9346), .C2(n10530), .A(n9345), .B(n9344), .ZN(n9367)
         );
  MUX2_X1 U10257 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9367), .S(n10657), .Z(
        P2_U3536) );
  AOI22_X1 U10258 ( .A1(n9348), .A2(n10629), .B1(n10628), .B2(n9347), .ZN(
        n9349) );
  OAI211_X1 U10259 ( .C1(n9351), .C2(n10530), .A(n9350), .B(n9349), .ZN(n9368)
         );
  MUX2_X1 U10260 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9368), .S(n10657), .Z(
        P2_U3535) );
  MUX2_X1 U10261 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9352), .S(n10660), .Z(
        P2_U3519) );
  MUX2_X1 U10262 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9353), .S(n10660), .Z(
        P2_U3518) );
  MUX2_X1 U10263 ( .A(n9354), .B(P2_REG0_REG_29__SCAN_IN), .S(n10658), .Z(
        P2_U3517) );
  MUX2_X1 U10264 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9355), .S(n10660), .Z(
        P2_U3516) );
  MUX2_X1 U10265 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9356), .S(n10660), .Z(
        P2_U3515) );
  MUX2_X1 U10266 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9357), .S(n10660), .Z(
        P2_U3514) );
  MUX2_X1 U10267 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9358), .S(n10660), .Z(
        P2_U3513) );
  MUX2_X1 U10268 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9359), .S(n10660), .Z(
        P2_U3512) );
  MUX2_X1 U10269 ( .A(n9360), .B(P2_REG0_REG_23__SCAN_IN), .S(n10658), .Z(
        P2_U3511) );
  MUX2_X1 U10270 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9361), .S(n10660), .Z(
        P2_U3510) );
  MUX2_X1 U10271 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9362), .S(n10660), .Z(
        P2_U3509) );
  MUX2_X1 U10272 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9363), .S(n10660), .Z(
        P2_U3508) );
  MUX2_X1 U10273 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9364), .S(n10660), .Z(
        P2_U3507) );
  MUX2_X1 U10274 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9365), .S(n10660), .Z(
        P2_U3505) );
  MUX2_X1 U10275 ( .A(n9366), .B(P2_REG0_REG_17__SCAN_IN), .S(n10658), .Z(
        P2_U3502) );
  MUX2_X1 U10276 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9367), .S(n10660), .Z(
        P2_U3499) );
  MUX2_X1 U10277 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9368), .S(n10660), .Z(
        P2_U3496) );
  INV_X1 U10278 ( .A(n9955), .ZN(n9372) );
  NOR4_X1 U10279 ( .A1(n4870), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3152), .A4(
        n9369), .ZN(n9370) );
  AOI21_X1 U10280 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n9373), .A(n9370), .ZN(
        n9371) );
  OAI21_X1 U10281 ( .B1(n9372), .B2(n9380), .A(n9371), .ZN(P2_U3327) );
  AOI22_X1 U10282 ( .A1(n9374), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9373), .ZN(n9375) );
  OAI21_X1 U10283 ( .B1(n9376), .B2(n9380), .A(n9375), .ZN(P2_U3328) );
  OAI222_X1 U10284 ( .A1(n9380), .A2(n9379), .B1(n9385), .B2(n9378), .C1(
        P2_U3152), .C2(n9377), .ZN(P2_U3329) );
  OAI222_X1 U10285 ( .A1(n9385), .A2(n7021), .B1(n9380), .B2(n9381), .C1(
        P2_U3152), .C2(n6125), .ZN(P2_U3330) );
  INV_X1 U10286 ( .A(n9382), .ZN(n9960) );
  OAI222_X1 U10287 ( .A1(n9380), .A2(n9960), .B1(n9383), .B2(P2_U3152), .C1(
        n7000), .C2(n9385), .ZN(P2_U3331) );
  INV_X1 U10288 ( .A(n9384), .ZN(n9963) );
  INV_X1 U10289 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9386) );
  OAI222_X1 U10290 ( .A1(n9380), .A2(n9963), .B1(P2_U3152), .B2(n9387), .C1(
        n9386), .C2(n9385), .ZN(P2_U3332) );
  MUX2_X1 U10291 ( .A(n9389), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10292 ( .A(n9391), .ZN(n9392) );
  NOR2_X1 U10293 ( .A1(n9393), .A2(n9392), .ZN(n9394) );
  XNOR2_X1 U10294 ( .A(n9390), .B(n9394), .ZN(n9400) );
  OAI22_X1 U10295 ( .A1(n9647), .A2(n9521), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9395), .ZN(n9397) );
  NOR2_X1 U10296 ( .A1(n9648), .A2(n9507), .ZN(n9396) );
  AOI211_X1 U10297 ( .C1(n9643), .C2(n9510), .A(n9397), .B(n9396), .ZN(n9399)
         );
  NAND2_X1 U10298 ( .A1(n9848), .A2(n9528), .ZN(n9398) );
  OAI211_X1 U10299 ( .C1(n9400), .C2(n9530), .A(n9399), .B(n9398), .ZN(
        P1_U3212) );
  XNOR2_X1 U10300 ( .A(n9403), .B(n9402), .ZN(n9404) );
  XNOR2_X1 U10301 ( .A(n9401), .B(n9404), .ZN(n9409) );
  NOR2_X1 U10302 ( .A1(n9526), .A2(n9702), .ZN(n9407) );
  AOI22_X1 U10303 ( .A1(n9710), .A2(n9523), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n9405) );
  OAI21_X1 U10304 ( .B1(n9742), .B2(n9521), .A(n9405), .ZN(n9406) );
  AOI211_X1 U10305 ( .C1(n9869), .C2(n9528), .A(n9407), .B(n9406), .ZN(n9408)
         );
  OAI21_X1 U10306 ( .B1(n9409), .B2(n9530), .A(n9408), .ZN(P1_U3214) );
  XOR2_X1 U10307 ( .A(n9410), .B(n9411), .Z(n9416) );
  NOR2_X1 U10308 ( .A1(n9526), .A2(n9772), .ZN(n9414) );
  NAND2_X1 U10309 ( .A1(n9523), .A2(n9534), .ZN(n9412) );
  NAND2_X1 U10310 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9601) );
  OAI211_X1 U10311 ( .C1(n9809), .C2(n9521), .A(n9412), .B(n9601), .ZN(n9413)
         );
  AOI211_X1 U10312 ( .C1(n9892), .C2(n9528), .A(n9414), .B(n9413), .ZN(n9415)
         );
  OAI21_X1 U10313 ( .B1(n9416), .B2(n9530), .A(n9415), .ZN(P1_U3217) );
  INV_X1 U10314 ( .A(n9417), .ZN(n9421) );
  OAI21_X1 U10315 ( .B1(n9419), .B2(n9421), .A(n9418), .ZN(n9420) );
  OAI21_X1 U10316 ( .B1(n5471), .B2(n9421), .A(n9420), .ZN(n9422) );
  NAND2_X1 U10317 ( .A1(n9422), .A2(n9485), .ZN(n9426) );
  AOI22_X1 U10318 ( .A1(n9523), .A2(n9709), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n9423) );
  OAI21_X1 U10319 ( .B1(n9780), .B2(n9521), .A(n9423), .ZN(n9424) );
  AOI21_X1 U10320 ( .B1(n9746), .B2(n9510), .A(n9424), .ZN(n9425) );
  OAI211_X1 U10321 ( .C1(n8800), .C2(n9513), .A(n9426), .B(n9425), .ZN(
        P1_U3221) );
  XOR2_X1 U10322 ( .A(n9428), .B(n9427), .Z(n9434) );
  NOR2_X1 U10323 ( .A1(n9526), .A2(n9670), .ZN(n9432) );
  AOI22_X1 U10324 ( .A1(n9677), .A2(n9523), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9429) );
  OAI21_X1 U10325 ( .B1(n9430), .B2(n9521), .A(n9429), .ZN(n9431) );
  AOI211_X1 U10326 ( .C1(n9859), .C2(n9528), .A(n9432), .B(n9431), .ZN(n9433)
         );
  OAI21_X1 U10327 ( .B1(n9434), .B2(n9530), .A(n9433), .ZN(P1_U3223) );
  INV_X1 U10328 ( .A(n9436), .ZN(n9437) );
  AOI21_X1 U10329 ( .B1(n9438), .B2(n9435), .A(n9437), .ZN(n9445) );
  NOR2_X1 U10330 ( .A1(n9526), .A2(n9439), .ZN(n9443) );
  NAND2_X1 U10331 ( .A1(n9523), .A2(n9799), .ZN(n9440) );
  NAND2_X1 U10332 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9558) );
  OAI211_X1 U10333 ( .C1(n9441), .C2(n9521), .A(n9440), .B(n9558), .ZN(n9442)
         );
  AOI211_X1 U10334 ( .C1(n9908), .C2(n9528), .A(n9443), .B(n9442), .ZN(n9444)
         );
  OAI21_X1 U10335 ( .B1(n9445), .B2(n9530), .A(n9444), .ZN(P1_U3224) );
  NAND2_X1 U10336 ( .A1(n4934), .A2(n9446), .ZN(n9447) );
  XNOR2_X1 U10337 ( .A(n9448), .B(n9447), .ZN(n9455) );
  NOR2_X1 U10338 ( .A1(n9449), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9573) );
  NOR2_X1 U10339 ( .A1(n9521), .A2(n9450), .ZN(n9451) );
  AOI211_X1 U10340 ( .C1(n9523), .C2(n9535), .A(n9573), .B(n9451), .ZN(n9452)
         );
  OAI21_X1 U10341 ( .B1(n9526), .B2(n9820), .A(n9452), .ZN(n9453) );
  AOI21_X1 U10342 ( .B1(n9901), .B2(n9528), .A(n9453), .ZN(n9454) );
  OAI21_X1 U10343 ( .B1(n9455), .B2(n9530), .A(n9454), .ZN(P1_U3226) );
  XOR2_X1 U10344 ( .A(n9457), .B(n9456), .Z(n9463) );
  AOI22_X1 U10345 ( .A1(n9533), .A2(n9523), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9459) );
  NAND2_X1 U10346 ( .A1(n9510), .A2(n9692), .ZN(n9458) );
  OAI211_X1 U10347 ( .C1(n9460), .C2(n9521), .A(n9459), .B(n9458), .ZN(n9461)
         );
  AOI21_X1 U10348 ( .B1(n9866), .B2(n9528), .A(n9461), .ZN(n9462) );
  OAI21_X1 U10349 ( .B1(n9463), .B2(n9530), .A(n9462), .ZN(P1_U3227) );
  XNOR2_X1 U10350 ( .A(n9465), .B(n9464), .ZN(n9466) );
  XNOR2_X1 U10351 ( .A(n9467), .B(n9466), .ZN(n9472) );
  NOR2_X1 U10352 ( .A1(n9526), .A2(n9765), .ZN(n9470) );
  AOI22_X1 U10353 ( .A1(n9523), .A2(n9720), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9468) );
  OAI21_X1 U10354 ( .B1(n9754), .B2(n9521), .A(n9468), .ZN(n9469) );
  AOI211_X1 U10355 ( .C1(n9885), .C2(n9528), .A(n9470), .B(n9469), .ZN(n9471)
         );
  OAI21_X1 U10356 ( .B1(n9472), .B2(n9530), .A(n9471), .ZN(P1_U3231) );
  INV_X1 U10357 ( .A(n9874), .ZN(n9482) );
  OAI21_X1 U10358 ( .B1(n9475), .B2(n9474), .A(n9473), .ZN(n9476) );
  NAND2_X1 U10359 ( .A1(n9476), .A2(n9485), .ZN(n9481) );
  INV_X1 U10360 ( .A(n9724), .ZN(n9479) );
  AOI22_X1 U10361 ( .A1(n9523), .A2(n9721), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9477) );
  OAI21_X1 U10362 ( .B1(n9755), .B2(n9521), .A(n9477), .ZN(n9478) );
  AOI21_X1 U10363 ( .B1(n9479), .B2(n9510), .A(n9478), .ZN(n9480) );
  OAI211_X1 U10364 ( .C1(n9482), .C2(n9513), .A(n9481), .B(n9480), .ZN(
        P1_U3233) );
  OAI21_X1 U10365 ( .B1(n6818), .B2(n9484), .A(n9483), .ZN(n9486) );
  NAND2_X1 U10366 ( .A1(n9486), .A2(n9485), .ZN(n9491) );
  AOI22_X1 U10367 ( .A1(n9487), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n9528), .B2(
        n10426), .ZN(n9490) );
  AOI22_X1 U10368 ( .A1(n9488), .A2(n9544), .B1(n9523), .B2(n6954), .ZN(n9489)
         );
  NAND3_X1 U10369 ( .A1(n9491), .A2(n9490), .A3(n9489), .ZN(P1_U3235) );
  NAND2_X1 U10370 ( .A1(n9493), .A2(n9492), .ZN(n9495) );
  XNOR2_X1 U10371 ( .A(n9495), .B(n9494), .ZN(n9501) );
  NOR2_X1 U10372 ( .A1(n9526), .A2(n9792), .ZN(n9499) );
  NAND2_X1 U10373 ( .A1(n9523), .A2(n9798), .ZN(n9496) );
  NAND2_X1 U10374 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9578) );
  OAI211_X1 U10375 ( .C1(n9497), .C2(n9521), .A(n9496), .B(n9578), .ZN(n9498)
         );
  AOI211_X1 U10376 ( .C1(n9895), .C2(n9528), .A(n9499), .B(n9498), .ZN(n9500)
         );
  OAI21_X1 U10377 ( .B1(n9501), .B2(n9530), .A(n9500), .ZN(P1_U3236) );
  AOI21_X1 U10378 ( .B1(n9502), .B2(n9503), .A(n9530), .ZN(n9505) );
  NAND2_X1 U10379 ( .A1(n9505), .A2(n9504), .ZN(n9512) );
  OAI22_X1 U10380 ( .A1(n9690), .A2(n9521), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9506), .ZN(n9509) );
  NOR2_X1 U10381 ( .A1(n9659), .A2(n9507), .ZN(n9508) );
  AOI211_X1 U10382 ( .C1(n9662), .C2(n9510), .A(n9509), .B(n9508), .ZN(n9511)
         );
  OAI211_X1 U10383 ( .C1(n9665), .C2(n9513), .A(n9512), .B(n9511), .ZN(
        P1_U3238) );
  INV_X1 U10384 ( .A(n9514), .ZN(n9516) );
  NAND2_X1 U10385 ( .A1(n9516), .A2(n9515), .ZN(n9518) );
  XNOR2_X1 U10386 ( .A(n9518), .B(n9517), .ZN(n9531) );
  OAI21_X1 U10387 ( .B1(n9521), .B2(n9520), .A(n9519), .ZN(n9522) );
  AOI21_X1 U10388 ( .B1(n9523), .B2(n9806), .A(n9522), .ZN(n9524) );
  OAI21_X1 U10389 ( .B1(n9526), .B2(n9525), .A(n9524), .ZN(n9527) );
  AOI21_X1 U10390 ( .B1(n9912), .B2(n9528), .A(n9527), .ZN(n9529) );
  OAI21_X1 U10391 ( .B1(n9531), .B2(n9530), .A(n9529), .ZN(P1_U3239) );
  MUX2_X1 U10392 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9608), .S(P1_U4006), .Z(
        P1_U3586) );
  MUX2_X1 U10393 ( .A(n9532), .B(P1_DATAO_REG_30__SCAN_IN), .S(n10340), .Z(
        P1_U3585) );
  MUX2_X1 U10394 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9677), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10395 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9533), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10396 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9710), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10397 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9721), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10398 ( .A(n9709), .B(P1_DATAO_REG_22__SCAN_IN), .S(n10340), .Z(
        P1_U3577) );
  MUX2_X1 U10399 ( .A(n9720), .B(P1_DATAO_REG_21__SCAN_IN), .S(n10340), .Z(
        P1_U3576) );
  MUX2_X1 U10400 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9534), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10401 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9798), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10402 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9535), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10403 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9799), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10404 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9806), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10405 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9536), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10406 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9537), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10407 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9538), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10408 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9539), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10409 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9540), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10410 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9541), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10411 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9542), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10412 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9543), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10413 ( .A(n6954), .B(P1_DATAO_REG_3__SCAN_IN), .S(n10340), .Z(
        P1_U3558) );
  MUX2_X1 U10414 ( .A(n6813), .B(P1_DATAO_REG_2__SCAN_IN), .S(n10340), .Z(
        P1_U3557) );
  MUX2_X1 U10415 ( .A(n9544), .B(P1_DATAO_REG_1__SCAN_IN), .S(n10340), .Z(
        P1_U3556) );
  MUX2_X1 U10416 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6676), .S(P1_U4006), .Z(
        P1_U3555) );
  NOR2_X1 U10417 ( .A1(n9553), .A2(n9546), .ZN(n9548) );
  NOR2_X1 U10418 ( .A1(n9548), .A2(n9547), .ZN(n9551) );
  NAND2_X1 U10419 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9570), .ZN(n9549) );
  OAI21_X1 U10420 ( .B1(n9570), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9549), .ZN(
        n9550) );
  NOR2_X1 U10421 ( .A1(n9551), .A2(n9550), .ZN(n9564) );
  AOI211_X1 U10422 ( .C1(n9551), .C2(n9550), .A(n9564), .B(n10370), .ZN(n9563)
         );
  NOR2_X1 U10423 ( .A1(n9553), .A2(n9552), .ZN(n9555) );
  NOR2_X1 U10424 ( .A1(n9555), .A2(n9554), .ZN(n9557) );
  XNOR2_X1 U10425 ( .A(n9570), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9556) );
  NOR2_X1 U10426 ( .A1(n9557), .A2(n9556), .ZN(n9569) );
  AOI211_X1 U10427 ( .C1(n9557), .C2(n9556), .A(n9569), .B(n10333), .ZN(n9562)
         );
  NAND2_X1 U10428 ( .A1(n10290), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9559) );
  OAI211_X1 U10429 ( .C1(n9560), .C2(n10364), .A(n9559), .B(n9558), .ZN(n9561)
         );
  OR3_X1 U10430 ( .A1(n9563), .A2(n9562), .A3(n9561), .ZN(P1_U3257) );
  INV_X1 U10431 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9577) );
  AOI21_X1 U10432 ( .B1(n9570), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9564), .ZN(
        n9567) );
  NAND2_X1 U10433 ( .A1(n9588), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9565) );
  OAI21_X1 U10434 ( .B1(n9588), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9565), .ZN(
        n9566) );
  NOR2_X1 U10435 ( .A1(n9567), .A2(n9566), .ZN(n9581) );
  AOI211_X1 U10436 ( .C1(n9567), .C2(n9566), .A(n9581), .B(n10370), .ZN(n9568)
         );
  AOI21_X1 U10437 ( .B1(n10288), .B2(n9588), .A(n9568), .ZN(n9576) );
  AOI21_X1 U10438 ( .B1(n9570), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9569), .ZN(
        n9572) );
  XNOR2_X1 U10439 ( .A(n9588), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9571) );
  NOR2_X1 U10440 ( .A1(n9572), .A2(n9571), .ZN(n9587) );
  AOI211_X1 U10441 ( .C1(n9572), .C2(n9571), .A(n9587), .B(n10333), .ZN(n9574)
         );
  NOR2_X1 U10442 ( .A1(n9574), .A2(n9573), .ZN(n9575) );
  OAI211_X1 U10443 ( .C1(n10376), .C2(n9577), .A(n9576), .B(n9575), .ZN(
        P1_U3258) );
  INV_X1 U10444 ( .A(n9598), .ZN(n9579) );
  OAI21_X1 U10445 ( .B1(n10364), .B2(n9579), .A(n9578), .ZN(n9585) );
  MUX2_X1 U10446 ( .A(P1_REG2_REG_18__SCAN_IN), .B(n8036), .S(n9598), .Z(n9580) );
  INV_X1 U10447 ( .A(n9580), .ZN(n9583) );
  AOI21_X1 U10448 ( .B1(n9588), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9581), .ZN(
        n9582) );
  NOR2_X1 U10449 ( .A1(n9582), .A2(n9583), .ZN(n9594) );
  AOI211_X1 U10450 ( .C1(n9583), .C2(n9582), .A(n9594), .B(n10370), .ZN(n9584)
         );
  AOI211_X1 U10451 ( .C1(n10290), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9585), .B(
        n9584), .ZN(n9593) );
  XNOR2_X1 U10452 ( .A(n9598), .B(n9586), .ZN(n9590) );
  AOI21_X1 U10453 ( .B1(n9588), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9587), .ZN(
        n9589) );
  NAND2_X1 U10454 ( .A1(n9589), .A2(n9590), .ZN(n9597) );
  OAI21_X1 U10455 ( .B1(n9590), .B2(n9589), .A(n9597), .ZN(n9591) );
  NAND2_X1 U10456 ( .A1(n9591), .A2(n10368), .ZN(n9592) );
  NAND2_X1 U10457 ( .A1(n9593), .A2(n9592), .ZN(P1_U3259) );
  AOI21_X1 U10458 ( .B1(n9598), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9594), .ZN(
        n9596) );
  XNOR2_X1 U10459 ( .A(n9781), .B(n9773), .ZN(n9595) );
  XNOR2_X1 U10460 ( .A(n9596), .B(n9595), .ZN(n9606) );
  OAI21_X1 U10461 ( .B1(n9598), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9597), .ZN(
        n9600) );
  XNOR2_X1 U10462 ( .A(n9781), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9599) );
  XNOR2_X1 U10463 ( .A(n9600), .B(n9599), .ZN(n9604) );
  NAND2_X1 U10464 ( .A1(n10290), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n9602) );
  OAI211_X1 U10465 ( .C1(n9781), .C2(n10364), .A(n9602), .B(n9601), .ZN(n9603)
         );
  AOI21_X1 U10466 ( .B1(n10368), .B2(n9604), .A(n9603), .ZN(n9605) );
  OAI21_X1 U10467 ( .B1(n9606), .B2(n10370), .A(n9605), .ZN(P1_U3260) );
  XNOR2_X1 U10468 ( .A(n9831), .B(n9611), .ZN(n9829) );
  NAND2_X1 U10469 ( .A1(n9829), .A2(n9825), .ZN(n9610) );
  NAND2_X1 U10470 ( .A1(n9608), .A2(n9607), .ZN(n9834) );
  NOR2_X1 U10471 ( .A1(n10425), .A2(n9834), .ZN(n9615) );
  AOI21_X1 U10472 ( .B1(n10425), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9615), .ZN(
        n9609) );
  OAI211_X1 U10473 ( .C1(n9831), .C2(n9818), .A(n9610), .B(n9609), .ZN(
        P1_U3261) );
  OAI21_X1 U10474 ( .B1(n9613), .B2(n9612), .A(n9611), .ZN(n9835) );
  NOR2_X1 U10475 ( .A1(n9822), .A2(n9614), .ZN(n9616) );
  AOI211_X1 U10476 ( .C1(n9832), .C2(n9785), .A(n9616), .B(n9615), .ZN(n9617)
         );
  OAI21_X1 U10477 ( .B1(n9835), .B2(n9728), .A(n9617), .ZN(P1_U3262) );
  NAND2_X1 U10478 ( .A1(n9618), .A2(n9624), .ZN(n9619) );
  NAND2_X1 U10479 ( .A1(n9620), .A2(n9619), .ZN(n9847) );
  AOI22_X1 U10480 ( .A1(n9622), .A2(n10393), .B1(n9621), .B2(n10392), .ZN(
        n9627) );
  OAI211_X1 U10481 ( .C1(n9625), .C2(n9624), .A(n9623), .B(n10397), .ZN(n9626)
         );
  OAI211_X1 U10482 ( .C1(n9847), .C2(n9836), .A(n9627), .B(n9626), .ZN(n9842)
         );
  OAI22_X1 U10483 ( .A1(n9629), .A2(n9819), .B1(n9628), .B2(n9822), .ZN(n9630)
         );
  AOI21_X1 U10484 ( .B1(n9843), .B2(n9785), .A(n9630), .ZN(n9634) );
  NAND2_X1 U10485 ( .A1(n9640), .A2(n9843), .ZN(n9631) );
  AND2_X1 U10486 ( .A1(n9632), .A2(n9631), .ZN(n9844) );
  NAND2_X1 U10487 ( .A1(n9844), .A2(n9825), .ZN(n9633) );
  OAI211_X1 U10488 ( .C1(n9847), .C2(n9635), .A(n9634), .B(n9633), .ZN(n9636)
         );
  AOI21_X1 U10489 ( .B1(n9842), .B2(n9822), .A(n9636), .ZN(n9637) );
  INV_X1 U10490 ( .A(n9637), .ZN(P1_U3263) );
  XOR2_X1 U10491 ( .A(n9639), .B(n9638), .Z(n9852) );
  INV_X1 U10492 ( .A(n9660), .ZN(n9642) );
  INV_X1 U10493 ( .A(n9640), .ZN(n9641) );
  AOI21_X1 U10494 ( .B1(n9848), .B2(n9642), .A(n9641), .ZN(n9849) );
  AOI22_X1 U10495 ( .A1(n9643), .A2(n10411), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n9684), .ZN(n9644) );
  OAI21_X1 U10496 ( .B1(n9645), .B2(n9818), .A(n9644), .ZN(n9653) );
  AOI21_X1 U10497 ( .B1(n4903), .B2(n9646), .A(n9811), .ZN(n9651) );
  OAI22_X1 U10498 ( .A1(n9648), .A2(n9808), .B1(n9647), .B2(n9779), .ZN(n9649)
         );
  AOI21_X1 U10499 ( .B1(n9651), .B2(n9650), .A(n9649), .ZN(n9851) );
  NOR2_X1 U10500 ( .A1(n9851), .A2(n10425), .ZN(n9652) );
  AOI211_X1 U10501 ( .C1(n9825), .C2(n9849), .A(n9653), .B(n9652), .ZN(n9654)
         );
  OAI21_X1 U10502 ( .B1(n9852), .B2(n9804), .A(n9654), .ZN(P1_U3264) );
  XOR2_X1 U10503 ( .A(n9657), .B(n9655), .Z(n9858) );
  INV_X1 U10504 ( .A(n9669), .ZN(n9661) );
  AOI21_X1 U10505 ( .B1(n9854), .B2(n9661), .A(n9660), .ZN(n9855) );
  NAND2_X1 U10506 ( .A1(n9855), .A2(n9825), .ZN(n9664) );
  AOI22_X1 U10507 ( .A1(n9662), .A2(n10411), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n9684), .ZN(n9663) );
  OAI211_X1 U10508 ( .C1(n9665), .C2(n9818), .A(n9664), .B(n9663), .ZN(n9666)
         );
  AOI21_X1 U10509 ( .B1(n9853), .B2(n9822), .A(n9666), .ZN(n9667) );
  OAI21_X1 U10510 ( .B1(n9858), .B2(n9804), .A(n9667), .ZN(P1_U3265) );
  XNOR2_X1 U10511 ( .A(n9668), .B(n9675), .ZN(n9863) );
  AOI21_X1 U10512 ( .B1(n9859), .B2(n9691), .A(n9669), .ZN(n9860) );
  INV_X1 U10513 ( .A(n9859), .ZN(n9673) );
  INV_X1 U10514 ( .A(n9670), .ZN(n9671) );
  AOI22_X1 U10515 ( .A1(n9671), .A2(n10411), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n9684), .ZN(n9672) );
  OAI21_X1 U10516 ( .B1(n9673), .B2(n9818), .A(n9672), .ZN(n9681) );
  OAI211_X1 U10517 ( .C1(n9676), .C2(n9675), .A(n9674), .B(n10397), .ZN(n9679)
         );
  AOI22_X1 U10518 ( .A1(n9677), .A2(n10392), .B1(n10393), .B2(n9710), .ZN(
        n9678) );
  AND2_X1 U10519 ( .A1(n9679), .A2(n9678), .ZN(n9862) );
  NOR2_X1 U10520 ( .A1(n9862), .A2(n10425), .ZN(n9680) );
  AOI211_X1 U10521 ( .C1(n9860), .C2(n9825), .A(n9681), .B(n9680), .ZN(n9682)
         );
  OAI21_X1 U10522 ( .B1(n9863), .B2(n9804), .A(n9682), .ZN(P1_U3266) );
  XOR2_X1 U10523 ( .A(n9686), .B(n9683), .Z(n9868) );
  AOI22_X1 U10524 ( .A1(n9866), .A2(n9785), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9684), .ZN(n9697) );
  OAI211_X1 U10525 ( .C1(n9687), .C2(n9686), .A(n9685), .B(n10397), .ZN(n9689)
         );
  NAND2_X1 U10526 ( .A1(n9721), .A2(n10393), .ZN(n9688) );
  OAI211_X1 U10527 ( .C1(n9690), .C2(n9808), .A(n9689), .B(n9688), .ZN(n9864)
         );
  AOI211_X1 U10528 ( .C1(n9866), .C2(n9699), .A(n10548), .B(n5138), .ZN(n9865)
         );
  INV_X1 U10529 ( .A(n9865), .ZN(n9694) );
  INV_X1 U10530 ( .A(n9692), .ZN(n9693) );
  OAI22_X1 U10531 ( .A1(n9694), .A2(n10415), .B1(n9693), .B2(n9819), .ZN(n9695) );
  OAI21_X1 U10532 ( .B1(n9864), .B2(n9695), .A(n9822), .ZN(n9696) );
  OAI211_X1 U10533 ( .C1(n9868), .C2(n9804), .A(n9697), .B(n9696), .ZN(
        P1_U3267) );
  XNOR2_X1 U10534 ( .A(n9698), .B(n9707), .ZN(n9873) );
  INV_X1 U10535 ( .A(n9726), .ZN(n9701) );
  INV_X1 U10536 ( .A(n9699), .ZN(n9700) );
  AOI21_X1 U10537 ( .B1(n9869), .B2(n9701), .A(n9700), .ZN(n9870) );
  INV_X1 U10538 ( .A(n9702), .ZN(n9703) );
  AOI22_X1 U10539 ( .A1(n10425), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9703), 
        .B2(n10411), .ZN(n9704) );
  OAI21_X1 U10540 ( .B1(n9705), .B2(n9818), .A(n9704), .ZN(n9714) );
  OAI211_X1 U10541 ( .C1(n9708), .C2(n9707), .A(n9706), .B(n10397), .ZN(n9712)
         );
  AOI22_X1 U10542 ( .A1(n9710), .A2(n10392), .B1(n10393), .B2(n9709), .ZN(
        n9711) );
  AND2_X1 U10543 ( .A1(n9712), .A2(n9711), .ZN(n9872) );
  NOR2_X1 U10544 ( .A1(n9872), .A2(n10425), .ZN(n9713) );
  AOI211_X1 U10545 ( .C1(n9870), .C2(n9825), .A(n9714), .B(n9713), .ZN(n9715)
         );
  OAI21_X1 U10546 ( .B1(n9873), .B2(n9804), .A(n9715), .ZN(P1_U3268) );
  XOR2_X1 U10547 ( .A(n9718), .B(n9716), .Z(n9878) );
  OAI211_X1 U10548 ( .C1(n9719), .C2(n9718), .A(n9717), .B(n10397), .ZN(n9723)
         );
  AOI22_X1 U10549 ( .A1(n9721), .A2(n10392), .B1(n10393), .B2(n9720), .ZN(
        n9722) );
  AND2_X1 U10550 ( .A1(n9723), .A2(n9722), .ZN(n9877) );
  OAI21_X1 U10551 ( .B1(n9724), .B2(n9819), .A(n9877), .ZN(n9731) );
  AND2_X1 U10552 ( .A1(n9874), .A2(n9744), .ZN(n9725) );
  NOR2_X1 U10553 ( .A1(n9726), .A2(n9725), .ZN(n9875) );
  INV_X1 U10554 ( .A(n9875), .ZN(n9729) );
  AOI22_X1 U10555 ( .A1(n9874), .A2(n9785), .B1(n10425), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9727) );
  OAI21_X1 U10556 ( .B1(n9729), .B2(n9728), .A(n9727), .ZN(n9730) );
  AOI21_X1 U10557 ( .B1(n9731), .B2(n9822), .A(n9730), .ZN(n9732) );
  OAI21_X1 U10558 ( .B1(n9878), .B2(n9804), .A(n9732), .ZN(P1_U3269) );
  NAND2_X1 U10559 ( .A1(n9734), .A2(n9733), .ZN(n9753) );
  NAND2_X1 U10560 ( .A1(n9753), .A2(n9760), .ZN(n9736) );
  NAND2_X1 U10561 ( .A1(n9736), .A2(n9735), .ZN(n9737) );
  XNOR2_X1 U10562 ( .A(n9740), .B(n9737), .ZN(n9883) );
  NAND2_X1 U10563 ( .A1(n9757), .A2(n9738), .ZN(n9739) );
  XOR2_X1 U10564 ( .A(n9740), .B(n9739), .Z(n9741) );
  OAI222_X1 U10565 ( .A1(n9808), .A2(n9742), .B1(n9779), .B2(n9780), .C1(n9811), .C2(n9741), .ZN(n9879) );
  INV_X1 U10566 ( .A(n9744), .ZN(n9745) );
  AOI211_X1 U10567 ( .C1(n9881), .C2(n9763), .A(n10548), .B(n9745), .ZN(n9880)
         );
  INV_X1 U10568 ( .A(n9880), .ZN(n9748) );
  INV_X1 U10569 ( .A(n9746), .ZN(n9747) );
  OAI22_X1 U10570 ( .A1(n9748), .A2(n10415), .B1(n9747), .B2(n9819), .ZN(n9749) );
  OAI21_X1 U10571 ( .B1(n9879), .B2(n9749), .A(n9822), .ZN(n9751) );
  AOI22_X1 U10572 ( .A1(n9881), .A2(n9785), .B1(n10425), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9750) );
  OAI211_X1 U10573 ( .C1(n9883), .C2(n9804), .A(n9751), .B(n9750), .ZN(
        P1_U3270) );
  XNOR2_X1 U10574 ( .A(n9753), .B(n9752), .ZN(n9884) );
  OAI22_X1 U10575 ( .A1(n9755), .A2(n9808), .B1(n9754), .B2(n9779), .ZN(n9762)
         );
  INV_X1 U10576 ( .A(n9756), .ZN(n9759) );
  INV_X1 U10577 ( .A(n9757), .ZN(n9758) );
  AOI211_X1 U10578 ( .C1(n9760), .C2(n9759), .A(n9811), .B(n9758), .ZN(n9761)
         );
  AOI211_X1 U10579 ( .C1(n9884), .C2(n9816), .A(n9762), .B(n9761), .ZN(n9888)
         );
  AOI21_X1 U10580 ( .B1(n9885), .B2(n9774), .A(n9743), .ZN(n9886) );
  INV_X1 U10581 ( .A(n9885), .ZN(n9764) );
  NOR2_X1 U10582 ( .A1(n9764), .A2(n9818), .ZN(n9768) );
  OAI22_X1 U10583 ( .A1(n9822), .A2(n9766), .B1(n9765), .B2(n9819), .ZN(n9767)
         );
  AOI211_X1 U10584 ( .C1(n9886), .C2(n9825), .A(n9768), .B(n9767), .ZN(n9770)
         );
  NAND2_X1 U10585 ( .A1(n9884), .A2(n9826), .ZN(n9769) );
  OAI211_X1 U10586 ( .C1(n9888), .C2(n10425), .A(n9770), .B(n9769), .ZN(
        P1_U3271) );
  XOR2_X1 U10587 ( .A(n9771), .B(n9777), .Z(n9894) );
  OAI22_X1 U10588 ( .A1(n9822), .A2(n9773), .B1(n9772), .B2(n9819), .ZN(n9784)
         );
  INV_X1 U10589 ( .A(n9774), .ZN(n9775) );
  AOI211_X1 U10590 ( .C1(n9892), .C2(n9790), .A(n10548), .B(n9775), .ZN(n9891)
         );
  XOR2_X1 U10591 ( .A(n9777), .B(n9776), .Z(n9778) );
  OAI222_X1 U10592 ( .A1(n9808), .A2(n9780), .B1(n9779), .B2(n9809), .C1(n9778), .C2(n9811), .ZN(n9890) );
  AOI21_X1 U10593 ( .B1(n9891), .B2(n9781), .A(n9890), .ZN(n9782) );
  NOR2_X1 U10594 ( .A1(n9782), .A2(n10425), .ZN(n9783) );
  AOI211_X1 U10595 ( .C1(n9785), .C2(n9892), .A(n9784), .B(n9783), .ZN(n9786)
         );
  OAI21_X1 U10596 ( .B1(n9804), .B2(n9894), .A(n9786), .ZN(P1_U3272) );
  OAI21_X1 U10597 ( .B1(n9789), .B2(n9788), .A(n9787), .ZN(n9899) );
  INV_X1 U10598 ( .A(n9790), .ZN(n9791) );
  AOI21_X1 U10599 ( .B1(n9895), .B2(n5142), .A(n9791), .ZN(n9896) );
  INV_X1 U10600 ( .A(n9792), .ZN(n9793) );
  AOI22_X1 U10601 ( .A1(n10425), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9793), 
        .B2(n10411), .ZN(n9794) );
  OAI21_X1 U10602 ( .B1(n9795), .B2(n9818), .A(n9794), .ZN(n9802) );
  OAI21_X1 U10603 ( .B1(n9797), .B2(n4939), .A(n9796), .ZN(n9800) );
  AOI222_X1 U10604 ( .A1(n10397), .A2(n9800), .B1(n9799), .B2(n10393), .C1(
        n9798), .C2(n10392), .ZN(n9898) );
  NOR2_X1 U10605 ( .A1(n9898), .A2(n10425), .ZN(n9801) );
  AOI211_X1 U10606 ( .C1(n9896), .C2(n9825), .A(n9802), .B(n9801), .ZN(n9803)
         );
  OAI21_X1 U10607 ( .B1(n9804), .B2(n9899), .A(n9803), .ZN(P1_U3273) );
  OAI21_X1 U10608 ( .B1(n5457), .B2(n9812), .A(n9805), .ZN(n9900) );
  NAND2_X1 U10609 ( .A1(n9806), .A2(n10393), .ZN(n9807) );
  OAI21_X1 U10610 ( .B1(n9809), .B2(n9808), .A(n9807), .ZN(n9815) );
  AOI211_X1 U10611 ( .C1(n9813), .C2(n9812), .A(n9811), .B(n9810), .ZN(n9814)
         );
  AOI211_X1 U10612 ( .C1(n9816), .C2(n9900), .A(n9815), .B(n9814), .ZN(n9904)
         );
  AOI21_X1 U10613 ( .B1(n9901), .B2(n9817), .A(n4863), .ZN(n9902) );
  NOR2_X1 U10614 ( .A1(n5140), .A2(n9818), .ZN(n9824) );
  OAI22_X1 U10615 ( .A1(n9822), .A2(n9821), .B1(n9820), .B2(n9819), .ZN(n9823)
         );
  AOI211_X1 U10616 ( .C1(n9902), .C2(n9825), .A(n9824), .B(n9823), .ZN(n9828)
         );
  NAND2_X1 U10617 ( .A1(n9900), .A2(n9826), .ZN(n9827) );
  OAI211_X1 U10618 ( .C1(n9904), .C2(n10425), .A(n9828), .B(n9827), .ZN(
        P1_U3274) );
  NAND2_X1 U10619 ( .A1(n9829), .A2(n10482), .ZN(n9830) );
  OAI211_X1 U10620 ( .C1(n9831), .C2(n10637), .A(n9830), .B(n9834), .ZN(n9930)
         );
  MUX2_X1 U10621 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9930), .S(n10644), .Z(
        P1_U3554) );
  NAND2_X1 U10622 ( .A1(n9832), .A2(n10501), .ZN(n9833) );
  OAI211_X1 U10623 ( .C1(n9835), .C2(n10548), .A(n9834), .B(n9833), .ZN(n9931)
         );
  INV_X2 U10624 ( .A(n10642), .ZN(n10644) );
  MUX2_X1 U10625 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9931), .S(n10644), .Z(
        P1_U3553) );
  AOI22_X1 U10626 ( .A1(n9838), .A2(n10482), .B1(n10501), .B2(n9837), .ZN(
        n9839) );
  INV_X1 U10627 ( .A(n9842), .ZN(n9846) );
  AOI22_X1 U10628 ( .A1(n9844), .A2(n10482), .B1(n10501), .B2(n9843), .ZN(
        n9845) );
  OAI211_X1 U10629 ( .C1(n10504), .C2(n9847), .A(n9846), .B(n9845), .ZN(n9932)
         );
  MUX2_X1 U10630 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9932), .S(n10644), .Z(
        P1_U3551) );
  AOI22_X1 U10631 ( .A1(n9849), .A2(n10482), .B1(n10501), .B2(n9848), .ZN(
        n9850) );
  OAI211_X1 U10632 ( .C1(n9852), .C2(n10406), .A(n9851), .B(n9850), .ZN(n9933)
         );
  MUX2_X1 U10633 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9933), .S(n10644), .Z(
        P1_U3550) );
  INV_X1 U10634 ( .A(n9853), .ZN(n9857) );
  AOI22_X1 U10635 ( .A1(n9855), .A2(n10482), .B1(n10501), .B2(n9854), .ZN(
        n9856) );
  OAI211_X1 U10636 ( .C1(n10406), .C2(n9858), .A(n9857), .B(n9856), .ZN(n9934)
         );
  MUX2_X1 U10637 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9934), .S(n10644), .Z(
        P1_U3549) );
  AOI22_X1 U10638 ( .A1(n9860), .A2(n10482), .B1(n10501), .B2(n9859), .ZN(
        n9861) );
  OAI211_X1 U10639 ( .C1(n9863), .C2(n10406), .A(n9862), .B(n9861), .ZN(n9935)
         );
  MUX2_X1 U10640 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9935), .S(n10644), .Z(
        P1_U3548) );
  AOI211_X1 U10641 ( .C1(n10501), .C2(n9866), .A(n9865), .B(n9864), .ZN(n9867)
         );
  OAI21_X1 U10642 ( .B1(n9868), .B2(n10406), .A(n9867), .ZN(n9936) );
  MUX2_X1 U10643 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9936), .S(n10644), .Z(
        P1_U3547) );
  AOI22_X1 U10644 ( .A1(n9870), .A2(n10482), .B1(n10501), .B2(n9869), .ZN(
        n9871) );
  OAI211_X1 U10645 ( .C1(n9873), .C2(n10406), .A(n9872), .B(n9871), .ZN(n9937)
         );
  MUX2_X1 U10646 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9937), .S(n10644), .Z(
        P1_U3546) );
  AOI22_X1 U10647 ( .A1(n9875), .A2(n10482), .B1(n10501), .B2(n9874), .ZN(
        n9876) );
  OAI211_X1 U10648 ( .C1(n9878), .C2(n10406), .A(n9877), .B(n9876), .ZN(n9938)
         );
  MUX2_X1 U10649 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9938), .S(n10644), .Z(
        P1_U3545) );
  AOI211_X1 U10650 ( .C1(n10501), .C2(n9881), .A(n9880), .B(n9879), .ZN(n9882)
         );
  OAI21_X1 U10651 ( .B1(n10406), .B2(n9883), .A(n9882), .ZN(n9939) );
  MUX2_X1 U10652 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9939), .S(n10644), .Z(
        P1_U3544) );
  INV_X1 U10653 ( .A(n9884), .ZN(n9889) );
  AOI22_X1 U10654 ( .A1(n9886), .A2(n10482), .B1(n10501), .B2(n9885), .ZN(
        n9887) );
  OAI211_X1 U10655 ( .C1(n10504), .C2(n9889), .A(n9888), .B(n9887), .ZN(n9940)
         );
  MUX2_X1 U10656 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9940), .S(n10644), .Z(
        P1_U3543) );
  AOI211_X1 U10657 ( .C1(n10501), .C2(n9892), .A(n9891), .B(n9890), .ZN(n9893)
         );
  OAI21_X1 U10658 ( .B1(n10406), .B2(n9894), .A(n9893), .ZN(n9941) );
  MUX2_X1 U10659 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9941), .S(n10644), .Z(
        P1_U3542) );
  AOI22_X1 U10660 ( .A1(n9896), .A2(n10482), .B1(n10501), .B2(n9895), .ZN(
        n9897) );
  OAI211_X1 U10661 ( .C1(n10406), .C2(n9899), .A(n9898), .B(n9897), .ZN(n9942)
         );
  MUX2_X1 U10662 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9942), .S(n10644), .Z(
        P1_U3541) );
  INV_X1 U10663 ( .A(n9900), .ZN(n9905) );
  AOI22_X1 U10664 ( .A1(n9902), .A2(n10482), .B1(n10501), .B2(n9901), .ZN(
        n9903) );
  OAI211_X1 U10665 ( .C1(n9905), .C2(n10504), .A(n9904), .B(n9903), .ZN(n9943)
         );
  MUX2_X1 U10666 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9943), .S(n10644), .Z(
        P1_U3540) );
  AOI211_X1 U10667 ( .C1(n10501), .C2(n9908), .A(n9907), .B(n9906), .ZN(n9909)
         );
  OAI21_X1 U10668 ( .B1(n10406), .B2(n9910), .A(n9909), .ZN(n9944) );
  MUX2_X1 U10669 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9944), .S(n10644), .Z(
        P1_U3539) );
  INV_X1 U10670 ( .A(n9911), .ZN(n9916) );
  AOI22_X1 U10671 ( .A1(n9913), .A2(n10482), .B1(n10501), .B2(n9912), .ZN(
        n9914) );
  OAI211_X1 U10672 ( .C1(n10504), .C2(n9916), .A(n9915), .B(n9914), .ZN(n9945)
         );
  MUX2_X1 U10673 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9945), .S(n10644), .Z(
        P1_U3538) );
  INV_X1 U10674 ( .A(n10504), .ZN(n10617) );
  INV_X1 U10675 ( .A(n9917), .ZN(n9918) );
  OAI22_X1 U10676 ( .A1(n9919), .A2(n10548), .B1(n9918), .B2(n10637), .ZN(
        n9920) );
  AOI21_X1 U10677 ( .B1(n9921), .B2(n10617), .A(n9920), .ZN(n9922) );
  NAND2_X1 U10678 ( .A1(n9923), .A2(n9922), .ZN(n9946) );
  MUX2_X1 U10679 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9946), .S(n10644), .Z(
        P1_U3536) );
  INV_X1 U10680 ( .A(n9924), .ZN(n9929) );
  AOI22_X1 U10681 ( .A1(n9926), .A2(n10482), .B1(n10501), .B2(n9925), .ZN(
        n9927) );
  OAI211_X1 U10682 ( .C1(n9929), .C2(n10504), .A(n9928), .B(n9927), .ZN(n9947)
         );
  MUX2_X1 U10683 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9947), .S(n10644), .Z(
        P1_U3534) );
  MUX2_X1 U10684 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9930), .S(n10491), .Z(
        P1_U3522) );
  MUX2_X1 U10685 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9931), .S(n10491), .Z(
        P1_U3521) );
  MUX2_X1 U10686 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9932), .S(n10491), .Z(
        P1_U3519) );
  MUX2_X1 U10687 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9933), .S(n10491), .Z(
        P1_U3518) );
  MUX2_X1 U10688 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9934), .S(n10491), .Z(
        P1_U3517) );
  MUX2_X1 U10689 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9935), .S(n10491), .Z(
        P1_U3516) );
  MUX2_X1 U10690 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9936), .S(n10491), .Z(
        P1_U3515) );
  MUX2_X1 U10691 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9937), .S(n10491), .Z(
        P1_U3514) );
  MUX2_X1 U10692 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9938), .S(n10491), .Z(
        P1_U3513) );
  MUX2_X1 U10693 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9939), .S(n10491), .Z(
        P1_U3512) );
  MUX2_X1 U10694 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9940), .S(n10491), .Z(
        P1_U3511) );
  MUX2_X1 U10695 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9941), .S(n10491), .Z(
        P1_U3510) );
  MUX2_X1 U10696 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9942), .S(n10491), .Z(
        P1_U3508) );
  MUX2_X1 U10697 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9943), .S(n10491), .Z(
        P1_U3505) );
  MUX2_X1 U10698 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9944), .S(n10491), .Z(
        P1_U3502) );
  MUX2_X1 U10699 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9945), .S(n10491), .Z(
        P1_U3499) );
  MUX2_X1 U10700 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9946), .S(n10491), .Z(
        P1_U3493) );
  MUX2_X1 U10701 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n9947), .S(n10491), .Z(
        P1_U3487) );
  MUX2_X1 U10702 ( .A(n9948), .B(P1_D_REG_0__SCAN_IN), .S(n9967), .Z(P1_U3440)
         );
  NAND3_X1 U10703 ( .A1(n9950), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n9952) );
  OAI22_X1 U10704 ( .A1(n9949), .A2(n9952), .B1(n9951), .B2(n9961), .ZN(n9953)
         );
  AOI21_X1 U10705 ( .B1(n9955), .B2(n9954), .A(n9953), .ZN(n9956) );
  INV_X1 U10706 ( .A(n9956), .ZN(P1_U3322) );
  AOI21_X1 U10707 ( .B1(n9958), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n9957), .ZN(
        n9959) );
  OAI21_X1 U10708 ( .B1(n9960), .B2(n8830), .A(n9959), .ZN(P1_U3326) );
  OAI222_X1 U10709 ( .A1(P1_U3084), .A2(n9964), .B1(n8830), .B2(n9963), .C1(
        n9962), .C2(n9961), .ZN(P1_U3327) );
  INV_X1 U10710 ( .A(n9965), .ZN(n9966) );
  MUX2_X1 U10711 ( .A(n9966), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AND2_X1 U10712 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9967), .ZN(P1_U3321) );
  AND2_X1 U10713 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9967), .ZN(P1_U3320) );
  AND2_X1 U10714 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9967), .ZN(P1_U3319) );
  AND2_X1 U10715 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9967), .ZN(P1_U3318) );
  AND2_X1 U10716 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9967), .ZN(P1_U3317) );
  AND2_X1 U10717 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9967), .ZN(P1_U3316) );
  AND2_X1 U10718 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9967), .ZN(P1_U3315) );
  AND2_X1 U10719 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9967), .ZN(P1_U3314) );
  AND2_X1 U10720 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9967), .ZN(P1_U3313) );
  AND2_X1 U10721 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9967), .ZN(P1_U3312) );
  AND2_X1 U10722 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9967), .ZN(P1_U3311) );
  AND2_X1 U10723 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9967), .ZN(P1_U3310) );
  AND2_X1 U10724 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9967), .ZN(P1_U3309) );
  AND2_X1 U10725 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9967), .ZN(P1_U3308) );
  AND2_X1 U10726 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9967), .ZN(P1_U3307) );
  AND2_X1 U10727 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9967), .ZN(P1_U3306) );
  AND2_X1 U10728 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9967), .ZN(P1_U3305) );
  AND2_X1 U10729 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9967), .ZN(P1_U3304) );
  AND2_X1 U10730 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9967), .ZN(P1_U3303) );
  AND2_X1 U10731 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9967), .ZN(P1_U3302) );
  AND2_X1 U10732 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9967), .ZN(P1_U3301) );
  AND2_X1 U10733 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9967), .ZN(P1_U3300) );
  AND2_X1 U10734 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9967), .ZN(P1_U3299) );
  AND2_X1 U10735 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9967), .ZN(P1_U3298) );
  AND2_X1 U10736 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9967), .ZN(P1_U3297) );
  AND2_X1 U10737 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9967), .ZN(P1_U3296) );
  AND2_X1 U10738 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9967), .ZN(P1_U3295) );
  AND2_X1 U10739 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9967), .ZN(P1_U3294) );
  AND2_X1 U10740 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9967), .ZN(P1_U3293) );
  AND2_X1 U10741 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9967), .ZN(P1_U3292) );
  INV_X1 U10742 ( .A(n9968), .ZN(n9972) );
  INV_X1 U10743 ( .A(n9969), .ZN(n9970) );
  AOI22_X1 U10744 ( .A1(n10300), .A2(n9972), .B1(n6079), .B2(n4857), .ZN(
        P2_U3438) );
  AND2_X1 U10745 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n4857), .ZN(P2_U3326) );
  AND2_X1 U10746 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n4857), .ZN(P2_U3325) );
  AND2_X1 U10747 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n4857), .ZN(P2_U3323) );
  AND2_X1 U10748 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n4857), .ZN(P2_U3322) );
  AND2_X1 U10749 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n4857), .ZN(P2_U3321) );
  AND2_X1 U10750 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n4857), .ZN(P2_U3320) );
  AND2_X1 U10751 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n4857), .ZN(P2_U3319) );
  AND2_X1 U10752 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n4857), .ZN(P2_U3318) );
  AND2_X1 U10753 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n4857), .ZN(P2_U3317) );
  AND2_X1 U10754 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n4857), .ZN(P2_U3316) );
  AND2_X1 U10755 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n4857), .ZN(P2_U3315) );
  AND2_X1 U10756 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n4857), .ZN(P2_U3314) );
  AND2_X1 U10757 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n4857), .ZN(P2_U3313) );
  AND2_X1 U10758 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n4857), .ZN(P2_U3312) );
  AND2_X1 U10759 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n4857), .ZN(P2_U3311) );
  AND2_X1 U10760 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n4857), .ZN(P2_U3310) );
  AND2_X1 U10761 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n4857), .ZN(P2_U3309) );
  AND2_X1 U10762 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n4857), .ZN(P2_U3308) );
  AND2_X1 U10763 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n4857), .ZN(P2_U3307) );
  AND2_X1 U10764 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n4857), .ZN(P2_U3306) );
  AND2_X1 U10765 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n4857), .ZN(P2_U3305) );
  AND2_X1 U10766 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n4857), .ZN(P2_U3304) );
  AND2_X1 U10767 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n4857), .ZN(P2_U3303) );
  AND2_X1 U10768 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n4857), .ZN(P2_U3302) );
  AND2_X1 U10769 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n4857), .ZN(P2_U3301) );
  AND2_X1 U10770 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n4857), .ZN(P2_U3300) );
  AND2_X1 U10771 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n4857), .ZN(P2_U3299) );
  AND2_X1 U10772 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n4857), .ZN(P2_U3298) );
  AND2_X1 U10773 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n4857), .ZN(P2_U3297) );
  NAND2_X1 U10774 ( .A1(n4857), .A2(P2_D_REG_4__SCAN_IN), .ZN(n10202) );
  AOI22_X1 U10775 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_62), .B1(n5595), 
        .B2(keyinput_61), .ZN(n9974) );
  OAI221_X1 U10776 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_62), .C1(n5595), .C2(keyinput_61), .A(n9974), .ZN(n10075) );
  AOI22_X1 U10777 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_59), .B1(n10078), 
        .B2(keyinput_58), .ZN(n9975) );
  OAI221_X1 U10778 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_59), .C1(n10078), .C2(keyinput_58), .A(n9975), .ZN(n10072) );
  INV_X1 U10779 ( .A(keyinput_57), .ZN(n10070) );
  INV_X1 U10780 ( .A(keyinput_56), .ZN(n10068) );
  AOI22_X1 U10781 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_54), .B1(n5740), 
        .B2(keyinput_53), .ZN(n9976) );
  OAI221_X1 U10782 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_54), .C1(n5740), 
        .C2(keyinput_53), .A(n9976), .ZN(n10065) );
  INV_X1 U10783 ( .A(keyinput_52), .ZN(n10063) );
  OAI22_X1 U10784 ( .A1(n10181), .A2(keyinput_49), .B1(keyinput_50), .B2(
        P2_REG3_REG_17__SCAN_IN), .ZN(n9977) );
  AOI221_X1 U10785 ( .B1(n10181), .B2(keyinput_49), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput_50), .A(n9977), .ZN(n10060) );
  OAI22_X1 U10786 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_46), .B1(
        P2_REG3_REG_25__SCAN_IN), .B2(keyinput_47), .ZN(n9978) );
  AOI221_X1 U10787 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_46), .C1(
        keyinput_47), .C2(P2_REG3_REG_25__SCAN_IN), .A(n9978), .ZN(n10057) );
  INV_X1 U10788 ( .A(keyinput_45), .ZN(n10055) );
  OAI22_X1 U10789 ( .A1(n5666), .A2(keyinput_40), .B1(keyinput_42), .B2(
        P2_REG3_REG_28__SCAN_IN), .ZN(n9979) );
  AOI221_X1 U10790 ( .B1(n5666), .B2(keyinput_40), .C1(P2_REG3_REG_28__SCAN_IN), .C2(keyinput_42), .A(n9979), .ZN(n10053) );
  INV_X1 U10791 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9981) );
  OAI22_X1 U10792 ( .A1(n9981), .A2(keyinput_43), .B1(keyinput_39), .B2(
        P2_REG3_REG_10__SCAN_IN), .ZN(n9980) );
  AOI221_X1 U10793 ( .B1(n9981), .B2(keyinput_43), .C1(P2_REG3_REG_10__SCAN_IN), .C2(keyinput_39), .A(n9980), .ZN(n10052) );
  OAI22_X1 U10794 ( .A1(n5902), .A2(keyinput_41), .B1(n9983), .B2(keyinput_44), 
        .ZN(n9982) );
  AOI221_X1 U10795 ( .B1(n5902), .B2(keyinput_41), .C1(keyinput_44), .C2(n9983), .A(n9982), .ZN(n10051) );
  INV_X1 U10796 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10515) );
  AOI22_X1 U10797 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput_33), .B1(n10515), 
        .B2(keyinput_35), .ZN(n9984) );
  OAI221_X1 U10798 ( .B1(P2_RD_REG_SCAN_IN), .B2(keyinput_33), .C1(n10515), 
        .C2(keyinput_35), .A(n9984), .ZN(n9988) );
  AOI22_X1 U10799 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_34), .B1(n9986), 
        .B2(keyinput_36), .ZN(n9985) );
  OAI221_X1 U10800 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_34), .C1(n9986), 
        .C2(keyinput_36), .A(n9985), .ZN(n9987) );
  AOI211_X1 U10801 ( .C1(keyinput_37), .C2(P2_REG3_REG_14__SCAN_IN), .A(n9988), 
        .B(n9987), .ZN(n9989) );
  OAI21_X1 U10802 ( .B1(keyinput_37), .B2(P2_REG3_REG_14__SCAN_IN), .A(n9989), 
        .ZN(n10049) );
  INV_X1 U10803 ( .A(keyinput_31), .ZN(n9990) );
  MUX2_X1 U10804 ( .A(keyinput_31), .B(n9990), .S(SI_1_), .Z(n9991) );
  INV_X1 U10805 ( .A(n9991), .ZN(n10046) );
  INV_X1 U10806 ( .A(keyinput_29), .ZN(n10040) );
  INV_X1 U10807 ( .A(keyinput_24), .ZN(n10032) );
  AOI22_X1 U10808 ( .A1(SI_11_), .A2(keyinput_21), .B1(n9993), .B2(keyinput_22), .ZN(n9992) );
  OAI221_X1 U10809 ( .B1(SI_11_), .B2(keyinput_21), .C1(n9993), .C2(
        keyinput_22), .A(n9992), .ZN(n10029) );
  OAI22_X1 U10810 ( .A1(SI_16_), .A2(keyinput_16), .B1(keyinput_17), .B2(
        SI_15_), .ZN(n9994) );
  AOI221_X1 U10811 ( .B1(SI_16_), .B2(keyinput_16), .C1(SI_15_), .C2(
        keyinput_17), .A(n9994), .ZN(n10027) );
  OAI22_X1 U10812 ( .A1(n9996), .A2(keyinput_13), .B1(n10099), .B2(keyinput_14), .ZN(n9995) );
  AOI221_X1 U10813 ( .B1(n9996), .B2(keyinput_13), .C1(keyinput_14), .C2(
        n10099), .A(n9995), .ZN(n10019) );
  INV_X1 U10814 ( .A(keyinput_12), .ZN(n10017) );
  INV_X1 U10815 ( .A(keyinput_11), .ZN(n10015) );
  INV_X1 U10816 ( .A(SI_21_), .ZN(n10124) );
  INV_X1 U10817 ( .A(keyinput_10), .ZN(n10013) );
  INV_X1 U10818 ( .A(keyinput_9), .ZN(n10011) );
  INV_X1 U10819 ( .A(keyinput_8), .ZN(n10009) );
  INV_X1 U10820 ( .A(keyinput_7), .ZN(n10007) );
  INV_X1 U10821 ( .A(keyinput_6), .ZN(n10005) );
  OAI22_X1 U10822 ( .A1(SI_31_), .A2(keyinput_1), .B1(P2_WR_REG_SCAN_IN), .B2(
        keyinput_0), .ZN(n9997) );
  AOI221_X1 U10823 ( .B1(SI_31_), .B2(keyinput_1), .C1(keyinput_0), .C2(
        P2_WR_REG_SCAN_IN), .A(n9997), .ZN(n10003) );
  AOI22_X1 U10824 ( .A1(SI_30_), .A2(keyinput_2), .B1(n10102), .B2(keyinput_3), 
        .ZN(n9998) );
  OAI221_X1 U10825 ( .B1(SI_30_), .B2(keyinput_2), .C1(n10102), .C2(keyinput_3), .A(n9998), .ZN(n10002) );
  OAI22_X1 U10826 ( .A1(n10000), .A2(keyinput_5), .B1(keyinput_4), .B2(SI_28_), 
        .ZN(n9999) );
  AOI221_X1 U10827 ( .B1(n10000), .B2(keyinput_5), .C1(SI_28_), .C2(keyinput_4), .A(n9999), .ZN(n10001) );
  OAI21_X1 U10828 ( .B1(n10003), .B2(n10002), .A(n10001), .ZN(n10004) );
  OAI221_X1 U10829 ( .B1(SI_26_), .B2(n10005), .C1(n10109), .C2(keyinput_6), 
        .A(n10004), .ZN(n10006) );
  OAI221_X1 U10830 ( .B1(SI_25_), .B2(keyinput_7), .C1(n10113), .C2(n10007), 
        .A(n10006), .ZN(n10008) );
  OAI221_X1 U10831 ( .B1(SI_24_), .B2(keyinput_8), .C1(n10116), .C2(n10009), 
        .A(n10008), .ZN(n10010) );
  OAI221_X1 U10832 ( .B1(SI_23_), .B2(keyinput_9), .C1(n10118), .C2(n10011), 
        .A(n10010), .ZN(n10012) );
  OAI221_X1 U10833 ( .B1(SI_22_), .B2(keyinput_10), .C1(n10122), .C2(n10013), 
        .A(n10012), .ZN(n10014) );
  OAI221_X1 U10834 ( .B1(SI_21_), .B2(n10015), .C1(n10124), .C2(keyinput_11), 
        .A(n10014), .ZN(n10016) );
  OAI221_X1 U10835 ( .B1(SI_20_), .B2(n10017), .C1(n10127), .C2(keyinput_12), 
        .A(n10016), .ZN(n10018) );
  AOI22_X1 U10836 ( .A1(keyinput_15), .A2(n10021), .B1(n10019), .B2(n10018), 
        .ZN(n10020) );
  OAI21_X1 U10837 ( .B1(n10021), .B2(keyinput_15), .A(n10020), .ZN(n10026) );
  XOR2_X1 U10838 ( .A(keyinput_18), .B(SI_14_), .Z(n10025) );
  INV_X1 U10839 ( .A(SI_12_), .ZN(n10023) );
  AOI22_X1 U10840 ( .A1(SI_13_), .A2(keyinput_19), .B1(n10023), .B2(
        keyinput_20), .ZN(n10022) );
  OAI221_X1 U10841 ( .B1(SI_13_), .B2(keyinput_19), .C1(n10023), .C2(
        keyinput_20), .A(n10022), .ZN(n10024) );
  AOI211_X1 U10842 ( .C1(n10027), .C2(n10026), .A(n10025), .B(n10024), .ZN(
        n10028) );
  OAI22_X1 U10843 ( .A1(n10029), .A2(n10028), .B1(keyinput_23), .B2(SI_9_), 
        .ZN(n10030) );
  AOI21_X1 U10844 ( .B1(keyinput_23), .B2(SI_9_), .A(n10030), .ZN(n10031) );
  AOI221_X1 U10845 ( .B1(SI_8_), .B2(n10032), .C1(n10093), .C2(keyinput_24), 
        .A(n10031), .ZN(n10038) );
  INV_X1 U10846 ( .A(SI_7_), .ZN(n10144) );
  AOI22_X1 U10847 ( .A1(n10034), .A2(keyinput_27), .B1(n10144), .B2(
        keyinput_25), .ZN(n10033) );
  OAI221_X1 U10848 ( .B1(n10034), .B2(keyinput_27), .C1(n10144), .C2(
        keyinput_25), .A(n10033), .ZN(n10037) );
  AOI22_X1 U10849 ( .A1(SI_4_), .A2(keyinput_28), .B1(SI_6_), .B2(keyinput_26), 
        .ZN(n10035) );
  OAI221_X1 U10850 ( .B1(SI_4_), .B2(keyinput_28), .C1(SI_6_), .C2(keyinput_26), .A(n10035), .ZN(n10036) );
  NOR3_X1 U10851 ( .A1(n10038), .A2(n10037), .A3(n10036), .ZN(n10039) );
  AOI221_X1 U10852 ( .B1(SI_3_), .B2(keyinput_29), .C1(n10151), .C2(n10040), 
        .A(n10039), .ZN(n10043) );
  INV_X1 U10853 ( .A(keyinput_30), .ZN(n10041) );
  MUX2_X1 U10854 ( .A(keyinput_30), .B(n10041), .S(SI_2_), .Z(n10042) );
  OR2_X1 U10855 ( .A1(n10043), .A2(n10042), .ZN(n10045) );
  INV_X1 U10856 ( .A(SI_0_), .ZN(n10157) );
  INV_X1 U10857 ( .A(keyinput_32), .ZN(n10044) );
  AOI222_X1 U10858 ( .A1(n10046), .A2(n10045), .B1(keyinput_32), .B2(n10157), 
        .C1(SI_0_), .C2(n10044), .ZN(n10048) );
  NAND2_X1 U10859 ( .A1(n10166), .A2(keyinput_38), .ZN(n10047) );
  OAI221_X1 U10860 ( .B1(n10049), .B2(n10048), .C1(n10166), .C2(keyinput_38), 
        .A(n10047), .ZN(n10050) );
  NAND4_X1 U10861 ( .A1(n10053), .A2(n10052), .A3(n10051), .A4(n10050), .ZN(
        n10054) );
  OAI221_X1 U10862 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_45), .C1(
        n10172), .C2(n10055), .A(n10054), .ZN(n10056) );
  AOI22_X1 U10863 ( .A1(keyinput_48), .A2(n10177), .B1(n10057), .B2(n10056), 
        .ZN(n10058) );
  OAI21_X1 U10864 ( .B1(n10177), .B2(keyinput_48), .A(n10058), .ZN(n10059) );
  OAI211_X1 U10865 ( .C1(P2_REG3_REG_24__SCAN_IN), .C2(keyinput_51), .A(n10060), .B(n10059), .ZN(n10061) );
  AOI21_X1 U10866 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_51), .A(n10061), 
        .ZN(n10062) );
  AOI221_X1 U10867 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(n10063), .C1(n5665), 
        .C2(keyinput_52), .A(n10062), .ZN(n10064) );
  OAI22_X1 U10868 ( .A1(n10065), .A2(n10064), .B1(keyinput_55), .B2(
        P2_REG3_REG_20__SCAN_IN), .ZN(n10066) );
  AOI21_X1 U10869 ( .B1(keyinput_55), .B2(P2_REG3_REG_20__SCAN_IN), .A(n10066), 
        .ZN(n10067) );
  AOI221_X1 U10870 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_56), .C1(n5791), .C2(n10068), .A(n10067), .ZN(n10069) );
  AOI221_X1 U10871 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(n10070), .C1(n10192), 
        .C2(keyinput_57), .A(n10069), .ZN(n10071) );
  OAI22_X1 U10872 ( .A1(n10072), .A2(n10071), .B1(keyinput_60), .B2(
        P2_REG3_REG_18__SCAN_IN), .ZN(n10073) );
  AOI21_X1 U10873 ( .B1(keyinput_60), .B2(P2_REG3_REG_18__SCAN_IN), .A(n10073), 
        .ZN(n10074) );
  OAI22_X1 U10874 ( .A1(keyinput_63), .A2(n5833), .B1(n10075), .B2(n10074), 
        .ZN(n10076) );
  AOI21_X1 U10875 ( .B1(keyinput_63), .B2(n5833), .A(n10076), .ZN(n10200) );
  AOI22_X1 U10876 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_123), .B1(n10078), .B2(keyinput_122), .ZN(n10077) );
  OAI221_X1 U10877 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_123), .C1(
        n10078), .C2(keyinput_122), .A(n10077), .ZN(n10194) );
  INV_X1 U10878 ( .A(keyinput_121), .ZN(n10191) );
  INV_X1 U10879 ( .A(keyinput_120), .ZN(n10189) );
  AOI22_X1 U10880 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_118), .B1(n5740), 
        .B2(keyinput_117), .ZN(n10079) );
  OAI221_X1 U10881 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_118), .C1(n5740), .C2(keyinput_117), .A(n10079), .ZN(n10185) );
  INV_X1 U10882 ( .A(keyinput_116), .ZN(n10183) );
  OAI22_X1 U10883 ( .A1(n5867), .A2(keyinput_114), .B1(n10081), .B2(
        keyinput_115), .ZN(n10080) );
  AOI221_X1 U10884 ( .B1(n5867), .B2(keyinput_114), .C1(keyinput_115), .C2(
        n10081), .A(n10080), .ZN(n10179) );
  OAI22_X1 U10885 ( .A1(n10083), .A2(keyinput_111), .B1(keyinput_110), .B2(
        P2_REG3_REG_12__SCAN_IN), .ZN(n10082) );
  AOI221_X1 U10886 ( .B1(n10083), .B2(keyinput_111), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_110), .A(n10082), .ZN(n10175)
         );
  INV_X1 U10887 ( .A(keyinput_109), .ZN(n10173) );
  OAI22_X1 U10888 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_107), .B1(
        P2_REG3_REG_10__SCAN_IN), .B2(keyinput_103), .ZN(n10084) );
  AOI221_X1 U10889 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_107), .C1(
        keyinput_103), .C2(P2_REG3_REG_10__SCAN_IN), .A(n10084), .ZN(n10170)
         );
  OAI22_X1 U10890 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_104), .B1(
        keyinput_108), .B2(P2_REG3_REG_1__SCAN_IN), .ZN(n10085) );
  AOI221_X1 U10891 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_104), .C1(
        P2_REG3_REG_1__SCAN_IN), .C2(keyinput_108), .A(n10085), .ZN(n10169) );
  OAI22_X1 U10892 ( .A1(n5902), .A2(keyinput_105), .B1(keyinput_106), .B2(
        P2_REG3_REG_28__SCAN_IN), .ZN(n10086) );
  AOI221_X1 U10893 ( .B1(n5902), .B2(keyinput_105), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_106), .A(n10086), .ZN(n10168)
         );
  AOI22_X1 U10894 ( .A1(n10515), .A2(keyinput_99), .B1(n5518), .B2(keyinput_97), .ZN(n10087) );
  OAI221_X1 U10895 ( .B1(n10515), .B2(keyinput_99), .C1(n5518), .C2(
        keyinput_97), .A(n10087), .ZN(n10092) );
  OAI22_X1 U10896 ( .A1(n10089), .A2(keyinput_101), .B1(P2_STATE_REG_SCAN_IN), 
        .B2(keyinput_98), .ZN(n10088) );
  AOI221_X1 U10897 ( .B1(n10089), .B2(keyinput_101), .C1(keyinput_98), .C2(
        P2_STATE_REG_SCAN_IN), .A(n10088), .ZN(n10090) );
  OAI21_X1 U10898 ( .B1(keyinput_100), .B2(P2_REG3_REG_27__SCAN_IN), .A(n10090), .ZN(n10091) );
  AOI211_X1 U10899 ( .C1(keyinput_100), .C2(P2_REG3_REG_27__SCAN_IN), .A(
        n10092), .B(n10091), .ZN(n10164) );
  INV_X1 U10900 ( .A(keyinput_93), .ZN(n10152) );
  XOR2_X1 U10901 ( .A(n10093), .B(keyinput_88), .Z(n10149) );
  INV_X1 U10902 ( .A(SI_11_), .ZN(n10095) );
  AOI22_X1 U10903 ( .A1(SI_10_), .A2(keyinput_86), .B1(n10095), .B2(
        keyinput_85), .ZN(n10094) );
  OAI221_X1 U10904 ( .B1(SI_10_), .B2(keyinput_86), .C1(n10095), .C2(
        keyinput_85), .A(n10094), .ZN(n10140) );
  OAI22_X1 U10905 ( .A1(n10097), .A2(keyinput_81), .B1(SI_16_), .B2(
        keyinput_80), .ZN(n10096) );
  AOI221_X1 U10906 ( .B1(n10097), .B2(keyinput_81), .C1(keyinput_80), .C2(
        SI_16_), .A(n10096), .ZN(n10138) );
  OAI22_X1 U10907 ( .A1(n10099), .A2(keyinput_78), .B1(keyinput_77), .B2(
        SI_19_), .ZN(n10098) );
  AOI221_X1 U10908 ( .B1(n10099), .B2(keyinput_78), .C1(SI_19_), .C2(
        keyinput_77), .A(n10098), .ZN(n10130) );
  INV_X1 U10909 ( .A(keyinput_76), .ZN(n10128) );
  INV_X1 U10910 ( .A(keyinput_75), .ZN(n10125) );
  INV_X1 U10911 ( .A(keyinput_74), .ZN(n10121) );
  INV_X1 U10912 ( .A(keyinput_73), .ZN(n10119) );
  INV_X1 U10913 ( .A(keyinput_72), .ZN(n10115) );
  INV_X1 U10914 ( .A(keyinput_71), .ZN(n10112) );
  INV_X1 U10915 ( .A(keyinput_70), .ZN(n10110) );
  OAI22_X1 U10916 ( .A1(SI_31_), .A2(keyinput_65), .B1(P2_WR_REG_SCAN_IN), 
        .B2(keyinput_64), .ZN(n10100) );
  AOI221_X1 U10917 ( .B1(SI_31_), .B2(keyinput_65), .C1(keyinput_64), .C2(
        P2_WR_REG_SCAN_IN), .A(n10100), .ZN(n10107) );
  AOI22_X1 U10918 ( .A1(SI_30_), .A2(keyinput_66), .B1(n10102), .B2(
        keyinput_67), .ZN(n10101) );
  OAI221_X1 U10919 ( .B1(SI_30_), .B2(keyinput_66), .C1(n10102), .C2(
        keyinput_67), .A(n10101), .ZN(n10106) );
  OAI22_X1 U10920 ( .A1(n10104), .A2(keyinput_68), .B1(keyinput_69), .B2(
        SI_27_), .ZN(n10103) );
  AOI221_X1 U10921 ( .B1(n10104), .B2(keyinput_68), .C1(SI_27_), .C2(
        keyinput_69), .A(n10103), .ZN(n10105) );
  OAI21_X1 U10922 ( .B1(n10107), .B2(n10106), .A(n10105), .ZN(n10108) );
  OAI221_X1 U10923 ( .B1(SI_26_), .B2(n10110), .C1(n10109), .C2(keyinput_70), 
        .A(n10108), .ZN(n10111) );
  OAI221_X1 U10924 ( .B1(SI_25_), .B2(keyinput_71), .C1(n10113), .C2(n10112), 
        .A(n10111), .ZN(n10114) );
  OAI221_X1 U10925 ( .B1(SI_24_), .B2(keyinput_72), .C1(n10116), .C2(n10115), 
        .A(n10114), .ZN(n10117) );
  OAI221_X1 U10926 ( .B1(SI_23_), .B2(n10119), .C1(n10118), .C2(keyinput_73), 
        .A(n10117), .ZN(n10120) );
  OAI221_X1 U10927 ( .B1(SI_22_), .B2(keyinput_74), .C1(n10122), .C2(n10121), 
        .A(n10120), .ZN(n10123) );
  OAI221_X1 U10928 ( .B1(SI_21_), .B2(n10125), .C1(n10124), .C2(keyinput_75), 
        .A(n10123), .ZN(n10126) );
  OAI221_X1 U10929 ( .B1(SI_20_), .B2(n10128), .C1(n10127), .C2(keyinput_76), 
        .A(n10126), .ZN(n10129) );
  AOI22_X1 U10930 ( .A1(n10130), .A2(n10129), .B1(keyinput_79), .B2(SI_17_), 
        .ZN(n10131) );
  OAI21_X1 U10931 ( .B1(keyinput_79), .B2(SI_17_), .A(n10131), .ZN(n10137) );
  INV_X1 U10932 ( .A(SI_14_), .ZN(n10132) );
  XOR2_X1 U10933 ( .A(n10132), .B(keyinput_82), .Z(n10136) );
  AOI22_X1 U10934 ( .A1(SI_12_), .A2(keyinput_84), .B1(n10134), .B2(
        keyinput_83), .ZN(n10133) );
  OAI221_X1 U10935 ( .B1(SI_12_), .B2(keyinput_84), .C1(n10134), .C2(
        keyinput_83), .A(n10133), .ZN(n10135) );
  AOI211_X1 U10936 ( .C1(n10138), .C2(n10137), .A(n10136), .B(n10135), .ZN(
        n10139) );
  OAI22_X1 U10937 ( .A1(keyinput_87), .A2(n10142), .B1(n10140), .B2(n10139), 
        .ZN(n10141) );
  AOI21_X1 U10938 ( .B1(keyinput_87), .B2(n10142), .A(n10141), .ZN(n10148) );
  OAI22_X1 U10939 ( .A1(n10144), .A2(keyinput_89), .B1(keyinput_90), .B2(SI_6_), .ZN(n10143) );
  AOI221_X1 U10940 ( .B1(n10144), .B2(keyinput_89), .C1(SI_6_), .C2(
        keyinput_90), .A(n10143), .ZN(n10147) );
  OAI22_X1 U10941 ( .A1(SI_5_), .A2(keyinput_91), .B1(SI_4_), .B2(keyinput_92), 
        .ZN(n10145) );
  AOI221_X1 U10942 ( .B1(SI_5_), .B2(keyinput_91), .C1(keyinput_92), .C2(SI_4_), .A(n10145), .ZN(n10146) );
  OAI211_X1 U10943 ( .C1(n10149), .C2(n10148), .A(n10147), .B(n10146), .ZN(
        n10150) );
  OAI221_X1 U10944 ( .B1(SI_3_), .B2(n10152), .C1(n10151), .C2(keyinput_93), 
        .A(n10150), .ZN(n10155) );
  INV_X1 U10945 ( .A(keyinput_94), .ZN(n10153) );
  MUX2_X1 U10946 ( .A(n10153), .B(keyinput_94), .S(SI_2_), .Z(n10154) );
  NAND2_X1 U10947 ( .A1(n10155), .A2(n10154), .ZN(n10161) );
  INV_X1 U10948 ( .A(keyinput_95), .ZN(n10156) );
  MUX2_X1 U10949 ( .A(n10156), .B(keyinput_95), .S(SI_1_), .Z(n10160) );
  INV_X1 U10950 ( .A(keyinput_96), .ZN(n10158) );
  OAI22_X1 U10951 ( .A1(SI_0_), .A2(n10158), .B1(keyinput_96), .B2(n10157), 
        .ZN(n10159) );
  AOI21_X1 U10952 ( .B1(n10161), .B2(n10160), .A(n10159), .ZN(n10162) );
  INV_X1 U10953 ( .A(n10162), .ZN(n10163) );
  AOI22_X1 U10954 ( .A1(keyinput_102), .A2(n10166), .B1(n10164), .B2(n10163), 
        .ZN(n10165) );
  OAI21_X1 U10955 ( .B1(n10166), .B2(keyinput_102), .A(n10165), .ZN(n10167) );
  NAND4_X1 U10956 ( .A1(n10170), .A2(n10169), .A3(n10168), .A4(n10167), .ZN(
        n10171) );
  OAI221_X1 U10957 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(n10173), .C1(n10172), 
        .C2(keyinput_109), .A(n10171), .ZN(n10174) );
  AOI22_X1 U10958 ( .A1(keyinput_112), .A2(n10177), .B1(n10175), .B2(n10174), 
        .ZN(n10176) );
  OAI21_X1 U10959 ( .B1(n10177), .B2(keyinput_112), .A(n10176), .ZN(n10178) );
  OAI211_X1 U10960 ( .C1(n10181), .C2(keyinput_113), .A(n10179), .B(n10178), 
        .ZN(n10180) );
  AOI21_X1 U10961 ( .B1(n10181), .B2(keyinput_113), .A(n10180), .ZN(n10182) );
  AOI221_X1 U10962 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(n10183), .C1(n5665), 
        .C2(keyinput_116), .A(n10182), .ZN(n10184) );
  OAI22_X1 U10963 ( .A1(keyinput_119), .A2(n10187), .B1(n10185), .B2(n10184), 
        .ZN(n10186) );
  AOI21_X1 U10964 ( .B1(keyinput_119), .B2(n10187), .A(n10186), .ZN(n10188) );
  AOI221_X1 U10965 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_120), .C1(
        n5791), .C2(n10189), .A(n10188), .ZN(n10190) );
  AOI221_X1 U10966 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_121), .C1(
        n10192), .C2(n10191), .A(n10190), .ZN(n10193) );
  OAI22_X1 U10967 ( .A1(n10194), .A2(n10193), .B1(keyinput_124), .B2(
        P2_REG3_REG_18__SCAN_IN), .ZN(n10195) );
  AOI21_X1 U10968 ( .B1(keyinput_124), .B2(P2_REG3_REG_18__SCAN_IN), .A(n10195), .ZN(n10198) );
  AOI22_X1 U10969 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_126), .B1(n5595), .B2(keyinput_125), .ZN(n10196) );
  OAI221_X1 U10970 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_126), .C1(
        n5595), .C2(keyinput_125), .A(n10196), .ZN(n10197) );
  OAI22_X1 U10971 ( .A1(n10198), .A2(n10197), .B1(keyinput_127), .B2(n5833), 
        .ZN(n10199) );
  AOI211_X1 U10972 ( .C1(keyinput_127), .C2(n5833), .A(n10200), .B(n10199), 
        .ZN(n10201) );
  XNOR2_X1 U10973 ( .A(n10202), .B(n10201), .ZN(P2_U3324) );
  XOR2_X1 U10974 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  INV_X1 U10975 ( .A(n10203), .ZN(n10204) );
  NAND2_X1 U10976 ( .A1(n10205), .A2(n10204), .ZN(n10206) );
  XOR2_X1 U10977 ( .A(n10207), .B(n10206), .Z(ADD_1071_U5) );
  XOR2_X1 U10978 ( .A(n10209), .B(n10208), .Z(ADD_1071_U54) );
  XOR2_X1 U10979 ( .A(n10211), .B(n10210), .Z(ADD_1071_U53) );
  XNOR2_X1 U10980 ( .A(n10213), .B(n10212), .ZN(ADD_1071_U52) );
  NOR2_X1 U10981 ( .A1(n10215), .A2(n10214), .ZN(n10216) );
  XOR2_X1 U10982 ( .A(n10216), .B(P2_ADDR_REG_5__SCAN_IN), .Z(ADD_1071_U51) );
  XOR2_X1 U10983 ( .A(n10217), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  XOR2_X1 U10984 ( .A(n10218), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U10985 ( .A(n10219), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  XOR2_X1 U10986 ( .A(n10220), .B(P2_ADDR_REG_9__SCAN_IN), .Z(ADD_1071_U47) );
  XOR2_X1 U10987 ( .A(n10222), .B(n10221), .Z(ADD_1071_U63) );
  XOR2_X1 U10988 ( .A(n10224), .B(n10223), .Z(ADD_1071_U62) );
  XNOR2_X1 U10989 ( .A(n10226), .B(n10225), .ZN(ADD_1071_U61) );
  XNOR2_X1 U10990 ( .A(n10228), .B(n10227), .ZN(ADD_1071_U60) );
  XNOR2_X1 U10991 ( .A(n10230), .B(n10229), .ZN(ADD_1071_U59) );
  XNOR2_X1 U10992 ( .A(n10232), .B(n10231), .ZN(ADD_1071_U58) );
  XNOR2_X1 U10993 ( .A(n10234), .B(n10233), .ZN(ADD_1071_U57) );
  XNOR2_X1 U10994 ( .A(n10236), .B(n10235), .ZN(ADD_1071_U56) );
  NOR2_X1 U10995 ( .A1(n10238), .A2(n10237), .ZN(n10239) );
  XOR2_X1 U10996 ( .A(P1_ADDR_REG_18__SCAN_IN), .B(n10239), .Z(ADD_1071_U55)
         );
  AOI22_X1 U10997 ( .A1(n10290), .A2(P1_ADDR_REG_10__SCAN_IN), .B1(n10240), 
        .B2(n10288), .ZN(n10251) );
  OAI21_X1 U10998 ( .B1(n10243), .B2(n10242), .A(n10241), .ZN(n10244) );
  NAND2_X1 U10999 ( .A1(n10244), .A2(n10368), .ZN(n10249) );
  OAI211_X1 U11000 ( .C1(n10247), .C2(n10246), .A(n10245), .B(n10348), .ZN(
        n10248) );
  NAND4_X1 U11001 ( .A1(n10251), .A2(n10250), .A3(n10249), .A4(n10248), .ZN(
        P1_U3251) );
  INV_X1 U11002 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10264) );
  AOI21_X1 U11003 ( .B1(n10288), .B2(n10253), .A(n10252), .ZN(n10263) );
  OAI21_X1 U11004 ( .B1(n10256), .B2(n10255), .A(n10254), .ZN(n10261) );
  OAI21_X1 U11005 ( .B1(n10259), .B2(n10258), .A(n10257), .ZN(n10260) );
  AOI22_X1 U11006 ( .A1(n10261), .A2(n10348), .B1(n10260), .B2(n10368), .ZN(
        n10262) );
  OAI211_X1 U11007 ( .C1(n10264), .C2(n10376), .A(n10263), .B(n10262), .ZN(
        P1_U3255) );
  INV_X1 U11008 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10282) );
  NAND2_X1 U11009 ( .A1(n10266), .A2(n10265), .ZN(n10269) );
  INV_X1 U11010 ( .A(n10267), .ZN(n10268) );
  NAND2_X1 U11011 ( .A1(n10269), .A2(n10268), .ZN(n10270) );
  OR2_X1 U11012 ( .A1(n10333), .A2(n10270), .ZN(n10273) );
  INV_X1 U11013 ( .A(n10271), .ZN(n10272) );
  OAI211_X1 U11014 ( .C1(n10364), .C2(n10274), .A(n10273), .B(n10272), .ZN(
        n10275) );
  INV_X1 U11015 ( .A(n10275), .ZN(n10281) );
  AOI21_X1 U11016 ( .B1(n10278), .B2(n10277), .A(n10276), .ZN(n10279) );
  OR2_X1 U11017 ( .A1(n10370), .A2(n10279), .ZN(n10280) );
  OAI211_X1 U11018 ( .C1(n10376), .C2(n10282), .A(n10281), .B(n10280), .ZN(
        P1_U3246) );
  NAND2_X1 U11019 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n10285) );
  AOI211_X1 U11020 ( .C1(n10285), .C2(n10284), .A(n10283), .B(n10333), .ZN(
        n10286) );
  AOI21_X1 U11021 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(P1_U3084), .A(n10286), 
        .ZN(n10296) );
  INV_X1 U11022 ( .A(n10287), .ZN(n10289) );
  AOI22_X1 U11023 ( .A1(n10290), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(n10289), 
        .B2(n10288), .ZN(n10295) );
  NOR2_X1 U11024 ( .A1(n10342), .A2(n10291), .ZN(n10337) );
  OAI211_X1 U11025 ( .C1(n10337), .C2(n10293), .A(n10348), .B(n10292), .ZN(
        n10294) );
  NAND3_X1 U11026 ( .A1(n10296), .A2(n10295), .A3(n10294), .ZN(P1_U3242) );
  INV_X1 U11027 ( .A(n10297), .ZN(n10299) );
  AOI22_X1 U11028 ( .A1(n10300), .A2(n10299), .B1(n10298), .B2(n4857), .ZN(
        P2_U3437) );
  OAI22_X1 U11029 ( .A1(n4946), .A2(n10303), .B1(n10380), .B2(n10320), .ZN(
        n10302) );
  AOI22_X1 U11030 ( .A1(n10302), .A2(n10301), .B1(P2_ADDR_REG_0__SCAN_IN), 
        .B2(n10319), .ZN(n10307) );
  AOI21_X1 U11031 ( .B1(n4948), .B2(n10303), .A(n10330), .ZN(n10304) );
  OAI21_X1 U11032 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n10320), .A(n10304), .ZN(
        n10305) );
  NAND2_X1 U11033 ( .A1(n10305), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n10306) );
  OAI211_X1 U11034 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10388), .A(n10307), .B(
        n10306), .ZN(P2_U3245) );
  AOI22_X1 U11035 ( .A1(n10319), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n10318) );
  NAND2_X1 U11036 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10310) );
  AOI211_X1 U11037 ( .C1(n10310), .C2(n10309), .A(n10308), .B(n10320), .ZN(
        n10315) );
  NAND2_X1 U11038 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n10313) );
  AOI211_X1 U11039 ( .C1(n10313), .C2(n10312), .A(n10311), .B(n4946), .ZN(
        n10314) );
  AOI211_X1 U11040 ( .C1(n10330), .C2(n10316), .A(n10315), .B(n10314), .ZN(
        n10317) );
  NAND2_X1 U11041 ( .A1(n10318), .A2(n10317), .ZN(P2_U3246) );
  AOI22_X1 U11042 ( .A1(n10319), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n10332) );
  AOI211_X1 U11043 ( .C1(n10323), .C2(n10322), .A(n10321), .B(n10320), .ZN(
        n10328) );
  AOI211_X1 U11044 ( .C1(n10326), .C2(n10325), .A(n10324), .B(n4946), .ZN(
        n10327) );
  AOI211_X1 U11045 ( .C1(n10330), .C2(n10329), .A(n10328), .B(n10327), .ZN(
        n10331) );
  NAND2_X1 U11046 ( .A1(n10332), .A2(n10331), .ZN(P2_U3247) );
  XOR2_X1 U11047 ( .A(P1_RD_REG_SCAN_IN), .B(n5518), .Z(U126) );
  AOI211_X1 U11048 ( .C1(n10336), .C2(n10335), .A(n10334), .B(n10333), .ZN(
        n10354) );
  AND3_X1 U11049 ( .A1(n10339), .A2(n10338), .A3(n10337), .ZN(n10341) );
  AOI211_X1 U11050 ( .C1(n10343), .C2(n10342), .A(n10341), .B(n10340), .ZN(
        n10344) );
  OAI21_X1 U11051 ( .B1(n10346), .B2(n10345), .A(n10344), .ZN(n10373) );
  OAI211_X1 U11052 ( .C1(n10350), .C2(n10349), .A(n10348), .B(n10347), .ZN(
        n10351) );
  OAI211_X1 U11053 ( .C1(n10364), .C2(n10352), .A(n10373), .B(n10351), .ZN(
        n10353) );
  AOI211_X1 U11054 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(P1_U3084), .A(n10354), 
        .B(n10353), .ZN(n10355) );
  OAI21_X1 U11055 ( .B1(n10356), .B2(n10376), .A(n10355), .ZN(P1_U3243) );
  AOI21_X1 U11056 ( .B1(n10359), .B2(n10358), .A(n10357), .ZN(n10371) );
  OAI21_X1 U11057 ( .B1(n10362), .B2(n10361), .A(n10360), .ZN(n10367) );
  NOR2_X1 U11058 ( .A1(n10364), .A2(n10363), .ZN(n10365) );
  AOI211_X1 U11059 ( .C1(n10368), .C2(n10367), .A(n10366), .B(n10365), .ZN(
        n10369) );
  OAI21_X1 U11060 ( .B1(n10371), .B2(n10370), .A(n10369), .ZN(n10372) );
  INV_X1 U11061 ( .A(n10372), .ZN(n10374) );
  OAI211_X1 U11062 ( .C1(n10376), .C2(n10375), .A(n10374), .B(n10373), .ZN(
        P1_U3245) );
  OAI21_X1 U11063 ( .B1(n9234), .B2(n10596), .A(n10377), .ZN(n10379) );
  NAND2_X1 U11064 ( .A1(n10379), .A2(n10378), .ZN(n10386) );
  NOR2_X1 U11065 ( .A1(n10605), .A2(n10380), .ZN(n10385) );
  AOI21_X1 U11066 ( .B1(n10383), .B2(n10382), .A(n10381), .ZN(n10384) );
  AOI211_X1 U11067 ( .C1(n10605), .C2(n10386), .A(n10385), .B(n10384), .ZN(
        n10387) );
  OAI21_X1 U11068 ( .B1(n10388), .B2(n10609), .A(n10387), .ZN(P2_U3296) );
  OR2_X1 U11069 ( .A1(n10405), .A2(n10389), .ZN(n10390) );
  NAND2_X1 U11070 ( .A1(n10391), .A2(n10390), .ZN(n10398) );
  NAND2_X1 U11071 ( .A1(n6813), .A2(n10392), .ZN(n10395) );
  NAND2_X1 U11072 ( .A1(n6676), .A2(n10393), .ZN(n10394) );
  NAND2_X1 U11073 ( .A1(n10395), .A2(n10394), .ZN(n10396) );
  AOI21_X1 U11074 ( .B1(n10398), .B2(n10397), .A(n10396), .ZN(n10422) );
  NAND2_X1 U11075 ( .A1(n10399), .A2(n10413), .ZN(n10401) );
  NAND3_X1 U11076 ( .A1(n10401), .A2(n10482), .A3(n10400), .ZN(n10416) );
  NAND2_X1 U11077 ( .A1(n10413), .A2(n10501), .ZN(n10402) );
  AND2_X1 U11078 ( .A1(n10416), .A2(n10402), .ZN(n10408) );
  INV_X1 U11079 ( .A(n10403), .ZN(n10404) );
  XNOR2_X1 U11080 ( .A(n10405), .B(n10404), .ZN(n10419) );
  NAND2_X1 U11081 ( .A1(n10419), .A2(n10640), .ZN(n10407) );
  AND3_X1 U11082 ( .A1(n10422), .A2(n10408), .A3(n10407), .ZN(n10410) );
  AOI22_X1 U11083 ( .A1(n10644), .A2(n10410), .B1(n6638), .B2(n10642), .ZN(
        P1_U3524) );
  INV_X1 U11084 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10409) );
  AOI22_X1 U11085 ( .A1(n10491), .A2(n10410), .B1(n10409), .B2(n10645), .ZN(
        P1_U3457) );
  AOI22_X1 U11086 ( .A1(n10413), .A2(n10412), .B1(n10411), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n10414) );
  OAI21_X1 U11087 ( .B1(n10416), .B2(n10415), .A(n10414), .ZN(n10417) );
  INV_X1 U11088 ( .A(n10417), .ZN(n10421) );
  NAND2_X1 U11089 ( .A1(n10419), .A2(n10418), .ZN(n10420) );
  AND3_X1 U11090 ( .A1(n10422), .A2(n10421), .A3(n10420), .ZN(n10423) );
  AOI22_X1 U11091 ( .A1(n10425), .A2(n10424), .B1(n10423), .B2(n9822), .ZN(
        P1_U3290) );
  AOI22_X1 U11092 ( .A1(n10427), .A2(n10482), .B1(n10501), .B2(n10426), .ZN(
        n10428) );
  OAI211_X1 U11093 ( .C1(n10430), .C2(n10504), .A(n10429), .B(n10428), .ZN(
        n10431) );
  INV_X1 U11094 ( .A(n10431), .ZN(n10434) );
  INV_X1 U11095 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10432) );
  AOI22_X1 U11096 ( .A1(n10644), .A2(n10434), .B1(n10432), .B2(n10642), .ZN(
        P1_U3525) );
  INV_X1 U11097 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10433) );
  AOI22_X1 U11098 ( .A1(n10491), .A2(n10434), .B1(n10433), .B2(n10645), .ZN(
        P1_U3460) );
  INV_X1 U11099 ( .A(n10435), .ZN(n10576) );
  OAI22_X1 U11100 ( .A1(n10437), .A2(n10650), .B1(n10436), .B2(n10648), .ZN(
        n10439) );
  AOI211_X1 U11101 ( .C1(n10576), .C2(n10440), .A(n10439), .B(n10438), .ZN(
        n10442) );
  AOI22_X1 U11102 ( .A1(n10657), .A2(n10442), .B1(n5630), .B2(n10656), .ZN(
        P2_U3522) );
  INV_X1 U11103 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10441) );
  AOI22_X1 U11104 ( .A1(n10660), .A2(n10442), .B1(n10441), .B2(n10658), .ZN(
        P2_U3457) );
  OAI22_X1 U11105 ( .A1(n10444), .A2(n10548), .B1(n10443), .B2(n10637), .ZN(
        n10445) );
  AOI21_X1 U11106 ( .B1(n10446), .B2(n10617), .A(n10445), .ZN(n10447) );
  AND2_X1 U11107 ( .A1(n10448), .A2(n10447), .ZN(n10451) );
  INV_X1 U11108 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10449) );
  AOI22_X1 U11109 ( .A1(n10644), .A2(n10451), .B1(n10449), .B2(n10642), .ZN(
        P1_U3526) );
  INV_X1 U11110 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10450) );
  AOI22_X1 U11111 ( .A1(n10491), .A2(n10451), .B1(n10450), .B2(n10645), .ZN(
        P1_U3463) );
  OAI22_X1 U11112 ( .A1(n10453), .A2(n10548), .B1(n10452), .B2(n10637), .ZN(
        n10454) );
  AOI21_X1 U11113 ( .B1(n10455), .B2(n10640), .A(n10454), .ZN(n10456) );
  AOI22_X1 U11114 ( .A1(n10644), .A2(n10459), .B1(n6419), .B2(n10642), .ZN(
        P1_U3527) );
  INV_X1 U11115 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10458) );
  AOI22_X1 U11116 ( .A1(n10491), .A2(n10459), .B1(n10458), .B2(n10645), .ZN(
        P1_U3466) );
  OAI22_X1 U11117 ( .A1(n10461), .A2(n10650), .B1(n10460), .B2(n10648), .ZN(
        n10463) );
  AOI211_X1 U11118 ( .C1(n10464), .C2(n10654), .A(n10463), .B(n10462), .ZN(
        n10465) );
  AOI22_X1 U11119 ( .A1(n10657), .A2(n10465), .B1(n6182), .B2(n10656), .ZN(
        P2_U3524) );
  AOI22_X1 U11120 ( .A1(n10660), .A2(n10465), .B1(n5669), .B2(n10658), .ZN(
        P2_U3463) );
  INV_X1 U11121 ( .A(n10466), .ZN(n10467) );
  OAI21_X1 U11122 ( .B1(n10468), .B2(n10637), .A(n10467), .ZN(n10470) );
  AOI211_X1 U11123 ( .C1(n10471), .C2(n10640), .A(n10470), .B(n10469), .ZN(
        n10473) );
  AOI22_X1 U11124 ( .A1(n10644), .A2(n10473), .B1(n6436), .B2(n10642), .ZN(
        P1_U3528) );
  INV_X1 U11125 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U11126 ( .A1(n10491), .A2(n10473), .B1(n10472), .B2(n10645), .ZN(
        P1_U3469) );
  AOI21_X1 U11127 ( .B1(n10628), .B2(n10475), .A(n10474), .ZN(n10476) );
  OAI211_X1 U11128 ( .C1(n10478), .C2(n10530), .A(n10477), .B(n10476), .ZN(
        n10479) );
  INV_X1 U11129 ( .A(n10479), .ZN(n10480) );
  AOI22_X1 U11130 ( .A1(n10657), .A2(n10480), .B1(n6183), .B2(n10656), .ZN(
        P2_U3525) );
  AOI22_X1 U11131 ( .A1(n10660), .A2(n10480), .B1(n5680), .B2(n10658), .ZN(
        P2_U3466) );
  INV_X1 U11132 ( .A(n10481), .ZN(n10488) );
  NAND2_X1 U11133 ( .A1(n10483), .A2(n10482), .ZN(n10484) );
  OAI21_X1 U11134 ( .B1(n10485), .B2(n10637), .A(n10484), .ZN(n10487) );
  AOI211_X1 U11135 ( .C1(n10488), .C2(n10640), .A(n10487), .B(n10486), .ZN(
        n10490) );
  AOI22_X1 U11136 ( .A1(n10644), .A2(n10490), .B1(n6429), .B2(n10642), .ZN(
        P1_U3529) );
  INV_X1 U11137 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10489) );
  AOI22_X1 U11138 ( .A1(n10491), .A2(n10490), .B1(n10489), .B2(n10645), .ZN(
        P1_U3472) );
  AOI22_X1 U11139 ( .A1(n10493), .A2(n10629), .B1(n10628), .B2(n10492), .ZN(
        n10497) );
  NAND3_X1 U11140 ( .A1(n10495), .A2(n10494), .A3(n10654), .ZN(n10496) );
  AND3_X1 U11141 ( .A1(n10498), .A2(n10497), .A3(n10496), .ZN(n10499) );
  AOI22_X1 U11142 ( .A1(n10657), .A2(n10499), .B1(n6184), .B2(n10656), .ZN(
        P2_U3526) );
  AOI22_X1 U11143 ( .A1(n10660), .A2(n10499), .B1(n5596), .B2(n10658), .ZN(
        P2_U3469) );
  AOI21_X1 U11144 ( .B1(n10501), .B2(n5131), .A(n10500), .ZN(n10502) );
  OAI211_X1 U11145 ( .C1(n10505), .C2(n10504), .A(n10503), .B(n10502), .ZN(
        n10506) );
  INV_X1 U11146 ( .A(n10506), .ZN(n10508) );
  AOI22_X1 U11147 ( .A1(n10644), .A2(n10508), .B1(n6412), .B2(n10642), .ZN(
        P1_U3530) );
  INV_X1 U11148 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10507) );
  AOI22_X1 U11149 ( .A1(n10491), .A2(n10508), .B1(n10507), .B2(n10645), .ZN(
        P1_U3475) );
  AOI211_X1 U11150 ( .C1(n10512), .C2(n10511), .A(n10510), .B(n10509), .ZN(
        n10521) );
  AND2_X1 U11151 ( .A1(n8918), .A2(n10525), .ZN(n10520) );
  NOR2_X1 U11152 ( .A1(n10514), .A2(n10513), .ZN(n10519) );
  OAI22_X1 U11153 ( .A1(n10517), .A2(n10516), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10515), .ZN(n10518) );
  NOR4_X1 U11154 ( .A1(n10521), .A2(n10520), .A3(n10519), .A4(n10518), .ZN(
        n10522) );
  OAI21_X1 U11155 ( .B1(n10524), .B2(n10523), .A(n10522), .ZN(P2_U3215) );
  AOI22_X1 U11156 ( .A1(n10526), .A2(n10629), .B1(n10628), .B2(n10525), .ZN(
        n10527) );
  OAI211_X1 U11157 ( .C1(n10530), .C2(n10529), .A(n10528), .B(n10527), .ZN(
        n10531) );
  INV_X1 U11158 ( .A(n10531), .ZN(n10533) );
  AOI22_X1 U11159 ( .A1(n10657), .A2(n10533), .B1(n6185), .B2(n10656), .ZN(
        P2_U3527) );
  INV_X1 U11160 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10532) );
  AOI22_X1 U11161 ( .A1(n10660), .A2(n10533), .B1(n10532), .B2(n10658), .ZN(
        P2_U3472) );
  INV_X1 U11162 ( .A(n10534), .ZN(n10535) );
  OAI22_X1 U11163 ( .A1(n10536), .A2(n10548), .B1(n10535), .B2(n10637), .ZN(
        n10538) );
  AOI211_X1 U11164 ( .C1(n10539), .C2(n10640), .A(n10538), .B(n10537), .ZN(
        n10541) );
  AOI22_X1 U11165 ( .A1(n10644), .A2(n10541), .B1(n7148), .B2(n10642), .ZN(
        P1_U3531) );
  INV_X1 U11166 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10540) );
  AOI22_X1 U11167 ( .A1(n10491), .A2(n10541), .B1(n10540), .B2(n10645), .ZN(
        P1_U3478) );
  OAI21_X1 U11168 ( .B1(n5286), .B2(n10648), .A(n10542), .ZN(n10544) );
  AOI211_X1 U11169 ( .C1(n10545), .C2(n10654), .A(n10544), .B(n10543), .ZN(
        n10546) );
  AOI22_X1 U11170 ( .A1(n10657), .A2(n10546), .B1(n6186), .B2(n10656), .ZN(
        P2_U3528) );
  AOI22_X1 U11171 ( .A1(n10660), .A2(n10546), .B1(n5713), .B2(n10658), .ZN(
        P2_U3475) );
  OAI22_X1 U11172 ( .A1(n10549), .A2(n10548), .B1(n5145), .B2(n10637), .ZN(
        n10551) );
  AOI211_X1 U11173 ( .C1(n10617), .C2(n10552), .A(n10551), .B(n10550), .ZN(
        n10554) );
  AOI22_X1 U11174 ( .A1(n10644), .A2(n10554), .B1(n7275), .B2(n10642), .ZN(
        P1_U3532) );
  INV_X1 U11175 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10553) );
  AOI22_X1 U11176 ( .A1(n10491), .A2(n10554), .B1(n10553), .B2(n10645), .ZN(
        P1_U3481) );
  OAI22_X1 U11177 ( .A1(n10556), .A2(n10650), .B1(n10555), .B2(n10648), .ZN(
        n10558) );
  AOI211_X1 U11178 ( .C1(n10654), .C2(n10559), .A(n10558), .B(n10557), .ZN(
        n10560) );
  AOI22_X1 U11179 ( .A1(n10657), .A2(n10560), .B1(n6187), .B2(n10656), .ZN(
        P2_U3529) );
  AOI22_X1 U11180 ( .A1(n10660), .A2(n10560), .B1(n5585), .B2(n10658), .ZN(
        P2_U3478) );
  OAI21_X1 U11181 ( .B1(n10562), .B2(n10637), .A(n10561), .ZN(n10563) );
  AOI21_X1 U11182 ( .B1(n10564), .B2(n10617), .A(n10563), .ZN(n10565) );
  AND2_X1 U11183 ( .A1(n10566), .A2(n10565), .ZN(n10569) );
  AOI22_X1 U11184 ( .A1(n10644), .A2(n10569), .B1(n10567), .B2(n10642), .ZN(
        P1_U3533) );
  INV_X1 U11185 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U11186 ( .A1(n10491), .A2(n10569), .B1(n10568), .B2(n10645), .ZN(
        P1_U3484) );
  INV_X1 U11187 ( .A(n10570), .ZN(n10575) );
  OAI22_X1 U11188 ( .A1(n10572), .A2(n10650), .B1(n10571), .B2(n10648), .ZN(
        n10574) );
  AOI211_X1 U11189 ( .C1(n10576), .C2(n10575), .A(n10574), .B(n10573), .ZN(
        n10578) );
  AOI22_X1 U11190 ( .A1(n10657), .A2(n10578), .B1(n6188), .B2(n10656), .ZN(
        P2_U3530) );
  INV_X1 U11191 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10577) );
  AOI22_X1 U11192 ( .A1(n10660), .A2(n10578), .B1(n10577), .B2(n10658), .ZN(
        P2_U3481) );
  OAI21_X1 U11193 ( .B1(n10580), .B2(n10581), .A(n10579), .ZN(n10603) );
  INV_X1 U11194 ( .A(n10603), .ZN(n10593) );
  NAND3_X1 U11195 ( .A1(n10583), .A2(n10582), .A3(n10581), .ZN(n10584) );
  NAND2_X1 U11196 ( .A1(n10585), .A2(n10584), .ZN(n10589) );
  AOI222_X1 U11197 ( .A1(n9234), .A2(n10589), .B1(n10588), .B2(n10587), .C1(
        n10586), .C2(n9230), .ZN(n10602) );
  OAI211_X1 U11198 ( .C1(n4975), .C2(n4974), .A(n10629), .B(n10591), .ZN(
        n10597) );
  OAI211_X1 U11199 ( .C1(n4974), .C2(n10648), .A(n10602), .B(n10597), .ZN(
        n10592) );
  AOI21_X1 U11200 ( .B1(n10593), .B2(n10654), .A(n10592), .ZN(n10595) );
  AOI22_X1 U11201 ( .A1(n10657), .A2(n10595), .B1(n6189), .B2(n10656), .ZN(
        P2_U3531) );
  INV_X1 U11202 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10594) );
  AOI22_X1 U11203 ( .A1(n10660), .A2(n10595), .B1(n10594), .B2(n10658), .ZN(
        P2_U3484) );
  INV_X1 U11204 ( .A(n10596), .ZN(n10604) );
  INV_X1 U11205 ( .A(n10597), .ZN(n10600) );
  AOI22_X1 U11206 ( .A1(n10600), .A2(n5582), .B1(n10599), .B2(n10598), .ZN(
        n10601) );
  OAI211_X1 U11207 ( .C1(n10604), .C2(n10603), .A(n10602), .B(n10601), .ZN(
        n10606) );
  AOI22_X1 U11208 ( .A1(n10607), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n10606), 
        .B2(n10605), .ZN(n10608) );
  OAI21_X1 U11209 ( .B1(n10610), .B2(n10609), .A(n10608), .ZN(P2_U3285) );
  INV_X1 U11210 ( .A(n10611), .ZN(n10616) );
  OAI21_X1 U11211 ( .B1(n10613), .B2(n10637), .A(n10612), .ZN(n10615) );
  AOI211_X1 U11212 ( .C1(n10617), .C2(n10616), .A(n10615), .B(n10614), .ZN(
        n10619) );
  AOI22_X1 U11213 ( .A1(n10644), .A2(n10619), .B1(n7559), .B2(n10642), .ZN(
        P1_U3535) );
  INV_X1 U11214 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10618) );
  AOI22_X1 U11215 ( .A1(n10491), .A2(n10619), .B1(n10618), .B2(n10645), .ZN(
        P1_U3490) );
  OAI22_X1 U11216 ( .A1(n10621), .A2(n10650), .B1(n4972), .B2(n10648), .ZN(
        n10623) );
  AOI211_X1 U11217 ( .C1(n10624), .C2(n10654), .A(n10623), .B(n10622), .ZN(
        n10625) );
  AOI22_X1 U11218 ( .A1(n10657), .A2(n10625), .B1(n6177), .B2(n10656), .ZN(
        P2_U3532) );
  AOI22_X1 U11219 ( .A1(n10660), .A2(n10625), .B1(n5775), .B2(n10658), .ZN(
        P2_U3487) );
  NAND3_X1 U11220 ( .A1(n4932), .A2(n10626), .A3(n10654), .ZN(n10633) );
  AOI22_X1 U11221 ( .A1(n10630), .A2(n10629), .B1(n10628), .B2(n10627), .ZN(
        n10631) );
  AOI22_X1 U11222 ( .A1(n10657), .A2(n10634), .B1(n6175), .B2(n10656), .ZN(
        P2_U3533) );
  AOI22_X1 U11223 ( .A1(n10660), .A2(n10634), .B1(n5790), .B2(n10658), .ZN(
        P2_U3490) );
  OAI211_X1 U11224 ( .C1(n10638), .C2(n10637), .A(n10636), .B(n10635), .ZN(
        n10639) );
  AOI21_X1 U11225 ( .B1(n10641), .B2(n10640), .A(n10639), .ZN(n10647) );
  AOI22_X1 U11226 ( .A1(n10644), .A2(n10647), .B1(n10643), .B2(n10642), .ZN(
        P1_U3537) );
  INV_X1 U11227 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10646) );
  AOI22_X1 U11228 ( .A1(n10491), .A2(n10647), .B1(n10646), .B2(n10645), .ZN(
        P1_U3496) );
  OAI22_X1 U11229 ( .A1(n10651), .A2(n10650), .B1(n10649), .B2(n10648), .ZN(
        n10652) );
  AOI211_X1 U11230 ( .C1(n10655), .C2(n10654), .A(n10653), .B(n10652), .ZN(
        n10659) );
  AOI22_X1 U11231 ( .A1(n10657), .A2(n10659), .B1(n6174), .B2(n10656), .ZN(
        P2_U3534) );
  AOI22_X1 U11232 ( .A1(n10660), .A2(n10659), .B1(n5803), .B2(n10658), .ZN(
        P2_U3493) );
  XNOR2_X1 U11233 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  AND2_X1 U4926 ( .A1(n6727), .A2(n7116), .ZN(n8188) );
  CLKBUF_X1 U4935 ( .A(n6788), .Z(n8145) );
  AND2_X1 U4965 ( .A1(n9971), .A2(n9970), .ZN(n10662) );
endmodule

