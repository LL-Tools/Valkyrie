

module b17_C_gen_AntiSAT_k_128_7 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput_f0, keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, 
        keyinput_f5, keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, 
        keyinput_f10, keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, 
        keyinput_f15, keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, 
        keyinput_f20, keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, 
        keyinput_f25, keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, 
        keyinput_f30, keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, 
        keyinput_f35, keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, 
        keyinput_f40, keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, 
        keyinput_f45, keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, 
        keyinput_f50, keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, 
        keyinput_f55, keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, 
        keyinput_f60, keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, 
        keyinput_g1, keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, 
        keyinput_g6, keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, 
        keyinput_g11, keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, 
        keyinput_g16, keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, 
        keyinput_g21, keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, 
        keyinput_g26, keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, 
        keyinput_g31, keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, 
        keyinput_g36, keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, 
        keyinput_g41, keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, 
        keyinput_g46, keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, 
        keyinput_g51, keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, 
        keyinput_g56, keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, 
        keyinput_g61, keyinput_g62, keyinput_g63, U355, U356, U357, U358, U359, 
        U360, U361, U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, 
        U373, U374, U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, 
        U376, U247, U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, 
        U236, U235, U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, 
        U224, U223, U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, 
        U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, 
        U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, 
        U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274, 
        P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, 
        P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, 
        P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, 
        P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, 
        P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, 
        P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, 
        P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, 
        P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, 
        P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, 
        P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, 
        P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, 
        P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, 
        P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, 
        P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, 
        P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, 
        P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, 
        P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, 
        P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, 
        P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, 
        P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, 
        P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, 
        P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, 
        P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, 
        P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, 
        P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, 
        P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, 
        P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, 
        P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, 
        P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, 
        P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, 
        P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, 
        P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, 
        P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, 
        P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, 
        P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, 
        P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, 
        P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, 
        P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, 
        P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, 
        P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, 
        P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, 
        P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, 
        P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, 
        P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, 
        P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, 
        P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, 
        P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, 
        P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, 
        P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, 
        P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, 
        P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, 
        P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, 
        P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, 
        P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, 
        P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, 
        P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, 
        P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, 
        P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, 
        P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, 
        P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, 
        P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, 
        P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, 
        P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, 
        P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, 
        P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, 
        P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, 
        P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, 
        P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, 
        P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, 
        P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, 
        P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, 
        P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, 
        P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, 
        P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, 
        P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, 
        P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, 
        P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, 
        P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, 
        P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, 
        P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, 
        P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, 
        P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, 
        P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, 
        P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, 
        P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, 
        P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, 
        P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, 
        P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, 
        P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, 
        P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, 
        P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, 
        P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, 
        P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, 
        P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, 
        P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, 
        P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, 
        P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, 
        P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, 
        P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, 
        P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, 
        P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, 
        P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, 
        P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, 
        P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, 
        P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, 
        P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, 
        P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, 
        P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, 
        P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, 
        P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, 
        P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, 
        P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, 
        P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, 
        P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, 
        P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, 
        P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, 
        P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, 
        P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, 
        P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, 
        P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, 
        P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, 
        P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, 
        P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, 
        P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, 
        P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, 
        P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, 
        P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, 
        P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, 
        P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, 
        P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, 
        P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, 
        P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, 
        P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, 
        P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, 
        P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, 
        P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, 
        P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, 
        P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, 
        P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, 
        P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, 
        P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, 
        P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, 
        P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, 
        P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, 
        P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, 
        P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, 
        P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, 
        P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, 
        P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, 
        P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, 
        P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, 
        P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, 
        P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, 
        P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, 
        P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, 
        P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, 
        P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, 
        P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, 
        P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, 
        P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, 
        P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, 
        P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, 
        P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, 
        P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, 
        P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, 
        P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, 
        P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, 
        P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, 
        P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, 
        P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, 
        P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, 
        P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, 
        P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, 
        P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, 
        P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, 
        P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, 
        P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, 
        P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, 
        P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, 
        P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, 
        P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9649, n9650, n9652, n9653, n9654, n9655, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
         n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
         n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
         n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
         n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,
         n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
         n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
         n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,
         n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
         n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,
         n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
         n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,
         n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
         n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,
         n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,
         n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16681, n16682, n16683, n16684, n16685,
         n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693,
         n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701,
         n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
         n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717,
         n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725,
         n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733,
         n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741,
         n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749,
         n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757,
         n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765,
         n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773,
         n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781,
         n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789,
         n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797,
         n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805,
         n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813,
         n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
         n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829,
         n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837,
         n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845,
         n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
         n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861,
         n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869,
         n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877,
         n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
         n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
         n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
         n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909,
         n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917,
         n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925,
         n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933,
         n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941,
         n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
         n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
         n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
         n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
         n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
         n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
         n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
         n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
         n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013,
         n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
         n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
         n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
         n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
         n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
         n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
         n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
         n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
         n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
         n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
         n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
         n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
         n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
         n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
         n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
         n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
         n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
         n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
         n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
         n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
         n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
         n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
         n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349,
         n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
         n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
         n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
         n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
         n17382, n17384, n17385, n17386, n17387, n17388, n17389, n17390,
         n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398,
         n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406,
         n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
         n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422,
         n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430,
         n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438,
         n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
         n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454,
         n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462,
         n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470,
         n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478,
         n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
         n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494,
         n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502,
         n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510,
         n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
         n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526,
         n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534,
         n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542,
         n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550,
         n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
         n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566,
         n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574,
         n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
         n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
         n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
         n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
         n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
         n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
         n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
         n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638,
         n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646,
         n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
         n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
         n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
         n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
         n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
         n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
         n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782,
         n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
         n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
         n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
         n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
         n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
         n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
         n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
         n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
         n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854,
         n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
         n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
         n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
         n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886,
         n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
         n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
         n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
         n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
         n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006,
         n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
         n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
         n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
         n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
         n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
         n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
         n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
         n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
         n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
         n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
         n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142,
         n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150,
         n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
         n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
         n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
         n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
         n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
         n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
         n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
         n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
         n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
         n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
         n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278,
         n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286,
         n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
         n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
         n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
         n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
         n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342,
         n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
         n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358,
         n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366,
         n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374,
         n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
         n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
         n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398,
         n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
         n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414,
         n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422,
         n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430,
         n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438,
         n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446,
         n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454,
         n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462,
         n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470,
         n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
         n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486,
         n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494,
         n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502,
         n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510,
         n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518,
         n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526,
         n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534,
         n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542,
         n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
         n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558,
         n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566,
         n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574,
         n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582,
         n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
         n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
         n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
         n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614,
         n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
         n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630,
         n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638,
         n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
         n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654,
         n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662,
         n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
         n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678,
         n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686,
         n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694,
         n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702,
         n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
         n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718,
         n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726,
         n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734,
         n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
         n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750,
         n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758,
         n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766,
         n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774,
         n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782,
         n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790,
         n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798,
         n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806,
         n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814,
         n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822,
         n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830,
         n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838,
         n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846,
         n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
         n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862,
         n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870,
         n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878,
         n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
         n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894,
         n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902,
         n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
         n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918,
         n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926,
         n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934,
         n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942,
         n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950,
         n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
         n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966,
         n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974,
         n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
         n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990,
         n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
         n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006,
         n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014,
         n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022,
         n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030,
         n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038,
         n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046,
         n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
         n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062,
         n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070,
         n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078,
         n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086,
         n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094,
         n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
         n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110,
         n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118,
         n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
         n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134,
         n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142,
         n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150,
         n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158,
         n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166,
         n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
         n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182,
         n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190,
         n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198,
         n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206,
         n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214,
         n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222,
         n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230,
         n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238,
         n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
         n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254,
         n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262,
         n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
         n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278,
         n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286,
         n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294,
         n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302,
         n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310,
         n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
         n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326,
         n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334,
         n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342,
         n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350,
         n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358,
         n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366,
         n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374,
         n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382,
         n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
         n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398,
         n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406,
         n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
         n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422,
         n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430,
         n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438,
         n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446,
         n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454,
         n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
         n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470,
         n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478,
         n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486,
         n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494,
         n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502,
         n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510,
         n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518,
         n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526,
         n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
         n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542,
         n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550,
         n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
         n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566,
         n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574,
         n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582,
         n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590,
         n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598,
         n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
         n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614,
         n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622,
         n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
         n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638,
         n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
         n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
         n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
         n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
         n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710,
         n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
         n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726,
         n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734,
         n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
         n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
         n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758,
         n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766,
         n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
         n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
         n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
         n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
         n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806,
         n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
         n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
         n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830,
         n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838,
         n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
         n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
         n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
         n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870,
         n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
         n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
         n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902,
         n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
         n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
         n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926,
         n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934,
         n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
         n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
         n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
         n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
         n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
         n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982,
         n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
         n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014,
         n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
         n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
         n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
         n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
         n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
         n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142,
         n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
         n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158,
         n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
         n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
         n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
         n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190,
         n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198,
         n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
         n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
         n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
         n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
         n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
         n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246,
         n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
         n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262,
         n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270,
         n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
         n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
         n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
         n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342,
         n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
         n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
         n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
         n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
         n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
         n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
         n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
         n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
         n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
         n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
         n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
         n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
         n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574,
         n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
         n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590,
         n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
         n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
         n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718,
         n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
         n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734,
         n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742,
         n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
         n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
         n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766,
         n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774,
         n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
         n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790,
         n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
         n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806,
         n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814,
         n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822,
         n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
         n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838,
         n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846,
         n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854,
         n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862,
         n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
         n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878,
         n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886,
         n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894,
         n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
         n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910,
         n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918,
         n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
         n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934,
         n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942,
         n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950,
         n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958,
         n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966,
         n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
         n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982,
         n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990,
         n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998,
         n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006,
         n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014,
         n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022,
         n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030,
         n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038,
         n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
         n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054,
         n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062,
         n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070,
         n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078,
         n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086,
         n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094,
         n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102,
         n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110,
         n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118,
         n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126,
         n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134,
         n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142,
         n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150,
         n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158,
         n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166,
         n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174,
         n21175, n21176;

  INV_X1 U11093 ( .A(n17984), .ZN(n17996) );
  OR2_X1 U11094 ( .A1(n10047), .A2(n16133), .ZN(n9988) );
  XNOR2_X1 U11095 ( .A(n11709), .B(n12872), .ZN(n16133) );
  INV_X1 U11096 ( .A(n18449), .ZN(n17527) );
  AND2_X1 U11097 ( .A1(n10441), .A2(n13743), .ZN(n10648) );
  AND2_X1 U11098 ( .A1(n10148), .A2(n11603), .ZN(n9957) );
  XNOR2_X1 U11100 ( .A(n10434), .B(n10433), .ZN(n10435) );
  AOI21_X1 U11101 ( .B1(n11598), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11599), .ZN(n11606) );
  CLKBUF_X3 U11102 ( .A(n10871), .Z(n9659) );
  AND2_X1 U11104 ( .A1(n12587), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10534) );
  AOI21_X1 U11105 ( .B1(n11525), .B2(n11512), .A(n11527), .ZN(n12867) );
  INV_X1 U11106 ( .A(n12918), .ZN(n17382) );
  CLKBUF_X2 U11107 ( .A(n11430), .Z(n12206) );
  INV_X2 U11108 ( .A(n17355), .ZN(n17376) );
  INV_X4 U11109 ( .A(n17358), .ZN(n17392) );
  NAND2_X1 U11110 ( .A1(n12742), .A2(n12864), .ZN(n14486) );
  CLKBUF_X1 U11111 ( .A(n11505), .Z(n20347) );
  NOR2_X2 U11112 ( .A1(n11499), .A2(n11588), .ZN(n11511) );
  INV_X1 U11113 ( .A(n11494), .ZN(n11510) );
  INV_X1 U11114 ( .A(n10361), .ZN(n19416) );
  NAND2_X1 U11115 ( .A1(n10264), .A2(n10263), .ZN(n10361) );
  AND2_X1 U11116 ( .A1(n11360), .A2(n11365), .ZN(n11414) );
  AND2_X1 U11117 ( .A1(n13681), .A2(n11366), .ZN(n11430) );
  AND2_X1 U11118 ( .A1(n13702), .A2(n11355), .ZN(n11569) );
  AND2_X1 U11119 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11365) );
  NOR2_X1 U11121 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10252) );
  AND2_X1 U11123 ( .A1(n11366), .A2(n11360), .ZN(n11399) );
  AND2_X1 U11125 ( .A1(n13702), .A2(n13704), .ZN(n11413) );
  AND2_X1 U11126 ( .A1(n11507), .A2(n11506), .ZN(n11509) );
  NAND2_X1 U11127 ( .A1(n13361), .A2(n13357), .ZN(n12840) );
  NAND4_X1 U11128 ( .A1(n11394), .A2(n11393), .A3(n11392), .A4(n11391), .ZN(
        n11437) );
  AND2_X1 U11129 ( .A1(n9683), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12563) );
  OR2_X1 U11130 ( .A1(n9671), .A2(n14458), .ZN(n10419) );
  NOR2_X1 U11131 ( .A1(n9832), .A2(n14800), .ZN(n14793) );
  BUF_X1 U11133 ( .A(n10578), .Z(n10974) );
  INV_X1 U11134 ( .A(n17585), .ZN(n13160) );
  NAND4_X1 U11135 ( .A1(n11492), .A2(n11491), .A3(n11490), .A4(n11489), .ZN(
        n11498) );
  NAND2_X1 U11136 ( .A1(n14372), .A2(n12019), .ZN(n14564) );
  INV_X2 U11137 ( .A(n13918), .ZN(n20316) );
  INV_X1 U11138 ( .A(n11498), .ZN(n20326) );
  NAND2_X1 U11140 ( .A1(n9649), .A2(n14045), .ZN(n13749) );
  INV_X2 U11141 ( .A(n17287), .ZN(n17320) );
  INV_X1 U11142 ( .A(n17396), .ZN(n9662) );
  INV_X1 U11143 ( .A(n18444), .ZN(n17436) );
  NAND2_X1 U11144 ( .A1(n17045), .A2(n19031), .ZN(n12896) );
  NAND2_X1 U11145 ( .A1(n13036), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17735) );
  INV_X1 U11146 ( .A(n13357), .ZN(n14485) );
  NOR2_X1 U11147 ( .A1(n14448), .A2(n14447), .ZN(n14449) );
  OR2_X1 U11149 ( .A1(n15429), .A2(n15428), .ZN(n15430) );
  CLKBUF_X2 U11150 ( .A(n10384), .Z(n9666) );
  OR2_X1 U11152 ( .A1(n9980), .A2(n13088), .ZN(n18449) );
  INV_X1 U11153 ( .A(n20165), .ZN(n20148) );
  AOI211_X1 U11154 ( .C1(n17217), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n12911), .B(n12910), .ZN(n17563) );
  INV_X1 U11155 ( .A(n18073), .ZN(n18065) );
  INV_X1 U11156 ( .A(n11281), .ZN(n9655) );
  AND2_X4 U11157 ( .A1(n10872), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9649) );
  INV_X1 U11158 ( .A(n13117), .ZN(n17268) );
  OR2_X2 U11160 ( .A1(n9994), .A2(n9991), .ZN(n9990) );
  XNOR2_X2 U11161 ( .A(n14488), .B(n14487), .ZN(n14826) );
  AND2_X4 U11162 ( .A1(n11734), .A2(n11745), .ZN(n16086) );
  OAI21_X2 U11163 ( .B1(n15227), .B2(n10130), .A(n10129), .ZN(n15165) );
  XNOR2_X2 U11164 ( .A(n12577), .B(n12600), .ZN(n15227) );
  XNOR2_X2 U11165 ( .A(n10677), .B(n14305), .ZN(n14298) );
  NAND2_X2 U11166 ( .A1(n10676), .A2(n19217), .ZN(n10677) );
  BUF_X2 U11167 ( .A(n10852), .Z(n9650) );
  BUF_X8 U11169 ( .A(n10484), .Z(n9652) );
  AND2_X2 U11170 ( .A1(n10252), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10484) );
  INV_X1 U11171 ( .A(n12938), .ZN(n14414) );
  NOR2_X2 U11172 ( .A1(n12899), .A2(n12896), .ZN(n12938) );
  AND2_X4 U11173 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10872) );
  BUF_X4 U11174 ( .A(n12968), .Z(n9653) );
  INV_X1 U11175 ( .A(n17367), .ZN(n12968) );
  NOR2_X4 U11176 ( .A1(n10768), .A2(n10766), .ZN(n10761) );
  OAI211_X2 U11177 ( .C1(n9994), .C2(n9992), .A(n9990), .B(n9993), .ZN(n10768)
         );
  INV_X1 U11178 ( .A(n9649), .ZN(n9654) );
  INV_X2 U11180 ( .A(n9655), .ZN(n9657) );
  NOR2_X2 U11181 ( .A1(n15041), .A2(n11067), .ZN(n15044) );
  AND2_X1 U11182 ( .A1(n9961), .A2(n9960), .ZN(n14717) );
  NAND2_X1 U11183 ( .A1(n15302), .A2(n15301), .ZN(n15303) );
  NAND2_X2 U11184 ( .A1(n11752), .A2(n9732), .ZN(n14815) );
  NAND2_X1 U11185 ( .A1(n13790), .A2(n13789), .ZN(n13791) );
  AND2_X1 U11187 ( .A1(n14536), .A2(n14522), .ZN(n14524) );
  INV_X4 U11188 ( .A(n18080), .ZN(n18039) );
  AND2_X1 U11189 ( .A1(n10446), .A2(n13743), .ZN(n10649) );
  NAND2_X1 U11190 ( .A1(n10800), .A2(n10820), .ZN(n10799) );
  NOR2_X1 U11191 ( .A1(n10459), .A2(n10445), .ZN(n10464) );
  AND2_X1 U11192 ( .A1(n18272), .A2(n17959), .ZN(n17995) );
  INV_X2 U11193 ( .A(n18843), .ZN(n18252) );
  OAI21_X1 U11194 ( .B1(n11840), .B2(n9837), .A(n9835), .ZN(n9838) );
  NAND2_X1 U11195 ( .A1(n10374), .A2(n10373), .ZN(n10410) );
  OAI21_X1 U11196 ( .B1(n11304), .B2(n10401), .A(n14901), .ZN(n10392) );
  AND2_X1 U11197 ( .A1(n13325), .A2(n13323), .ZN(n12739) );
  AND2_X1 U11198 ( .A1(n10364), .A2(n10363), .ZN(n11180) );
  INV_X1 U11199 ( .A(n10415), .ZN(n10427) );
  AND2_X1 U11200 ( .A1(n10390), .A2(n10880), .ZN(n11179) );
  INV_X2 U11201 ( .A(n11526), .ZN(n11512) );
  AND2_X1 U11202 ( .A1(n10356), .A2(n19411), .ZN(n11314) );
  INV_X1 U11205 ( .A(n11437), .ZN(n11505) );
  BUF_X2 U11206 ( .A(n11508), .Z(n14479) );
  INV_X1 U11207 ( .A(n10366), .ZN(n9658) );
  AND3_X1 U11208 ( .A1(n11412), .A2(n11411), .A3(n10249), .ZN(n10251) );
  INV_X1 U11209 ( .A(n13080), .ZN(n17303) );
  BUF_X2 U11210 ( .A(n11569), .Z(n12300) );
  CLKBUF_X2 U11211 ( .A(n11414), .Z(n12295) );
  AND2_X2 U11212 ( .A1(n11360), .A2(n13707), .ZN(n11612) );
  AND2_X4 U11213 ( .A1(n13681), .A2(n11365), .ZN(n11422) );
  INV_X2 U11214 ( .A(n13246), .ZN(n9660) );
  INV_X4 U11215 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17045) );
  INV_X2 U11216 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14069) );
  AND2_X1 U11217 ( .A1(n13320), .A2(n13321), .ZN(n9913) );
  OAI21_X1 U11218 ( .B1(n12339), .B2(n10207), .A(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10204) );
  AND2_X1 U11219 ( .A1(n14728), .A2(n10041), .ZN(n12387) );
  AND2_X1 U11220 ( .A1(n14738), .A2(n9745), .ZN(n9960) );
  NOR2_X1 U11221 ( .A1(n14755), .A2(n12707), .ZN(n12711) );
  OR2_X1 U11222 ( .A1(n14748), .A2(n16143), .ZN(n14756) );
  XNOR2_X1 U11223 ( .A(n12395), .B(n12394), .ZN(n14489) );
  NOR2_X1 U11224 ( .A1(n15320), .A2(n15555), .ZN(n15560) );
  NOR2_X1 U11225 ( .A1(n15354), .A2(n15351), .ZN(n15344) );
  NAND2_X1 U11226 ( .A1(n15303), .A2(n10197), .ZN(n10196) );
  AND2_X1 U11227 ( .A1(n15929), .A2(n15928), .ZN(n16068) );
  INV_X1 U11228 ( .A(n9901), .ZN(n15354) );
  AOI21_X1 U11229 ( .B1(n19189), .B2(n14933), .A(n14932), .ZN(n14934) );
  AND2_X1 U11230 ( .A1(n15412), .A2(n15411), .ZN(n10246) );
  NAND2_X1 U11231 ( .A1(n10804), .A2(n15513), .ZN(n15302) );
  OAI21_X1 U11232 ( .B1(n16391), .B2(n15306), .A(n16389), .ZN(n15382) );
  CLKBUF_X1 U11233 ( .A(n14768), .Z(n16163) );
  NAND2_X1 U11234 ( .A1(n14606), .A2(n14607), .ZN(n14604) );
  AND2_X1 U11235 ( .A1(n13266), .A2(n13265), .ZN(n15407) );
  XNOR2_X1 U11236 ( .A(n13265), .B(n11177), .ZN(n16306) );
  OR2_X1 U11237 ( .A1(n14450), .A2(n14449), .ZN(n16317) );
  NAND2_X1 U11238 ( .A1(n14448), .A2(n12364), .ZN(n15197) );
  OR2_X1 U11239 ( .A1(n10608), .A2(n9919), .ZN(n9916) );
  NOR2_X1 U11240 ( .A1(n9710), .A2(n9822), .ZN(n9821) );
  OR2_X1 U11241 ( .A1(n17765), .A2(n13034), .ZN(n13035) );
  OAI21_X1 U11242 ( .B1(n10926), .B2(n11014), .A(n15111), .ZN(n10608) );
  NAND2_X1 U11243 ( .A1(n10209), .A2(n9716), .ZN(n10952) );
  NOR2_X1 U11244 ( .A1(n10016), .A2(n9723), .ZN(n10015) );
  AND2_X1 U11245 ( .A1(n14793), .A2(n10012), .ZN(n11759) );
  XNOR2_X1 U11246 ( .A(n10845), .B(n10844), .ZN(n14933) );
  NOR2_X1 U11247 ( .A1(n19859), .A2(n20071), .ZN(n19795) );
  NAND2_X1 U11248 ( .A1(n10714), .A2(n10713), .ZN(n10953) );
  OAI21_X1 U11249 ( .B1(n9844), .B2(n9846), .A(n10557), .ZN(n10560) );
  OR3_X1 U11250 ( .A1(n10698), .A2(n10697), .A3(n10696), .ZN(n10714) );
  NOR2_X1 U11251 ( .A1(n16568), .A2(n17887), .ZN(n17742) );
  NAND2_X1 U11252 ( .A1(n17980), .A2(n18187), .ZN(n17887) );
  NOR2_X1 U11253 ( .A1(n13025), .A2(n17873), .ZN(n17869) );
  XNOR2_X1 U11254 ( .A(n11734), .B(n11733), .ZN(n11885) );
  NOR2_X1 U11255 ( .A1(n10797), .A2(n9924), .ZN(n9923) );
  NOR2_X1 U11256 ( .A1(n13832), .A2(n13833), .ZN(n15047) );
  AND2_X1 U11257 ( .A1(n14589), .A2(n14534), .ZN(n14536) );
  NAND2_X1 U11258 ( .A1(n9839), .A2(n11723), .ZN(n11734) );
  AOI22_X1 U11259 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10637), .B1(
        n10511), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10518) );
  NAND2_X1 U11260 ( .A1(n17559), .A2(n18074), .ZN(n17999) );
  NAND2_X1 U11261 ( .A1(n10820), .A2(n9707), .ZN(n10850) );
  INV_X1 U11262 ( .A(n11725), .ZN(n9839) );
  NAND2_X1 U11263 ( .A1(n17757), .A2(n18080), .ZN(n17830) );
  AND2_X1 U11264 ( .A1(n19800), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n9849) );
  INV_X1 U11265 ( .A(n13026), .ZN(n17798) );
  INV_X1 U11266 ( .A(n18070), .ZN(n18084) );
  INV_X1 U11267 ( .A(n11662), .ZN(n11636) );
  NOR3_X1 U11268 ( .A1(n10808), .A2(n10807), .A3(P2_EBX_REG_24__SCAN_IN), .ZN(
        n10822) );
  OR2_X1 U11269 ( .A1(n10808), .A2(n10807), .ZN(n10810) );
  CLKBUF_X1 U11270 ( .A(n13344), .Z(n14708) );
  NOR2_X1 U11271 ( .A1(n10470), .A2(n10473), .ZN(n19800) );
  NOR2_X2 U11272 ( .A1(n10472), .A2(n10473), .ZN(n10637) );
  INV_X1 U11273 ( .A(n19666), .ZN(n19663) );
  OR2_X1 U11274 ( .A1(n10456), .A2(n13653), .ZN(n10650) );
  AND2_X1 U11275 ( .A1(n10464), .A2(n10461), .ZN(n19666) );
  NOR2_X1 U11276 ( .A1(n20475), .A2(n20327), .ZN(n20834) );
  NOR2_X1 U11277 ( .A1(n20475), .A2(n20332), .ZN(n20840) );
  AND2_X1 U11278 ( .A1(n10450), .A2(n15129), .ZN(n19704) );
  NOR2_X1 U11279 ( .A1(n20475), .A2(n20317), .ZN(n20821) );
  AND2_X1 U11280 ( .A1(n10450), .A2(n13653), .ZN(n19829) );
  OR2_X2 U11281 ( .A1(n18848), .A2(n18904), .ZN(n16696) );
  NOR2_X1 U11282 ( .A1(n20475), .A2(n20340), .ZN(n20846) );
  AND2_X1 U11283 ( .A1(n13743), .A2(n10447), .ZN(n19446) );
  NAND2_X1 U11284 ( .A1(n17994), .A2(n17959), .ZN(n17931) );
  NAND2_X1 U11285 ( .A1(n10799), .A2(n10798), .ZN(n10808) );
  OAI21_X1 U11286 ( .B1(n10459), .B2(n12426), .A(n12425), .ZN(n13737) );
  OR2_X1 U11287 ( .A1(n10459), .A2(n10455), .ZN(n10456) );
  NAND2_X2 U11288 ( .A1(n14711), .A2(n13816), .ZN(n14715) );
  CLKBUF_X1 U11289 ( .A(n13866), .Z(n9675) );
  NAND2_X1 U11290 ( .A1(n11661), .A2(n11660), .ZN(n13874) );
  NAND2_X1 U11291 ( .A1(n17995), .A2(n10059), .ZN(n17994) );
  NAND2_X1 U11292 ( .A1(n9864), .A2(n9863), .ZN(n10459) );
  NAND2_X1 U11293 ( .A1(n17658), .A2(n18233), .ZN(n18843) );
  INV_X1 U11294 ( .A(n10460), .ZN(n10473) );
  OR2_X1 U11295 ( .A1(n15033), .A2(n10961), .ZN(n10792) );
  AND2_X1 U11296 ( .A1(n9824), .A2(n9734), .ZN(n11833) );
  NAND2_X1 U11297 ( .A1(n12416), .A2(n12415), .ZN(n13601) );
  CLKBUF_X1 U11298 ( .A(n14642), .Z(n14633) );
  NAND2_X1 U11299 ( .A1(n9862), .A2(n11183), .ZN(n9863) );
  OR2_X2 U11300 ( .A1(n14011), .A2(n13943), .ZN(n14193) );
  OAI21_X1 U11301 ( .B1(n11838), .B2(n11743), .A(n11591), .ZN(n13665) );
  AND2_X1 U11302 ( .A1(n10757), .A2(n10753), .ZN(n10782) );
  INV_X2 U11303 ( .A(n19252), .ZN(n19259) );
  CLKBUF_X1 U11304 ( .A(n12408), .Z(n15129) );
  NAND2_X1 U11305 ( .A1(n9838), .A2(n11744), .ZN(n11629) );
  NAND2_X1 U11306 ( .A1(n18387), .A2(n18859), .ZN(n18309) );
  NAND2_X1 U11307 ( .A1(n9955), .A2(n9954), .ZN(n11607) );
  NOR2_X1 U11308 ( .A1(n18007), .A2(n18324), .ZN(n18006) );
  NAND2_X1 U11309 ( .A1(n10009), .A2(n11537), .ZN(n11538) );
  OAI211_X1 U11310 ( .C1(n18017), .C2(n10074), .A(n10072), .B(n10069), .ZN(
        n18007) );
  NOR2_X1 U11311 ( .A1(n10992), .A2(n10991), .ZN(n10998) );
  NOR2_X1 U11312 ( .A1(n18017), .A2(n18016), .ZN(n18015) );
  INV_X1 U11313 ( .A(n10820), .ZN(n9994) );
  NAND2_X1 U11314 ( .A1(n10422), .A2(n10421), .ZN(n10433) );
  OR2_X1 U11315 ( .A1(n10732), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10736) );
  AND2_X1 U11316 ( .A1(n13605), .A2(n13604), .ZN(n13607) );
  AND2_X1 U11317 ( .A1(n10071), .A2(n10070), .ZN(n10069) );
  NAND2_X1 U11318 ( .A1(n10982), .A2(n10981), .ZN(n13605) );
  AOI21_X1 U11319 ( .B1(n10407), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10406), 
        .ZN(n10408) );
  AND3_X1 U11320 ( .A1(n11536), .A2(n12867), .A3(n11535), .ZN(n11568) );
  NOR2_X1 U11321 ( .A1(n12594), .A2(n14114), .ZN(n12419) );
  INV_X4 U11322 ( .A(n10427), .ZN(n11188) );
  NAND2_X1 U11323 ( .A1(n11180), .A2(n11314), .ZN(n13752) );
  AND2_X1 U11324 ( .A1(n10417), .A2(n10416), .ZN(n10418) );
  NAND2_X1 U11325 ( .A1(n10378), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10400) );
  AND2_X1 U11326 ( .A1(n11623), .A2(n9836), .ZN(n9835) );
  AND2_X2 U11327 ( .A1(n10389), .A2(n10369), .ZN(n11281) );
  AND2_X1 U11328 ( .A1(n10370), .A2(n10369), .ZN(n10415) );
  INV_X1 U11329 ( .A(n11581), .ZN(n9837) );
  INV_X1 U11330 ( .A(n11724), .ZN(n11723) );
  AND2_X1 U11331 ( .A1(n14899), .A2(n10983), .ZN(n10369) );
  AND2_X1 U11332 ( .A1(n10723), .A2(n10007), .ZN(n10006) );
  XNOR2_X1 U11333 ( .A(n13010), .B(n13009), .ZN(n13011) );
  OR2_X1 U11334 ( .A1(n13357), .A2(n12742), .ZN(n12820) );
  NOR2_X1 U11335 ( .A1(n18424), .A2(n13150), .ZN(n13134) );
  NOR2_X1 U11336 ( .A1(n18444), .A2(n17446), .ZN(n18858) );
  OR2_X1 U11337 ( .A1(n13496), .A2(n10988), .ZN(n10982) );
  AND2_X1 U11338 ( .A1(n11493), .A2(n13959), .ZN(n11528) );
  AND2_X1 U11339 ( .A1(n10896), .A2(n11314), .ZN(n11311) );
  NOR2_X1 U11340 ( .A1(n10385), .A2(n10375), .ZN(n10389) );
  AND2_X1 U11341 ( .A1(n9861), .A2(n9859), .ZN(n10380) );
  AND2_X1 U11342 ( .A1(n11449), .A2(n11530), .ZN(n11450) );
  INV_X1 U11343 ( .A(n10591), .ZN(n13414) );
  NAND2_X2 U11344 ( .A1(n13267), .A2(n10975), .ZN(n11175) );
  NAND2_X1 U11345 ( .A1(n13115), .A2(n13114), .ZN(n18411) );
  OR2_X1 U11346 ( .A1(n12856), .A2(n11497), .ZN(n15877) );
  OAI211_X1 U11347 ( .C1(n17367), .C2(n17232), .A(n13079), .B(n13078), .ZN(
        n18424) );
  NAND4_X1 U11348 ( .A1(n10367), .A2(n9658), .A3(n19416), .A4(n13764), .ZN(
        n11318) );
  OAI211_X1 U11349 ( .C1(n17120), .C2(n15832), .A(n13069), .B(n13068), .ZN(
        n18439) );
  OAI211_X1 U11350 ( .C1(n17287), .C2(n17172), .A(n13059), .B(n13058), .ZN(
        n18444) );
  AND2_X1 U11351 ( .A1(n10367), .A2(n13279), .ZN(n13267) );
  INV_X2 U11352 ( .A(n10974), .ZN(n19422) );
  OAI211_X1 U11353 ( .C1(n17367), .C2(n17319), .A(n12936), .B(n12935), .ZN(
        n13155) );
  AOI211_X1 U11354 ( .C1(n17321), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n13077), .B(n13076), .ZN(n13078) );
  OAI211_X1 U11355 ( .C1(n15784), .C2(n17420), .A(n13101), .B(n13100), .ZN(
        n18429) );
  OR2_X1 U11356 ( .A1(n10556), .A2(n10555), .ZN(n10993) );
  NAND2_X1 U11357 ( .A1(n11498), .A2(n11588), .ZN(n12864) );
  AND2_X1 U11358 ( .A1(n12953), .A2(n12952), .ZN(n17578) );
  INV_X1 U11359 ( .A(n10917), .ZN(n19411) );
  AND2_X1 U11360 ( .A1(n9860), .A2(n10366), .ZN(n10883) );
  AND2_X1 U11361 ( .A1(n12925), .A2(n12924), .ZN(n17571) );
  OR2_X1 U11362 ( .A1(n10626), .A2(n10625), .ZN(n10976) );
  NAND2_X1 U11363 ( .A1(n9805), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18079) );
  INV_X1 U11364 ( .A(n10384), .ZN(n10973) );
  CLKBUF_X3 U11365 ( .A(n11498), .Z(n13943) );
  OR2_X1 U11366 ( .A1(n10669), .A2(n10668), .ZN(n11006) );
  NAND2_X1 U11367 ( .A1(n9857), .A2(n9856), .ZN(n10578) );
  AND2_X1 U11368 ( .A1(n10352), .A2(n10351), .ZN(n10384) );
  NAND2_X1 U11369 ( .A1(n10275), .A2(n10276), .ZN(n10917) );
  NAND2_X1 U11370 ( .A1(n10304), .A2(n10305), .ZN(n10366) );
  OR2_X1 U11371 ( .A1(n11448), .A2(n11447), .ZN(n11588) );
  AND4_X1 U11372 ( .A1(n11479), .A2(n11478), .A3(n11477), .A4(n11476), .ZN(
        n11491) );
  AND4_X1 U11373 ( .A1(n11455), .A2(n11454), .A3(n11453), .A4(n11452), .ZN(
        n11471) );
  OR2_X2 U11374 ( .A1(n16645), .A2(n16600), .ZN(n16647) );
  AND4_X1 U11375 ( .A1(n11378), .A2(n11377), .A3(n11376), .A4(n11375), .ZN(
        n11394) );
  INV_X2 U11376 ( .A(U212), .ZN(n16630) );
  AND4_X1 U11377 ( .A1(n11364), .A2(n11363), .A3(n11362), .A4(n11361), .ZN(
        n11372) );
  AND4_X1 U11378 ( .A1(n11354), .A2(n11353), .A3(n11352), .A4(n11351), .ZN(
        n11374) );
  AND4_X1 U11379 ( .A1(n11459), .A2(n11458), .A3(n11457), .A4(n11456), .ZN(
        n11470) );
  AND4_X1 U11380 ( .A1(n11463), .A2(n11462), .A3(n11461), .A4(n11460), .ZN(
        n11469) );
  CLKBUF_X3 U11381 ( .A(n13039), .Z(n17374) );
  AND4_X1 U11382 ( .A1(n11475), .A2(n11474), .A3(n11473), .A4(n11472), .ZN(
        n11492) );
  AND4_X1 U11383 ( .A1(n11467), .A2(n11466), .A3(n11465), .A4(n11464), .ZN(
        n11468) );
  AND4_X1 U11384 ( .A1(n11386), .A2(n11385), .A3(n11384), .A4(n11383), .ZN(
        n11392) );
  AND4_X1 U11385 ( .A1(n11390), .A2(n11389), .A3(n11388), .A4(n11387), .ZN(
        n11391) );
  AND4_X1 U11386 ( .A1(n11359), .A2(n11358), .A3(n11357), .A4(n11356), .ZN(
        n11373) );
  INV_X4 U11387 ( .A(n14414), .ZN(n17336) );
  AND4_X1 U11388 ( .A1(n11382), .A2(n11381), .A3(n11380), .A4(n11379), .ZN(
        n11393) );
  INV_X2 U11389 ( .A(n19198), .ZN(n19214) );
  BUF_X2 U11390 ( .A(n11413), .Z(n12120) );
  NAND2_X2 U11391 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20108), .ZN(n20058) );
  INV_X2 U11392 ( .A(n15833), .ZN(n17385) );
  NAND2_X2 U11393 ( .A1(n20108), .A2(n20011), .ZN(n20061) );
  NAND2_X2 U11394 ( .A1(n19070), .A2(n19059), .ZN(n18380) );
  INV_X2 U11395 ( .A(n17355), .ZN(n17306) );
  AND2_X1 U11396 ( .A1(n10481), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10871) );
  NAND2_X2 U11397 ( .A1(n19000), .A2(n18933), .ZN(n18985) );
  AND2_X2 U11398 ( .A1(n9677), .A2(n10588), .ZN(n13249) );
  OR2_X2 U11399 ( .A1(n20980), .A2(n20894), .ZN(n20884) );
  BUF_X2 U11400 ( .A(n11399), .Z(n11480) );
  CLKBUF_X1 U11401 ( .A(n15220), .Z(n14107) );
  AND2_X1 U11402 ( .A1(n10278), .A2(n10277), .ZN(n10279) );
  INV_X1 U11403 ( .A(n9678), .ZN(n9682) );
  AND2_X2 U11404 ( .A1(n10481), .A2(n14045), .ZN(n12556) );
  OR2_X1 U11405 ( .A1(n12896), .A2(n12900), .ZN(n15833) );
  NOR2_X1 U11406 ( .A1(n17060), .A2(n12900), .ZN(n12990) );
  OR2_X2 U11407 ( .A1(n12899), .A2(n12901), .ZN(n17396) );
  OR3_X2 U11408 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n12901), .ZN(n17355) );
  INV_X2 U11409 ( .A(n16686), .ZN(n16688) );
  NAND2_X1 U11410 ( .A1(n12897), .A2(n19014), .ZN(n17287) );
  CLKBUF_X2 U11411 ( .A(n10490), .Z(n9677) );
  NAND2_X2 U11412 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12897), .ZN(
        n17367) );
  NAND4_X2 U11413 ( .A1(n19025), .A2(n19031), .A3(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A4(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17358) );
  AND3_X1 U11414 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n12895), .ZN(n12897) );
  NAND2_X1 U11415 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19025), .ZN(
        n12899) );
  AND2_X2 U11416 ( .A1(n13704), .A2(n11365), .ZN(n12267) );
  AND2_X2 U11417 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13704) );
  INV_X2 U11418 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n19025) );
  AND2_X1 U11419 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17078) );
  BUF_X1 U11420 ( .A(n17657), .Z(n9661) );
  NOR4_X1 U11421 ( .A1(n14411), .A2(n13135), .A3(n18439), .A4(n13138), .ZN(
        n17657) );
  INV_X1 U11422 ( .A(n9678), .ZN(n9681) );
  INV_X1 U11423 ( .A(n9678), .ZN(n9680) );
  XNOR2_X1 U11424 ( .A(n13608), .B(n12419), .ZN(n13602) );
  AND2_X1 U11425 ( .A1(n9677), .A2(n10588), .ZN(n9663) );
  AND2_X1 U11426 ( .A1(n9677), .A2(n10588), .ZN(n9664) );
  AND2_X1 U11427 ( .A1(n10761), .A2(n9766), .ZN(n10757) );
  NAND2_X1 U11428 ( .A1(n12409), .A2(n10357), .ZN(n12594) );
  INV_X1 U11429 ( .A(n17120), .ZN(n9665) );
  OR2_X1 U11430 ( .A1(n12901), .A2(n12900), .ZN(n17120) );
  NAND2_X1 U11431 ( .A1(n10578), .A2(n10354), .ZN(n10386) );
  AND4_X1 U11432 ( .A1(n9858), .A2(n10354), .A3(n10578), .A4(n10917), .ZN(
        n9859) );
  NOR2_X2 U11433 ( .A1(n14564), .A2(n10158), .ZN(n14617) );
  AND2_X1 U11434 ( .A1(n10459), .A2(n15709), .ZN(n10462) );
  NOR2_X2 U11435 ( .A1(n14321), .A2(n12789), .ZN(n14404) );
  NOR2_X1 U11436 ( .A1(n12899), .A2(n17060), .ZN(n9667) );
  NAND2_X1 U11437 ( .A1(n10436), .A2(n10423), .ZN(n10185) );
  NAND2_X2 U11438 ( .A1(n10414), .A2(n10413), .ZN(n10436) );
  INV_X1 U11439 ( .A(n10560), .ZN(n10558) );
  NOR2_X2 U11440 ( .A1(n14604), .A2(n10150), .ZN(n14584) );
  NOR2_X2 U11441 ( .A1(n15154), .A2(n12642), .ZN(n12664) );
  NOR2_X2 U11442 ( .A1(n15156), .A2(n15155), .ZN(n15154) );
  OR2_X2 U11443 ( .A1(n12664), .A2(n12663), .ZN(n15138) );
  INV_X1 U11444 ( .A(n11034), .ZN(n9668) );
  INV_X1 U11445 ( .A(n11034), .ZN(n9669) );
  NAND2_X1 U11446 ( .A1(n10983), .A2(n13484), .ZN(n11034) );
  AND2_X2 U11447 ( .A1(n14519), .A2(n12246), .ZN(n13306) );
  NOR2_X4 U11448 ( .A1(n14537), .A2(n14538), .ZN(n14519) );
  NAND2_X2 U11449 ( .A1(n15395), .A2(n10191), .ZN(n10190) );
  NAND2_X2 U11450 ( .A1(n10717), .A2(n10716), .ZN(n15395) );
  NAND2_X2 U11451 ( .A1(n11636), .A2(n11635), .ZN(n11830) );
  OAI211_X1 U11452 ( .C1(n11840), .C2(n10052), .A(n10050), .B(n10048), .ZN(
        n11838) );
  NAND3_X2 U11453 ( .A1(n10199), .A2(n10558), .A3(n10976), .ZN(n10937) );
  XNOR2_X2 U11454 ( .A(n10411), .B(n10410), .ZN(n10437) );
  NAND2_X1 U11455 ( .A1(n11300), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9671) );
  NAND2_X1 U11456 ( .A1(n11300), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9672) );
  NAND2_X1 U11457 ( .A1(n11300), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11286) );
  AND2_X1 U11458 ( .A1(n12336), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14899) );
  NOR2_X2 U11459 ( .A1(n14003), .A2(n14120), .ZN(n14119) );
  OAI21_X2 U11460 ( .B1(n12329), .B2(n15285), .A(n12328), .ZN(n12331) );
  NOR2_X2 U11461 ( .A1(n15165), .A2(n12601), .ZN(n12621) );
  INV_X1 U11462 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9673) );
  OAI21_X2 U11463 ( .B1(n10400), .B2(n10591), .A(n10396), .ZN(n10420) );
  NOR2_X2 U11464 ( .A1(n12699), .A2(n12698), .ZN(n13238) );
  NOR2_X4 U11465 ( .A1(n13909), .A2(n19236), .ZN(n14028) );
  NOR2_X2 U11466 ( .A1(n15171), .A2(n16339), .ZN(n12577) );
  INV_X1 U11467 ( .A(n10321), .ZN(n9678) );
  INV_X1 U11468 ( .A(n10321), .ZN(n9679) );
  INV_X1 U11469 ( .A(n9679), .ZN(n9683) );
  INV_X1 U11470 ( .A(n9679), .ZN(n9684) );
  AND3_X1 U11471 ( .A1(n14074), .A2(n9673), .A3(n14069), .ZN(n10321) );
  AND2_X1 U11472 ( .A1(n9677), .A2(n10588), .ZN(n9685) );
  OAI211_X2 U11473 ( .C1(n13735), .C2(n12428), .A(n12427), .B(n13738), .ZN(
        n13759) );
  OAI21_X2 U11474 ( .B1(n13669), .B2(n13670), .A(n12420), .ZN(n13735) );
  INV_X1 U11475 ( .A(n11710), .ZN(n10047) );
  NAND2_X1 U11476 ( .A1(n10367), .A2(n10357), .ZN(n10375) );
  NOR2_X1 U11477 ( .A1(n15877), .A2(n20971), .ZN(n12312) );
  NAND2_X1 U11478 ( .A1(n20245), .A2(n11594), .ZN(n11642) );
  NAND2_X1 U11479 ( .A1(n16127), .A2(n16126), .ZN(n9989) );
  NAND2_X1 U11480 ( .A1(n10430), .A2(n10429), .ZN(n11184) );
  INV_X1 U11481 ( .A(n11014), .ZN(n10961) );
  INV_X1 U11482 ( .A(n18429), .ZN(n13149) );
  NAND2_X1 U11483 ( .A1(n9661), .A2(n9969), .ZN(n9979) );
  NOR2_X1 U11484 ( .A1(n16082), .A2(n11762), .ZN(n9953) );
  NAND2_X1 U11485 ( .A1(n14815), .A2(n9821), .ZN(n9823) );
  INV_X1 U11486 ( .A(n11286), .ZN(n11298) );
  NOR2_X1 U11487 ( .A1(n19014), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12902) );
  INV_X2 U11488 ( .A(n17380), .ZN(n17321) );
  OR2_X1 U11489 ( .A1(n11549), .A2(n11548), .ZN(n11562) );
  INV_X1 U11490 ( .A(n10017), .ZN(n10016) );
  NAND2_X1 U11491 ( .A1(n9834), .A2(n11662), .ZN(n11711) );
  AND2_X1 U11492 ( .A1(n13874), .A2(n9952), .ZN(n9834) );
  OR2_X1 U11493 ( .A1(n11580), .A2(n11579), .ZN(n11747) );
  NAND2_X1 U11494 ( .A1(n9727), .A2(n11662), .ZN(n11725) );
  AND2_X1 U11495 ( .A1(n9986), .A2(n9952), .ZN(n9833) );
  NAND2_X1 U11496 ( .A1(n10377), .A2(n10376), .ZN(n10378) );
  NAND2_X1 U11497 ( .A1(n10169), .A2(n10375), .ZN(n10887) );
  AND2_X1 U11498 ( .A1(n19416), .A2(n10386), .ZN(n10169) );
  AND2_X1 U11499 ( .A1(n10375), .A2(n10386), .ZN(n10882) );
  NAND2_X1 U11500 ( .A1(n13155), .A2(n13005), .ZN(n13010) );
  NOR2_X1 U11501 ( .A1(n17578), .A2(n13160), .ZN(n13005) );
  NAND2_X1 U11502 ( .A1(n9805), .A2(n17585), .ZN(n13157) );
  NAND2_X1 U11503 ( .A1(n10154), .A2(n9781), .ZN(n10153) );
  INV_X1 U11504 ( .A(n14550), .ZN(n10154) );
  INV_X1 U11505 ( .A(n14374), .ZN(n10155) );
  NAND2_X1 U11506 ( .A1(n11531), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12016) );
  NAND2_X1 U11507 ( .A1(n16110), .A2(n10013), .ZN(n10012) );
  AOI21_X1 U11508 ( .B1(n20081), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10611), .ZN(n10854) );
  NOR2_X1 U11509 ( .A1(n10610), .A2(n10609), .ZN(n10611) );
  NAND2_X1 U11510 ( .A1(n10675), .A2(n10006), .ZN(n10733) );
  OAI21_X1 U11511 ( .B1(n9672), .B2(n16534), .A(n9853), .ZN(n11185) );
  AOI21_X1 U11512 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n11188), .A(n9854), .ZN(
        n9853) );
  NAND2_X1 U11513 ( .A1(n10428), .A2(n9855), .ZN(n9854) );
  NAND2_X1 U11514 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n9855) );
  INV_X1 U11515 ( .A(n10578), .ZN(n10367) );
  NAND2_X1 U11516 ( .A1(n10196), .A2(n9927), .ZN(n12329) );
  AND2_X1 U11517 ( .A1(n15469), .A2(n9995), .ZN(n9927) );
  INV_X1 U11518 ( .A(n15277), .ZN(n9995) );
  NOR2_X1 U11519 ( .A1(n10193), .A2(n15647), .ZN(n10191) );
  OR2_X1 U11520 ( .A1(n19174), .A2(n10961), .ZN(n10748) );
  NAND2_X1 U11521 ( .A1(n10955), .A2(n10954), .ZN(n10962) );
  AND2_X1 U11522 ( .A1(n11309), .A2(n10362), .ZN(n10363) );
  NOR2_X1 U11523 ( .A1(n18411), .A2(n17658), .ZN(n13142) );
  NAND2_X1 U11524 ( .A1(n13012), .A2(n17566), .ZN(n12987) );
  CLKBUF_X1 U11525 ( .A(n12912), .Z(n15784) );
  OR2_X1 U11526 ( .A1(n14470), .A2(n14477), .ZN(n13627) );
  NAND2_X1 U11527 ( .A1(n13329), .A2(n13328), .ZN(n13631) );
  INV_X1 U11528 ( .A(n12321), .ZN(n12392) );
  AND2_X1 U11529 ( .A1(n12391), .A2(n10167), .ZN(n10165) );
  AOI21_X1 U11530 ( .B1(n12264), .B2(n12263), .A(n12262), .ZN(n13307) );
  AND2_X1 U11531 ( .A1(n14435), .A2(n12289), .ZN(n12262) );
  NAND2_X1 U11532 ( .A1(n9961), .A2(n14738), .ZN(n14728) );
  NAND2_X1 U11533 ( .A1(n14331), .A2(n11749), .ZN(n11752) );
  NOR2_X1 U11534 ( .A1(n16127), .A2(n16126), .ZN(n9987) );
  NAND2_X1 U11535 ( .A1(n13791), .A2(n11643), .ZN(n11670) );
  INV_X1 U11536 ( .A(n20702), .ZN(n20824) );
  NAND2_X1 U11537 ( .A1(n10973), .A2(n12336), .ZN(n10591) );
  NAND2_X1 U11538 ( .A1(n10093), .A2(n16375), .ZN(n10092) );
  INV_X1 U11539 ( .A(n10095), .ZN(n10093) );
  AOI21_X1 U11540 ( .B1(n10085), .B2(n13435), .A(n10105), .ZN(n10095) );
  NAND2_X1 U11541 ( .A1(n11293), .A2(n11292), .ZN(n12381) );
  OR2_X1 U11542 ( .A1(n13737), .A2(n13736), .ZN(n13738) );
  AOI21_X1 U11543 ( .B1(n9897), .B2(n15307), .A(n9895), .ZN(n9894) );
  INV_X1 U11544 ( .A(n15309), .ZN(n9895) );
  NAND2_X1 U11545 ( .A1(n19926), .A2(n13484), .ZN(n19860) );
  AND2_X1 U11546 ( .A1(n12353), .A2(n14091), .ZN(n19936) );
  NOR2_X1 U11547 ( .A1(n15848), .A2(n14410), .ZN(n15939) );
  INV_X2 U11548 ( .A(n12928), .ZN(n17352) );
  INV_X1 U11549 ( .A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17302) );
  NAND2_X1 U11550 ( .A1(n15862), .A2(n16586), .ZN(n15917) );
  NOR2_X1 U11551 ( .A1(n17563), .A2(n12987), .ZN(n13228) );
  NAND2_X1 U11552 ( .A1(n17798), .A2(n17774), .ZN(n13028) );
  OAI211_X1 U11553 ( .C1(n17268), .C2(n17406), .A(n12986), .B(n12985), .ZN(
        n16559) );
  NAND2_X1 U11554 ( .A1(n15846), .A2(n15845), .ZN(n15852) );
  INV_X1 U11555 ( .A(n10472), .ZN(n10474) );
  AOI22_X1 U11556 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n11510), .B1(n11792), 
        .B2(n13943), .ZN(n11798) );
  INV_X1 U11557 ( .A(n10510), .ZN(n9850) );
  AND4_X1 U11558 ( .A1(n10469), .A2(n10468), .A3(n10467), .A4(n10466), .ZN(
        n10479) );
  AOI22_X1 U11559 ( .A1(n13249), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10284), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10286) );
  OR2_X1 U11560 ( .A1(n11682), .A2(n11681), .ZN(n11701) );
  NAND2_X1 U11561 ( .A1(n20347), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11649) );
  NAND2_X1 U11562 ( .A1(n11771), .A2(n20347), .ZN(n12859) );
  NAND2_X1 U11563 ( .A1(n11597), .A2(n11519), .ZN(n9827) );
  NOR2_X1 U11564 ( .A1(n11518), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9828) );
  NAND2_X1 U11565 ( .A1(n10590), .A2(n10589), .ZN(n10610) );
  INV_X1 U11566 ( .A(n10596), .ZN(n10867) );
  NAND3_X1 U11567 ( .A1(n14069), .A2(n14074), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13246) );
  AND2_X1 U11568 ( .A1(n9676), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12409) );
  INV_X1 U11569 ( .A(n13486), .ZN(n10896) );
  NAND2_X1 U11570 ( .A1(n13018), .A2(n10077), .ZN(n10076) );
  OAI21_X1 U11571 ( .B1(n13228), .B2(n16559), .A(n17819), .ZN(n13018) );
  NOR2_X1 U11572 ( .A1(n17571), .A2(n13167), .ZN(n13169) );
  INV_X1 U11573 ( .A(n13008), .ZN(n10058) );
  NOR2_X1 U11574 ( .A1(n17571), .A2(n13010), .ZN(n13012) );
  NOR2_X1 U11575 ( .A1(n14507), .A2(n10168), .ZN(n10167) );
  INV_X1 U11576 ( .A(n12312), .ZN(n12284) );
  NOR2_X1 U11577 ( .A1(n10161), .A2(n14630), .ZN(n10160) );
  INV_X1 U11578 ( .A(n10163), .ZN(n10161) );
  AND2_X1 U11579 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n11878), .ZN(
        n11886) );
  INV_X1 U11580 ( .A(n11879), .ZN(n11878) );
  AND2_X1 U11581 ( .A1(n16110), .A2(n14735), .ZN(n12707) );
  NAND3_X1 U11582 ( .A1(n9816), .A2(n9962), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n9961) );
  AND2_X1 U11583 ( .A1(n11758), .A2(n16095), .ZN(n10017) );
  NAND2_X1 U11584 ( .A1(n14404), .A2(n9756), .ZN(n9975) );
  INV_X1 U11585 ( .A(n14573), .ZN(n9973) );
  AND2_X1 U11586 ( .A1(n14804), .A2(n14802), .ZN(n14791) );
  NAND2_X1 U11587 ( .A1(n16110), .A2(n9748), .ZN(n11750) );
  NOR2_X1 U11588 ( .A1(n12766), .A2(n13926), .ZN(n9966) );
  INV_X1 U11589 ( .A(n11643), .ZN(n9820) );
  NAND2_X1 U11590 ( .A1(n11833), .A2(n13943), .ZN(n11567) );
  AOI21_X1 U11591 ( .B1(n11480), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A(
        n11484), .ZN(n11490) );
  AND2_X1 U11592 ( .A1(n11509), .A2(n14479), .ZN(n13676) );
  NAND2_X1 U11593 ( .A1(n10388), .A2(n10387), .ZN(n10863) );
  INV_X1 U11594 ( .A(n10386), .ZN(n10387) );
  AND2_X1 U11595 ( .A1(n9698), .A2(n9998), .ZN(n9997) );
  INV_X1 U11596 ( .A(n10770), .ZN(n9998) );
  NOR2_X1 U11597 ( .A1(n10008), .A2(n10718), .ZN(n10007) );
  INV_X1 U11598 ( .A(n10674), .ZN(n10008) );
  NAND2_X1 U11599 ( .A1(n10593), .A2(n10592), .ZN(n10594) );
  NAND2_X1 U11600 ( .A1(n10856), .A2(n10974), .ZN(n10593) );
  INV_X1 U11601 ( .A(n14964), .ZN(n10034) );
  INV_X1 U11602 ( .A(n15166), .ZN(n10132) );
  AND2_X1 U11603 ( .A1(n15505), .A2(n14983), .ZN(n10035) );
  NAND2_X1 U11604 ( .A1(n10143), .A2(n10139), .ZN(n15171) );
  NOR2_X1 U11605 ( .A1(n10140), .A2(n10146), .ZN(n10139) );
  INV_X1 U11606 ( .A(n15173), .ZN(n10146) );
  INV_X1 U11607 ( .A(n10141), .ZN(n10140) );
  INV_X1 U11608 ( .A(n15180), .ZN(n10145) );
  INV_X1 U11609 ( .A(n12568), .ZN(n12529) );
  INV_X1 U11610 ( .A(n15151), .ZN(n10187) );
  AND2_X1 U11611 ( .A1(n14954), .A2(n14968), .ZN(n10188) );
  INV_X1 U11612 ( .A(n13906), .ZN(n10174) );
  NOR2_X1 U11613 ( .A1(n10176), .A2(n13883), .ZN(n10175) );
  INV_X1 U11614 ( .A(n15633), .ZN(n10176) );
  OR2_X1 U11615 ( .A1(n10128), .A2(n16445), .ZN(n10127) );
  NAND2_X1 U11616 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10128) );
  NOR2_X1 U11617 ( .A1(n11318), .A2(n10368), .ZN(n10370) );
  NAND2_X1 U11618 ( .A1(n10402), .A2(n10401), .ZN(n10403) );
  NOR2_X1 U11619 ( .A1(n10973), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10975) );
  AND2_X1 U11620 ( .A1(n12330), .A2(n15267), .ZN(n10826) );
  OR2_X1 U11621 ( .A1(n16318), .A2(n10816), .ZN(n10836) );
  INV_X1 U11622 ( .A(n15363), .ZN(n9892) );
  OR2_X1 U11623 ( .A1(n10792), .A2(n11230), .ZN(n16389) );
  AOI21_X1 U11624 ( .B1(n9871), .B2(n9924), .A(n9869), .ZN(n9868) );
  INV_X1 U11625 ( .A(n15620), .ZN(n9869) );
  NOR2_X1 U11626 ( .A1(n15079), .A2(n10029), .ZN(n10028) );
  INV_X1 U11627 ( .A(n14273), .ZN(n10029) );
  NAND2_X1 U11628 ( .A1(n10182), .A2(n10181), .ZN(n10180) );
  INV_X1 U11629 ( .A(n13760), .ZN(n10181) );
  INV_X1 U11630 ( .A(n10183), .ZN(n10182) );
  INV_X1 U11631 ( .A(n14203), .ZN(n9915) );
  NAND2_X1 U11632 ( .A1(n16480), .A2(n10933), .ZN(n10940) );
  AND3_X1 U11633 ( .A1(n11307), .A2(n10892), .A3(n10891), .ZN(n11303) );
  NAND2_X1 U11634 ( .A1(n12412), .A2(n12411), .ZN(n12420) );
  AND2_X1 U11635 ( .A1(n13476), .A2(n13475), .ZN(n13540) );
  AOI22_X1 U11636 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12945), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13123) );
  NAND2_X1 U11637 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18000), .ZN(
        n13182) );
  INV_X1 U11638 ( .A(n10076), .ZN(n10073) );
  OR2_X1 U11639 ( .A1(n10076), .A2(n10075), .ZN(n10071) );
  NAND2_X1 U11640 ( .A1(n10078), .A2(n13017), .ZN(n10070) );
  INV_X1 U11641 ( .A(n18016), .ZN(n10075) );
  INV_X1 U11642 ( .A(n13018), .ZN(n10078) );
  NOR2_X1 U11643 ( .A1(n13176), .A2(n18011), .ZN(n13179) );
  NOR2_X1 U11644 ( .A1(n18036), .A2(n13168), .ZN(n13170) );
  INV_X1 U11645 ( .A(n9803), .ZN(n13166) );
  INV_X1 U11646 ( .A(n17571), .ZN(n13009) );
  NOR2_X1 U11647 ( .A1(n13004), .A2(n13003), .ZN(n13007) );
  XNOR2_X1 U11648 ( .A(n13160), .B(n17578), .ZN(n13002) );
  OR3_X1 U11649 ( .A1(n13135), .A2(n13151), .A3(n17446), .ZN(n14406) );
  NAND2_X1 U11650 ( .A1(n18434), .A2(n17436), .ZN(n13151) );
  INV_X1 U11651 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17232) );
  AOI21_X1 U11652 ( .B1(n18434), .B2(n15943), .A(n13129), .ZN(n16551) );
  NAND2_X1 U11653 ( .A1(n19055), .A2(n15844), .ZN(n17594) );
  NAND2_X1 U11654 ( .A1(n11647), .A2(n11646), .ZN(n20469) );
  OR2_X1 U11655 ( .A1(n13360), .A2(n14508), .ZN(n14510) );
  OR2_X1 U11656 ( .A1(n15913), .A2(n20971), .ZN(n13355) );
  NAND2_X2 U11657 ( .A1(n13331), .A2(n11508), .ZN(n13821) );
  AND2_X1 U11658 ( .A1(n14500), .A2(n12289), .ZN(n12317) );
  OR2_X1 U11659 ( .A1(n12286), .A2(n13311), .ZN(n12287) );
  INV_X1 U11660 ( .A(n10168), .ZN(n10166) );
  NAND2_X1 U11661 ( .A1(n12241), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12286) );
  NAND2_X1 U11662 ( .A1(n12198), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12239) );
  NAND2_X1 U11663 ( .A1(n10151), .A2(n14594), .ZN(n10150) );
  INV_X1 U11664 ( .A(n10153), .ZN(n10151) );
  AND2_X1 U11665 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n12112), .ZN(
        n12113) );
  INV_X1 U11666 ( .A(n12111), .ZN(n12112) );
  INV_X1 U11667 ( .A(n14645), .ZN(n12019) );
  AOI21_X1 U11668 ( .B1(n11875), .B2(n11967), .A(n11874), .ZN(n13931) );
  NAND2_X1 U11669 ( .A1(n11867), .A2(n11866), .ZN(n10147) );
  NAND2_X1 U11670 ( .A1(n14524), .A2(n12843), .ZN(n13360) );
  NOR2_X1 U11671 ( .A1(n12708), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10054) );
  NAND2_X1 U11672 ( .A1(n14404), .A2(n9974), .ZN(n14650) );
  AND2_X1 U11673 ( .A1(n16086), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14792) );
  OR2_X1 U11674 ( .A1(n14801), .A2(n16102), .ZN(n9832) );
  INV_X1 U11675 ( .A(n16120), .ZN(n9810) );
  NAND2_X1 U11676 ( .A1(n9809), .A2(n16120), .ZN(n9808) );
  INV_X1 U11677 ( .A(n10044), .ZN(n9809) );
  AND2_X1 U11678 ( .A1(n11730), .A2(n11729), .ZN(n16127) );
  NOR2_X1 U11679 ( .A1(n20958), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12324) );
  NAND2_X1 U11680 ( .A1(n16134), .A2(n16133), .ZN(n16132) );
  OR2_X1 U11681 ( .A1(n20305), .A2(n11743), .ZN(n11669) );
  AND2_X1 U11682 ( .A1(n12735), .A2(n14483), .ZN(n12874) );
  INV_X1 U11683 ( .A(n11538), .ZN(n9954) );
  AOI21_X1 U11684 ( .B1(n11833), .B2(n11832), .A(n11632), .ZN(n11634) );
  NOR2_X1 U11685 ( .A1(n11629), .A2(n11631), .ZN(n11632) );
  INV_X1 U11686 ( .A(n20553), .ZN(n20549) );
  NOR2_X1 U11687 ( .A1(n20475), .A2(n20709), .ZN(n20640) );
  OR2_X1 U11688 ( .A1(n11830), .A2(n13875), .ZN(n20702) );
  AOI21_X1 U11689 ( .B1(n20751), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20475), 
        .ZN(n20827) );
  NAND2_X1 U11690 ( .A1(n11823), .A2(n11822), .ZN(n14477) );
  OR2_X1 U11691 ( .A1(n11810), .A2(n11781), .ZN(n11823) );
  AOI221_X1 U11692 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n10854), 
        .C1(n13490), .C2(n10854), .A(n10853), .ZN(n10915) );
  NAND2_X2 U11693 ( .A1(n10340), .A2(n10339), .ZN(n12336) );
  NAND2_X1 U11694 ( .A1(n10333), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10340) );
  NAND2_X1 U11695 ( .A1(n13433), .A2(n10121), .ZN(n13442) );
  AND2_X1 U11696 ( .A1(n9703), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10121) );
  AND2_X1 U11697 ( .A1(n16375), .A2(n13435), .ZN(n10094) );
  AOI21_X1 U11699 ( .B1(n13426), .B2(n10104), .A(n10103), .ZN(n10102) );
  INV_X1 U11700 ( .A(n19113), .ZN(n10103) );
  INV_X1 U11701 ( .A(n19131), .ZN(n10104) );
  NOR2_X1 U11702 ( .A1(n14091), .A2(n10970), .ZN(n13387) );
  NAND2_X1 U11703 ( .A1(n10761), .A2(n9997), .ZN(n10773) );
  INV_X1 U11704 ( .A(n10736), .ZN(n9992) );
  AOI21_X1 U11705 ( .B1(n10820), .B2(P2_EBX_REG_11__SCAN_IN), .A(n9689), .ZN(
        n9993) );
  NOR2_X1 U11706 ( .A1(n10736), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10737) );
  NAND2_X1 U11707 ( .A1(n10737), .A2(n13886), .ZN(n10746) );
  INV_X1 U11708 ( .A(n13911), .ZN(n10137) );
  AND2_X1 U11709 ( .A1(n9652), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12562) );
  AND2_X1 U11710 ( .A1(n9652), .A2(n14045), .ZN(n12569) );
  NAND2_X1 U11711 ( .A1(n19253), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10138) );
  NAND2_X1 U11712 ( .A1(n10185), .A2(n10426), .ZN(n9862) );
  INV_X1 U11713 ( .A(n15220), .ZN(n14108) );
  INV_X1 U11714 ( .A(n9887), .ZN(n9883) );
  NOR2_X1 U11715 ( .A1(n13382), .A2(n19187), .ZN(n13385) );
  INV_X1 U11716 ( .A(n10236), .ZN(n9910) );
  NOR2_X1 U11717 ( .A1(n15422), .A2(n12341), .ZN(n9842) );
  INV_X1 U11718 ( .A(n15380), .ZN(n9898) );
  NOR2_X1 U11719 ( .A1(n9926), .A2(n15626), .ZN(n9925) );
  INV_X1 U11720 ( .A(n15680), .ZN(n10194) );
  OR2_X1 U11721 ( .A1(n15395), .A2(n10730), .ZN(n10195) );
  OR3_X1 U11722 ( .A1(n10962), .A2(n10961), .A3(n11205), .ZN(n10963) );
  NAND2_X1 U11723 ( .A1(n10607), .A2(n16534), .ZN(n9918) );
  NOR2_X1 U11724 ( .A1(n10607), .A2(n16534), .ZN(n9919) );
  AND2_X1 U11725 ( .A1(n13618), .A2(n14057), .ZN(n10971) );
  INV_X1 U11726 ( .A(n10608), .ZN(n9917) );
  NAND2_X1 U11727 ( .A1(n14068), .A2(n12414), .ZN(n12416) );
  AND3_X1 U11728 ( .A1(n11317), .A2(n11316), .A3(n11315), .ZN(n14066) );
  OR2_X1 U11729 ( .A1(n20074), .A2(n19541), .ZN(n19634) );
  OR2_X1 U11730 ( .A1(n20074), .A2(n20101), .ZN(n19627) );
  NAND2_X1 U11731 ( .A1(n19540), .A2(n20091), .ZN(n19836) );
  NAND2_X1 U11732 ( .A1(n20074), .A2(n20101), .ZN(n19859) );
  NAND2_X1 U11733 ( .A1(n20074), .A2(n14097), .ZN(n19837) );
  NAND2_X1 U11734 ( .A1(n19540), .A2(n20094), .ZN(n19931) );
  OR2_X1 U11735 ( .A1(n16745), .A2(n16746), .ZN(n16743) );
  AOI21_X1 U11736 ( .B1(n17018), .B2(n16785), .A(n17751), .ZN(n9942) );
  OR2_X1 U11737 ( .A1(n16784), .A2(n16785), .ZN(n9943) );
  OR2_X1 U11738 ( .A1(n16796), .A2(n17769), .ZN(n16794) );
  OR2_X1 U11739 ( .A1(n17018), .A2(n16821), .ZN(n9931) );
  OR2_X1 U11740 ( .A1(n16831), .A2(n9932), .ZN(n9930) );
  NAND2_X1 U11741 ( .A1(n17807), .A2(n17813), .ZN(n9932) );
  OR2_X1 U11742 ( .A1(n16831), .A2(n16832), .ZN(n9933) );
  NOR2_X1 U11743 ( .A1(n9983), .A2(n9982), .ZN(n9981) );
  OAI22_X1 U11744 ( .A1(n17380), .A2(n13090), .B1(n17367), .B2(n17127), .ZN(
        n9982) );
  INV_X1 U11745 ( .A(n13091), .ZN(n9983) );
  NAND2_X1 U11746 ( .A1(n12898), .A2(n19014), .ZN(n17249) );
  NOR3_X1 U11747 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(n17045), .ZN(n12898) );
  NAND2_X1 U11748 ( .A1(n17384), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12920) );
  AOI21_X1 U11749 ( .B1(n13080), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n12939), .ZN(n12940) );
  NAND2_X1 U11750 ( .A1(n12956), .A2(n12955), .ZN(n12960) );
  AOI21_X1 U11751 ( .B1(n17392), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n12954), .ZN(n12955) );
  INV_X1 U11752 ( .A(n18858), .ZN(n15943) );
  NOR3_X1 U11753 ( .A1(n15939), .A2(n18411), .A3(n9969), .ZN(n15940) );
  AND2_X1 U11754 ( .A1(n17713), .A2(n9948), .ZN(n16591) );
  AND2_X1 U11755 ( .A1(n9699), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9948) );
  AND3_X1 U11756 ( .A1(n9747), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17923) );
  AND2_X1 U11757 ( .A1(n9944), .A2(n9945), .ZN(n17985) );
  NAND2_X1 U11758 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18040) );
  NAND2_X1 U11759 ( .A1(n13227), .A2(n10065), .ZN(n15916) );
  NOR2_X1 U11760 ( .A1(n13036), .A2(n10064), .ZN(n15862) );
  NAND2_X1 U11761 ( .A1(n10221), .A2(n17727), .ZN(n10064) );
  AND2_X1 U11762 ( .A1(n13029), .A2(n10067), .ZN(n10066) );
  NAND2_X1 U11763 ( .A1(n17781), .A2(n17818), .ZN(n17820) );
  NOR2_X1 U11764 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n13027), .ZN(
        n17821) );
  NOR2_X1 U11765 ( .A1(n10059), .A2(n9782), .ZN(n10082) );
  NAND2_X1 U11766 ( .A1(n13140), .A2(n13149), .ZN(n14408) );
  AND2_X1 U11767 ( .A1(n13150), .A2(n9969), .ZN(n9968) );
  XNOR2_X1 U11768 ( .A(n13002), .B(n13001), .ZN(n18063) );
  INV_X1 U11769 ( .A(n18880), .ZN(n18844) );
  XNOR2_X1 U11770 ( .A(n19020), .B(n17585), .ZN(n18072) );
  OAI21_X1 U11771 ( .B1(n13206), .B2(n13205), .A(n13204), .ZN(n16690) );
  AND2_X1 U11772 ( .A1(n13049), .A2(n10228), .ZN(n13199) );
  NOR2_X1 U11773 ( .A1(n19068), .A2(n14406), .ZN(n18880) );
  INV_X1 U11774 ( .A(n18881), .ZN(n18882) );
  AOI22_X1 U11775 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17320), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13069) );
  AOI211_X1 U11776 ( .C1(n17374), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n13067), .B(n13066), .ZN(n13068) );
  AND2_X1 U11777 ( .A1(n20144), .A2(n13949), .ZN(n20171) );
  INV_X1 U11778 ( .A(n20190), .ZN(n20173) );
  AND2_X1 U11779 ( .A1(n14711), .A2(n13820), .ZN(n14707) );
  INV_X1 U11780 ( .A(n14711), .ZN(n16057) );
  AND2_X1 U11781 ( .A1(n13878), .A2(n16289), .ZN(n20313) );
  XNOR2_X1 U11782 ( .A(n11770), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14842) );
  INV_X1 U11783 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20751) );
  NOR2_X1 U11784 ( .A1(n9692), .A2(n10049), .ZN(n10048) );
  INV_X1 U11785 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20638) );
  OAI211_X1 U11786 ( .C1(n20809), .C2(n20788), .A(n20787), .B(n20786), .ZN(
        n20812) );
  XNOR2_X1 U11787 ( .A(n12381), .B(n10177), .ZN(n16302) );
  INV_X1 U11788 ( .A(n11299), .ZN(n10177) );
  NAND2_X1 U11789 ( .A1(n14931), .A2(n14930), .ZN(n14932) );
  AOI21_X1 U11790 ( .B1(n14929), .B2(n19226), .A(n14928), .ZN(n14930) );
  NAND2_X1 U11791 ( .A1(n15407), .A2(n19209), .ZN(n14931) );
  AOI21_X1 U11792 ( .B1(n16315), .B2(n19189), .A(n16314), .ZN(n10113) );
  NOR2_X1 U11793 ( .A1(n16311), .A2(n10105), .ZN(n10117) );
  INV_X1 U11794 ( .A(n16310), .ZN(n10115) );
  NAND2_X1 U11795 ( .A1(n10116), .A2(n16310), .ZN(n14922) );
  INV_X1 U11796 ( .A(n10117), .ZN(n10116) );
  OR2_X1 U11797 ( .A1(n19390), .A2(n14092), .ZN(n19231) );
  OR2_X1 U11798 ( .A1(n13426), .A2(n16312), .ZN(n19151) );
  NAND2_X1 U11799 ( .A1(n13426), .A2(n19227), .ZN(n15103) );
  NAND2_X1 U11800 ( .A1(n9881), .A2(n9880), .ZN(n9878) );
  NAND2_X1 U11801 ( .A1(n15319), .A2(n9885), .ZN(n9880) );
  NAND2_X1 U11802 ( .A1(n9884), .A2(n9882), .ZN(n9881) );
  NAND2_X1 U11803 ( .A1(n9885), .A2(n9883), .ZN(n9882) );
  INV_X1 U11804 ( .A(n19405), .ZN(n16473) );
  NAND2_X1 U11805 ( .A1(n19394), .A2(n13498), .ZN(n19405) );
  NAND2_X1 U11806 ( .A1(n19936), .A2(n12354), .ZN(n16414) );
  INV_X1 U11807 ( .A(n16465), .ZN(n19397) );
  AND2_X1 U11808 ( .A1(n15410), .A2(n15409), .ZN(n15411) );
  NAND2_X1 U11809 ( .A1(n15407), .A2(n16502), .ZN(n15412) );
  OR2_X1 U11810 ( .A1(n15408), .A2(n15710), .ZN(n15410) );
  XNOR2_X1 U11811 ( .A(n9843), .B(n11342), .ZN(n15416) );
  INV_X1 U11812 ( .A(n10037), .ZN(n10036) );
  OAI211_X1 U11813 ( .C1(n15197), .C2(n16522), .A(n10039), .B(n10038), .ZN(
        n10037) );
  NOR2_X1 U11814 ( .A1(n12368), .A2(n10040), .ZN(n10039) );
  NAND2_X1 U11815 ( .A1(n14936), .A2(n16525), .ZN(n10038) );
  NAND2_X1 U11816 ( .A1(n9875), .A2(n9753), .ZN(n9874) );
  INV_X1 U11817 ( .A(n15344), .ZN(n9875) );
  NAND2_X1 U11818 ( .A1(n15344), .A2(n9750), .ZN(n9879) );
  AND2_X1 U11819 ( .A1(n9878), .A2(n16530), .ZN(n9877) );
  INV_X1 U11820 ( .A(n19540), .ZN(n20084) );
  NOR2_X1 U11821 ( .A1(n18909), .A2(n19056), .ZN(n19054) );
  AND2_X1 U11822 ( .A1(n16731), .A2(n9938), .ZN(n9937) );
  OR2_X1 U11823 ( .A1(n16733), .A2(n16732), .ZN(n9938) );
  INV_X1 U11824 ( .A(n16730), .ZN(n9936) );
  AND2_X1 U11825 ( .A1(n16743), .A2(n17018), .ZN(n16734) );
  NAND2_X1 U11826 ( .A1(n18449), .A2(n17593), .ZN(n17577) );
  OR3_X1 U11827 ( .A1(n12997), .A2(n12999), .A3(n12998), .ZN(n9805) );
  NAND2_X1 U11828 ( .A1(n16559), .A2(n18074), .ZN(n17984) );
  NAND2_X1 U11829 ( .A1(n13224), .A2(n13223), .ZN(n13226) );
  OR2_X1 U11830 ( .A1(n13230), .A2(n13229), .ZN(n13233) );
  INV_X1 U11831 ( .A(n18302), .ZN(n18315) );
  AOI22_X1 U11832 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10502), .B1(
        n19666), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10467) );
  INV_X1 U11833 ( .A(n11683), .ZN(n9952) );
  NAND2_X1 U11834 ( .A1(n12856), .A2(n11588), .ZN(n11530) );
  AND2_X2 U11835 ( .A1(n10010), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11355) );
  NAND2_X1 U11836 ( .A1(n10474), .A2(n9717), .ZN(n10654) );
  NAND2_X1 U11837 ( .A1(n10516), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n9845) );
  NOR2_X1 U11838 ( .A1(n10509), .A2(n9849), .ZN(n9848) );
  AOI21_X1 U11839 ( .B1(n10648), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A(n9666), .ZN(n10504) );
  NOR2_X1 U11840 ( .A1(n19863), .A2(n10471), .ZN(n10477) );
  AND4_X1 U11841 ( .A1(n10454), .A2(n10453), .A3(n10452), .A4(n10451), .ZN(
        n10480) );
  NAND2_X1 U11842 ( .A1(n9712), .A2(n11683), .ZN(n11684) );
  NAND2_X1 U11843 ( .A1(n11581), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9836) );
  OR2_X1 U11844 ( .A1(n12856), .A2(n12845), .ZN(n11496) );
  OR2_X1 U11845 ( .A1(n11659), .A2(n11658), .ZN(n11702) );
  AOI22_X1 U11846 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n11612), .ZN(n11418) );
  AOI21_X1 U11847 ( .B1(n11785), .B2(n11784), .A(n11779), .ZN(n11783) );
  OR3_X1 U11848 ( .A1(n11806), .A2(n11805), .A3(n12718), .ZN(n11807) );
  NAND2_X1 U11849 ( .A1(n11649), .A2(n11648), .ZN(n11792) );
  NOR2_X1 U11850 ( .A1(n10361), .A2(n10917), .ZN(n9914) );
  NOR2_X1 U11851 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(P2_EBX_REG_24__SCAN_IN), 
        .ZN(n10002) );
  NOR2_X1 U11852 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10491) );
  INV_X1 U11853 ( .A(n9872), .ZN(n9871) );
  OAI21_X1 U11854 ( .B1(n9925), .B2(n9924), .A(n15619), .ZN(n9872) );
  INV_X1 U11855 ( .A(n10937), .ZN(n10209) );
  AND2_X1 U11856 ( .A1(n10361), .A2(n13279), .ZN(n10362) );
  AND2_X1 U11857 ( .A1(n10358), .A2(n10384), .ZN(n11310) );
  INV_X1 U11858 ( .A(n9860), .ZN(n9858) );
  INV_X1 U11859 ( .A(n10455), .ZN(n10442) );
  AOI22_X1 U11860 ( .A1(n10284), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10273) );
  NAND2_X1 U11861 ( .A1(n10484), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10278) );
  AOI22_X1 U11862 ( .A1(n10284), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10282) );
  AOI22_X1 U11863 ( .A1(n9649), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10285) );
  NAND2_X1 U11864 ( .A1(n10582), .A2(n10581), .ZN(n10585) );
  NOR2_X1 U11865 ( .A1(n17527), .A2(n18411), .ZN(n13139) );
  NAND2_X1 U11866 ( .A1(n13307), .A2(n12246), .ZN(n10168) );
  INV_X1 U11867 ( .A(n11753), .ZN(n9822) );
  NOR2_X1 U11868 ( .A1(n10164), .A2(n14566), .ZN(n10163) );
  INV_X1 U11869 ( .A(n14638), .ZN(n10164) );
  AND2_X1 U11870 ( .A1(n11986), .A2(n10157), .ZN(n10156) );
  OR2_X1 U11871 ( .A1(n14362), .A2(n14380), .ZN(n10157) );
  AND2_X1 U11872 ( .A1(n14383), .A2(n14382), .ZN(n11986) );
  NOR2_X2 U11873 ( .A1(n14264), .A2(n11939), .ZN(n14319) );
  INV_X1 U11874 ( .A(n14556), .ZN(n9978) );
  AND2_X1 U11875 ( .A1(n9764), .A2(n12797), .ZN(n9974) );
  INV_X1 U11876 ( .A(n12832), .ZN(n12835) );
  AND2_X1 U11877 ( .A1(n14402), .A2(n14384), .ZN(n12797) );
  AND2_X1 U11878 ( .A1(n11494), .A2(n13943), .ZN(n11773) );
  MUX2_X1 U11879 ( .A(n12840), .B(n9674), .S(P1_EBX_REG_1__SCAN_IN), .Z(n12745) );
  OR2_X1 U11880 ( .A1(n11561), .A2(n11560), .ZN(n11589) );
  NAND2_X1 U11881 ( .A1(n11598), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9811) );
  AND3_X1 U11882 ( .A1(n11628), .A2(n11627), .A3(n11626), .ZN(n11630) );
  NAND2_X1 U11883 ( .A1(n20316), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11648) );
  OR2_X1 U11884 ( .A1(n11618), .A2(n11617), .ZN(n11619) );
  AND3_X1 U11885 ( .A1(n12845), .A2(n13918), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11813) );
  NAND2_X1 U11886 ( .A1(n11538), .A2(n11605), .ZN(n10148) );
  OAI21_X1 U11887 ( .B1(n11597), .B2(n9828), .A(n9827), .ZN(n9826) );
  AOI21_X1 U11888 ( .B1(n20970), .B2(n16295), .A(n13861), .ZN(n20315) );
  NAND2_X1 U11889 ( .A1(n11813), .A2(n11773), .ZN(n11810) );
  INV_X1 U11890 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13845) );
  NAND2_X1 U11891 ( .A1(n10799), .A2(n9999), .ZN(n10814) );
  NOR2_X1 U11892 ( .A1(n10001), .A2(n10000), .ZN(n9999) );
  NAND2_X1 U11893 ( .A1(n10003), .A2(n10002), .ZN(n10001) );
  INV_X1 U11894 ( .A(n10798), .ZN(n10000) );
  AND2_X1 U11895 ( .A1(n10092), .A2(n13426), .ZN(n10090) );
  AND2_X1 U11896 ( .A1(n19422), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10721) );
  NAND2_X1 U11897 ( .A1(n10604), .A2(n10603), .ZN(n10602) );
  NOR2_X1 U11898 ( .A1(n10142), .A2(n16342), .ZN(n10141) );
  INV_X1 U11899 ( .A(n10144), .ZN(n10142) );
  NOR2_X1 U11900 ( .A1(n10712), .A2(n10711), .ZN(n11009) );
  NAND2_X1 U11901 ( .A1(n10310), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9857) );
  NOR2_X1 U11902 ( .A1(n13436), .A2(n10123), .ZN(n10122) );
  INV_X1 U11903 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10123) );
  NOR2_X1 U11904 ( .A1(n16409), .A2(n10120), .ZN(n10119) );
  NOR2_X1 U11905 ( .A1(n15446), .A2(n15456), .ZN(n10200) );
  AND2_X1 U11906 ( .A1(n14947), .A2(n11014), .ZN(n10834) );
  NOR2_X1 U11907 ( .A1(n15471), .A2(n10198), .ZN(n10197) );
  INV_X1 U11908 ( .A(n10806), .ZN(n10198) );
  OR2_X1 U11909 ( .A1(n15867), .A2(n10961), .ZN(n10802) );
  NOR2_X1 U11910 ( .A1(n10966), .A2(n10203), .ZN(n10202) );
  INV_X1 U11911 ( .A(n10232), .ZN(n10203) );
  INV_X1 U11912 ( .A(n15188), .ZN(n10170) );
  INV_X1 U11913 ( .A(n16493), .ZN(n9841) );
  AND2_X1 U11914 ( .A1(n10025), .A2(n15612), .ZN(n10024) );
  INV_X1 U11915 ( .A(n11175), .ZN(n11170) );
  NOR2_X1 U11916 ( .A1(n15674), .A2(n15691), .ZN(n10208) );
  NAND2_X1 U11917 ( .A1(n10184), .A2(n13780), .ZN(n10183) );
  INV_X1 U11918 ( .A(n13773), .ZN(n10184) );
  OAI222_X1 U11919 ( .A1(n11034), .A2(n13550), .B1(n9736), .B2(n19354), .C1(
        n11175), .C2(n20013), .ZN(n10990) );
  NOR2_X1 U11920 ( .A1(n10540), .A2(n10539), .ZN(n10989) );
  NAND2_X1 U11921 ( .A1(n10975), .A2(n10974), .ZN(n10988) );
  INV_X1 U11922 ( .A(n10988), .ZN(n11147) );
  NAND2_X1 U11923 ( .A1(n12403), .A2(n13484), .ZN(n12424) );
  NOR2_X1 U11924 ( .A1(n12594), .A2(n12410), .ZN(n12411) );
  AND2_X2 U11925 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13747) );
  NAND2_X1 U11926 ( .A1(n10462), .A2(n13653), .ZN(n10472) );
  AND2_X1 U11927 ( .A1(n12408), .A2(n10460), .ZN(n10461) );
  NAND2_X1 U11928 ( .A1(n10464), .A2(n13653), .ZN(n10470) );
  NAND2_X1 U11929 ( .A1(n10457), .A2(n13653), .ZN(n19924) );
  NAND2_X1 U11930 ( .A1(n10866), .A2(n10865), .ZN(n10912) );
  NAND2_X1 U11931 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19014), .ZN(
        n12900) );
  NAND2_X1 U11932 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n17045), .ZN(
        n12901) );
  INV_X1 U11933 ( .A(n13134), .ZN(n13135) );
  INV_X1 U11934 ( .A(n17831), .ZN(n16723) );
  NOR2_X1 U11935 ( .A1(n18040), .A2(n18042), .ZN(n9944) );
  NOR2_X1 U11936 ( .A1(n18019), .A2(n9946), .ZN(n9945) );
  OAI22_X1 U11937 ( .A1(n10065), .A2(n17819), .B1(n19019), .B2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10062) );
  NOR2_X1 U11938 ( .A1(n10211), .A2(n16586), .ZN(n10065) );
  AND3_X1 U11939 ( .A1(n17820), .A2(n10068), .A3(n9704), .ZN(n13032) );
  NOR2_X1 U11940 ( .A1(n18027), .A2(n13172), .ZN(n13174) );
  OAI21_X1 U11941 ( .B1(n18048), .B2(n10057), .A(n10056), .ZN(n13014) );
  NAND2_X1 U11942 ( .A1(n10058), .A2(n9713), .ZN(n10057) );
  OR2_X1 U11943 ( .A1(n18051), .A2(n13165), .ZN(n9803) );
  INV_X1 U11944 ( .A(n15852), .ZN(n18870) );
  NOR2_X1 U11945 ( .A1(n19032), .A2(n18914), .ZN(n18410) );
  OR2_X1 U11946 ( .A1(n20973), .A2(n13939), .ZN(n20144) );
  NAND2_X1 U11947 ( .A1(n20144), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13960) );
  AND2_X1 U11948 ( .A1(n13917), .A2(n13916), .ZN(n20201) );
  OR2_X1 U11949 ( .A1(n14731), .A2(n12315), .ZN(n12244) );
  AND2_X1 U11950 ( .A1(n12203), .A2(n12202), .ZN(n14585) );
  OR2_X1 U11951 ( .A1(n15946), .A2(n12315), .ZN(n12202) );
  NOR2_X1 U11952 ( .A1(n12157), .A2(n15974), .ZN(n12158) );
  OR2_X1 U11953 ( .A1(n16067), .A2(n12315), .ZN(n12160) );
  AND2_X1 U11954 ( .A1(n12115), .A2(n12114), .ZN(n14607) );
  AND2_X1 U11955 ( .A1(n12096), .A2(n12095), .ZN(n14619) );
  NOR2_X1 U11956 ( .A1(n12077), .A2(n16011), .ZN(n12078) );
  NAND2_X1 U11957 ( .A1(n10160), .A2(n10159), .ZN(n10158) );
  INV_X1 U11958 ( .A(n14620), .ZN(n10159) );
  NAND2_X1 U11959 ( .A1(n12047), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12077) );
  NAND2_X1 U11960 ( .A1(n14778), .A2(n14777), .ZN(n14768) );
  AND2_X1 U11961 ( .A1(n12034), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12047) );
  AND2_X1 U11962 ( .A1(n12002), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12020) );
  NOR2_X1 U11963 ( .A1(n11987), .A2(n14809), .ZN(n12002) );
  NAND2_X1 U11964 ( .A1(n11970), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11987) );
  NAND2_X1 U11965 ( .A1(n14319), .A2(n10156), .ZN(n14373) );
  INV_X1 U11966 ( .A(n11955), .ZN(n11970) );
  AND2_X1 U11967 ( .A1(n11940), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11941) );
  NAND2_X1 U11968 ( .A1(n11941), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11955) );
  CLKBUF_X1 U11969 ( .A(n14319), .Z(n14320) );
  NAND2_X1 U11970 ( .A1(n11907), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11935) );
  AND3_X1 U11971 ( .A1(n11906), .A2(n11905), .A3(n11904), .ZN(n14120) );
  AND2_X1 U11972 ( .A1(n11886), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11907) );
  CLKBUF_X1 U11973 ( .A(n14003), .Z(n14004) );
  AOI21_X1 U11974 ( .B1(n11884), .B2(n11967), .A(n11883), .ZN(n13996) );
  CLKBUF_X1 U11975 ( .A(n13994), .Z(n13995) );
  INV_X1 U11976 ( .A(n11869), .ZN(n11870) );
  INV_X1 U11977 ( .A(n13931), .ZN(n11876) );
  INV_X1 U11978 ( .A(n13932), .ZN(n11877) );
  NAND2_X1 U11979 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11851) );
  NOR2_X1 U11980 ( .A1(n11851), .A2(n11850), .ZN(n11861) );
  INV_X1 U11981 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11850) );
  OAI21_X1 U11982 ( .B1(n11830), .B2(n12016), .A(n11829), .ZN(n11831) );
  NOR2_X1 U11983 ( .A1(n11828), .A2(n10250), .ZN(n11829) );
  NOR2_X1 U11984 ( .A1(n11768), .A2(n10042), .ZN(n10041) );
  NAND2_X1 U11985 ( .A1(n12711), .A2(n10229), .ZN(n10022) );
  OAI21_X1 U11986 ( .B1(n14764), .B2(n9813), .A(n9812), .ZN(n9962) );
  NOR2_X1 U11987 ( .A1(n14598), .A2(n14587), .ZN(n14589) );
  AND2_X1 U11988 ( .A1(n14881), .A2(n12880), .ZN(n14869) );
  NAND2_X1 U11989 ( .A1(n14611), .A2(n9976), .ZN(n14598) );
  AND2_X1 U11990 ( .A1(n9777), .A2(n9977), .ZN(n9976) );
  INV_X1 U11991 ( .A(n14595), .ZN(n9977) );
  NAND2_X1 U11992 ( .A1(n14611), .A2(n9777), .ZN(n14596) );
  NAND2_X1 U11993 ( .A1(n14611), .A2(n14601), .ZN(n14603) );
  AND2_X1 U11994 ( .A1(n14615), .A2(n14609), .ZN(n14611) );
  NOR2_X1 U11995 ( .A1(n14624), .A2(n14614), .ZN(n14615) );
  OR2_X1 U11996 ( .A1(n14628), .A2(n14622), .ZN(n14624) );
  NOR2_X1 U11997 ( .A1(n9975), .A2(n12806), .ZN(n14637) );
  NAND2_X1 U11998 ( .A1(n14637), .A2(n14626), .ZN(n14628) );
  OR2_X1 U11999 ( .A1(n11759), .A2(n16082), .ZN(n10018) );
  AND3_X1 U12000 ( .A1(n12804), .A2(n12820), .A3(n12803), .ZN(n14573) );
  INV_X1 U12001 ( .A(n11759), .ZN(n14782) );
  NAND2_X1 U12002 ( .A1(n14404), .A2(n12797), .ZN(n14646) );
  NAND2_X1 U12003 ( .A1(n11757), .A2(n10014), .ZN(n14800) );
  NAND2_X1 U12004 ( .A1(n16110), .A2(n16213), .ZN(n10014) );
  OR2_X1 U12005 ( .A1(n14268), .A2(n14269), .ZN(n14321) );
  INV_X1 U12006 ( .A(n11750), .ZN(n14333) );
  NAND2_X1 U12007 ( .A1(n9965), .A2(n9691), .ZN(n14123) );
  AND2_X1 U12008 ( .A1(n12779), .A2(n12778), .ZN(n14124) );
  OR2_X1 U12009 ( .A1(n14123), .A2(n14124), .ZN(n14268) );
  NOR2_X1 U12010 ( .A1(n13927), .A2(n9964), .ZN(n14096) );
  NAND2_X1 U12011 ( .A1(n9966), .A2(n13997), .ZN(n9964) );
  NAND2_X1 U12012 ( .A1(n9820), .A2(n11644), .ZN(n9819) );
  NAND2_X1 U12013 ( .A1(n13791), .A2(n9690), .ZN(n9817) );
  NAND2_X1 U12014 ( .A1(n13895), .A2(n13894), .ZN(n13893) );
  NAND2_X1 U12015 ( .A1(n9965), .A2(n9967), .ZN(n13964) );
  XNOR2_X1 U12016 ( .A(n11592), .B(n13664), .ZN(n20246) );
  NAND2_X1 U12017 ( .A1(n11584), .A2(n11581), .ZN(n10052) );
  NOR2_X1 U12018 ( .A1(n11584), .A2(n11581), .ZN(n10053) );
  NAND2_X1 U12019 ( .A1(n10149), .A2(n11607), .ZN(n9958) );
  NAND2_X1 U12020 ( .A1(n9712), .A2(n11663), .ZN(n20305) );
  CLKBUF_X1 U12021 ( .A(n13681), .Z(n13859) );
  NOR2_X1 U12022 ( .A1(n14472), .A2(n20326), .ZN(n15880) );
  CLKBUF_X1 U12023 ( .A(n13325), .Z(n13326) );
  INV_X1 U12024 ( .A(n20548), .ZN(n20674) );
  NOR2_X1 U12025 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20315), .ZN(n20377) );
  OR2_X1 U12026 ( .A1(n20675), .A2(n20674), .ZN(n20703) );
  AND2_X1 U12027 ( .A1(n9675), .A2(n20306), .ZN(n20548) );
  NAND2_X1 U12028 ( .A1(n20313), .A2(n20311), .ZN(n20370) );
  AND2_X1 U12029 ( .A1(n12736), .A2(n14477), .ZN(n15898) );
  INV_X1 U12030 ( .A(n11281), .ZN(n11296) );
  AOI21_X1 U12031 ( .B1(n10086), .B2(n10084), .A(n10083), .ZN(n16324) );
  NOR2_X1 U12032 ( .A1(n10089), .A2(n10085), .ZN(n10084) );
  OAI21_X1 U12033 ( .B1(n10087), .B2(n10085), .A(n15281), .ZN(n10083) );
  AOI21_X1 U12034 ( .B1(n10090), .B2(n10088), .A(n15290), .ZN(n10087) );
  INV_X1 U12035 ( .A(n10094), .ZN(n10088) );
  INV_X1 U12036 ( .A(n10090), .ZN(n10089) );
  NOR2_X1 U12037 ( .A1(n19132), .A2(n10085), .ZN(n10098) );
  INV_X1 U12039 ( .A(n10756), .ZN(n9996) );
  AND2_X1 U12040 ( .A1(n13385), .A2(n10118), .ZN(n13420) );
  AND2_X1 U12041 ( .A1(n9700), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10118) );
  NAND2_X1 U12042 ( .A1(n10004), .A2(n10675), .ZN(n10732) );
  AND2_X1 U12043 ( .A1(n10006), .A2(n10005), .ZN(n10004) );
  INV_X1 U12044 ( .A(n10721), .ZN(n10005) );
  AND2_X1 U12045 ( .A1(n10675), .A2(n10007), .ZN(n10725) );
  OR2_X1 U12046 ( .A1(n11064), .A2(n11063), .ZN(n13882) );
  NAND2_X1 U12047 ( .A1(n10185), .A2(n10426), .ZN(n9866) );
  AND2_X1 U12048 ( .A1(n11192), .A2(n11191), .ZN(n14218) );
  NAND2_X1 U12049 ( .A1(n10135), .A2(n10133), .ZN(n12699) );
  INV_X1 U12050 ( .A(n15141), .ZN(n10134) );
  INV_X1 U12051 ( .A(n14949), .ZN(n10033) );
  NAND2_X1 U12052 ( .A1(n15504), .A2(n9774), .ZN(n14966) );
  NAND2_X1 U12053 ( .A1(n10132), .A2(n10131), .ZN(n10130) );
  NAND2_X1 U12054 ( .A1(n16338), .A2(n9779), .ZN(n10129) );
  INV_X1 U12055 ( .A(n15229), .ZN(n10131) );
  NOR2_X1 U12056 ( .A1(n15227), .A2(n15229), .ZN(n15228) );
  OR4_X1 U12057 ( .A1(n12519), .A2(n12518), .A3(n12517), .A4(n12516), .ZN(
        n15173) );
  CLKBUF_X1 U12058 ( .A(n15171), .Z(n15172) );
  OR4_X1 U12059 ( .A1(n12489), .A2(n12488), .A3(n12487), .A4(n12486), .ZN(
        n15180) );
  OR4_X1 U12060 ( .A1(n12459), .A2(n12458), .A3(n12457), .A4(n12456), .ZN(
        n14350) );
  CLKBUF_X1 U12061 ( .A(n14348), .Z(n14349) );
  CLKBUF_X1 U12062 ( .A(n14346), .Z(n14347) );
  AND2_X1 U12063 ( .A1(n10028), .A2(n15065), .ZN(n10027) );
  INV_X1 U12064 ( .A(n15109), .ZN(n10032) );
  AND2_X1 U12065 ( .A1(n13542), .A2(n19996), .ZN(n19331) );
  NAND2_X1 U12066 ( .A1(n10111), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10108) );
  NOR2_X1 U12067 ( .A1(n13442), .A2(n12356), .ZN(n14920) );
  AND2_X1 U12068 ( .A1(n14981), .A2(n9788), .ZN(n13447) );
  INV_X1 U12069 ( .A(n13448), .ZN(n10186) );
  NAND2_X1 U12070 ( .A1(n14981), .A2(n9775), .ZN(n15153) );
  NAND2_X1 U12071 ( .A1(n13433), .A2(n9703), .ZN(n13440) );
  NAND2_X1 U12072 ( .A1(n13433), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13437) );
  NAND2_X1 U12073 ( .A1(n13430), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13434) );
  OR2_X1 U12074 ( .A1(n15181), .A2(n15334), .ZN(n15336) );
  NAND2_X1 U12075 ( .A1(n13424), .A2(n9701), .ZN(n13431) );
  AND2_X1 U12076 ( .A1(n13424), .A2(n9778), .ZN(n13429) );
  AND2_X1 U12077 ( .A1(n13424), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13427) );
  AND2_X1 U12078 ( .A1(n13411), .A2(n9744), .ZN(n15183) );
  NAND2_X1 U12079 ( .A1(n13420), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13421) );
  NOR2_X1 U12080 ( .A1(n13421), .A2(n19141), .ZN(n13424) );
  NOR2_X1 U12081 ( .A1(n9740), .A2(n10173), .ZN(n10172) );
  INV_X1 U12082 ( .A(n15026), .ZN(n10173) );
  AND2_X1 U12083 ( .A1(n11238), .A2(n11237), .ZN(n13412) );
  NAND2_X1 U12084 ( .A1(n13385), .A2(n9700), .ZN(n13386) );
  AND2_X1 U12085 ( .A1(n11229), .A2(n11228), .ZN(n13906) );
  NOR2_X1 U12086 ( .A1(n15049), .A2(n9740), .ZN(n15025) );
  NAND2_X1 U12087 ( .A1(n13385), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13384) );
  AND2_X1 U12088 ( .A1(n11221), .A2(n11220), .ZN(n13883) );
  NOR2_X1 U12089 ( .A1(n15049), .A2(n13883), .ZN(n15632) );
  NOR2_X1 U12090 ( .A1(n10127), .A2(n10126), .ZN(n10125) );
  INV_X1 U12091 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10126) );
  NOR2_X1 U12092 ( .A1(n13380), .A2(n10127), .ZN(n13383) );
  INV_X1 U12093 ( .A(n10180), .ZN(n10179) );
  NOR2_X1 U12094 ( .A1(n13378), .A2(n16470), .ZN(n13381) );
  NAND2_X1 U12095 ( .A1(n13381), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13380) );
  NOR2_X1 U12096 ( .A1(n13772), .A2(n13773), .ZN(n13781) );
  NOR2_X1 U12097 ( .A1(n13377), .A2(n16484), .ZN(n13379) );
  NAND2_X1 U12098 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13377) );
  NAND2_X1 U12099 ( .A1(n10409), .A2(n10408), .ZN(n10432) );
  NAND2_X1 U12100 ( .A1(n11300), .A2(n9758), .ZN(n10404) );
  NAND2_X1 U12101 ( .A1(n10431), .A2(n10432), .ZN(n10439) );
  NOR2_X1 U12102 ( .A1(n10529), .A2(n10528), .ZN(n13496) );
  NAND2_X1 U12103 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10207) );
  NAND2_X1 U12104 ( .A1(n9650), .A2(n9912), .ZN(n9911) );
  INV_X1 U12105 ( .A(n12376), .ZN(n9912) );
  NAND2_X1 U12106 ( .A1(n9908), .A2(n9905), .ZN(n9903) );
  OR2_X1 U12107 ( .A1(n9650), .A2(n9731), .ZN(n9907) );
  NAND2_X1 U12108 ( .A1(n9650), .A2(n10236), .ZN(n9906) );
  INV_X1 U12109 ( .A(n12365), .ZN(n10040) );
  OR2_X1 U12110 ( .A1(n13445), .A2(n10961), .ZN(n12330) );
  NAND2_X1 U12111 ( .A1(n10817), .A2(n10836), .ZN(n15277) );
  NOR2_X1 U12112 ( .A1(n10834), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15285) );
  NAND2_X1 U12113 ( .A1(n10196), .A2(n15469), .ZN(n15286) );
  AND2_X1 U12114 ( .A1(n15502), .A2(n14979), .ZN(n14981) );
  AND2_X1 U12115 ( .A1(n10201), .A2(n9796), .ZN(n9840) );
  AND2_X1 U12116 ( .A1(n10202), .A2(n11335), .ZN(n10201) );
  AOI21_X1 U12117 ( .B1(n9923), .B2(n9921), .A(n9725), .ZN(n9920) );
  INV_X1 U12118 ( .A(n9923), .ZN(n9922) );
  INV_X1 U12119 ( .A(n9925), .ZN(n9921) );
  OR2_X1 U12120 ( .A1(n15336), .A2(n15174), .ZN(n15501) );
  NOR2_X1 U12121 ( .A1(n15501), .A2(n15500), .ZN(n15502) );
  AOI21_X1 U12122 ( .B1(n15327), .B2(n15314), .A(n9886), .ZN(n9885) );
  INV_X1 U12123 ( .A(n15328), .ZN(n9886) );
  INV_X1 U12124 ( .A(n15319), .ZN(n9884) );
  NOR2_X1 U12125 ( .A1(n15315), .A2(n9888), .ZN(n9887) );
  INV_X1 U12126 ( .A(n15342), .ZN(n9888) );
  OAI21_X1 U12127 ( .B1(n15382), .B2(n9891), .A(n9889), .ZN(n9901) );
  AOI21_X1 U12128 ( .B1(n9890), .B2(n9896), .A(n15312), .ZN(n9889) );
  NOR2_X1 U12129 ( .A1(n10026), .A2(n15631), .ZN(n10025) );
  INV_X1 U12130 ( .A(n15650), .ZN(n10026) );
  AOI21_X1 U12131 ( .B1(n10191), .B2(n10730), .A(n9759), .ZN(n10189) );
  NAND2_X1 U12132 ( .A1(n10195), .A2(n10192), .ZN(n15645) );
  INV_X1 U12133 ( .A(n15683), .ZN(n15608) );
  OR2_X1 U12134 ( .A1(n10962), .A2(n10961), .ZN(n10960) );
  AND2_X1 U12135 ( .A1(n11204), .A2(n11203), .ZN(n13760) );
  OR2_X1 U12136 ( .A1(n13772), .A2(n10183), .ZN(n13779) );
  XNOR2_X1 U12137 ( .A(n10962), .B(n10961), .ZN(n15390) );
  OAI21_X1 U12138 ( .B1(n10949), .B2(n9718), .A(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n9851) );
  XNOR2_X1 U12139 ( .A(n10715), .B(n15695), .ZN(n15402) );
  NAND2_X1 U12140 ( .A1(n9916), .A2(n9754), .ZN(n10636) );
  AND2_X1 U12141 ( .A1(n10943), .A2(n10942), .ZN(n14312) );
  NAND2_X1 U12142 ( .A1(n14312), .A2(n14309), .ZN(n14314) );
  NOR2_X1 U12143 ( .A1(n13805), .A2(n10030), .ZN(n14300) );
  NAND2_X1 U12144 ( .A1(n10031), .A2(n14214), .ZN(n10030) );
  NAND2_X1 U12145 ( .A1(n16480), .A2(n16479), .ZN(n16478) );
  AND2_X1 U12146 ( .A1(n11303), .A2(n11302), .ZN(n14054) );
  OAI211_X1 U12147 ( .C1(n11175), .C2(n19091), .A(n10985), .B(n10984), .ZN(
        n13604) );
  NAND3_X1 U12148 ( .A1(n11311), .A2(n13267), .A3(n13764), .ZN(n10355) );
  NAND2_X1 U12149 ( .A1(n10918), .A2(n10916), .ZN(n13261) );
  NAND2_X1 U12150 ( .A1(n10353), .A2(n10384), .ZN(n13486) );
  NAND2_X1 U12151 ( .A1(n20084), .A2(n20091), .ZN(n19700) );
  INV_X1 U12152 ( .A(n19436), .ZN(n19428) );
  NAND2_X1 U12153 ( .A1(n19936), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19438) );
  INV_X1 U12154 ( .A(n19936), .ZN(n19865) );
  NOR2_X2 U12155 ( .A1(n14107), .A2(n16414), .ZN(n19437) );
  OR3_X1 U12156 ( .A1(n9661), .A2(n16713), .A3(n18870), .ZN(n18840) );
  AND2_X1 U12157 ( .A1(n9940), .A2(n17018), .ZN(n16764) );
  OR2_X1 U12158 ( .A1(n16784), .A2(n9941), .ZN(n9940) );
  INV_X1 U12159 ( .A(n9942), .ZN(n9941) );
  AND2_X1 U12160 ( .A1(n9930), .A2(n9767), .ZN(n16809) );
  INV_X1 U12161 ( .A(n16885), .ZN(n16897) );
  INV_X1 U12162 ( .A(n18411), .ZN(n14411) );
  NOR2_X1 U12163 ( .A1(n17604), .A2(n9972), .ZN(n9971) );
  NOR2_X1 U12164 ( .A1(n19014), .A2(n19025), .ZN(n9984) );
  INV_X1 U12165 ( .A(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15832) );
  NOR2_X1 U12166 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9807) );
  INV_X1 U12167 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15825) );
  NAND2_X1 U12168 ( .A1(n17374), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12995) );
  NOR2_X1 U12169 ( .A1(n17659), .A2(n17594), .ZN(n17624) );
  INV_X1 U12170 ( .A(n17659), .ZN(n17656) );
  NAND2_X1 U12171 ( .A1(n17713), .A2(n9699), .ZN(n16554) );
  NOR2_X1 U12172 ( .A1(n17711), .A2(n9950), .ZN(n9949) );
  INV_X1 U12173 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n9950) );
  NAND2_X1 U12174 ( .A1(n17713), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17719) );
  NOR2_X1 U12175 ( .A1(n17749), .A2(n17748), .ZN(n17713) );
  NOR2_X1 U12176 ( .A1(n18227), .A2(n16568), .ZN(n17726) );
  NAND2_X1 U12177 ( .A1(n9714), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17770) );
  AND2_X1 U12178 ( .A1(n17831), .A2(n9928), .ZN(n17802) );
  NOR2_X1 U12179 ( .A1(n17834), .A2(n17833), .ZN(n9928) );
  INV_X1 U12180 ( .A(n17770), .ZN(n17759) );
  NOR2_X1 U12181 ( .A1(n17875), .A2(n9929), .ZN(n17831) );
  NAND2_X1 U12182 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n9929) );
  INV_X1 U12183 ( .A(n17999), .ZN(n17809) );
  INV_X1 U12184 ( .A(n17918), .ZN(n17879) );
  OR2_X1 U12185 ( .A1(n17877), .A2(n17878), .ZN(n17875) );
  OR2_X1 U12186 ( .A1(n13126), .A2(n13125), .ZN(n13127) );
  NAND2_X1 U12187 ( .A1(n15916), .A2(n10059), .ZN(n13285) );
  NAND2_X1 U12188 ( .A1(n10063), .A2(n10060), .ZN(n13284) );
  NAND2_X1 U12189 ( .A1(n17735), .A2(n10059), .ZN(n10063) );
  AND2_X1 U12190 ( .A1(n15917), .A2(n10061), .ZN(n10060) );
  INV_X1 U12191 ( .A(n10062), .ZN(n10061) );
  OAI21_X1 U12192 ( .B1(n17710), .B2(n13037), .A(n16559), .ZN(n13133) );
  AND2_X1 U12193 ( .A1(n13227), .A2(n13228), .ZN(n13037) );
  NOR2_X1 U12194 ( .A1(n16568), .A2(n18218), .ZN(n18090) );
  NOR2_X1 U12195 ( .A1(n17746), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17745) );
  NOR2_X1 U12196 ( .A1(n13032), .A2(n17819), .ZN(n17765) );
  NOR2_X1 U12197 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n10059), .ZN(
        n17858) );
  OR2_X1 U12198 ( .A1(n17959), .A2(n10079), .ZN(n17891) );
  NAND2_X1 U12199 ( .A1(n9687), .A2(n17933), .ZN(n10079) );
  NOR2_X1 U12200 ( .A1(n17891), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17907) );
  INV_X1 U12201 ( .A(n18309), .ZN(n18233) );
  OR2_X1 U12202 ( .A1(n17992), .A2(n13184), .ZN(n18277) );
  INV_X1 U12203 ( .A(n18277), .ZN(n18244) );
  NOR2_X1 U12204 ( .A1(n13181), .A2(n9806), .ZN(n17993) );
  AND2_X1 U12205 ( .A1(n13182), .A2(n13183), .ZN(n9806) );
  NOR2_X1 U12206 ( .A1(n17993), .A2(n18312), .ZN(n17992) );
  NAND2_X1 U12207 ( .A1(n10078), .A2(n10075), .ZN(n10074) );
  NOR2_X1 U12208 ( .A1(n18012), .A2(n18336), .ZN(n18011) );
  XNOR2_X1 U12209 ( .A(n13170), .B(n13171), .ZN(n18028) );
  NOR2_X1 U12210 ( .A1(n18028), .A2(n18344), .ZN(n18027) );
  XNOR2_X1 U12211 ( .A(n13014), .B(n13013), .ZN(n18026) );
  XNOR2_X1 U12212 ( .A(n9803), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18038) );
  NOR2_X1 U12213 ( .A1(n18038), .A2(n18037), .ZN(n18036) );
  XNOR2_X1 U12214 ( .A(n13164), .B(n18050), .ZN(n18052) );
  NOR2_X1 U12215 ( .A1(n18059), .A2(n13163), .ZN(n18053) );
  NOR2_X1 U12216 ( .A1(n18053), .A2(n18052), .ZN(n18051) );
  INV_X1 U12217 ( .A(n9805), .ZN(n13161) );
  NOR2_X1 U12218 ( .A1(n13130), .A2(n13209), .ZN(n18839) );
  NOR2_X1 U12219 ( .A1(n9805), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18069) );
  NAND2_X1 U12220 ( .A1(n13152), .A2(n9755), .ZN(n18868) );
  NOR2_X2 U12221 ( .A1(n19031), .A2(n19025), .ZN(n18850) );
  NOR2_X1 U12222 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18410), .ZN(n18758) );
  AOI211_X1 U12223 ( .C1(n17374), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n13099), .B(n13098), .ZN(n13100) );
  INV_X1 U12224 ( .A(n13199), .ZN(n18434) );
  AOI211_X1 U12225 ( .C1(n17321), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n13057), .B(n13056), .ZN(n13058) );
  NOR2_X2 U12226 ( .A1(n18755), .A2(n18525), .ZN(n18786) );
  INV_X1 U12227 ( .A(n18758), .ZN(n18525) );
  AOI22_X1 U12228 ( .A1(n18845), .A2(n18252), .B1(n16551), .B2(n16550), .ZN(
        n18848) );
  OAI21_X1 U12229 ( .B1(n15850), .B2(n17594), .A(n15849), .ZN(n18881) );
  OAI21_X1 U12230 ( .B1(n13276), .B2(n13275), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n15220) );
  NAND3_X1 U12231 ( .A1(n13501), .A2(n14483), .A3(n14477), .ZN(n14011) );
  NAND2_X1 U12232 ( .A1(n13504), .A2(n14011), .ZN(n20973) );
  INV_X1 U12233 ( .A(n20175), .ZN(n20146) );
  INV_X1 U12234 ( .A(n20171), .ZN(n20189) );
  INV_X1 U12235 ( .A(n20187), .ZN(n20177) );
  AND2_X1 U12236 ( .A1(n20144), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20186) );
  NAND2_X1 U12237 ( .A1(n13947), .A2(n13946), .ZN(n20190) );
  AND2_X1 U12238 ( .A1(n14510), .A2(n14509), .ZN(n14844) );
  OAI21_X1 U12239 ( .B1(n13627), .B2(n13355), .A(n13354), .ZN(n14642) );
  INV_X1 U12240 ( .A(n14496), .ZN(n14659) );
  INV_X1 U12241 ( .A(n14691), .ZN(n14705) );
  NAND2_X1 U12242 ( .A1(n13333), .A2(n13332), .ZN(n14711) );
  NAND2_X1 U12243 ( .A1(n13631), .A2(n14483), .ZN(n13333) );
  INV_X1 U12244 ( .A(n16059), .ZN(n14713) );
  NOR2_X1 U12245 ( .A1(n20201), .A2(n20231), .ZN(n20218) );
  BUF_X1 U12246 ( .A(n20218), .Z(n20230) );
  BUF_X1 U12247 ( .A(n14243), .Z(n20231) );
  INV_X1 U12248 ( .A(n14187), .ZN(n14012) );
  NOR2_X1 U12249 ( .A1(n12397), .A2(n12396), .ZN(n12398) );
  INV_X1 U12250 ( .A(n12393), .ZN(n12394) );
  AND2_X1 U12251 ( .A1(n12397), .A2(n12288), .ZN(n14719) );
  OR2_X1 U12252 ( .A1(n13306), .A2(n13307), .ZN(n13309) );
  INV_X1 U12253 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n16011) );
  INV_X1 U12254 ( .A(n10147), .ZN(n13890) );
  INV_X1 U12255 ( .A(n16074), .ZN(n20244) );
  NAND2_X1 U12256 ( .A1(n14728), .A2(n14846), .ZN(n10043) );
  AND2_X1 U12257 ( .A1(n12844), .A2(n13360), .ZN(n14440) );
  XNOR2_X1 U12258 ( .A(n10020), .B(n10019), .ZN(n13314) );
  INV_X1 U12259 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10019) );
  NAND2_X1 U12260 ( .A1(n10023), .A2(n10021), .ZN(n10020) );
  NAND2_X1 U12261 ( .A1(n10022), .A2(n16110), .ZN(n10021) );
  AND2_X1 U12262 ( .A1(n16138), .A2(n12886), .ZN(n14858) );
  NAND2_X1 U12263 ( .A1(n20260), .A2(n20294), .ZN(n20279) );
  NOR3_X1 U12264 ( .A1(n16273), .A2(n12883), .A3(n16213), .ZN(n16205) );
  NAND2_X1 U12265 ( .A1(n11752), .A2(n11751), .ZN(n14342) );
  NAND2_X1 U12266 ( .A1(n10045), .A2(n10044), .ZN(n16122) );
  NAND2_X1 U12267 ( .A1(n16132), .A2(n11710), .ZN(n16129) );
  AND2_X1 U12268 ( .A1(n12874), .A2(n12854), .ZN(n20276) );
  AND2_X1 U12269 ( .A1(n12874), .A2(n12740), .ZN(n20296) );
  AND2_X1 U12270 ( .A1(n12874), .A2(n12847), .ZN(n20292) );
  INV_X1 U12271 ( .A(n20296), .ZN(n16225) );
  INV_X1 U12272 ( .A(n20823), .ZN(n20817) );
  NAND2_X1 U12273 ( .A1(n14477), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20950) );
  OR2_X1 U12274 ( .A1(n20448), .A2(n20701), .ZN(n20382) );
  INV_X1 U12275 ( .A(n20447), .ZN(n20465) );
  OAI21_X1 U12276 ( .B1(n20492), .B2(n20476), .A(n20787), .ZN(n20494) );
  NOR2_X1 U12277 ( .A1(n20751), .A2(n20551), .ZN(n20571) );
  OAI211_X1 U12278 ( .C1(n20603), .C2(n11516), .A(n20640), .B(n20587), .ZN(
        n20605) );
  INV_X1 U12279 ( .A(n20644), .ZN(n20662) );
  INV_X1 U12280 ( .A(n20700), .ZN(n20660) );
  INV_X1 U12281 ( .A(n20737), .ZN(n20857) );
  INV_X1 U12282 ( .A(n20741), .ZN(n20863) );
  NOR2_X1 U12283 ( .A1(n20751), .A2(n20825), .ZN(n20873) );
  NAND2_X1 U12284 ( .A1(n20824), .A2(n20779), .ZN(n20880) );
  INV_X1 U12285 ( .A(n20747), .ZN(n20871) );
  NAND2_X1 U12286 ( .A1(n16292), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15913) );
  INV_X1 U12287 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16292) );
  OR2_X1 U12288 ( .A1(n13472), .A2(n13398), .ZN(n13464) );
  OAI21_X1 U12289 ( .B1(n14976), .B2(n10089), .A(n10087), .ZN(n16326) );
  NAND2_X1 U12290 ( .A1(n14976), .A2(n10094), .ZN(n10091) );
  NAND2_X1 U12291 ( .A1(n10099), .A2(n10096), .ZN(n19100) );
  INV_X1 U12292 ( .A(n10100), .ZN(n10099) );
  NAND2_X1 U12293 ( .A1(n10098), .A2(n13426), .ZN(n10096) );
  OAI21_X1 U12294 ( .B1(n10102), .B2(n10085), .A(n13432), .ZN(n10100) );
  OR2_X1 U12295 ( .A1(n19132), .A2(n10105), .ZN(n10101) );
  OAI21_X1 U12296 ( .B1(n19132), .B2(n10085), .A(n19131), .ZN(n19112) );
  NAND2_X1 U12297 ( .A1(n10761), .A2(n9698), .ZN(n10771) );
  NAND2_X1 U12298 ( .A1(n10746), .A2(n10820), .ZN(n10745) );
  NAND2_X1 U12299 ( .A1(n16297), .A2(n13397), .ZN(n19183) );
  INV_X1 U12300 ( .A(n16302), .ZN(n16334) );
  NAND2_X1 U12301 ( .A1(n12381), .A2(n12380), .ZN(n15408) );
  OR2_X1 U12302 ( .A1(n11146), .A2(n11145), .ZN(n14029) );
  OR2_X1 U12303 ( .A1(n11113), .A2(n11112), .ZN(n13911) );
  CLKBUF_X1 U12304 ( .A(n13909), .Z(n13910) );
  OR2_X1 U12305 ( .A1(n11081), .A2(n11080), .ZN(n19241) );
  OR2_X1 U12306 ( .A1(n11029), .A2(n11028), .ZN(n19253) );
  AND4_X1 U12307 ( .A1(n9676), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A3(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .A4(P2_INSTQUEUE_REG_0__4__SCAN_IN), 
        .ZN(n12427) );
  AND2_X1 U12308 ( .A1(n13737), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12428) );
  AND2_X1 U12309 ( .A1(n12701), .A2(n13539), .ZN(n19252) );
  AND3_X1 U12310 ( .A1(n15138), .A2(n10136), .A3(n10135), .ZN(n15145) );
  CLKBUF_X1 U12311 ( .A(n15159), .Z(n15160) );
  NOR2_X1 U12312 ( .A1(n19308), .A2(n19321), .ZN(n19304) );
  INV_X1 U12313 ( .A(n19325), .ZN(n19308) );
  AND2_X1 U12314 ( .A1(n19293), .A2(n9658), .ZN(n19321) );
  NOR2_X1 U12315 ( .A1(n19331), .A2(n19356), .ZN(n19339) );
  BUF_X1 U12317 ( .A(n13728), .Z(n19356) );
  INV_X1 U12318 ( .A(n19359), .ZN(n19376) );
  INV_X1 U12319 ( .A(n15569), .ZN(n19143) );
  INV_X1 U12320 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n19187) );
  INV_X1 U12321 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16470) );
  INV_X1 U12322 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16484) );
  INV_X1 U12323 ( .A(n16414), .ZN(n19399) );
  INV_X1 U12324 ( .A(n19394), .ZN(n16447) );
  AOI21_X1 U12325 ( .B1(n16302), .B2(n16525), .A(n9726), .ZN(n10214) );
  NAND2_X1 U12326 ( .A1(n15421), .A2(n16525), .ZN(n15427) );
  INV_X1 U12327 ( .A(n9843), .ZN(n15260) );
  NAND2_X1 U12328 ( .A1(n15303), .A2(n10806), .ZN(n15473) );
  OR2_X1 U12329 ( .A1(n15499), .A2(n15498), .ZN(n16382) );
  NAND2_X1 U12330 ( .A1(n9893), .A2(n9894), .ZN(n15362) );
  AND2_X1 U12331 ( .A1(n9893), .A2(n9890), .ZN(n15361) );
  NAND2_X1 U12332 ( .A1(n15382), .A2(n9897), .ZN(n9893) );
  NAND2_X1 U12333 ( .A1(n9899), .A2(n15380), .ZN(n15370) );
  NAND2_X1 U12334 ( .A1(n9900), .A2(n15379), .ZN(n9899) );
  INV_X1 U12335 ( .A(n15382), .ZN(n9900) );
  NAND2_X1 U12336 ( .A1(n10190), .A2(n9925), .ZN(n9870) );
  AND2_X1 U12337 ( .A1(n10195), .A2(n9741), .ZN(n15663) );
  NAND2_X1 U12338 ( .A1(n10195), .A2(n10729), .ZN(n15682) );
  NAND2_X1 U12339 ( .A1(n9916), .A2(n9918), .ZN(n14204) );
  NAND2_X1 U12340 ( .A1(n10608), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n16474) );
  NAND2_X1 U12341 ( .A1(n9917), .A2(n16534), .ZN(n16475) );
  NAND2_X1 U12342 ( .A1(n13618), .A2(n11182), .ZN(n16522) );
  INV_X1 U12343 ( .A(n16522), .ZN(n16502) );
  AND2_X1 U12344 ( .A1(n15575), .A2(n15581), .ZN(n16501) );
  INV_X1 U12345 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20106) );
  INV_X1 U12346 ( .A(n20094), .ZN(n20091) );
  INV_X1 U12347 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20088) );
  XNOR2_X1 U12348 ( .A(n13669), .B(n13671), .ZN(n19540) );
  AND2_X1 U12349 ( .A1(n13742), .A2(n13768), .ZN(n20074) );
  AND2_X1 U12350 ( .A1(n13261), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16543) );
  NOR2_X1 U12351 ( .A1(n19700), .A2(n19597), .ZN(n19465) );
  INV_X1 U12352 ( .A(n19564), .ZN(n19557) );
  NOR2_X1 U12353 ( .A1(n19931), .A2(n19597), .ZN(n19649) );
  OAI21_X1 U12354 ( .B1(n19664), .B2(n19672), .A(n19936), .ZN(n19696) );
  INV_X1 U12355 ( .A(n19747), .ZN(n19762) );
  NOR2_X1 U12356 ( .A1(n19837), .A2(n20071), .ZN(n19825) );
  OAI22_X1 U12357 ( .A1(n20338), .A2(n19427), .B1(n18430), .B2(n19428), .ZN(
        n19892) );
  OAI21_X1 U12358 ( .B1(n19874), .B2(n19873), .A(n19872), .ZN(n19919) );
  INV_X1 U12359 ( .A(n19779), .ZN(n19938) );
  INV_X1 U12360 ( .A(n19869), .ZN(n19928) );
  INV_X1 U12361 ( .A(n19882), .ZN(n19948) );
  INV_X1 U12362 ( .A(n19889), .ZN(n19954) );
  INV_X1 U12363 ( .A(n19895), .ZN(n19960) );
  INV_X1 U12364 ( .A(n19688), .ZN(n19972) );
  OR2_X1 U12365 ( .A1(n19837), .A2(n19931), .ZN(n19989) );
  INV_X1 U12366 ( .A(n19978), .ZN(n19985) );
  INV_X1 U12367 ( .A(n19069), .ZN(n19073) );
  NAND2_X1 U12368 ( .A1(n18840), .A2(n17656), .ZN(n19069) );
  NOR2_X1 U12369 ( .A1(n9661), .A2(n13213), .ZN(n16695) );
  NAND2_X1 U12370 ( .A1(n19054), .A2(n16690), .ZN(n17659) );
  AND2_X1 U12371 ( .A1(n9943), .A2(n17018), .ZN(n16774) );
  NAND2_X1 U12372 ( .A1(n16784), .A2(n17018), .ZN(n9939) );
  AND2_X1 U12373 ( .A1(n16794), .A2(n17018), .ZN(n16784) );
  INV_X1 U12374 ( .A(n17086), .ZN(n17065) );
  AND2_X1 U12375 ( .A1(n9933), .A2(n17018), .ZN(n16820) );
  INV_X1 U12376 ( .A(n17093), .ZN(n17083) );
  NOR2_X2 U12377 ( .A1(n19071), .A2(n18897), .ZN(n17086) );
  OAI211_X1 U12378 ( .C1(n18909), .C2(n18780), .A(n19069), .B(n16986), .ZN(
        n17094) );
  NOR2_X1 U12379 ( .A1(n16806), .A2(n17163), .ZN(n17169) );
  NOR4_X1 U12380 ( .A1(n16867), .A2(n17260), .A3(n17263), .A4(n17262), .ZN(
        n17246) );
  NAND2_X1 U12381 ( .A1(n13089), .A2(n9981), .ZN(n9980) );
  NOR2_X1 U12382 ( .A1(n17397), .A2(n17373), .ZN(n17371) );
  NOR2_X1 U12383 ( .A1(n17263), .A2(n15820), .ZN(n17416) );
  NAND2_X1 U12384 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17416), .ZN(n17415) );
  NOR4_X1 U12385 ( .A1(n17658), .A2(n14411), .A3(n15939), .A4(n18904), .ZN(
        n17435) );
  NAND2_X1 U12386 ( .A1(n17452), .A2(n17577), .ZN(n17450) );
  NAND2_X1 U12387 ( .A1(n17453), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n17452) );
  NAND2_X1 U12388 ( .A1(n17442), .A2(n9706), .ZN(n17456) );
  NAND2_X1 U12389 ( .A1(n17442), .A2(n9971), .ZN(n17464) );
  NOR2_X1 U12390 ( .A1(n17474), .A2(n17604), .ZN(n17469) );
  NOR2_X1 U12391 ( .A1(n17480), .A2(n17608), .ZN(n17479) );
  NOR4_X1 U12392 ( .A1(n17519), .A2(n17489), .A3(n17612), .A4(n17662), .ZN(
        n10240) );
  NAND2_X1 U12393 ( .A1(n17518), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n17519) );
  INV_X1 U12394 ( .A(n17577), .ZN(n17555) );
  NOR2_X1 U12395 ( .A1(n12923), .A2(n12922), .ZN(n12924) );
  NOR2_X1 U12396 ( .A1(n12943), .A2(n12942), .ZN(n12953) );
  NAND2_X1 U12397 ( .A1(n12941), .A2(n12940), .ZN(n12942) );
  INV_X1 U12398 ( .A(n17586), .ZN(n17579) );
  INV_X1 U12399 ( .A(n17587), .ZN(n17580) );
  NOR2_X1 U12400 ( .A1(n12960), .A2(n12959), .ZN(n12965) );
  OAI211_X1 U12401 ( .C1(n19050), .C2(n17658), .A(n9661), .B(n17656), .ZN(
        n17692) );
  BUF_X1 U12402 ( .A(n17692), .Z(n17703) );
  NOR2_X1 U12403 ( .A1(n17703), .A2(n17658), .ZN(n17704) );
  AND2_X1 U12404 ( .A1(n17809), .A2(n16560), .ZN(n16561) );
  INV_X1 U12405 ( .A(n17887), .ZN(n17812) );
  NOR2_X1 U12406 ( .A1(n17939), .A2(n17927), .ZN(n17920) );
  INV_X1 U12407 ( .A(n17926), .ZN(n17943) );
  INV_X1 U12408 ( .A(n17923), .ZN(n17905) );
  AND2_X1 U12409 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17986) );
  INV_X1 U12410 ( .A(n18040), .ZN(n9947) );
  INV_X1 U12411 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18019) );
  NOR2_X1 U12412 ( .A1(n18040), .A2(n18042), .ZN(n18024) );
  XNOR2_X1 U12413 ( .A(n15918), .B(n16579), .ZN(n16577) );
  NOR2_X1 U12414 ( .A1(n17735), .A2(n10211), .ZN(n15861) );
  NAND2_X1 U12415 ( .A1(n17781), .A2(n13029), .ZN(n17776) );
  NAND2_X1 U12416 ( .A1(n17820), .A2(n13030), .ZN(n17782) );
  NOR2_X1 U12417 ( .A1(n18880), .A2(n18857), .ZN(n18387) );
  NOR2_X1 U12418 ( .A1(n18209), .A2(n9801), .ZN(n18201) );
  OR2_X1 U12419 ( .A1(n18194), .A2(n9802), .ZN(n9801) );
  NOR2_X1 U12420 ( .A1(n9752), .A2(n18367), .ZN(n9802) );
  NAND2_X1 U12421 ( .A1(n18277), .A2(n18187), .ZN(n18227) );
  NAND2_X1 U12422 ( .A1(n10081), .A2(n10082), .ZN(n17948) );
  OAI21_X2 U12423 ( .B1(n14408), .B2(n18872), .A(n13152), .ZN(n18857) );
  NOR2_X1 U12424 ( .A1(n18048), .A2(n13008), .ZN(n18035) );
  INV_X1 U12425 ( .A(n18378), .ZN(n18388) );
  NOR2_X1 U12426 ( .A1(n15845), .A2(n18872), .ZN(n18859) );
  AOI21_X2 U12427 ( .B1(n13220), .B2(n13219), .A(n18904), .ZN(n18394) );
  NOR2_X1 U12428 ( .A1(n18843), .A2(n18386), .ZN(n18397) );
  OR2_X1 U12429 ( .A1(n9804), .A2(n18069), .ZN(n18400) );
  INV_X1 U12430 ( .A(n18079), .ZN(n9804) );
  INV_X1 U12431 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18864) );
  INV_X1 U12432 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18884) );
  INV_X1 U12433 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18887) );
  NOR2_X1 U12434 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19008), .ZN(
        n19032) );
  INV_X1 U12435 ( .A(n19036), .ZN(n19038) );
  INV_X1 U12436 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18849) );
  OAI211_X1 U12437 ( .C1(n18904), .C2(n18882), .A(n18409), .B(n15851), .ZN(
        n19036) );
  AND2_X1 U12439 ( .A1(n13343), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20311)
         );
  CLKBUF_X1 U12440 ( .A(n16676), .Z(n16682) );
  OAI21_X1 U12441 ( .B1(n14842), .B2(n20115), .A(n12327), .ZN(P1_U2969) );
  INV_X1 U12442 ( .A(n14922), .ZN(n16313) );
  AOI21_X1 U12443 ( .B1(n14922), .B2(n10114), .A(n10112), .ZN(n16316) );
  AOI21_X1 U12444 ( .B1(n10117), .B2(n10115), .A(n16312), .ZN(n10114) );
  INV_X1 U12445 ( .A(n10113), .ZN(n10112) );
  AND2_X1 U12446 ( .A1(n12385), .A2(n10243), .ZN(n12386) );
  INV_X1 U12447 ( .A(n12359), .ZN(n12360) );
  OAI21_X1 U12448 ( .B1(n12369), .B2(n16463), .A(n12358), .ZN(n12359) );
  NAND2_X1 U12449 ( .A1(n9728), .A2(n9874), .ZN(n15527) );
  OAI21_X1 U12450 ( .B1(n12369), .B2(n16527), .A(n10036), .ZN(n12370) );
  OAI21_X1 U12451 ( .B1(n9876), .B2(n9873), .A(n15526), .ZN(P2_U3025) );
  NAND2_X1 U12452 ( .A1(n9879), .A2(n9877), .ZN(n9876) );
  INV_X1 U12453 ( .A(n9874), .ZN(n9873) );
  OAI21_X1 U12454 ( .B1(n16734), .B2(n9791), .A(n9934), .ZN(P3_U2640) );
  AOI21_X1 U12455 ( .B1(n16739), .B2(n17104), .A(n9935), .ZN(n9934) );
  NAND2_X1 U12456 ( .A1(n9937), .A2(n9936), .ZN(n9935) );
  AOI22_X1 U12457 ( .A1(n17587), .A2(BUF2_REG_0__SCAN_IN), .B1(n17586), .B2(
        n9805), .ZN(n15944) );
  AOI21_X1 U12458 ( .B1(n17725), .B2(n17724), .A(n17723), .ZN(n17730) );
  AND2_X1 U12459 ( .A1(n13303), .A2(n10227), .ZN(n13304) );
  NAND2_X1 U12460 ( .A1(n13226), .A2(n13225), .ZN(n13235) );
  OAI211_X1 U12461 ( .C1(n18214), .C2(n18204), .A(n9799), .B(n9798), .ZN(
        P3_U2845) );
  AOI21_X1 U12462 ( .B1(n18203), .B2(n18315), .A(n18202), .ZN(n9798) );
  OR2_X1 U12463 ( .A1(n18201), .A2(n9800), .ZN(n9799) );
  NAND2_X1 U12464 ( .A1(n18380), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9800) );
  OR3_X1 U12465 ( .A1(n18909), .A2(n18908), .A3(n18907), .ZN(n18910) );
  NAND3_X2 U12466 ( .A1(n10055), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12918) );
  INV_X1 U12467 ( .A(n11407), .ZN(n11427) );
  NAND2_X1 U12468 ( .A1(n10152), .A2(n9781), .ZN(n14548) );
  INV_X1 U12469 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17988) );
  AND2_X1 U12470 ( .A1(n10179), .A2(n15077), .ZN(n9686) );
  INV_X1 U12471 ( .A(n17819), .ZN(n10059) );
  AND2_X1 U12472 ( .A1(n9649), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10612) );
  NAND2_X1 U12473 ( .A1(n15688), .A2(n9795), .ZN(n15607) );
  NAND2_X1 U12474 ( .A1(n10968), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15278) );
  AND2_X1 U12475 ( .A1(n15688), .A2(n9796), .ZN(n15366) );
  NOR2_X1 U12476 ( .A1(n14564), .A2(n14566), .ZN(n14565) );
  NOR2_X1 U12477 ( .A1(n15369), .A2(n9898), .ZN(n9897) );
  AND2_X1 U12478 ( .A1(n10082), .A2(n10080), .ZN(n9687) );
  NOR2_X1 U12479 ( .A1(n15228), .A2(n9761), .ZN(n9688) );
  OR2_X1 U12480 ( .A1(n11405), .A2(n11404), .ZN(n11499) );
  AND2_X1 U12481 ( .A1(n19422), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n9689) );
  AND2_X1 U12482 ( .A1(n11643), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9690) );
  AND2_X1 U12483 ( .A1(n9966), .A2(n9722), .ZN(n9691) );
  INV_X1 U12484 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18004) );
  OR2_X1 U12485 ( .A1(n10053), .A2(n9724), .ZN(n9692) );
  AND2_X1 U12486 ( .A1(n11563), .A2(n11588), .ZN(n11506) );
  AND2_X1 U12487 ( .A1(n10031), .A2(n9751), .ZN(n9693) );
  AND3_X1 U12488 ( .A1(n10367), .A2(n10357), .A3(n12336), .ZN(n9694) );
  INV_X1 U12489 ( .A(n12896), .ZN(n10055) );
  AND2_X1 U12490 ( .A1(n13789), .A2(n11644), .ZN(n9695) );
  AND2_X1 U12491 ( .A1(n9729), .A2(n9903), .ZN(n9696) );
  INV_X1 U12492 ( .A(n11712), .ZN(n9986) );
  NOR2_X1 U12493 ( .A1(n13759), .A2(n10138), .ZN(n9697) );
  NAND2_X1 U12494 ( .A1(n10143), .A2(n10144), .ZN(n15179) );
  NAND2_X1 U12495 ( .A1(n14274), .A2(n14273), .ZN(n14275) );
  AND2_X1 U12496 ( .A1(n15044), .A2(n9765), .ZN(n13408) );
  NAND2_X1 U12497 ( .A1(n9958), .A2(n13638), .ZN(n13690) );
  NOR2_X1 U12498 ( .A1(n13380), .A2(n15394), .ZN(n13376) );
  AND2_X1 U12499 ( .A1(n13411), .A2(n9743), .ZN(n14998) );
  AND2_X1 U12500 ( .A1(n9760), .A2(n10749), .ZN(n9698) );
  AND2_X1 U12501 ( .A1(n9949), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9699) );
  AND2_X1 U12502 ( .A1(n10119), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9700) );
  AND2_X1 U12503 ( .A1(n9778), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9701) );
  AND2_X1 U12504 ( .A1(n11153), .A2(n14353), .ZN(n9702) );
  INV_X1 U12505 ( .A(n13426), .ZN(n10085) );
  AND2_X1 U12506 ( .A1(n13424), .A2(n9787), .ZN(n13430) );
  AND2_X1 U12507 ( .A1(n10122), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9703) );
  AND2_X1 U12508 ( .A1(n13030), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9704) );
  AND2_X1 U12509 ( .A1(n9971), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n9705) );
  AND2_X1 U12510 ( .A1(n9705), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n9706) );
  NAND2_X1 U12512 ( .A1(n14815), .A2(n11753), .ZN(n14781) );
  NAND2_X1 U12513 ( .A1(n15366), .A2(n10232), .ZN(n15320) );
  INV_X1 U12514 ( .A(n9860), .ZN(n10356) );
  AND2_X1 U12515 ( .A1(n13918), .A2(n13943), .ZN(n12741) );
  CLKBUF_X3 U12516 ( .A(n12741), .Z(n13357) );
  OR2_X1 U12517 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n10814), .ZN(n9707) );
  NAND2_X1 U12518 ( .A1(n10964), .A2(n10963), .ZN(n15688) );
  AND2_X1 U12519 ( .A1(n15366), .A2(n10202), .ZN(n15295) );
  INV_X1 U12520 ( .A(n14068), .ZN(n10460) );
  NOR2_X1 U12521 ( .A1(n17473), .A2(n17606), .ZN(n17442) );
  AND2_X1 U12522 ( .A1(n10443), .A2(n10459), .ZN(n9708) );
  NAND2_X1 U12523 ( .A1(n10162), .A2(n10163), .ZN(n14629) );
  NOR2_X1 U12524 ( .A1(n14604), .A2(n10153), .ZN(n14549) );
  INV_X1 U12525 ( .A(n10068), .ZN(n17775) );
  NAND2_X1 U12526 ( .A1(n17781), .A2(n10066), .ZN(n10068) );
  AND2_X1 U12527 ( .A1(n17442), .A2(n9705), .ZN(n9709) );
  NAND2_X1 U12528 ( .A1(n10015), .A2(n11759), .ZN(n9710) );
  AND2_X1 U12529 ( .A1(n14617), .A2(n14619), .ZN(n14606) );
  AND2_X1 U12530 ( .A1(n15688), .A2(n10208), .ZN(n15657) );
  NAND2_X1 U12531 ( .A1(n14319), .A2(n14362), .ZN(n14361) );
  NAND2_X1 U12532 ( .A1(n15688), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15673) );
  AND2_X1 U12533 ( .A1(n10968), .A2(n10200), .ZN(n15265) );
  AND4_X1 U12534 ( .A1(n10396), .A2(n10399), .A3(n10247), .A4(n10403), .ZN(
        n9711) );
  NAND2_X1 U12535 ( .A1(n11662), .A2(n13874), .ZN(n9712) );
  INV_X1 U12536 ( .A(n16713), .ZN(n9970) );
  BUF_X1 U12537 ( .A(n10459), .Z(n13743) );
  NAND2_X1 U12538 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13011), .ZN(
        n9713) );
  NAND2_X1 U12539 ( .A1(n9870), .A2(n15627), .ZN(n15618) );
  NAND2_X1 U12540 ( .A1(n10959), .A2(n10958), .ZN(n16455) );
  AND2_X1 U12541 ( .A1(n17802), .A2(n16552), .ZN(n9714) );
  NAND2_X1 U12542 ( .A1(n9711), .A2(n10404), .ZN(n10431) );
  INV_X2 U12543 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14045) );
  AND4_X1 U12544 ( .A1(n11418), .A2(n11417), .A3(n11416), .A4(n11415), .ZN(
        n9715) );
  OAI21_X2 U12545 ( .B1(n10431), .B2(n10432), .A(n10439), .ZN(n15709) );
  NAND2_X1 U12546 ( .A1(n10761), .A2(n10749), .ZN(n10759) );
  XNOR2_X1 U12547 ( .A(n11185), .B(n11184), .ZN(n11183) );
  INV_X1 U12548 ( .A(n13926), .ZN(n9967) );
  AND2_X1 U12549 ( .A1(n10672), .A2(n10671), .ZN(n9716) );
  NAND2_X1 U12550 ( .A1(n10462), .A2(n10463), .ZN(n19479) );
  AND2_X1 U12551 ( .A1(n10473), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n9717) );
  INV_X1 U12552 ( .A(n14604), .ZN(n10152) );
  NAND2_X1 U12553 ( .A1(n16086), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9719) );
  AND2_X1 U12554 ( .A1(n10018), .A2(n10017), .ZN(n9720) );
  OR2_X1 U12555 ( .A1(n15285), .A2(n10826), .ZN(n9721) );
  AND2_X1 U12556 ( .A1(n13997), .A2(n14095), .ZN(n9722) );
  OR2_X1 U12557 ( .A1(n10470), .A2(n10460), .ZN(n19863) );
  NAND2_X1 U12558 ( .A1(n15688), .A2(n9840), .ZN(n15296) );
  NOR2_X1 U12559 ( .A1(n16086), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9723) );
  AND2_X1 U12560 ( .A1(n11587), .A2(n11586), .ZN(n9724) );
  OAI21_X1 U12561 ( .B1(n12339), .B2(n10205), .A(n10204), .ZN(n13319) );
  NAND2_X1 U12562 ( .A1(n9914), .A2(n10883), .ZN(n10385) );
  INV_X1 U12563 ( .A(n9891), .ZN(n9890) );
  NAND2_X1 U12564 ( .A1(n9894), .A2(n9892), .ZN(n9891) );
  NAND2_X1 U12565 ( .A1(n10796), .A2(n15327), .ZN(n9725) );
  NAND2_X1 U12566 ( .A1(n11346), .A2(n11345), .ZN(n9726) );
  AND2_X1 U12567 ( .A1(n13874), .A2(n9833), .ZN(n9727) );
  AND2_X1 U12568 ( .A1(n9879), .A2(n9878), .ZN(n9728) );
  NAND2_X1 U12569 ( .A1(n9907), .A2(n9906), .ZN(n9729) );
  NAND2_X1 U12570 ( .A1(n10162), .A2(n10160), .ZN(n9730) );
  AND2_X1 U12571 ( .A1(n14981), .A2(n14968), .ZN(n14953) );
  AND2_X1 U12572 ( .A1(n13447), .A2(n12346), .ZN(n12347) );
  AND2_X1 U12573 ( .A1(n10236), .A2(n12376), .ZN(n9731) );
  AND2_X1 U12574 ( .A1(n11751), .A2(n9719), .ZN(n9732) );
  OR2_X1 U12575 ( .A1(n11664), .A2(n11649), .ZN(n9733) );
  OR2_X1 U12576 ( .A1(n11649), .A2(n11625), .ZN(n9734) );
  AND2_X1 U12577 ( .A1(n11605), .A2(n11604), .ZN(n9735) );
  INV_X1 U12578 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14074) );
  INV_X2 U12579 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19014) );
  INV_X1 U12580 ( .A(n9909), .ZN(n9908) );
  OR2_X1 U12581 ( .A1(n9650), .A2(n9910), .ZN(n9909) );
  INV_X1 U12582 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n13484) );
  INV_X1 U12583 ( .A(n17658), .ZN(n9969) );
  BUF_X1 U12584 ( .A(n11429), .Z(n12266) );
  OR2_X1 U12585 ( .A1(n13279), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n9736) );
  NAND2_X1 U12586 ( .A1(n11607), .A2(n20753), .ZN(n13673) );
  NAND2_X1 U12587 ( .A1(n11016), .A2(n11015), .ZN(n14274) );
  NAND2_X1 U12588 ( .A1(n13841), .A2(n13840), .ZN(n13839) );
  NAND2_X1 U12589 ( .A1(n10675), .A2(n10674), .ZN(n10719) );
  INV_X1 U12590 ( .A(n17018), .ZN(n17048) );
  NOR2_X1 U12591 ( .A1(n17959), .A2(n10059), .ZN(n17960) );
  NAND2_X1 U12592 ( .A1(n15044), .A2(n10024), .ZN(n15029) );
  NAND2_X1 U12593 ( .A1(n10171), .A2(n10175), .ZN(n13905) );
  AND2_X1 U12594 ( .A1(n10143), .A2(n10141), .ZN(n9737) );
  NOR2_X1 U12595 ( .A1(n17532), .A2(n17707), .ZN(n17518) );
  AND2_X1 U12596 ( .A1(n10091), .A2(n10092), .ZN(n9738) );
  NAND2_X1 U12597 ( .A1(n14352), .A2(n14353), .ZN(n14351) );
  AOI21_X1 U12598 ( .B1(n19100), .B2(n13426), .A(n15871), .ZN(n14976) );
  AND2_X1 U12599 ( .A1(n10081), .A2(n9687), .ZN(n9739) );
  NAND2_X1 U12600 ( .A1(n10175), .A2(n10174), .ZN(n9740) );
  NOR2_X1 U12601 ( .A1(n15027), .A2(n13412), .ZN(n13411) );
  NOR2_X1 U12602 ( .A1(n15021), .A2(n15020), .ZN(n14352) );
  BUF_X1 U12603 ( .A(n10354), .Z(n13764) );
  NAND2_X1 U12604 ( .A1(n13411), .A2(n15008), .ZN(n15009) );
  NOR2_X1 U12605 ( .A1(n17439), .A2(n17438), .ZN(n17526) );
  AND2_X1 U12606 ( .A1(n14274), .A2(n10028), .ZN(n15064) );
  NAND2_X1 U12607 ( .A1(n14352), .A2(n9702), .ZN(n14994) );
  NAND2_X1 U12608 ( .A1(n15504), .A2(n10035), .ZN(n14963) );
  AND2_X1 U12609 ( .A1(n10729), .A2(n10194), .ZN(n9741) );
  INV_X1 U12610 ( .A(n11499), .ZN(n11563) );
  OR2_X1 U12611 ( .A1(n12430), .A2(n10138), .ZN(n9742) );
  OAI211_X1 U12612 ( .C1(n10045), .C2(n9810), .A(n9808), .B(n16119), .ZN(
        n14331) );
  NOR2_X1 U12613 ( .A1(n13805), .A2(n10999), .ZN(n15108) );
  NAND2_X1 U12614 ( .A1(n9851), .A2(n10951), .ZN(n15389) );
  NAND2_X1 U12615 ( .A1(n13486), .A2(n10591), .ZN(n11309) );
  AND2_X1 U12616 ( .A1(n10170), .A2(n15008), .ZN(n9743) );
  AND2_X1 U12617 ( .A1(n9743), .A2(n14999), .ZN(n9744) );
  INV_X1 U12618 ( .A(n15627), .ZN(n9924) );
  AND2_X1 U12619 ( .A1(n16086), .A2(n12887), .ZN(n9745) );
  INV_X1 U12620 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10588) );
  NOR2_X2 U12621 ( .A1(n14471), .A2(n20372), .ZN(n13501) );
  AND2_X1 U12622 ( .A1(n11496), .A2(n11529), .ZN(n11771) );
  OR2_X1 U12623 ( .A1(n13380), .A2(n10128), .ZN(n9746) );
  AND3_X1 U12624 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n9747) );
  OR2_X1 U12625 ( .A1(n14009), .A2(n11748), .ZN(n9748) );
  INV_X1 U12626 ( .A(n10105), .ZN(n13426) );
  AND2_X1 U12627 ( .A1(n10101), .A2(n10102), .ZN(n9749) );
  AND2_X1 U12628 ( .A1(n15319), .A2(n9887), .ZN(n9750) );
  AND2_X1 U12629 ( .A1(n14214), .A2(n14301), .ZN(n9751) );
  NOR2_X1 U12630 ( .A1(n18213), .A2(n18189), .ZN(n9752) );
  AND2_X1 U12631 ( .A1(n9884), .A2(n9885), .ZN(n9753) );
  AND2_X1 U12632 ( .A1(n9918), .A2(n9915), .ZN(n9754) );
  INV_X1 U12633 ( .A(n9897), .ZN(n9896) );
  OR2_X1 U12634 ( .A1(n14408), .A2(n13151), .ZN(n9755) );
  AND2_X1 U12635 ( .A1(n9974), .A2(n9973), .ZN(n9756) );
  AND2_X1 U12636 ( .A1(n9939), .A2(n9942), .ZN(n9757) );
  INV_X1 U12637 ( .A(n14564), .ZN(n10162) );
  AND2_X1 U12638 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n9758) );
  INV_X1 U12639 ( .A(n10193), .ZN(n10192) );
  NAND2_X1 U12640 ( .A1(n15665), .A2(n9741), .ZN(n10193) );
  OR2_X1 U12641 ( .A1(n15643), .A2(n15646), .ZN(n9759) );
  OR2_X1 U12642 ( .A1(n10974), .A2(n15014), .ZN(n9760) );
  AND2_X1 U12643 ( .A1(n16338), .A2(n12600), .ZN(n9761) );
  AND2_X1 U12644 ( .A1(n15504), .A2(n15505), .ZN(n14982) );
  AND2_X1 U12645 ( .A1(n15044), .A2(n10025), .ZN(n9762) );
  AND2_X1 U12646 ( .A1(n9744), .A2(n15182), .ZN(n9763) );
  AND2_X1 U12647 ( .A1(n14647), .A2(n14648), .ZN(n9764) );
  AND2_X1 U12648 ( .A1(n10024), .A2(n11132), .ZN(n9765) );
  AND2_X1 U12649 ( .A1(n9997), .A2(n9996), .ZN(n9766) );
  AND2_X1 U12650 ( .A1(n9931), .A2(n17018), .ZN(n9767) );
  AND2_X1 U12651 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n9768) );
  OR2_X1 U12652 ( .A1(n9742), .A2(n10137), .ZN(n9769) );
  NAND2_X2 U12653 ( .A1(n13228), .A2(n16559), .ZN(n17819) );
  NOR2_X1 U12654 ( .A1(n13427), .A2(n13425), .ZN(n9770) );
  NOR2_X1 U12655 ( .A1(n10999), .A2(n10032), .ZN(n10031) );
  NAND2_X1 U12656 ( .A1(n15044), .A2(n15650), .ZN(n15630) );
  INV_X1 U12657 ( .A(n13927), .ZN(n9965) );
  NOR2_X1 U12658 ( .A1(n13759), .A2(n9742), .ZN(n9771) );
  AND2_X1 U12659 ( .A1(n9965), .A2(n9966), .ZN(n9772) );
  AND2_X1 U12660 ( .A1(n13385), .A2(n10119), .ZN(n9773) );
  BUF_X1 U12661 ( .A(n9660), .Z(n12686) );
  NAND2_X1 U12662 ( .A1(n10971), .A2(n9676), .ZN(n16490) );
  AND2_X1 U12663 ( .A1(n10035), .A2(n10034), .ZN(n9774) );
  AND2_X1 U12664 ( .A1(n10188), .A2(n10187), .ZN(n9775) );
  NAND2_X1 U12665 ( .A1(n10388), .A2(n9694), .ZN(n13392) );
  AND2_X1 U12666 ( .A1(n13433), .A2(n10122), .ZN(n9776) );
  AND2_X1 U12667 ( .A1(n9978), .A2(n14601), .ZN(n9777) );
  NAND2_X1 U12668 ( .A1(n11012), .A2(n11011), .ZN(n15698) );
  AND2_X1 U12669 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n9778) );
  AOI21_X1 U12670 ( .B1(n13426), .B2(n19148), .A(n9770), .ZN(n19132) );
  NOR2_X1 U12671 ( .A1(n13434), .A2(n15297), .ZN(n13433) );
  AND2_X1 U12672 ( .A1(n14920), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13317) );
  AND2_X1 U12673 ( .A1(n10132), .A2(n12600), .ZN(n9779) );
  AND2_X1 U12674 ( .A1(n11831), .A2(n11848), .ZN(n10216) );
  OR2_X1 U12675 ( .A1(n13759), .A2(n12429), .ZN(n9780) );
  INV_X1 U12676 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9963) );
  AND2_X1 U12677 ( .A1(n12131), .A2(n12130), .ZN(n9781) );
  AND2_X1 U12678 ( .A1(n15898), .A2(n14483), .ZN(n20250) );
  INV_X1 U12679 ( .A(n20250), .ZN(n20115) );
  NAND2_X1 U12680 ( .A1(n17981), .A2(n18286), .ZN(n9782) );
  NAND3_X1 U12681 ( .A1(n9829), .A2(n9826), .A3(n9825), .ZN(n11539) );
  INV_X1 U12682 ( .A(n11539), .ZN(n9955) );
  NOR2_X1 U12683 ( .A1(n13772), .A2(n10180), .ZN(n9783) );
  AND2_X1 U12684 ( .A1(n13806), .A2(n10031), .ZN(n9784) );
  AND2_X1 U12685 ( .A1(n10156), .A2(n10155), .ZN(n9785) );
  AND2_X1 U12686 ( .A1(n9774), .A2(n10033), .ZN(n9786) );
  AND2_X1 U12687 ( .A1(n9701), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9787) );
  AND2_X1 U12688 ( .A1(n9775), .A2(n10186), .ZN(n9788) );
  AND2_X1 U12689 ( .A1(n9702), .A2(n11155), .ZN(n9789) );
  INV_X1 U12690 ( .A(n10807), .ZN(n10003) );
  INV_X1 U12691 ( .A(n17078), .ZN(n17060) );
  AND2_X1 U12692 ( .A1(n17713), .A2(n9949), .ZN(n9790) );
  OR3_X1 U12693 ( .A1(n17048), .A2(n16735), .A3(n18913), .ZN(n9791) );
  AND2_X2 U12694 ( .A1(n9985), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13702) );
  INV_X1 U12695 ( .A(n15146), .ZN(n10136) );
  NOR2_X1 U12696 ( .A1(n18035), .A2(n18034), .ZN(n9792) );
  AND2_X1 U12697 ( .A1(n11511), .A2(n11510), .ZN(n9793) );
  NOR2_X1 U12698 ( .A1(n14069), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10490) );
  INV_X1 U12699 ( .A(n10111), .ZN(n10110) );
  NAND2_X1 U12700 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10111) );
  INV_X1 U12701 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9985) );
  AND2_X1 U12702 ( .A1(n10110), .A2(n10109), .ZN(n9794) );
  AND2_X1 U12703 ( .A1(n10208), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9795) );
  AND2_X1 U12704 ( .A1(n9795), .A2(n9841), .ZN(n9796) );
  AND2_X1 U12705 ( .A1(n10200), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9797) );
  INV_X1 U12706 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18042) );
  INV_X1 U12707 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10013) );
  INV_X1 U12708 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10080) );
  INV_X1 U12709 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10067) );
  INV_X1 U12710 ( .A(n14735), .ZN(n9814) );
  INV_X1 U12711 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9946) );
  INV_X1 U12712 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n9815) );
  INV_X1 U12713 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10109) );
  INV_X1 U12714 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n9972) );
  INV_X1 U12715 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9951) );
  INV_X1 U12716 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10120) );
  INV_X1 U12717 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n9991) );
  NOR2_X1 U12718 ( .A1(n16344), .A2(n10145), .ZN(n10144) );
  NOR2_X1 U12719 ( .A1(n14348), .A2(n16344), .ZN(n15178) );
  OAI22_X2 U12720 ( .A1(n21027), .A2(n20368), .B1(n14356), .B2(n20370), .ZN(
        n20835) );
  NAND2_X1 U12721 ( .A1(n20313), .A2(n20312), .ZN(n20368) );
  AOI22_X2 U12722 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19437), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19436), .ZN(n19971) );
  OAI22_X2 U12723 ( .A1(n21108), .A2(n20368), .B1(n20333), .B2(n20370), .ZN(
        n20841) );
  AOI22_X2 U12724 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19437), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19436), .ZN(n19913) );
  NOR2_X2 U12725 ( .A1(n14108), .A2(n16414), .ZN(n19436) );
  NOR4_X4 U12726 ( .A1(n19018), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(
        P3_STATE2_REG_0__SCAN_IN), .A4(P3_STATEBS16_REG_SCAN_IN), .ZN(n17070)
         );
  INV_X1 U12727 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19018) );
  NOR2_X2 U12728 ( .A1(n20373), .A2(n11531), .ZN(n20864) );
  AND2_X2 U12729 ( .A1(n17078), .A2(n9807), .ZN(n14415) );
  NAND2_X2 U12730 ( .A1(n9811), .A2(n11522), .ZN(n10009) );
  NAND2_X2 U12731 ( .A1(n11515), .A2(n11520), .ZN(n11598) );
  AOI21_X1 U12732 ( .B1(n14763), .B2(n9815), .A(n9814), .ZN(n9812) );
  INV_X1 U12733 ( .A(n14763), .ZN(n9813) );
  INV_X1 U12734 ( .A(n9816), .ZN(n14748) );
  NAND2_X1 U12735 ( .A1(n14725), .A2(n16110), .ZN(n9816) );
  NAND2_X2 U12736 ( .A1(n14764), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14725) );
  NAND2_X1 U12737 ( .A1(n14725), .A2(n14763), .ZN(n16063) );
  NAND3_X1 U12738 ( .A1(n9818), .A2(n9817), .A3(n9819), .ZN(n13895) );
  NAND2_X1 U12739 ( .A1(n9695), .A2(n13790), .ZN(n9818) );
  NAND2_X2 U12740 ( .A1(n9823), .A2(n9953), .ZN(n14778) );
  NAND3_X1 U12741 ( .A1(n11607), .A2(n20971), .A3(n20753), .ZN(n9824) );
  NAND3_X1 U12743 ( .A1(n11597), .A2(n11598), .A3(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9825) );
  NAND3_X1 U12744 ( .A1(n9831), .A2(n9830), .A3(n11519), .ZN(n9829) );
  INV_X1 U12745 ( .A(n11597), .ZN(n9830) );
  INV_X1 U12746 ( .A(n11598), .ZN(n9831) );
  NAND2_X1 U12747 ( .A1(n12387), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12388) );
  NAND2_X1 U12748 ( .A1(n10969), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12339) );
  NAND2_X1 U12749 ( .A1(n10969), .A2(n9842), .ZN(n9843) );
  OR2_X1 U12750 ( .A1(n15416), .A2(n16463), .ZN(n10238) );
  NAND3_X1 U12751 ( .A1(n10517), .A2(n9845), .A3(n10518), .ZN(n9844) );
  NAND3_X1 U12752 ( .A1(n9850), .A2(n9848), .A3(n9847), .ZN(n9846) );
  INV_X1 U12753 ( .A(n10508), .ZN(n9847) );
  NAND2_X1 U12754 ( .A1(n9852), .A2(n10950), .ZN(n15400) );
  NAND2_X1 U12755 ( .A1(n10951), .A2(n10949), .ZN(n9852) );
  INV_X1 U12756 ( .A(n10950), .ZN(n9718) );
  NAND3_X1 U12757 ( .A1(n10462), .A2(n13653), .A3(n10473), .ZN(n19603) );
  AND2_X2 U12758 ( .A1(n10395), .A2(n10394), .ZN(n10411) );
  NAND2_X1 U12759 ( .A1(n10315), .A2(n14045), .ZN(n9856) );
  NAND2_X2 U12760 ( .A1(n10291), .A2(n10290), .ZN(n9860) );
  NOR2_X1 U12761 ( .A1(n9658), .A2(n10361), .ZN(n9861) );
  INV_X1 U12762 ( .A(n11183), .ZN(n9865) );
  NAND3_X1 U12763 ( .A1(n9865), .A2(n10185), .A3(n10426), .ZN(n9864) );
  NAND2_X1 U12764 ( .A1(n9865), .A2(n9866), .ZN(n11187) );
  XNOR2_X2 U12765 ( .A(n10952), .B(n10953), .ZN(n10948) );
  NAND2_X1 U12766 ( .A1(n10190), .A2(n9871), .ZN(n9867) );
  NAND2_X1 U12767 ( .A1(n9867), .A2(n9868), .ZN(n16391) );
  AOI21_X1 U12768 ( .B1(n15344), .B2(n15342), .A(n15314), .ZN(n15329) );
  NAND2_X1 U12769 ( .A1(n15258), .A2(n9904), .ZN(n9902) );
  OAI211_X1 U12770 ( .C1(n15258), .C2(n9909), .A(n9696), .B(n9902), .ZN(n13322) );
  NAND2_X1 U12771 ( .A1(n15258), .A2(n15256), .ZN(n12373) );
  OAI21_X1 U12772 ( .B1(n13322), .B2(n16465), .A(n9913), .ZN(P2_U2983) );
  NOR2_X1 U12773 ( .A1(n9911), .A2(n9905), .ZN(n9904) );
  INV_X1 U12774 ( .A(n15256), .ZN(n9905) );
  INV_X2 U12775 ( .A(n10354), .ZN(n10357) );
  OAI21_X2 U12776 ( .B1(n10190), .B2(n9922), .A(n9920), .ZN(n15515) );
  NAND2_X1 U12777 ( .A1(n10190), .A2(n10189), .ZN(n15625) );
  INV_X1 U12778 ( .A(n10189), .ZN(n9926) );
  NAND2_X1 U12779 ( .A1(n15515), .A2(n15512), .ZN(n10804) );
  NAND2_X2 U12780 ( .A1(n10365), .A2(n13752), .ZN(n11300) );
  NOR2_X2 U12781 ( .A1(n12329), .A2(n9721), .ZN(n10833) );
  NAND2_X1 U12782 ( .A1(n9930), .A2(n9931), .ZN(n16819) );
  INV_X1 U12783 ( .A(n9933), .ZN(n16830) );
  INV_X1 U12784 ( .A(n9943), .ZN(n16783) );
  NAND4_X1 U12785 ( .A1(n17986), .A2(n9945), .A3(n9944), .A4(n9747), .ZN(
        n17877) );
  NAND3_X1 U12786 ( .A1(n9947), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18014) );
  NAND2_X1 U12787 ( .A1(n9956), .A2(n9733), .ZN(n11622) );
  NAND3_X1 U12788 ( .A1(n9958), .A2(n20971), .A3(n13638), .ZN(n9956) );
  NAND2_X2 U12789 ( .A1(n9957), .A2(n9959), .ZN(n13638) );
  NAND2_X1 U12790 ( .A1(n11539), .A2(n11605), .ZN(n9959) );
  NAND2_X1 U12791 ( .A1(n9962), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14726) );
  AND2_X2 U12792 ( .A1(n9963), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11360) );
  NOR2_X4 U12793 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11366) );
  OAI21_X2 U12794 ( .B1(n18868), .B2(n18439), .A(n9970), .ZN(n18872) );
  AOI21_X2 U12795 ( .B1(n9970), .B2(n9968), .A(n13154), .ZN(n13152) );
  NAND2_X1 U12796 ( .A1(n17479), .A2(n17527), .ZN(n17473) );
  NAND2_X1 U12797 ( .A1(n10240), .A2(P3_EAX_REG_22__SCAN_IN), .ZN(n17480) );
  INV_X1 U12798 ( .A(n9975), .ZN(n14635) );
  AOI211_X2 U12799 ( .C1(n15852), .C2(n9979), .A(n19057), .B(n18841), .ZN(
        n15941) );
  AND2_X2 U12800 ( .A1(n17078), .A2(n9984), .ZN(n13117) );
  AOI21_X2 U12801 ( .B1(n10046), .B2(n10047), .A(n9987), .ZN(n10044) );
  NAND3_X1 U12802 ( .A1(n11734), .A2(n11884), .A3(n11773), .ZN(n11730) );
  AND2_X4 U12803 ( .A1(n13747), .A2(n9673), .ZN(n10485) );
  XNOR2_X2 U12804 ( .A(n10009), .B(n11568), .ZN(n11840) );
  INV_X1 U12805 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10010) );
  OAI21_X2 U12806 ( .B1(n14778), .B2(n10011), .A(n16086), .ZN(n14763) );
  NAND3_X1 U12807 ( .A1(n10217), .A2(n11766), .A3(n15934), .ZN(n10011) );
  NAND2_X1 U12808 ( .A1(n11765), .A2(n16110), .ZN(n14764) );
  NAND2_X1 U12809 ( .A1(n12712), .A2(n16086), .ZN(n10023) );
  NAND2_X1 U12810 ( .A1(n14274), .A2(n10027), .ZN(n15041) );
  NAND2_X1 U12811 ( .A1(n13806), .A2(n9693), .ZN(n11012) );
  NAND2_X1 U12812 ( .A1(n14352), .A2(n9789), .ZN(n15529) );
  AND2_X2 U12813 ( .A1(n15504), .A2(n9786), .ZN(n15209) );
  INV_X1 U12814 ( .A(n14846), .ZN(n10042) );
  MUX2_X1 U12815 ( .A(n16110), .B(n14717), .S(n10043), .Z(n14718) );
  NAND2_X1 U12816 ( .A1(n16134), .A2(n10046), .ZN(n10045) );
  NOR2_X1 U12817 ( .A1(n10052), .A2(n20971), .ZN(n10049) );
  NAND2_X1 U12818 ( .A1(n11840), .A2(n10051), .ZN(n10050) );
  NOR2_X1 U12819 ( .A1(n11584), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10051) );
  NAND3_X1 U12820 ( .A1(n14725), .A2(n14763), .A3(n16143), .ZN(n14746) );
  NAND3_X1 U12821 ( .A1(n14725), .A2(n14763), .A3(n10054), .ZN(n11767) );
  INV_X2 U12822 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19031) );
  NAND2_X1 U12823 ( .A1(n18034), .A2(n9713), .ZN(n10056) );
  NOR2_X1 U12824 ( .A1(n13036), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17733) );
  NAND2_X1 U12825 ( .A1(n18017), .A2(n10073), .ZN(n10072) );
  NOR2_X1 U12826 ( .A1(n18015), .A2(n13017), .ZN(n13019) );
  INV_X1 U12827 ( .A(n13017), .ZN(n10077) );
  INV_X1 U12828 ( .A(n17959), .ZN(n10081) );
  INV_X1 U12829 ( .A(n14976), .ZN(n10086) );
  OAI21_X1 U12830 ( .B1(n14976), .B2(n10105), .A(n13435), .ZN(n14977) );
  NAND3_X1 U12831 ( .A1(n10107), .A2(n10106), .A3(n10108), .ZN(n13388) );
  NAND2_X1 U12832 ( .A1(n14920), .A2(n9794), .ZN(n10106) );
  OR2_X1 U12833 ( .A1(n14920), .A2(n10109), .ZN(n10107) );
  AOI21_X1 U12834 ( .B1(n13388), .B2(n14091), .A(n13387), .ZN(n10105) );
  INV_X1 U12835 ( .A(n13380), .ZN(n10124) );
  NAND2_X1 U12836 ( .A1(n10124), .A2(n10125), .ZN(n13382) );
  NAND2_X1 U12837 ( .A1(n12664), .A2(n12663), .ZN(n10135) );
  AOI21_X2 U12838 ( .B1(n15138), .B2(n15146), .A(n10134), .ZN(n10133) );
  NAND2_X1 U12839 ( .A1(n15138), .A2(n10135), .ZN(n15147) );
  OR2_X2 U12840 ( .A1(n13759), .A2(n9769), .ZN(n13909) );
  INV_X1 U12841 ( .A(n14348), .ZN(n10143) );
  NAND2_X1 U12842 ( .A1(n11300), .A2(n9768), .ZN(n10374) );
  NAND3_X1 U12843 ( .A1(n11509), .A2(n14479), .A3(n12741), .ZN(n13323) );
  NAND3_X1 U12844 ( .A1(n10147), .A2(n13841), .A3(n13840), .ZN(n13932) );
  AND2_X1 U12845 ( .A1(n9735), .A2(n11606), .ZN(n10149) );
  AND2_X2 U12846 ( .A1(n14319), .A2(n9785), .ZN(n14372) );
  AND2_X1 U12847 ( .A1(n14519), .A2(n10167), .ZN(n14506) );
  NAND2_X1 U12848 ( .A1(n14519), .A2(n10166), .ZN(n13308) );
  NAND2_X1 U12849 ( .A1(n14519), .A2(n10165), .ZN(n12395) );
  NAND2_X1 U12850 ( .A1(n10358), .A2(n10361), .ZN(n10889) );
  NAND3_X1 U12851 ( .A1(n10889), .A2(n13279), .A3(n10887), .ZN(n11306) );
  NAND2_X1 U12852 ( .A1(n11306), .A2(n9860), .ZN(n10377) );
  NAND2_X1 U12853 ( .A1(n13411), .A2(n9763), .ZN(n15181) );
  INV_X1 U12854 ( .A(n15049), .ZN(n10171) );
  NAND2_X1 U12855 ( .A1(n10171), .A2(n10172), .ZN(n15027) );
  INV_X1 U12856 ( .A(n13772), .ZN(n10178) );
  NAND2_X1 U12857 ( .A1(n10178), .A2(n9686), .ZN(n13832) );
  NAND2_X1 U12858 ( .A1(n14981), .A2(n10188), .ZN(n14952) );
  OAI21_X2 U12859 ( .B1(n10948), .B2(n11014), .A(n19202), .ZN(n10715) );
  AND3_X2 U12860 ( .A1(n14074), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10284) );
  INV_X1 U12861 ( .A(n10559), .ZN(n10199) );
  NAND2_X1 U12862 ( .A1(n10199), .A2(n10558), .ZN(n10935) );
  NAND2_X1 U12863 ( .A1(n10968), .A2(n9797), .ZN(n12340) );
  INV_X1 U12864 ( .A(n12340), .ZN(n10969) );
  INV_X1 U12865 ( .A(n15296), .ZN(n10967) );
  NAND2_X1 U12866 ( .A1(n10206), .A2(n10970), .ZN(n10205) );
  INV_X1 U12867 ( .A(n10207), .ZN(n10206) );
  OR2_X1 U12868 ( .A1(n9675), .A2(n11838), .ZN(n20749) );
  AND2_X1 U12869 ( .A1(n12267), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11442) );
  CLKBUF_X1 U12870 ( .A(n12577), .Z(n16338) );
  AND3_X1 U12871 ( .A1(n11531), .A2(n11505), .A3(n11510), .ZN(n11507) );
  INV_X1 U12872 ( .A(n12370), .ZN(n12371) );
  NAND2_X1 U12873 ( .A1(n11860), .A2(n11967), .ZN(n11867) );
  AOI21_X1 U12874 ( .B1(n12302), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n11442), .ZN(n11443) );
  INV_X1 U12875 ( .A(n15408), .ZN(n14929) );
  INV_X1 U12876 ( .A(n10439), .ZN(n10440) );
  OR2_X1 U12877 ( .A1(n13871), .A2(n20305), .ZN(n20675) );
  NAND2_X1 U12878 ( .A1(n20305), .A2(n11830), .ZN(n20448) );
  NAND2_X1 U12879 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20106), .ZN(
        n10596) );
  NOR3_X2 U12880 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(n12539), .ZN(n11088) );
  INV_X1 U12881 ( .A(n10952), .ZN(n10955) );
  NAND2_X1 U12882 ( .A1(n10462), .A2(n10461), .ZN(n10641) );
  OR2_X2 U12883 ( .A1(n11436), .A2(n11435), .ZN(n11508) );
  OR2_X1 U12884 ( .A1(n11634), .A2(n11633), .ZN(n11635) );
  AND2_X4 U12885 ( .A1(n11366), .A2(n13704), .ZN(n12265) );
  INV_X1 U12886 ( .A(n15288), .ZN(n10968) );
  XNOR2_X1 U12887 ( .A(n11833), .B(n11832), .ZN(n13866) );
  OR2_X1 U12888 ( .A1(n11662), .A2(n13874), .ZN(n11663) );
  NAND2_X1 U12889 ( .A1(n10437), .A2(n10439), .ZN(n10414) );
  NOR2_X1 U12890 ( .A1(n20635), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10210) );
  OR2_X1 U12891 ( .A1(n17819), .A2(n15858), .ZN(n10211) );
  OR2_X1 U12892 ( .A1(n17819), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10212) );
  NAND2_X1 U12893 ( .A1(n14446), .A2(n19260), .ZN(n10213) );
  AND2_X1 U12894 ( .A1(n10386), .A2(n19411), .ZN(n10215) );
  INV_X1 U12895 ( .A(n11824), .ZN(n12315) );
  INV_X1 U12896 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20081) );
  INV_X1 U12897 ( .A(n12016), .ZN(n11967) );
  INV_X1 U12898 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11934) );
  AND2_X1 U12899 ( .A1(n16174), .A2(n14893), .ZN(n10217) );
  AND4_X1 U12900 ( .A1(n10647), .A2(n10646), .A3(n10645), .A4(n10644), .ZN(
        n10218) );
  OR2_X1 U12901 ( .A1(n14442), .A2(n20254), .ZN(n10219) );
  INV_X1 U12902 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11776) );
  INV_X1 U12903 ( .A(n14655), .ZN(n14001) );
  INV_X1 U12904 ( .A(n11843), .ZN(n11893) );
  NAND2_X1 U12905 ( .A1(n12343), .A2(n9666), .ZN(n16463) );
  AND2_X1 U12906 ( .A1(n13388), .A2(n16473), .ZN(n10220) );
  NOR2_X1 U12907 ( .A1(n10059), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10221) );
  OR2_X1 U12908 ( .A1(n17367), .A2(n17305), .ZN(n10222) );
  OR2_X1 U12909 ( .A1(n17303), .A2(n17395), .ZN(n10223) );
  OR2_X1 U12910 ( .A1(n17396), .A2(n17313), .ZN(n10224) );
  OR3_X1 U12911 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17797), .ZN(n10225) );
  AND2_X1 U12912 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_14__SCAN_IN), 
        .ZN(n10226) );
  INV_X1 U12913 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10970) );
  AND2_X1 U12914 ( .A1(n13302), .A2(n13301), .ZN(n10227) );
  NOR2_X1 U12915 ( .A1(n13048), .A2(n13047), .ZN(n10228) );
  INV_X1 U12916 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17427) );
  AND2_X1 U12917 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10229) );
  AND2_X1 U12918 ( .A1(n11763), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10230) );
  XOR2_X1 U12919 ( .A(n13366), .B(n13365), .Z(n10231) );
  INV_X1 U12920 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19926) );
  NAND2_X1 U12921 ( .A1(n14633), .A2(n20372), .ZN(n14643) );
  INV_X1 U12922 ( .A(n14643), .ZN(n13368) );
  AND3_X1 U12923 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10232) );
  AND2_X1 U12924 ( .A1(n12640), .A2(n13769), .ZN(n10233) );
  NAND2_X1 U12925 ( .A1(n12324), .A2(n20968), .ZN(n10234) );
  AND4_X1 U12926 ( .A1(n12964), .A2(n12963), .A3(n12962), .A4(n12961), .ZN(
        n10235) );
  INV_X1 U12927 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13001) );
  INV_X2 U12928 ( .A(n17432), .ZN(n17423) );
  INV_X1 U12929 ( .A(n19129), .ZN(n19226) );
  AND2_X1 U12930 ( .A1(n12374), .A2(n15257), .ZN(n10236) );
  NOR3_X1 U12931 ( .A1(n16105), .A2(n14805), .A3(n16102), .ZN(n10237) );
  AND2_X1 U12932 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10239) );
  OR3_X1 U12933 ( .A1(n15440), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15424), .ZN(n10241) );
  OR3_X1 U12934 ( .A1(n15440), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15413), .ZN(n10242) );
  OR2_X1 U12935 ( .A1(n12384), .A2(n19405), .ZN(n10243) );
  AND2_X1 U12936 ( .A1(n19183), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10244) );
  AND2_X1 U12937 ( .A1(n12706), .A2(n12705), .ZN(n10245) );
  NAND2_X1 U12938 ( .A1(n11281), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10247) );
  AND4_X1 U12939 ( .A1(n10654), .A2(n10653), .A3(n10652), .A4(n10651), .ZN(
        n10248) );
  INV_X1 U12940 ( .A(n15366), .ZN(n16393) );
  AND2_X1 U12941 ( .A1(n11410), .A2(n11409), .ZN(n10249) );
  AND2_X1 U12942 ( .A1(n11842), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10250) );
  OAI22_X1 U12943 ( .A1(n12485), .A2(n10650), .B1(n19924), .B2(n12482), .ZN(
        n10458) );
  NAND2_X1 U12944 ( .A1(n10649), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10507) );
  NOR2_X1 U12945 ( .A1(n19603), .A2(n10475), .ZN(n10476) );
  OAI22_X1 U12946 ( .A1(n11525), .A2(n11511), .B1(n20316), .B2(n13629), .ZN(
        n11501) );
  INV_X1 U12947 ( .A(n11792), .ZN(n11806) );
  OR2_X1 U12948 ( .A1(n11700), .A2(n11699), .ZN(n11726) );
  NAND2_X1 U12949 ( .A1(n10283), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10291) );
  INV_X1 U12950 ( .A(n11790), .ZN(n11787) );
  NAND2_X1 U12951 ( .A1(n11778), .A2(n11777), .ZN(n11785) );
  INV_X1 U12952 ( .A(n14265), .ZN(n11923) );
  NOR2_X1 U12953 ( .A1(n12849), .A2(n12864), .ZN(n12855) );
  NAND2_X1 U12954 ( .A1(n12856), .A2(n11494), .ZN(n11419) );
  NAND2_X1 U12955 ( .A1(n19422), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10592) );
  NAND2_X1 U12956 ( .A1(n11318), .A2(n10356), .ZN(n10376) );
  AND2_X1 U12957 ( .A1(n10372), .A2(n10371), .ZN(n10373) );
  NOR2_X1 U12958 ( .A1(n14414), .A2(n17348), .ZN(n12939) );
  NAND2_X1 U12959 ( .A1(n17321), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n13045) );
  AND2_X1 U12960 ( .A1(n11783), .A2(n11782), .ZN(n12721) );
  INV_X1 U12961 ( .A(n12196), .ZN(n12197) );
  INV_X1 U12962 ( .A(n14318), .ZN(n11939) );
  OR2_X1 U12963 ( .A1(n11722), .A2(n11721), .ZN(n11735) );
  INV_X1 U12964 ( .A(n11619), .ZN(n11664) );
  INV_X1 U12965 ( .A(n11747), .ZN(n11585) );
  AND4_X1 U12966 ( .A1(n11370), .A2(n11369), .A3(n11368), .A4(n11367), .ZN(
        n11371) );
  INV_X1 U12967 ( .A(n13749), .ZN(n12555) );
  OR2_X1 U12968 ( .A1(n12412), .A2(n12411), .ZN(n12413) );
  AND2_X1 U12969 ( .A1(n12641), .A2(n10233), .ZN(n12642) );
  INV_X1 U12970 ( .A(n12622), .ZN(n12623) );
  AND2_X1 U12971 ( .A1(n12600), .A2(n12599), .ZN(n12601) );
  INV_X1 U12972 ( .A(n10948), .ZN(n10946) );
  NAND2_X1 U12973 ( .A1(n14314), .A2(n10948), .ZN(n10949) );
  NAND2_X1 U12974 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12946) );
  NOR2_X1 U12975 ( .A1(n17396), .A2(n17359), .ZN(n12954) );
  AOI21_X1 U12976 ( .B1(n11783), .B2(n11780), .A(n11782), .ZN(n12723) );
  OR2_X1 U12977 ( .A1(n12287), .A2(n14721), .ZN(n12397) );
  AND2_X1 U12978 ( .A1(n12197), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12198) );
  OR2_X1 U12979 ( .A1(n11649), .A2(n11585), .ZN(n11744) );
  INV_X1 U12980 ( .A(n14792), .ZN(n11757) );
  NAND2_X1 U12981 ( .A1(n12624), .A2(n12623), .ZN(n12625) );
  INV_X1 U12982 ( .A(n13121), .ZN(n13122) );
  INV_X1 U12983 ( .A(n12944), .ZN(n12951) );
  NAND2_X1 U12984 ( .A1(n10059), .A2(n18213), .ZN(n13023) );
  AND2_X1 U12985 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13016), .ZN(
        n13017) );
  OAI21_X1 U12986 ( .B1(n13149), .B2(n13148), .A(n13212), .ZN(n13154) );
  AND4_X1 U12987 ( .A1(n11488), .A2(n11487), .A3(n11486), .A4(n11485), .ZN(
        n11489) );
  AND2_X1 U12988 ( .A1(n12240), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12241) );
  AND2_X1 U12989 ( .A1(n12020), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12034) );
  NAND2_X1 U12990 ( .A1(n13893), .A2(n11671), .ZN(n20237) );
  AND2_X1 U12991 ( .A1(n11247), .A2(n11246), .ZN(n15188) );
  AND2_X1 U12992 ( .A1(n11198), .A2(n11197), .ZN(n13773) );
  AND2_X1 U12993 ( .A1(n12554), .A2(n12553), .ZN(n12597) );
  INV_X1 U12994 ( .A(n12569), .ZN(n12531) );
  AND2_X1 U12995 ( .A1(n11213), .A2(n11212), .ZN(n13833) );
  AND2_X1 U12996 ( .A1(n15425), .A2(n10241), .ZN(n15426) );
  AND2_X1 U12997 ( .A1(n15692), .A2(n11338), .ZN(n15547) );
  OR3_X1 U12998 ( .A1(n13407), .A2(n10961), .A3(n15589), .ZN(n15379) );
  INV_X1 U12999 ( .A(n16543), .ZN(n12352) );
  INV_X1 U13000 ( .A(n18424), .ZN(n13140) );
  OAI21_X1 U13001 ( .B1(n18849), .B2(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n13195), .ZN(n13205) );
  NAND2_X1 U13002 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17805) );
  NAND2_X1 U13003 ( .A1(n16560), .A2(n15859), .ZN(n13301) );
  NOR2_X1 U13004 ( .A1(n13178), .A2(n13182), .ZN(n13184) );
  AND2_X1 U13005 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13112) );
  NOR2_X1 U13006 ( .A1(n13154), .A2(n13153), .ZN(n15845) );
  INV_X1 U13007 ( .A(n13956), .ZN(n13947) );
  INV_X1 U13008 ( .A(n15970), .ZN(n15968) );
  OR2_X1 U13009 ( .A1(n13960), .A2(n20316), .ZN(n13956) );
  AND2_X1 U13010 ( .A1(n15963), .A2(n11824), .ZN(n12178) );
  INV_X1 U13011 ( .A(n12391), .ZN(n12320) );
  NAND2_X1 U13012 ( .A1(n12113), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12157) );
  INV_X1 U13013 ( .A(n14372), .ZN(n14644) );
  NOR2_X1 U13014 ( .A1(n11935), .A2(n11934), .ZN(n11940) );
  INV_X1 U13015 ( .A(n14119), .ZN(n14266) );
  INV_X1 U13016 ( .A(n14800), .ZN(n14807) );
  AND2_X1 U13017 ( .A1(n16165), .A2(n12870), .ZN(n20293) );
  OR2_X1 U13018 ( .A1(n11830), .A2(n13874), .ZN(n20553) );
  OR2_X1 U13019 ( .A1(n20675), .A2(n20749), .ZN(n20633) );
  INV_X1 U13020 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20710) );
  NOR2_X1 U13021 ( .A1(n20637), .A2(n20475), .ZN(n20787) );
  OR3_X1 U13022 ( .A1(n11516), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n20315), 
        .ZN(n20373) );
  OR2_X1 U13023 ( .A1(n16309), .A2(n19259), .ZN(n12706) );
  INV_X1 U13024 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15394) );
  NAND2_X1 U13025 ( .A1(n15427), .A2(n15426), .ZN(n15428) );
  XNOR2_X1 U13026 ( .A(n10960), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16456) );
  OR2_X1 U13027 ( .A1(n15581), .A2(n11324), .ZN(n11336) );
  AND2_X1 U13028 ( .A1(n10925), .A2(n13539), .ZN(n13618) );
  OR3_X1 U13029 ( .A1(n19446), .A2(n19468), .A3(n19926), .ZN(n19451) );
  OR2_X1 U13030 ( .A1(n20074), .A2(n14097), .ZN(n19597) );
  NAND2_X1 U13031 ( .A1(n12352), .A2(n12351), .ZN(n12353) );
  NAND2_X1 U13032 ( .A1(n20084), .A2(n20094), .ZN(n20071) );
  OR3_X1 U13033 ( .A1(n19829), .A2(n19862), .A3(n19926), .ZN(n19834) );
  INV_X1 U13034 ( .A(n19437), .ZN(n19427) );
  INV_X1 U13035 ( .A(n20101), .ZN(n14097) );
  NOR2_X1 U13036 ( .A1(n18838), .A2(n13209), .ZN(n16550) );
  AOI21_X1 U13037 ( .B1(n17801), .B2(n16887), .A(n17048), .ZN(n16840) );
  INV_X1 U13038 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16891) );
  INV_X1 U13039 ( .A(n17092), .ZN(n17082) );
  NOR2_X1 U13040 ( .A1(n14407), .A2(n14406), .ZN(n15848) );
  INV_X1 U13041 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17267) );
  INV_X1 U13042 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17354) );
  NOR2_X1 U13043 ( .A1(n13221), .A2(n18272), .ZN(n17899) );
  INV_X1 U13044 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17927) );
  INV_X1 U13045 ( .A(n18272), .ZN(n17955) );
  NAND2_X1 U13046 ( .A1(n13133), .A2(n13132), .ZN(n13224) );
  NAND2_X1 U13047 ( .A1(n13028), .A2(n10225), .ZN(n13029) );
  NAND2_X1 U13048 ( .A1(n13179), .A2(n13180), .ZN(n18000) );
  INV_X1 U13049 ( .A(n18306), .ZN(n18367) );
  AOI211_X1 U13050 ( .C1(n18845), .C2(n13214), .A(n16550), .B(n15847), .ZN(
        n13220) );
  NOR2_X1 U13051 ( .A1(n13113), .A2(n13112), .ZN(n13114) );
  INV_X1 U13052 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17127) );
  INV_X1 U13053 ( .A(n13355), .ZN(n14483) );
  NAND2_X1 U13054 ( .A1(n13947), .A2(n15906), .ZN(n20175) );
  AND2_X1 U13055 ( .A1(n20144), .A2(n13940), .ZN(n20165) );
  NOR2_X2 U13056 ( .A1(n13956), .A2(n13955), .ZN(n20196) );
  INV_X1 U13057 ( .A(n14479), .ZN(n20372) );
  OAI211_X1 U13058 ( .C1(n11893), .C2(n11892), .A(n11891), .B(n11890), .ZN(
        n14005) );
  OR2_X1 U13059 ( .A1(n14707), .A2(n13823), .ZN(n16059) );
  INV_X1 U13060 ( .A(n14012), .ZN(n14190) );
  OR2_X1 U13061 ( .A1(n14011), .A2(n14010), .ZN(n14187) );
  NAND2_X1 U13062 ( .A1(n12158), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12196) );
  NAND2_X1 U13063 ( .A1(n12078), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12111) );
  NAND2_X1 U13064 ( .A1(n11870), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11879) );
  NAND2_X1 U13065 ( .A1(n11861), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11869) );
  AND2_X1 U13066 ( .A1(n16074), .A2(n12323), .ZN(n20249) );
  AND2_X1 U13067 ( .A1(n12890), .A2(n12889), .ZN(n12891) );
  AND2_X1 U13068 ( .A1(n16205), .A2(n12885), .ZN(n16138) );
  INV_X1 U13069 ( .A(n20293), .ZN(n16188) );
  NOR2_X1 U13070 ( .A1(n16244), .A2(n20279), .ZN(n16222) );
  INV_X1 U13071 ( .A(n20377), .ZN(n20475) );
  INV_X1 U13072 ( .A(n20950), .ZN(n13861) );
  OR2_X1 U13073 ( .A1(n9675), .A2(n20306), .ZN(n20701) );
  INV_X1 U13074 ( .A(n20382), .ZN(n20405) );
  INV_X1 U13075 ( .A(n20409), .ZN(n20433) );
  NOR2_X2 U13076 ( .A1(n20553), .A2(n20749), .ZN(n20543) );
  INV_X1 U13077 ( .A(n20583), .ZN(n20604) );
  INV_X1 U13078 ( .A(n20701), .ZN(n20576) );
  INV_X1 U13079 ( .A(n20633), .ZN(n20661) );
  NAND2_X1 U13080 ( .A1(n9675), .A2(n11838), .ZN(n20778) );
  INV_X1 U13081 ( .A(n20703), .ZN(n20743) );
  NOR2_X2 U13082 ( .A1(n20702), .A2(n20701), .ZN(n20774) );
  INV_X1 U13083 ( .A(n20789), .ZN(n20811) );
  INV_X1 U13084 ( .A(n20733), .ZN(n20851) );
  INV_X1 U13085 ( .A(n20869), .ZN(n20876) );
  INV_X1 U13086 ( .A(n20928), .ZN(n20939) );
  NAND2_X1 U13087 ( .A1(n13464), .A2(n13400), .ZN(n19215) );
  INV_X1 U13088 ( .A(n19215), .ZN(n19199) );
  INV_X1 U13089 ( .A(n19231), .ZN(n19209) );
  INV_X1 U13090 ( .A(n15103), .ZN(n15133) );
  INV_X1 U13091 ( .A(n19151), .ZN(n19167) );
  OR2_X1 U13092 ( .A1(n11048), .A2(n11047), .ZN(n13831) );
  INV_X1 U13093 ( .A(n19254), .ZN(n19260) );
  XNOR2_X1 U13094 ( .A(n13601), .B(n13602), .ZN(n20094) );
  INV_X1 U13095 ( .A(n19293), .ZN(n19320) );
  INV_X1 U13096 ( .A(n19390), .ZN(n13593) );
  INV_X1 U13097 ( .A(n13509), .ZN(n13508) );
  AND2_X1 U13098 ( .A1(n13835), .A2(n13834), .ZN(n16442) );
  INV_X1 U13099 ( .A(n16463), .ZN(n19400) );
  OAI21_X1 U13100 ( .B1(n16306), .B2(n16522), .A(n10214), .ZN(n11347) );
  AND2_X1 U13101 ( .A1(n14209), .A2(n11337), .ZN(n15692) );
  INV_X1 U13102 ( .A(n16490), .ZN(n16530) );
  INV_X1 U13103 ( .A(n16548), .ZN(n13539) );
  OAI21_X1 U13104 ( .B1(n14106), .B2(n14105), .A(n14104), .ZN(n19442) );
  NOR2_X1 U13105 ( .A1(n19700), .A2(n19627), .ZN(n19499) );
  NOR2_X1 U13106 ( .A1(n19597), .A2(n20071), .ZN(n19518) );
  NOR2_X1 U13107 ( .A1(n19627), .A2(n20071), .ZN(n19564) );
  NOR2_X1 U13108 ( .A1(n19597), .A2(n19836), .ZN(n19592) );
  NOR2_X1 U13109 ( .A1(n19627), .A2(n19836), .ZN(n19618) );
  INV_X1 U13110 ( .A(n19693), .ZN(n19673) );
  OAI21_X1 U13111 ( .B1(n19669), .B2(n19668), .A(n19667), .ZN(n19695) );
  INV_X1 U13112 ( .A(n19726), .ZN(n19722) );
  NOR2_X1 U13113 ( .A1(n19837), .A2(n19700), .ZN(n19761) );
  AND2_X1 U13114 ( .A1(n19774), .A2(n19770), .ZN(n19794) );
  NOR2_X1 U13115 ( .A1(n19859), .A2(n19836), .ZN(n19855) );
  INV_X1 U13116 ( .A(n19965), .ZN(n19898) );
  INV_X1 U13117 ( .A(n19917), .ZN(n19910) );
  INV_X1 U13118 ( .A(n19902), .ZN(n19966) );
  INV_X1 U13119 ( .A(n13142), .ZN(n13136) );
  NOR2_X1 U13120 ( .A1(n17065), .A2(n16908), .ZN(n16885) );
  OR2_X1 U13121 ( .A1(n16908), .A2(n17029), .ZN(n16915) );
  INV_X1 U13122 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17055) );
  INV_X1 U13123 ( .A(n17094), .ZN(n17029) );
  INV_X1 U13124 ( .A(n17050), .ZN(n17076) );
  NOR2_X1 U13125 ( .A1(n16836), .A2(n17201), .ZN(n17170) );
  NOR2_X1 U13126 ( .A1(n14412), .A2(n15836), .ZN(n17297) );
  NOR2_X1 U13127 ( .A1(n17026), .A2(n17415), .ZN(n17408) );
  INV_X1 U13128 ( .A(n17435), .ZN(n17263) );
  INV_X1 U13129 ( .A(n17456), .ZN(n17453) );
  NOR3_X1 U13130 ( .A1(n18449), .A2(n17662), .A3(n17519), .ZN(n17507) );
  INV_X1 U13131 ( .A(n17510), .ZN(n17517) );
  NOR2_X1 U13132 ( .A1(n18092), .A2(n13185), .ZN(n13298) );
  OR2_X1 U13133 ( .A1(n17722), .A2(n17721), .ZN(n17723) );
  INV_X1 U13134 ( .A(n17899), .ZN(n18218) );
  OAI21_X1 U13135 ( .B1(n18093), .B2(n17732), .A(n17716), .ZN(n13232) );
  NOR2_X1 U13136 ( .A1(n18136), .A2(n18386), .ZN(n18142) );
  INV_X1 U13137 ( .A(n18401), .ZN(n18384) );
  INV_X1 U13138 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19056) );
  INV_X1 U13139 ( .A(n18523), .ZN(n18584) );
  INV_X1 U13140 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19059) );
  INV_X1 U13141 ( .A(n20980), .ZN(n20979) );
  INV_X1 U13142 ( .A(n20186), .ZN(n20141) );
  INV_X1 U13143 ( .A(n20196), .ZN(n20162) );
  OR3_X1 U13144 ( .A1(n20175), .A2(n20134), .A3(n14569), .ZN(n16053) );
  INV_X1 U13145 ( .A(n20198), .ZN(n14024) );
  NAND2_X1 U13146 ( .A1(n14496), .A2(n14001), .ZN(n13370) );
  INV_X1 U13147 ( .A(n14001), .ZN(n14640) );
  NAND2_X1 U13148 ( .A1(n14633), .A2(n14479), .ZN(n14655) );
  INV_X1 U13149 ( .A(n20201), .ZN(n20233) );
  AOI21_X1 U13150 ( .B1(n20249), .B2(n14435), .A(n13312), .ZN(n13313) );
  OR2_X1 U13151 ( .A1(n20250), .A2(n12322), .ZN(n16074) );
  INV_X1 U13152 ( .A(n20249), .ZN(n20243) );
  AND2_X1 U13153 ( .A1(n12892), .A2(n12891), .ZN(n12893) );
  AOI21_X1 U13154 ( .B1(n12882), .B2(n20276), .A(n16222), .ZN(n16273) );
  INV_X1 U13155 ( .A(n20292), .ZN(n20288) );
  INV_X1 U13156 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20303) );
  INV_X1 U13157 ( .A(n20953), .ZN(n20955) );
  OR2_X1 U13158 ( .A1(n20448), .A2(n20749), .ZN(n20409) );
  AOI22_X1 U13159 ( .A1(n20412), .A2(n20416), .B1(n10210), .B2(n20637), .ZN(
        n20437) );
  NAND2_X1 U13160 ( .A1(n20549), .A2(n20576), .ZN(n20520) );
  AOI22_X1 U13161 ( .A1(n20526), .A2(n20523), .B1(n10210), .B2(n20709), .ZN(
        n20547) );
  NAND2_X1 U13162 ( .A1(n20549), .A2(n20548), .ZN(n20583) );
  NAND2_X1 U13163 ( .A1(n20577), .A2(n20576), .ZN(n20632) );
  AOI22_X1 U13164 ( .A1(n20643), .A2(n20639), .B1(n20637), .B2(n20636), .ZN(
        n20665) );
  OR2_X1 U13165 ( .A1(n20675), .A2(n20778), .ZN(n20700) );
  AOI22_X1 U13166 ( .A1(n20715), .A2(n20712), .B1(n20709), .B2(n20708), .ZN(
        n20748) );
  NAND2_X1 U13167 ( .A1(n20824), .A2(n20750), .ZN(n20789) );
  NAND2_X1 U13168 ( .A1(n20824), .A2(n20548), .ZN(n20869) );
  INV_X1 U13169 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20971) );
  INV_X1 U13170 ( .A(n20945), .ZN(n20980) );
  OR2_X1 U13171 ( .A1(n13472), .A2(n13394), .ZN(n13509) );
  INV_X1 U13172 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n14091) );
  INV_X1 U13173 ( .A(n19189), .ZN(n19216) );
  INV_X1 U13174 ( .A(n19183), .ZN(n19218) );
  NAND2_X1 U13175 ( .A1(n15722), .A2(n13610), .ZN(n20101) );
  AND2_X1 U13176 ( .A1(n13263), .A2(n13539), .ZN(n19293) );
  INV_X1 U13177 ( .A(n19295), .ZN(n19329) );
  INV_X1 U13178 ( .A(n19331), .ZN(n19358) );
  NAND2_X1 U13179 ( .A1(n13508), .A2(n9666), .ZN(n19390) );
  INV_X1 U13180 ( .A(n19388), .ZN(n13599) );
  NAND2_X1 U13181 ( .A1(n12343), .A2(n9676), .ZN(n16465) );
  INV_X1 U13182 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16409) );
  INV_X1 U13183 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16445) );
  NAND2_X1 U13184 ( .A1(n13473), .A2(n12344), .ZN(n19394) );
  NAND2_X1 U13185 ( .A1(n10971), .A2(n9666), .ZN(n16527) );
  INV_X1 U13186 ( .A(n16525), .ZN(n15710) );
  INV_X1 U13187 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20098) );
  INV_X1 U13188 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13490) );
  INV_X1 U13189 ( .A(n19443), .ZN(n19435) );
  INV_X1 U13190 ( .A(n19465), .ZN(n19473) );
  INV_X1 U13191 ( .A(n19499), .ZN(n19492) );
  INV_X1 U13192 ( .A(n19518), .ZN(n19534) );
  INV_X1 U13193 ( .A(n19592), .ZN(n19589) );
  INV_X1 U13194 ( .A(n19618), .ZN(n19626) );
  INV_X1 U13195 ( .A(n19649), .ZN(n19659) );
  NAND2_X1 U13196 ( .A1(n19629), .A2(n19628), .ZN(n19693) );
  OR2_X1 U13197 ( .A1(n19859), .A2(n19700), .ZN(n19726) );
  INV_X1 U13198 ( .A(n19761), .ZN(n19758) );
  INV_X1 U13199 ( .A(n19795), .ZN(n19790) );
  INV_X1 U13200 ( .A(n19825), .ZN(n19818) );
  INV_X1 U13201 ( .A(n19855), .ZN(n19851) );
  OR2_X1 U13202 ( .A1(n19837), .A2(n19836), .ZN(n19917) );
  AND2_X1 U13203 ( .A1(n19868), .A2(n19867), .ZN(n19905) );
  OR2_X1 U13204 ( .A1(n19859), .A2(n19931), .ZN(n19978) );
  INV_X1 U13205 ( .A(n20068), .ZN(n19991) );
  NAND2_X1 U13206 ( .A1(n19073), .A2(n18411), .ZN(n19071) );
  INV_X1 U13207 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17897) );
  NAND2_X1 U13208 ( .A1(n17094), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n17050) );
  NOR2_X1 U13209 ( .A1(n17099), .A2(n17153), .ZN(n17158) );
  AND2_X1 U13210 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17202), .ZN(n17216) );
  NOR2_X1 U13211 ( .A1(n16960), .A2(n17370), .ZN(n17351) );
  NOR2_X2 U13212 ( .A1(n17263), .A2(n17527), .ZN(n17432) );
  INV_X1 U13213 ( .A(n17516), .ZN(n17504) );
  NOR2_X1 U13214 ( .A1(n17528), .A2(n17550), .ZN(n17553) );
  NOR2_X1 U13215 ( .A1(n17558), .A2(n17589), .ZN(n17584) );
  NAND2_X1 U13216 ( .A1(n17624), .A2(n18411), .ZN(n17622) );
  INV_X1 U13217 ( .A(n17624), .ZN(n17654) );
  AOI21_X1 U13218 ( .B1(n13233), .B2(n18315), .A(n13232), .ZN(n13234) );
  INV_X1 U13219 ( .A(n18394), .ZN(n18386) );
  NAND2_X1 U13220 ( .A1(n16559), .A2(n18384), .ZN(n18302) );
  INV_X1 U13221 ( .A(n17995), .ZN(n18320) );
  INV_X1 U13222 ( .A(n18397), .ZN(n18391) );
  INV_X1 U13223 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18414) );
  INV_X1 U13224 ( .A(n19054), .ZN(n18904) );
  INV_X1 U13225 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19008) );
  INV_X1 U13226 ( .A(n19005), .ZN(n18918) );
  INV_X1 U13227 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18931) );
  NAND2_X1 U13228 ( .A1(n13370), .A2(n13369), .ZN(P1_U2842) );
  OAI211_X1 U13229 ( .C1(n20115), .C2(n13314), .A(n10219), .B(n13313), .ZN(
        P1_U2971) );
  OAI21_X1 U13230 ( .B1(n13314), .B2(n16225), .A(n12893), .ZN(P1_U3003) );
  OAI21_X1 U13231 ( .B1(n13238), .B2(n10213), .A(n10245), .ZN(P2_U2858) );
  NAND2_X1 U13232 ( .A1(n13235), .A2(n13234), .ZN(P3_U2834) );
  AND2_X4 U13233 ( .A1(n10872), .A2(n14069), .ZN(n12587) );
  AOI22_X1 U13234 ( .A1(n13249), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10256) );
  AOI22_X1 U13235 ( .A1(n10284), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10255) );
  AOI22_X1 U13236 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9660), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10254) );
  AOI22_X1 U13237 ( .A1(n9683), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10253) );
  NAND4_X1 U13238 ( .A1(n10256), .A2(n10255), .A3(n10254), .A4(n10253), .ZN(
        n10257) );
  NAND2_X1 U13239 ( .A1(n10257), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10264) );
  AOI22_X1 U13240 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10261) );
  AOI22_X1 U13241 ( .A1(n10284), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10260) );
  AOI22_X1 U13242 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(n9660), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10259) );
  AOI22_X1 U13243 ( .A1(n9681), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10258) );
  NAND4_X1 U13244 ( .A1(n10261), .A2(n10260), .A3(n10259), .A4(n10258), .ZN(
        n10262) );
  NAND2_X1 U13245 ( .A1(n10262), .A2(n14045), .ZN(n10263) );
  AOI22_X1 U13246 ( .A1(n10284), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10268) );
  AOI22_X1 U13247 ( .A1(n9664), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10267) );
  AOI22_X1 U13248 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9660), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10266) );
  AOI22_X1 U13249 ( .A1(n9682), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10265) );
  NAND4_X1 U13250 ( .A1(n10268), .A2(n10267), .A3(n10266), .A4(n10265), .ZN(
        n10269) );
  NAND2_X1 U13251 ( .A1(n10269), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10276) );
  AOI22_X1 U13252 ( .A1(n13249), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10272) );
  AOI22_X1 U13253 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(n9660), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10271) );
  AOI22_X1 U13254 ( .A1(n9684), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10270) );
  NAND4_X1 U13255 ( .A1(n10273), .A2(n10272), .A3(n10271), .A4(n10270), .ZN(
        n10274) );
  NAND2_X1 U13256 ( .A1(n10274), .A2(n14045), .ZN(n10275) );
  AOI22_X1 U13257 ( .A1(n13249), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10281) );
  AOI22_X1 U13258 ( .A1(n9680), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(n9660), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10280) );
  NAND2_X1 U13259 ( .A1(n10485), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10277) );
  NAND4_X1 U13260 ( .A1(n10282), .A2(n10281), .A3(n10280), .A4(n10279), .ZN(
        n10283) );
  AOI22_X1 U13261 ( .A1(n9680), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10288) );
  AOI22_X1 U13262 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n9660), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10287) );
  NAND4_X1 U13263 ( .A1(n10288), .A2(n10287), .A3(n10286), .A4(n10285), .ZN(
        n10289) );
  NAND2_X1 U13264 ( .A1(n10289), .A2(n14045), .ZN(n10290) );
  AOI22_X1 U13265 ( .A1(n10284), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10293) );
  AOI22_X1 U13266 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9660), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10292) );
  NAND2_X1 U13267 ( .A1(n10293), .A2(n10292), .ZN(n10297) );
  AOI22_X1 U13268 ( .A1(n9683), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10295) );
  AOI22_X1 U13269 ( .A1(n9664), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10294) );
  NAND2_X1 U13270 ( .A1(n10295), .A2(n10294), .ZN(n10296) );
  OAI21_X1 U13271 ( .B1(n10297), .B2(n10296), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10305) );
  AOI22_X1 U13272 ( .A1(n10284), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10299) );
  AOI22_X1 U13273 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(n9660), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10298) );
  NAND2_X1 U13274 ( .A1(n10299), .A2(n10298), .ZN(n10303) );
  AOI22_X1 U13275 ( .A1(n13249), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10301) );
  AOI22_X1 U13276 ( .A1(n9683), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10300) );
  NAND2_X1 U13277 ( .A1(n10301), .A2(n10300), .ZN(n10302) );
  OAI21_X1 U13278 ( .B1(n10303), .B2(n10302), .A(n14045), .ZN(n10304) );
  AOI22_X1 U13279 ( .A1(n10284), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10309) );
  AOI22_X1 U13280 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9660), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10308) );
  AOI22_X1 U13281 ( .A1(n9664), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10307) );
  AOI22_X1 U13282 ( .A1(n9682), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10306) );
  NAND4_X1 U13283 ( .A1(n10309), .A2(n10308), .A3(n10307), .A4(n10306), .ZN(
        n10310) );
  AOI22_X1 U13284 ( .A1(n10284), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10314) );
  AOI22_X1 U13285 ( .A1(n13249), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10313) );
  AOI22_X1 U13286 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(n9660), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10312) );
  AOI22_X1 U13287 ( .A1(n9684), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10311) );
  NAND4_X1 U13288 ( .A1(n10314), .A2(n10313), .A3(n10312), .A4(n10311), .ZN(
        n10315) );
  AOI22_X1 U13289 ( .A1(n10284), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10319) );
  AOI22_X1 U13290 ( .A1(n13249), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10318) );
  AOI22_X1 U13291 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9660), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10317) );
  AOI22_X1 U13292 ( .A1(n9682), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10316) );
  NAND4_X1 U13293 ( .A1(n10319), .A2(n10318), .A3(n10317), .A4(n10316), .ZN(
        n10320) );
  NAND2_X1 U13294 ( .A1(n10320), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10328) );
  AOI22_X1 U13295 ( .A1(n10284), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10325) );
  AOI22_X1 U13296 ( .A1(n9663), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10324) );
  AOI22_X1 U13297 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n9660), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10323) );
  AOI22_X1 U13298 ( .A1(n9684), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10322) );
  NAND4_X1 U13299 ( .A1(n10325), .A2(n10324), .A3(n10323), .A4(n10322), .ZN(
        n10326) );
  NAND2_X1 U13300 ( .A1(n10326), .A2(n14045), .ZN(n10327) );
  NAND2_X2 U13301 ( .A1(n10328), .A2(n10327), .ZN(n10354) );
  AOI22_X1 U13302 ( .A1(n10284), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10332) );
  AOI22_X1 U13303 ( .A1(n13249), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10331) );
  AOI22_X1 U13304 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9660), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10330) );
  AOI22_X1 U13305 ( .A1(n9681), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10329) );
  NAND4_X1 U13306 ( .A1(n10332), .A2(n10331), .A3(n10330), .A4(n10329), .ZN(
        n10333) );
  AOI22_X1 U13307 ( .A1(n10284), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10337) );
  AOI22_X1 U13308 ( .A1(n13249), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U13309 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(n9660), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10335) );
  AOI22_X1 U13310 ( .A1(n9680), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10334) );
  NAND4_X1 U13311 ( .A1(n10337), .A2(n10336), .A3(n10335), .A4(n10334), .ZN(
        n10338) );
  NAND2_X1 U13312 ( .A1(n10338), .A2(n14045), .ZN(n10339) );
  NAND2_X1 U13313 ( .A1(n10380), .A2(n10353), .ZN(n10888) );
  AND2_X2 U13314 ( .A1(n13392), .A2(n10888), .ZN(n11178) );
  INV_X2 U13315 ( .A(n12336), .ZN(n10353) );
  AOI22_X1 U13316 ( .A1(n13249), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10344) );
  AOI22_X1 U13317 ( .A1(n10284), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10343) );
  AOI22_X1 U13318 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9660), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10342) );
  AOI22_X1 U13319 ( .A1(n9684), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10341) );
  NAND4_X1 U13320 ( .A1(n10344), .A2(n10343), .A3(n10342), .A4(n10341), .ZN(
        n10345) );
  NAND2_X1 U13321 ( .A1(n10345), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10352) );
  AOI22_X1 U13322 ( .A1(n9664), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10349) );
  AOI22_X1 U13323 ( .A1(n10284), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10348) );
  AOI22_X1 U13324 ( .A1(n9682), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(n9660), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10347) );
  AOI22_X1 U13325 ( .A1(n9652), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10346) );
  NAND4_X1 U13326 ( .A1(n10349), .A2(n10348), .A3(n10347), .A4(n10346), .ZN(
        n10350) );
  NAND2_X1 U13327 ( .A1(n10350), .A2(n14045), .ZN(n10351) );
  NAND2_X2 U13328 ( .A1(n11178), .A2(n10355), .ZN(n10393) );
  NAND2_X1 U13329 ( .A1(n10393), .A2(n9666), .ZN(n10365) );
  NOR2_X1 U13330 ( .A1(n10375), .A2(n12336), .ZN(n10359) );
  AND2_X2 U13331 ( .A1(n10357), .A2(n10578), .ZN(n10979) );
  INV_X1 U13332 ( .A(n10979), .ZN(n10358) );
  NAND2_X1 U13333 ( .A1(n10358), .A2(n9860), .ZN(n10379) );
  OAI21_X1 U13334 ( .B1(n10359), .B2(n9860), .A(n10379), .ZN(n10360) );
  INV_X1 U13335 ( .A(n10360), .ZN(n10364) );
  INV_X1 U13336 ( .A(n10384), .ZN(n10983) );
  NAND2_X1 U13337 ( .A1(n11281), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10372) );
  INV_X1 U13338 ( .A(n11314), .ZN(n10368) );
  AOI22_X1 U13339 ( .A1(n10415), .A2(P2_EBX_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10371) );
  NAND2_X1 U13340 ( .A1(n10379), .A2(n10215), .ZN(n10381) );
  INV_X1 U13341 ( .A(n10380), .ZN(n13488) );
  NAND2_X1 U13342 ( .A1(n10381), .A2(n13488), .ZN(n10383) );
  MUX2_X1 U13343 ( .A(n13764), .B(n13279), .S(n10361), .Z(n10382) );
  NAND2_X1 U13344 ( .A1(n10383), .A2(n10382), .ZN(n11304) );
  NAND2_X1 U13345 ( .A1(n11310), .A2(n11318), .ZN(n10401) );
  NOR2_X1 U13346 ( .A1(n12336), .A2(n14091), .ZN(n14901) );
  INV_X1 U13347 ( .A(n10385), .ZN(n10388) );
  NAND3_X1 U13348 ( .A1(n10863), .A2(n19411), .A3(n10983), .ZN(n10390) );
  INV_X1 U13349 ( .A(n10389), .ZN(n10880) );
  NAND2_X1 U13350 ( .A1(n11179), .A2(n14899), .ZN(n10391) );
  AND2_X2 U13351 ( .A1(n10392), .A2(n10391), .ZN(n10396) );
  NAND2_X1 U13352 ( .A1(n10420), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10395) );
  NOR2_X1 U13353 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n14093) );
  AOI22_X1 U13354 ( .A1(n10393), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n14093), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10394) );
  INV_X1 U13355 ( .A(n14093), .ZN(n10405) );
  NAND2_X1 U13356 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10397) );
  NAND2_X1 U13357 ( .A1(n10405), .A2(n10397), .ZN(n10398) );
  AOI21_X1 U13358 ( .B1(n10415), .B2(P2_EBX_REG_0__SCAN_IN), .A(n10398), .ZN(
        n10399) );
  INV_X1 U13359 ( .A(n10400), .ZN(n10402) );
  NAND2_X1 U13360 ( .A1(n10420), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10409) );
  INV_X1 U13361 ( .A(n13752), .ZN(n10407) );
  OAI21_X1 U13362 ( .B1(n10405), .B2(n20106), .A(n10427), .ZN(n10406) );
  INV_X1 U13363 ( .A(n10410), .ZN(n10412) );
  NAND2_X1 U13364 ( .A1(n10412), .A2(n10411), .ZN(n10413) );
  INV_X1 U13365 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14458) );
  NAND2_X1 U13366 ( .A1(n9657), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10417) );
  AOI22_X1 U13367 ( .A1(n10415), .A2(P2_EBX_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10416) );
  NAND2_X2 U13368 ( .A1(n10419), .A2(n10418), .ZN(n10434) );
  NAND2_X1 U13369 ( .A1(n10420), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10422) );
  AOI21_X1 U13370 ( .B1(n14091), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10421) );
  NAND2_X1 U13371 ( .A1(n10434), .A2(n10433), .ZN(n10423) );
  INV_X1 U13372 ( .A(n10434), .ZN(n10425) );
  INV_X1 U13373 ( .A(n10433), .ZN(n10424) );
  NAND2_X1 U13374 ( .A1(n10425), .A2(n10424), .ZN(n10426) );
  INV_X1 U13375 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16534) );
  NAND2_X1 U13376 ( .A1(n9657), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10428) );
  NAND2_X1 U13377 ( .A1(n10420), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10430) );
  NAND2_X1 U13378 ( .A1(n14093), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10429) );
  XNOR2_X2 U13379 ( .A(n10436), .B(n10435), .ZN(n12408) );
  INV_X1 U13380 ( .A(n12408), .ZN(n13653) );
  INV_X1 U13382 ( .A(n10438), .ZN(n10444) );
  XNOR2_X2 U13383 ( .A(n10444), .B(n10440), .ZN(n14068) );
  NAND2_X1 U13384 ( .A1(n10637), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10454) );
  OR2_X1 U13385 ( .A1(n10444), .A2(n15709), .ZN(n10455) );
  AND2_X1 U13386 ( .A1(n15129), .A2(n10442), .ZN(n10441) );
  AND2_X1 U13387 ( .A1(n13653), .A2(n10442), .ZN(n10443) );
  AOI22_X1 U13388 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10648), .B1(
        n9708), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10453) );
  INV_X1 U13389 ( .A(n15709), .ZN(n10445) );
  AND2_X1 U13390 ( .A1(n10445), .A2(n10444), .ZN(n10448) );
  AND2_X1 U13391 ( .A1(n13653), .A2(n10448), .ZN(n10446) );
  AND2_X1 U13392 ( .A1(n12408), .A2(n10448), .ZN(n10447) );
  AOI22_X1 U13393 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10649), .B1(
        n19446), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10452) );
  INV_X1 U13394 ( .A(n10448), .ZN(n10449) );
  NOR2_X1 U13395 ( .A1(n10459), .A2(n10449), .ZN(n10450) );
  AOI22_X1 U13396 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19704), .B1(
        n19829), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10451) );
  INV_X1 U13397 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12485) );
  INV_X1 U13398 ( .A(n10456), .ZN(n10457) );
  INV_X1 U13399 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12482) );
  INV_X1 U13400 ( .A(n10458), .ZN(n10469) );
  NAND2_X1 U13401 ( .A1(n19800), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10468) );
  AND2_X1 U13402 ( .A1(n12408), .A2(n14068), .ZN(n10463) );
  INV_X1 U13403 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14118) );
  NAND2_X1 U13404 ( .A1(n10464), .A2(n10463), .ZN(n10682) );
  INV_X1 U13405 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12481) );
  OAI22_X1 U13406 ( .A1(n10641), .A2(n14118), .B1(n10682), .B2(n12481), .ZN(
        n10465) );
  INV_X1 U13407 ( .A(n10465), .ZN(n10466) );
  INV_X1 U13408 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10471) );
  INV_X1 U13409 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10475) );
  NOR2_X1 U13410 ( .A1(n10477), .A2(n10476), .ZN(n10478) );
  NAND3_X1 U13411 ( .A1(n10480), .A2(n10479), .A3(n10478), .ZN(n10501) );
  AND2_X1 U13412 ( .A1(n9663), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10519) );
  NAND2_X1 U13413 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10483) );
  BUF_X1 U13414 ( .A(n10284), .Z(n10481) );
  NAND2_X1 U13415 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10482) );
  AND2_X1 U13416 ( .A1(n10483), .A2(n10482), .ZN(n10489) );
  AOI22_X1 U13417 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10612), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10488) );
  AND2_X2 U13418 ( .A1(n10485), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10542) );
  AOI22_X1 U13419 ( .A1(n12562), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10487) );
  AND2_X2 U13420 ( .A1(n12587), .A2(n14045), .ZN(n10562) );
  AOI22_X1 U13421 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10562), .B1(
        n12555), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10486) );
  NAND4_X1 U13422 ( .A1(n10489), .A2(n10488), .A3(n10487), .A4(n10486), .ZN(
        n10499) );
  AND2_X2 U13423 ( .A1(n12686), .A2(n14045), .ZN(n12557) );
  AOI22_X1 U13424 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12557), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10497) );
  AND2_X2 U13425 ( .A1(n12686), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12568) );
  AOI22_X1 U13426 ( .A1(n12563), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12568), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10496) );
  INV_X1 U13427 ( .A(n10534), .ZN(n10570) );
  AND2_X2 U13428 ( .A1(n13747), .A2(n10491), .ZN(n12565) );
  INV_X1 U13429 ( .A(n10491), .ZN(n12539) );
  AOI22_X1 U13430 ( .A1(n12565), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n11088), .ZN(n10493) );
  AND2_X1 U13431 ( .A1(n9677), .A2(n10491), .ZN(n10547) );
  NAND2_X1 U13432 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n10492) );
  OAI211_X1 U13433 ( .C1(n10570), .C2(n12482), .A(n10493), .B(n10492), .ZN(
        n10494) );
  INV_X1 U13434 ( .A(n10494), .ZN(n10495) );
  NAND3_X1 U13435 ( .A1(n10497), .A2(n10496), .A3(n10495), .ZN(n10498) );
  NOR2_X1 U13436 ( .A1(n10499), .A2(n10498), .ZN(n11002) );
  NAND2_X1 U13437 ( .A1(n11002), .A2(n9666), .ZN(n10500) );
  NAND2_X1 U13438 ( .A1(n10501), .A2(n10500), .ZN(n10559) );
  INV_X1 U13439 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11041) );
  INV_X1 U13440 ( .A(n19704), .ZN(n19701) );
  INV_X1 U13441 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12453) );
  OAI22_X1 U13442 ( .A1(n11041), .A2(n19701), .B1(n19924), .B2(n12453), .ZN(
        n10510) );
  NAND2_X1 U13443 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10505) );
  INV_X1 U13444 ( .A(n19479), .ZN(n10502) );
  NAND2_X1 U13445 ( .A1(n10502), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10503) );
  NAND3_X1 U13446 ( .A1(n10505), .A2(n10504), .A3(n10503), .ZN(n10509) );
  INV_X1 U13447 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12455) );
  NAND2_X1 U13448 ( .A1(n19446), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10506) );
  OAI211_X1 U13449 ( .C1(n10650), .C2(n12455), .A(n10507), .B(n10506), .ZN(
        n10508) );
  INV_X1 U13450 ( .A(n19863), .ZN(n10511) );
  INV_X1 U13451 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14114) );
  INV_X1 U13452 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12451) );
  OAI22_X1 U13453 ( .A1(n14114), .A2(n10641), .B1(n10682), .B2(n12451), .ZN(
        n10515) );
  INV_X1 U13454 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10513) );
  INV_X1 U13455 ( .A(n19829), .ZN(n10512) );
  INV_X1 U13456 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12454) );
  OAI22_X1 U13457 ( .A1(n10513), .A2(n19663), .B1(n10512), .B2(n12454), .ZN(
        n10514) );
  NOR2_X1 U13458 ( .A1(n10515), .A2(n10514), .ZN(n10517) );
  INV_X1 U13459 ( .A(n19603), .ZN(n10516) );
  AOI22_X1 U13460 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n10562), .B1(
        n12568), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10523) );
  AOI22_X1 U13461 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12569), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10522) );
  AOI22_X1 U13462 ( .A1(n12563), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10521) );
  AOI22_X1 U13463 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10612), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10520) );
  NAND4_X1 U13464 ( .A1(n10523), .A2(n10522), .A3(n10521), .A4(n10520), .ZN(
        n10529) );
  AOI22_X1 U13465 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__0__SCAN_IN), .B2(n12564), .ZN(n10527) );
  AOI22_X1 U13466 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12565), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10526) );
  AOI22_X1 U13467 ( .A1(n12562), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10534), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10525) );
  AOI22_X1 U13468 ( .A1(n12555), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12557), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10524) );
  NAND4_X1 U13469 ( .A1(n10527), .A2(n10526), .A3(n10525), .A4(n10524), .ZN(
        n10528) );
  AOI22_X1 U13470 ( .A1(n12555), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12568), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10533) );
  AOI22_X1 U13471 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12562), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10532) );
  AOI22_X1 U13472 ( .A1(n12563), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10612), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10531) );
  AOI22_X1 U13473 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10530) );
  NAND4_X1 U13474 ( .A1(n10533), .A2(n10532), .A3(n10531), .A4(n10530), .ZN(
        n10540) );
  AOI22_X1 U13475 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n12565), .ZN(n10538) );
  AOI22_X1 U13476 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n11088), .ZN(n10537) );
  AOI22_X1 U13477 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10542), .B1(
        n12557), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U13478 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10534), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10535) );
  NAND4_X1 U13479 ( .A1(n10538), .A2(n10537), .A3(n10536), .A4(n10535), .ZN(
        n10539) );
  NOR2_X1 U13480 ( .A1(n13496), .A2(n10989), .ZN(n10541) );
  NAND2_X1 U13481 ( .A1(n9666), .A2(n10541), .ZN(n10930) );
  AOI22_X1 U13482 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10546) );
  AOI22_X1 U13483 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10534), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10545) );
  AOI22_X1 U13484 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10612), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10544) );
  AOI22_X1 U13485 ( .A1(n12562), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10542), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10543) );
  NAND4_X1 U13486 ( .A1(n10546), .A2(n10545), .A3(n10544), .A4(n10543), .ZN(
        n10556) );
  AOI22_X1 U13487 ( .A1(n12563), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12557), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10554) );
  AOI22_X1 U13488 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12568), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10553) );
  INV_X1 U13489 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10550) );
  AOI22_X1 U13490 ( .A1(n12565), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n11088), .ZN(n10549) );
  NAND2_X1 U13491 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n10548) );
  OAI211_X1 U13492 ( .C1(n13749), .C2(n10550), .A(n10549), .B(n10548), .ZN(
        n10551) );
  INV_X1 U13493 ( .A(n10551), .ZN(n10552) );
  NAND3_X1 U13494 ( .A1(n10554), .A2(n10553), .A3(n10552), .ZN(n10555) );
  INV_X1 U13495 ( .A(n10993), .ZN(n10929) );
  NAND2_X1 U13496 ( .A1(n10930), .A2(n10929), .ZN(n10557) );
  NAND2_X1 U13497 ( .A1(n10560), .A2(n10559), .ZN(n10561) );
  NAND2_X1 U13498 ( .A1(n10935), .A2(n10561), .ZN(n10926) );
  AOI22_X1 U13499 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10566) );
  AOI22_X1 U13500 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12555), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10565) );
  AOI22_X1 U13501 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10612), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10564) );
  AOI22_X1 U13502 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n10542), .B1(
        n12557), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10563) );
  NAND4_X1 U13503 ( .A1(n10566), .A2(n10565), .A3(n10564), .A4(n10563), .ZN(
        n10577) );
  AOI22_X1 U13504 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12568), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10575) );
  INV_X1 U13505 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10569) );
  AOI22_X1 U13506 ( .A1(n12565), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n11088), .ZN(n10568) );
  NAND2_X1 U13507 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10567) );
  OAI211_X1 U13508 ( .C1(n10570), .C2(n10569), .A(n10568), .B(n10567), .ZN(
        n10571) );
  INV_X1 U13509 ( .A(n10571), .ZN(n10574) );
  NAND2_X1 U13510 ( .A1(n12563), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10573) );
  NAND2_X1 U13511 ( .A1(n12562), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10572) );
  NAND4_X1 U13512 ( .A1(n10575), .A2(n10574), .A3(n10573), .A4(n10572), .ZN(
        n10576) );
  OR2_X2 U13513 ( .A1(n10577), .A2(n10576), .ZN(n11014) );
  OR2_X1 U13514 ( .A1(n10989), .A2(n19422), .ZN(n10580) );
  NOR2_X1 U13515 ( .A1(n10974), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10597) );
  INV_X1 U13516 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n14258) );
  NAND2_X1 U13517 ( .A1(n10597), .A2(n14258), .ZN(n10579) );
  NAND2_X1 U13518 ( .A1(n10580), .A2(n10579), .ZN(n10604) );
  INV_X1 U13519 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n15123) );
  NAND2_X1 U13520 ( .A1(n13414), .A2(n10993), .ZN(n10584) );
  MUX2_X1 U13521 ( .A(n20098), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n10868) );
  NAND2_X1 U13522 ( .A1(n10868), .A2(n10867), .ZN(n10582) );
  NAND2_X1 U13523 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20098), .ZN(
        n10581) );
  XNOR2_X1 U13524 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10583) );
  XNOR2_X1 U13525 ( .A(n10585), .B(n10583), .ZN(n10905) );
  INV_X1 U13526 ( .A(n10905), .ZN(n10895) );
  NAND2_X1 U13527 ( .A1(n10591), .A2(n10895), .ZN(n10906) );
  NAND2_X1 U13528 ( .A1(n10584), .A2(n10906), .ZN(n10858) );
  MUX2_X1 U13529 ( .A(n15123), .B(n10858), .S(n10974), .Z(n10603) );
  INV_X1 U13530 ( .A(n10585), .ZN(n10587) );
  NAND2_X1 U13531 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20088), .ZN(
        n10586) );
  NAND2_X1 U13532 ( .A1(n10587), .A2(n10586), .ZN(n10590) );
  NAND2_X1 U13533 ( .A1(n10588), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10589) );
  MUX2_X1 U13534 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n20081), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10609) );
  XNOR2_X1 U13535 ( .A(n10610), .B(n10609), .ZN(n10864) );
  MUX2_X1 U13536 ( .A(n11002), .B(n10864), .S(n10591), .Z(n10856) );
  NOR2_X2 U13537 ( .A1(n10602), .A2(n10594), .ZN(n10628) );
  INV_X1 U13538 ( .A(n10628), .ZN(n10631) );
  NAND2_X1 U13539 ( .A1(n10602), .A2(n10594), .ZN(n10595) );
  NAND2_X1 U13540 ( .A1(n10631), .A2(n10595), .ZN(n15111) );
  OAI21_X1 U13541 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20106), .A(
        n10596), .ZN(n10901) );
  MUX2_X1 U13542 ( .A(n10901), .B(n13496), .S(n13414), .Z(n10598) );
  AOI21_X1 U13543 ( .B1(n10598), .B2(n10974), .A(n10597), .ZN(n14289) );
  NAND2_X1 U13544 ( .A1(n14289), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13546) );
  INV_X1 U13545 ( .A(n10604), .ZN(n10600) );
  NAND3_X1 U13546 ( .A1(n19422), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n10599) );
  NAND2_X1 U13547 ( .A1(n10600), .A2(n10599), .ZN(n14255) );
  NOR2_X1 U13548 ( .A1(n13546), .A2(n14255), .ZN(n10601) );
  NAND2_X1 U13549 ( .A1(n13546), .A2(n14255), .ZN(n13545) );
  OAI21_X1 U13550 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10601), .A(
        n13545), .ZN(n13648) );
  OAI21_X1 U13551 ( .B1(n10604), .B2(n10603), .A(n10602), .ZN(n10605) );
  XNOR2_X1 U13552 ( .A(n10605), .B(n14458), .ZN(n13647) );
  OR2_X1 U13553 ( .A1(n13648), .A2(n13647), .ZN(n13650) );
  INV_X1 U13554 ( .A(n10605), .ZN(n15125) );
  NAND2_X1 U13555 ( .A1(n15125), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10606) );
  NAND2_X1 U13556 ( .A1(n13650), .A2(n10606), .ZN(n16476) );
  INV_X1 U13557 ( .A(n16476), .ZN(n10607) );
  INV_X1 U13558 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n10627) );
  NAND3_X1 U13559 ( .A1(n13490), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n10854), .ZN(n10866) );
  AOI22_X1 U13560 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10616) );
  AOI22_X1 U13561 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10612), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10615) );
  AOI22_X1 U13562 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10534), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10614) );
  AOI22_X1 U13563 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10542), .B1(
        n12557), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10613) );
  NAND4_X1 U13564 ( .A1(n10616), .A2(n10615), .A3(n10614), .A4(n10613), .ZN(
        n10626) );
  AOI22_X1 U13565 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12568), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10624) );
  INV_X1 U13566 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10619) );
  AOI22_X1 U13567 ( .A1(n12565), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n11088), .ZN(n10618) );
  NAND2_X1 U13568 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10617) );
  OAI211_X1 U13569 ( .C1(n13749), .C2(n10619), .A(n10618), .B(n10617), .ZN(
        n10620) );
  INV_X1 U13570 ( .A(n10620), .ZN(n10623) );
  NAND2_X1 U13571 ( .A1(n12563), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10622) );
  NAND2_X1 U13572 ( .A1(n12562), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10621) );
  NAND4_X1 U13573 ( .A1(n10624), .A2(n10623), .A3(n10622), .A4(n10621), .ZN(
        n10625) );
  MUX2_X1 U13574 ( .A(n10866), .B(n10976), .S(n13414), .Z(n10855) );
  MUX2_X1 U13575 ( .A(n10627), .B(n10855), .S(n10974), .Z(n10629) );
  AND2_X2 U13576 ( .A1(n10628), .A2(n10629), .ZN(n10675) );
  INV_X1 U13577 ( .A(n10675), .ZN(n10633) );
  INV_X1 U13578 ( .A(n10629), .ZN(n10630) );
  NAND2_X1 U13579 ( .A1(n10631), .A2(n10630), .ZN(n10632) );
  NAND2_X1 U13580 ( .A1(n10633), .A2(n10632), .ZN(n10634) );
  INV_X1 U13581 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14304) );
  XNOR2_X1 U13582 ( .A(n10634), .B(n14304), .ZN(n14203) );
  INV_X1 U13583 ( .A(n10634), .ZN(n15091) );
  NAND2_X1 U13584 ( .A1(n15091), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10635) );
  NAND2_X1 U13585 ( .A1(n10636), .A2(n10635), .ZN(n14297) );
  INV_X1 U13586 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10639) );
  INV_X1 U13587 ( .A(n10637), .ZN(n19543) );
  INV_X1 U13588 ( .A(n19800), .ZN(n19803) );
  INV_X1 U13589 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10638) );
  OAI22_X1 U13590 ( .A1(n10639), .A2(n19543), .B1(n19803), .B2(n10638), .ZN(
        n10640) );
  INV_X1 U13591 ( .A(n10640), .ZN(n10655) );
  INV_X1 U13592 ( .A(n10641), .ZN(n14103) );
  INV_X1 U13593 ( .A(n10682), .ZN(n19739) );
  AOI22_X1 U13594 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n14103), .B1(
        n19739), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10647) );
  INV_X1 U13595 ( .A(n19924), .ZN(n10690) );
  AOI22_X1 U13596 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19704), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10646) );
  INV_X1 U13597 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10642) );
  INV_X1 U13598 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10662) );
  OAI22_X1 U13599 ( .A1(n10642), .A2(n19479), .B1(n19663), .B2(n10662), .ZN(
        n10643) );
  INV_X1 U13600 ( .A(n10643), .ZN(n10645) );
  NAND2_X1 U13601 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10644) );
  AOI22_X1 U13602 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n10648), .B1(
        n10649), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10653) );
  INV_X1 U13603 ( .A(n10650), .ZN(n10691) );
  AOI22_X1 U13604 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n10691), .B1(
        n19829), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10652) );
  AOI22_X1 U13605 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19446), .B1(
        n9708), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10651) );
  NAND3_X1 U13606 ( .A1(n10655), .A2(n10218), .A3(n10248), .ZN(n10672) );
  AOI22_X1 U13607 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10659) );
  AOI22_X1 U13608 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10612), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10658) );
  AOI22_X1 U13609 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10534), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10657) );
  AOI22_X1 U13610 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n10542), .B1(
        n12557), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10656) );
  NAND4_X1 U13611 ( .A1(n10659), .A2(n10658), .A3(n10657), .A4(n10656), .ZN(
        n10669) );
  AOI22_X1 U13612 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12568), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10667) );
  AOI22_X1 U13613 ( .A1(n12565), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__5__SCAN_IN), .B2(n11088), .ZN(n10661) );
  NAND2_X1 U13614 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10660) );
  OAI211_X1 U13615 ( .C1(n13749), .C2(n10662), .A(n10661), .B(n10660), .ZN(
        n10663) );
  INV_X1 U13616 ( .A(n10663), .ZN(n10666) );
  NAND2_X1 U13617 ( .A1(n12563), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10665) );
  NAND2_X1 U13618 ( .A1(n12562), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10664) );
  NAND4_X1 U13619 ( .A1(n10667), .A2(n10666), .A3(n10665), .A4(n10664), .ZN(
        n10668) );
  INV_X1 U13620 ( .A(n11006), .ZN(n10670) );
  NAND2_X1 U13621 ( .A1(n10670), .A2(n9666), .ZN(n10671) );
  XNOR2_X2 U13622 ( .A(n10937), .B(n9716), .ZN(n10944) );
  NAND2_X1 U13623 ( .A1(n10944), .A2(n10961), .ZN(n10676) );
  INV_X1 U13624 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n10673) );
  MUX2_X1 U13625 ( .A(n10673), .B(n11006), .S(n10974), .Z(n10674) );
  OAI21_X1 U13626 ( .B1(n10675), .B2(n10674), .A(n10719), .ZN(n19217) );
  INV_X1 U13627 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14305) );
  NAND2_X1 U13628 ( .A1(n14297), .A2(n14298), .ZN(n10679) );
  NAND2_X1 U13629 ( .A1(n10677), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10678) );
  NAND2_X1 U13630 ( .A1(n10679), .A2(n10678), .ZN(n15401) );
  INV_X1 U13631 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10681) );
  INV_X1 U13632 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10680) );
  OAI22_X1 U13633 ( .A1(n10681), .A2(n19543), .B1(n19803), .B2(n10680), .ZN(
        n10698) );
  AOI22_X1 U13634 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19704), .B1(
        n19829), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10689) );
  INV_X1 U13635 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19434) );
  INV_X1 U13636 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12534) );
  OAI22_X1 U13637 ( .A1(n19434), .A2(n10641), .B1(n10682), .B2(n12534), .ZN(
        n10683) );
  INV_X1 U13638 ( .A(n10683), .ZN(n10688) );
  INV_X1 U13639 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10684) );
  INV_X1 U13640 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10705) );
  OAI22_X1 U13641 ( .A1(n10684), .A2(n19479), .B1(n19663), .B2(n10705), .ZN(
        n10685) );
  INV_X1 U13642 ( .A(n10685), .ZN(n10687) );
  NAND2_X1 U13643 ( .A1(n10511), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10686) );
  NAND4_X1 U13644 ( .A1(n10689), .A2(n10688), .A3(n10687), .A4(n10686), .ZN(
        n10697) );
  AOI22_X1 U13645 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10691), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10695) );
  AOI22_X1 U13646 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10648), .B1(
        n9708), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10694) );
  NAND2_X1 U13647 ( .A1(n10516), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10693) );
  AOI22_X1 U13648 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19446), .B1(
        n10649), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10692) );
  NAND4_X1 U13649 ( .A1(n10695), .A2(n10694), .A3(n10693), .A4(n10692), .ZN(
        n10696) );
  AOI22_X1 U13650 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10702) );
  AOI22_X1 U13651 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10612), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10701) );
  AOI22_X1 U13652 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10534), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10700) );
  AOI22_X1 U13653 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n10542), .B1(
        n12557), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10699) );
  NAND4_X1 U13654 ( .A1(n10702), .A2(n10701), .A3(n10700), .A4(n10699), .ZN(
        n10712) );
  AOI22_X1 U13655 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12568), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10710) );
  AOI22_X1 U13656 ( .A1(n12565), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n11088), .ZN(n10704) );
  NAND2_X1 U13657 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n10703) );
  OAI211_X1 U13658 ( .C1(n13749), .C2(n10705), .A(n10704), .B(n10703), .ZN(
        n10706) );
  INV_X1 U13659 ( .A(n10706), .ZN(n10709) );
  NAND2_X1 U13660 ( .A1(n12562), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10708) );
  NAND2_X1 U13661 ( .A1(n12563), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10707) );
  NAND4_X1 U13662 ( .A1(n10710), .A2(n10709), .A3(n10708), .A4(n10707), .ZN(
        n10711) );
  NAND2_X1 U13663 ( .A1(n11009), .A2(n9666), .ZN(n10713) );
  MUX2_X1 U13664 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n11009), .S(n10974), .Z(
        n10718) );
  XNOR2_X1 U13665 ( .A(n10719), .B(n10718), .ZN(n19202) );
  INV_X1 U13666 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15695) );
  NAND2_X1 U13667 ( .A1(n15401), .A2(n15402), .ZN(n10717) );
  NAND2_X1 U13668 ( .A1(n10715), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10716) );
  INV_X1 U13669 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n10720) );
  MUX2_X1 U13670 ( .A(n10720), .B(n11014), .S(n10974), .Z(n10723) );
  NAND2_X1 U13671 ( .A1(n10733), .A2(n10721), .ZN(n10722) );
  NAND2_X1 U13672 ( .A1(n10732), .A2(n10722), .ZN(n15082) );
  NOR2_X1 U13673 ( .A1(n15082), .A2(n10961), .ZN(n10726) );
  NAND2_X1 U13674 ( .A1(n10726), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16449) );
  INV_X1 U13675 ( .A(n10723), .ZN(n10724) );
  XNOR2_X1 U13676 ( .A(n10725), .B(n10724), .ZN(n14281) );
  NAND2_X1 U13677 ( .A1(n14281), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16450) );
  NAND2_X1 U13678 ( .A1(n16449), .A2(n16450), .ZN(n10730) );
  INV_X1 U13679 ( .A(n10726), .ZN(n10727) );
  INV_X1 U13680 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11205) );
  NAND2_X1 U13681 ( .A1(n10727), .A2(n11205), .ZN(n16448) );
  INV_X1 U13682 ( .A(n14281), .ZN(n10728) );
  INV_X1 U13683 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16514) );
  NAND2_X1 U13684 ( .A1(n10728), .A2(n16514), .ZN(n16452) );
  AND2_X1 U13685 ( .A1(n16448), .A2(n16452), .ZN(n10729) );
  NAND2_X1 U13686 ( .A1(n19422), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10731) );
  XNOR2_X1 U13687 ( .A(n10732), .B(n10731), .ZN(n15072) );
  AOI21_X1 U13688 ( .B1(n15072), .B2(n11014), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15680) );
  OR2_X2 U13689 ( .A1(n10733), .A2(n19422), .ZN(n10820) );
  AND2_X1 U13690 ( .A1(n19422), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10734) );
  NAND2_X1 U13691 ( .A1(n10736), .A2(n10734), .ZN(n10735) );
  OAI211_X1 U13692 ( .C1(n10736), .C2(P2_EBX_REG_10__SCAN_IN), .A(n10820), .B(
        n10735), .ZN(n15054) );
  INV_X1 U13693 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15674) );
  OAI21_X1 U13694 ( .B1(n15054), .B2(n10961), .A(n15674), .ZN(n15665) );
  INV_X1 U13695 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13886) );
  INV_X1 U13696 ( .A(n10737), .ZN(n10738) );
  AND3_X1 U13697 ( .A1(n19422), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n10738), .ZN(
        n10739) );
  NOR2_X1 U13698 ( .A1(n10745), .A2(n10739), .ZN(n19190) );
  AOI21_X1 U13699 ( .B1(n19190), .B2(n11014), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15647) );
  INV_X1 U13700 ( .A(n15054), .ZN(n10741) );
  AND2_X1 U13701 ( .A1(n11014), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10740) );
  NAND2_X1 U13702 ( .A1(n10741), .A2(n10740), .ZN(n15664) );
  AND2_X1 U13703 ( .A1(n11014), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10742) );
  NAND2_X1 U13704 ( .A1(n15072), .A2(n10742), .ZN(n15662) );
  NAND2_X1 U13705 ( .A1(n15664), .A2(n15662), .ZN(n15643) );
  INV_X1 U13706 ( .A(n19190), .ZN(n10744) );
  NAND2_X1 U13707 ( .A1(n11014), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10743) );
  NOR2_X1 U13708 ( .A1(n10744), .A2(n10743), .ZN(n15646) );
  NAND3_X1 U13709 ( .A1(n19422), .A2(P2_EBX_REG_12__SCAN_IN), .A3(n10746), 
        .ZN(n10747) );
  NAND2_X1 U13710 ( .A1(n10768), .A2(n10747), .ZN(n19174) );
  INV_X1 U13711 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15635) );
  NOR2_X1 U13712 ( .A1(n10748), .A2(n15635), .ZN(n15626) );
  NAND2_X1 U13713 ( .A1(n10748), .A2(n15635), .ZN(n15627) );
  INV_X1 U13714 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n19159) );
  NOR2_X1 U13715 ( .A1(n10974), .A2(n19159), .ZN(n10766) );
  OAI21_X1 U13716 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(P2_EBX_REG_14__SCAN_IN), 
        .A(n19422), .ZN(n10749) );
  INV_X1 U13717 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n15014) );
  INV_X1 U13718 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n19145) );
  NOR2_X1 U13719 ( .A1(n10974), .A2(n19145), .ZN(n10770) );
  INV_X1 U13720 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n15001) );
  NOR2_X1 U13721 ( .A1(n10974), .A2(n15001), .ZN(n10756) );
  NAND2_X1 U13722 ( .A1(n19422), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n10753) );
  INV_X1 U13723 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10750) );
  NAND2_X1 U13724 ( .A1(n10782), .A2(n10750), .ZN(n10751) );
  OR2_X2 U13725 ( .A1(n10751), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10800) );
  AND3_X1 U13726 ( .A1(n10751), .A2(n19422), .A3(P2_EBX_REG_21__SCAN_IN), .ZN(
        n10752) );
  OR2_X1 U13727 ( .A1(n10799), .A2(n10752), .ZN(n19102) );
  INV_X1 U13728 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15321) );
  OAI21_X1 U13729 ( .B1(n19102), .B2(n10961), .A(n15321), .ZN(n15317) );
  NOR2_X1 U13730 ( .A1(n10757), .A2(n10753), .ZN(n10754) );
  OR2_X1 U13731 ( .A1(n10782), .A2(n10754), .ZN(n19125) );
  NOR2_X1 U13732 ( .A1(n19125), .A2(n10961), .ZN(n10786) );
  INV_X1 U13733 ( .A(n10786), .ZN(n10755) );
  INV_X1 U13734 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15549) );
  NAND2_X1 U13735 ( .A1(n10755), .A2(n15549), .ZN(n15341) );
  AND2_X1 U13736 ( .A1(n10773), .A2(n10756), .ZN(n10758) );
  OR2_X1 U13737 ( .A1(n10758), .A2(n10757), .ZN(n15006) );
  INV_X1 U13738 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15555) );
  OAI21_X1 U13739 ( .B1(n15006), .B2(n10961), .A(n15555), .ZN(n15343) );
  NAND2_X1 U13740 ( .A1(n15341), .A2(n15343), .ZN(n15314) );
  NAND3_X1 U13741 ( .A1(n10759), .A2(n19422), .A3(P2_EBX_REG_16__SCAN_IN), 
        .ZN(n10760) );
  OAI211_X1 U13742 ( .C1(n10759), .C2(P2_EBX_REG_16__SCAN_IN), .A(n10820), .B(
        n10760), .ZN(n15007) );
  OR2_X1 U13743 ( .A1(n15007), .A2(n10961), .ZN(n10788) );
  XNOR2_X1 U13744 ( .A(n10788), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15308) );
  INV_X1 U13745 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n10762) );
  NAND2_X1 U13746 ( .A1(n10761), .A2(n10762), .ZN(n10777) );
  AND2_X1 U13747 ( .A1(n19422), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10763) );
  NAND2_X1 U13748 ( .A1(n10777), .A2(n10763), .ZN(n10764) );
  NAND2_X1 U13749 ( .A1(n10764), .A2(n10759), .ZN(n13407) );
  OR2_X1 U13750 ( .A1(n13407), .A2(n10961), .ZN(n10765) );
  INV_X1 U13751 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15589) );
  NAND2_X1 U13752 ( .A1(n10765), .A2(n15589), .ZN(n15380) );
  INV_X1 U13753 ( .A(n10766), .ZN(n10767) );
  XNOR2_X1 U13754 ( .A(n10768), .B(n10767), .ZN(n19164) );
  NAND2_X1 U13755 ( .A1(n19164), .A2(n11014), .ZN(n10769) );
  INV_X1 U13756 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16392) );
  NAND2_X1 U13757 ( .A1(n10769), .A2(n16392), .ZN(n15620) );
  AND2_X1 U13758 ( .A1(n15380), .A2(n15620), .ZN(n10779) );
  NAND2_X1 U13759 ( .A1(n10771), .A2(n10770), .ZN(n10772) );
  AND2_X1 U13760 ( .A1(n10773), .A2(n10772), .ZN(n19154) );
  INV_X1 U13761 ( .A(n19154), .ZN(n10775) );
  INV_X1 U13762 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10774) );
  OAI21_X1 U13763 ( .B1(n10775), .B2(n10961), .A(n10774), .ZN(n15311) );
  NAND2_X1 U13764 ( .A1(n19422), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10776) );
  MUX2_X1 U13765 ( .A(n10776), .B(n19422), .S(n10761), .Z(n10778) );
  NAND2_X1 U13766 ( .A1(n10778), .A2(n10777), .ZN(n15033) );
  INV_X1 U13767 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11230) );
  NAND2_X1 U13768 ( .A1(n10792), .A2(n11230), .ZN(n16388) );
  NAND4_X1 U13769 ( .A1(n15308), .A2(n10779), .A3(n15311), .A4(n16388), .ZN(
        n10780) );
  NOR2_X1 U13770 ( .A1(n15314), .A2(n10780), .ZN(n10784) );
  AND2_X1 U13771 ( .A1(n19422), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10781) );
  XNOR2_X1 U13772 ( .A(n10782), .B(n10781), .ZN(n19119) );
  NAND2_X1 U13773 ( .A1(n19119), .A2(n11014), .ZN(n10783) );
  INV_X1 U13774 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15538) );
  NAND2_X1 U13775 ( .A1(n10783), .A2(n15538), .ZN(n15328) );
  NAND3_X1 U13776 ( .A1(n15317), .A2(n10784), .A3(n15328), .ZN(n10797) );
  NAND2_X1 U13777 ( .A1(n11014), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10785) );
  NOR2_X1 U13778 ( .A1(n19102), .A2(n10785), .ZN(n15316) );
  NAND2_X1 U13779 ( .A1(n10786), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15342) );
  AND2_X1 U13780 ( .A1(n11014), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10787) );
  NAND2_X1 U13781 ( .A1(n19154), .A2(n10787), .ZN(n15310) );
  INV_X1 U13782 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11239) );
  OR2_X1 U13783 ( .A1(n10788), .A2(n11239), .ZN(n15309) );
  AND2_X1 U13784 ( .A1(n11014), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10789) );
  NAND2_X1 U13785 ( .A1(n19164), .A2(n10789), .ZN(n15619) );
  AND4_X1 U13786 ( .A1(n15310), .A2(n15309), .A3(n15379), .A4(n15619), .ZN(
        n10793) );
  INV_X1 U13787 ( .A(n15006), .ZN(n10791) );
  AND2_X1 U13788 ( .A1(n11014), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10790) );
  NAND2_X1 U13789 ( .A1(n10791), .A2(n10790), .ZN(n15313) );
  NAND4_X1 U13790 ( .A1(n15342), .A2(n10793), .A3(n15313), .A4(n16389), .ZN(
        n10794) );
  NOR2_X1 U13791 ( .A1(n15316), .A2(n10794), .ZN(n10796) );
  AND2_X1 U13792 ( .A1(n11014), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10795) );
  NAND2_X1 U13793 ( .A1(n19119), .A2(n10795), .ZN(n15327) );
  NAND2_X1 U13794 ( .A1(n19422), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10798) );
  NAND3_X1 U13795 ( .A1(n10800), .A2(n19422), .A3(P2_EBX_REG_22__SCAN_IN), 
        .ZN(n10801) );
  NAND2_X1 U13796 ( .A1(n10808), .A2(n10801), .ZN(n15867) );
  INV_X1 U13797 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15486) );
  NAND2_X1 U13798 ( .A1(n10802), .A2(n15486), .ZN(n15512) );
  INV_X1 U13799 ( .A(n10802), .ZN(n10803) );
  NAND2_X1 U13800 ( .A1(n10803), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15513) );
  INV_X1 U13801 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n14987) );
  NOR2_X1 U13802 ( .A1(n10974), .A2(n14987), .ZN(n10807) );
  XNOR2_X1 U13803 ( .A(n10808), .B(n10003), .ZN(n14975) );
  NAND2_X1 U13804 ( .A1(n14975), .A2(n11014), .ZN(n10805) );
  XNOR2_X1 U13805 ( .A(n10805), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15301) );
  INV_X1 U13806 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15485) );
  OR2_X1 U13807 ( .A1(n10805), .A2(n15485), .ZN(n10806) );
  NAND3_X1 U13808 ( .A1(n10810), .A2(n19422), .A3(P2_EBX_REG_24__SCAN_IN), 
        .ZN(n10809) );
  NAND2_X1 U13809 ( .A1(n10809), .A2(n10820), .ZN(n10811) );
  OR2_X1 U13810 ( .A1(n10811), .A2(n10822), .ZN(n14974) );
  NOR2_X1 U13811 ( .A1(n14974), .A2(n10961), .ZN(n10812) );
  AND2_X1 U13812 ( .A1(n10812), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15471) );
  INV_X1 U13813 ( .A(n10812), .ZN(n10813) );
  INV_X1 U13814 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15474) );
  NAND2_X1 U13815 ( .A1(n10813), .A2(n15474), .ZN(n15469) );
  INV_X1 U13816 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n15163) );
  AND3_X1 U13817 ( .A1(n19422), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n10814), .ZN(
        n10815) );
  OR2_X1 U13818 ( .A1(n10850), .A2(n10815), .ZN(n16318) );
  INV_X1 U13819 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15446) );
  OAI21_X1 U13820 ( .B1(n16318), .B2(n10961), .A(n15446), .ZN(n10817) );
  NAND2_X1 U13821 ( .A1(n11014), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10816) );
  NOR2_X1 U13822 ( .A1(n10822), .A2(n15163), .ZN(n10818) );
  NAND2_X1 U13823 ( .A1(n19422), .A2(n10818), .ZN(n10819) );
  NAND2_X1 U13824 ( .A1(n10820), .A2(n10819), .ZN(n10821) );
  AOI21_X1 U13825 ( .B1(n10822), .B2(n15163), .A(n10821), .ZN(n14947) );
  NAND2_X1 U13826 ( .A1(n19422), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10823) );
  NAND2_X1 U13827 ( .A1(n10850), .A2(n10823), .ZN(n10829) );
  INV_X1 U13828 ( .A(n10823), .ZN(n10824) );
  NAND2_X1 U13829 ( .A1(n10824), .A2(n9707), .ZN(n10825) );
  NAND2_X1 U13830 ( .A1(n10829), .A2(n10825), .ZN(n13445) );
  INV_X1 U13831 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15267) );
  NAND2_X1 U13832 ( .A1(n15267), .A2(n12341), .ZN(n10832) );
  INV_X1 U13833 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n10827) );
  NOR2_X1 U13834 ( .A1(n10974), .A2(n10827), .ZN(n10828) );
  OR2_X2 U13835 ( .A1(n10829), .A2(n10828), .ZN(n10843) );
  NAND2_X1 U13836 ( .A1(n10829), .A2(n10828), .ZN(n10830) );
  AND2_X1 U13837 ( .A1(n10843), .A2(n10830), .ZN(n14944) );
  NAND2_X1 U13838 ( .A1(n14944), .A2(n11014), .ZN(n12333) );
  INV_X1 U13839 ( .A(n12333), .ZN(n10831) );
  OAI21_X1 U13840 ( .B1(n10833), .B2(n10832), .A(n10831), .ZN(n10839) );
  NAND2_X1 U13841 ( .A1(n10833), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10838) );
  INV_X1 U13842 ( .A(n10834), .ZN(n10835) );
  INV_X1 U13843 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15456) );
  NOR2_X1 U13844 ( .A1(n10835), .A2(n15456), .ZN(n15284) );
  INV_X1 U13845 ( .A(n10836), .ZN(n10837) );
  NOR2_X1 U13846 ( .A1(n15284), .A2(n10837), .ZN(n12328) );
  NAND3_X1 U13847 ( .A1(n10839), .A2(n10838), .A3(n12328), .ZN(n15258) );
  INV_X1 U13848 ( .A(n10843), .ZN(n10840) );
  NAND2_X1 U13849 ( .A1(n19422), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n10841) );
  XNOR2_X1 U13850 ( .A(n10840), .B(n10841), .ZN(n10847) );
  INV_X1 U13851 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15422) );
  OAI21_X1 U13852 ( .B1(n10847), .B2(n10961), .A(n15422), .ZN(n15256) );
  INV_X1 U13853 ( .A(n10841), .ZN(n10842) );
  NOR2_X2 U13854 ( .A1(n10843), .A2(n10842), .ZN(n10848) );
  INV_X1 U13855 ( .A(n10848), .ZN(n10845) );
  NAND2_X1 U13856 ( .A1(n19422), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10844) );
  AOI21_X1 U13857 ( .B1(n14933), .B2(n11014), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12376) );
  AND2_X1 U13858 ( .A1(n11014), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10846) );
  NAND2_X1 U13859 ( .A1(n14933), .A2(n10846), .ZN(n12374) );
  INV_X1 U13860 ( .A(n10847), .ZN(n16315) );
  NAND3_X1 U13861 ( .A1(n16315), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11014), .ZN(n15257) );
  INV_X1 U13862 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n14443) );
  NAND2_X1 U13863 ( .A1(n10848), .A2(n14443), .ZN(n10849) );
  MUX2_X1 U13864 ( .A(n10850), .B(n10849), .S(n19422), .Z(n16300) );
  NOR2_X1 U13865 ( .A1(n16300), .A2(n10961), .ZN(n10851) );
  XOR2_X1 U13866 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n10851), .Z(
        n10852) );
  INV_X1 U13867 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15938) );
  NOR2_X1 U13868 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15938), .ZN(
        n10853) );
  INV_X1 U13869 ( .A(n10855), .ZN(n10861) );
  INV_X1 U13870 ( .A(n10868), .ZN(n10900) );
  NOR2_X1 U13871 ( .A1(n10900), .A2(n10901), .ZN(n10859) );
  INV_X1 U13872 ( .A(n10856), .ZN(n10857) );
  OAI21_X1 U13873 ( .B1(n10859), .B2(n10858), .A(n10857), .ZN(n10860) );
  NOR2_X1 U13874 ( .A1(n10861), .A2(n10860), .ZN(n10862) );
  OR2_X1 U13875 ( .A1(n10915), .A2(n10862), .ZN(n14912) );
  INV_X1 U13876 ( .A(n10863), .ZN(n10877) );
  NAND2_X1 U13877 ( .A1(n10877), .A2(n12336), .ZN(n14916) );
  NOR2_X1 U13878 ( .A1(n14912), .A2(n14916), .ZN(n10879) );
  INV_X1 U13879 ( .A(n10864), .ZN(n10865) );
  OR2_X1 U13880 ( .A1(n10912), .A2(n10905), .ZN(n10870) );
  XNOR2_X1 U13881 ( .A(n10868), .B(n10867), .ZN(n10897) );
  NOR2_X1 U13882 ( .A1(n10897), .A2(n10870), .ZN(n10869) );
  OR2_X1 U13883 ( .A1(n10915), .A2(n10869), .ZN(n13472) );
  INV_X1 U13884 ( .A(n13472), .ZN(n14051) );
  OAI21_X1 U13885 ( .B1(n10901), .B2(n10870), .A(n14051), .ZN(n10876) );
  INV_X1 U13886 ( .A(n10871), .ZN(n10873) );
  AOI21_X1 U13887 ( .B1(n10872), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13487) );
  NAND2_X1 U13888 ( .A1(n10873), .A2(n13487), .ZN(n10874) );
  INV_X1 U13889 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n15936) );
  NAND2_X1 U13890 ( .A1(n10874), .A2(n15936), .ZN(n10875) );
  NAND2_X1 U13891 ( .A1(n10875), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20099) );
  OAI21_X1 U13892 ( .B1(n10876), .B2(P2_STATE2_REG_1__SCAN_IN), .A(n20099), 
        .ZN(n16540) );
  AND2_X1 U13893 ( .A1(n16540), .A2(n10877), .ZN(n10878) );
  MUX2_X1 U13894 ( .A(n10879), .B(n10878), .S(n9676), .Z(n12338) );
  INV_X1 U13895 ( .A(n12338), .ZN(n10924) );
  MUX2_X1 U13896 ( .A(n10880), .B(n19411), .S(n9666), .Z(n10881) );
  NAND2_X1 U13897 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n14909) );
  INV_X1 U13898 ( .A(n14909), .ZN(n20003) );
  NOR2_X1 U13899 ( .A1(n10881), .A2(n20003), .ZN(n10894) );
  INV_X1 U13900 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19074) );
  INV_X1 U13901 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20011) );
  NOR2_X1 U13902 ( .A1(n19074), .A2(n20011), .ZN(n20002) );
  NOR2_X1 U13903 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20004) );
  NOR3_X1 U13904 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20002), .A3(n20004), 
        .ZN(n19996) );
  NAND2_X1 U13905 ( .A1(n14909), .A2(n19996), .ZN(n13395) );
  INV_X1 U13906 ( .A(n13395), .ZN(n13477) );
  NAND2_X1 U13907 ( .A1(n14051), .A2(n13477), .ZN(n10893) );
  OAI211_X1 U13908 ( .C1(n10882), .C2(n9658), .A(n9666), .B(n12336), .ZN(
        n11307) );
  NAND2_X1 U13909 ( .A1(n9666), .A2(n10361), .ZN(n11301) );
  NAND2_X1 U13910 ( .A1(n11301), .A2(n10353), .ZN(n10884) );
  NAND2_X1 U13911 ( .A1(n10884), .A2(n10883), .ZN(n10885) );
  NAND2_X1 U13912 ( .A1(n10885), .A2(n19411), .ZN(n10886) );
  AND2_X1 U13913 ( .A1(n10887), .A2(n10886), .ZN(n10892) );
  NAND2_X1 U13914 ( .A1(n10889), .A2(n19411), .ZN(n10890) );
  NAND2_X1 U13915 ( .A1(n10888), .A2(n10890), .ZN(n10891) );
  OAI21_X1 U13916 ( .B1(n10893), .B2(n10880), .A(n11303), .ZN(n13478) );
  AOI21_X1 U13917 ( .B1(n14051), .B2(n10894), .A(n13478), .ZN(n10923) );
  NAND2_X1 U13918 ( .A1(n10896), .A2(n10895), .ZN(n10904) );
  INV_X1 U13919 ( .A(n10901), .ZN(n10899) );
  INV_X1 U13920 ( .A(n10897), .ZN(n10898) );
  OAI211_X1 U13921 ( .C1(n9676), .C2(n10899), .A(n10353), .B(n10898), .ZN(
        n10903) );
  OAI21_X1 U13922 ( .B1(n10901), .B2(n10900), .A(n13414), .ZN(n10902) );
  NAND3_X1 U13923 ( .A1(n10904), .A2(n10903), .A3(n10902), .ZN(n10909) );
  OAI21_X1 U13924 ( .B1(n14899), .B2(n9666), .A(n10905), .ZN(n10907) );
  NAND2_X1 U13925 ( .A1(n10907), .A2(n10906), .ZN(n10908) );
  NAND2_X1 U13926 ( .A1(n10909), .A2(n10908), .ZN(n10911) );
  NAND2_X1 U13927 ( .A1(n10912), .A2(n13414), .ZN(n10910) );
  OAI21_X1 U13928 ( .B1(n10912), .B2(n10911), .A(n10910), .ZN(n10913) );
  OR2_X1 U13929 ( .A1(n10915), .A2(n10913), .ZN(n10914) );
  MUX2_X1 U13930 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n10914), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n10918) );
  NAND2_X1 U13931 ( .A1(n10915), .A2(n14899), .ZN(n10916) );
  AND2_X1 U13932 ( .A1(n13261), .A2(n9676), .ZN(n13476) );
  NAND3_X1 U13933 ( .A1(n13476), .A2(n10917), .A3(n13477), .ZN(n10922) );
  INV_X1 U13934 ( .A(n13476), .ZN(n10920) );
  AOI21_X1 U13935 ( .B1(n10918), .B2(n10353), .A(n19416), .ZN(n10919) );
  NAND2_X1 U13936 ( .A1(n10920), .A2(n10919), .ZN(n10921) );
  NAND4_X1 U13937 ( .A1(n10924), .A2(n10923), .A3(n10922), .A4(n10921), .ZN(
        n10925) );
  INV_X1 U13938 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n11320) );
  NAND3_X1 U13939 ( .A1(n11320), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n16548) );
  INV_X1 U13940 ( .A(n14916), .ZN(n14057) );
  INV_X1 U13941 ( .A(n10926), .ZN(n16480) );
  NAND2_X1 U13942 ( .A1(n13496), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13495) );
  NOR2_X1 U13943 ( .A1(n10989), .A2(n13495), .ZN(n10928) );
  INV_X1 U13944 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13550) );
  AND2_X1 U13945 ( .A1(n13496), .A2(n13494), .ZN(n10927) );
  XNOR2_X1 U13946 ( .A(n10927), .B(n10989), .ZN(n13549) );
  NOR2_X1 U13947 ( .A1(n13550), .A2(n13549), .ZN(n13548) );
  NOR2_X1 U13948 ( .A1(n10928), .A2(n13548), .ZN(n10931) );
  XNOR2_X1 U13949 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n10931), .ZN(
        n13645) );
  XNOR2_X1 U13950 ( .A(n10930), .B(n10929), .ZN(n13644) );
  NAND2_X1 U13951 ( .A1(n13645), .A2(n13644), .ZN(n13643) );
  OR2_X1 U13952 ( .A1(n10931), .A2(n14458), .ZN(n10932) );
  NAND2_X1 U13953 ( .A1(n13643), .A2(n10932), .ZN(n10938) );
  XNOR2_X1 U13954 ( .A(n10938), .B(n16534), .ZN(n16479) );
  AND2_X1 U13955 ( .A1(n16479), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10933) );
  INV_X1 U13956 ( .A(n10976), .ZN(n10934) );
  NAND2_X1 U13957 ( .A1(n10935), .A2(n10934), .ZN(n10936) );
  NAND2_X1 U13958 ( .A1(n10937), .A2(n10936), .ZN(n14205) );
  NAND2_X1 U13959 ( .A1(n10938), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14206) );
  OR2_X1 U13960 ( .A1(n14304), .A2(n14206), .ZN(n10939) );
  NAND3_X1 U13961 ( .A1(n10940), .A2(n14205), .A3(n10939), .ZN(n10943) );
  AND2_X1 U13962 ( .A1(n14304), .A2(n14206), .ZN(n10941) );
  NAND2_X1 U13963 ( .A1(n16478), .A2(n10941), .ZN(n10942) );
  INV_X1 U13964 ( .A(n10944), .ZN(n10945) );
  NAND2_X1 U13965 ( .A1(n10945), .A2(n14305), .ZN(n14309) );
  NAND2_X1 U13966 ( .A1(n10944), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14310) );
  NAND2_X1 U13967 ( .A1(n14314), .A2(n14310), .ZN(n10947) );
  NAND2_X1 U13968 ( .A1(n10947), .A2(n10946), .ZN(n10951) );
  INV_X1 U13969 ( .A(n14310), .ZN(n14313) );
  NAND2_X1 U13970 ( .A1(n14313), .A2(n10953), .ZN(n10950) );
  INV_X1 U13971 ( .A(n10953), .ZN(n10954) );
  NAND2_X1 U13972 ( .A1(n15390), .A2(n16514), .ZN(n10956) );
  NAND2_X1 U13973 ( .A1(n15389), .A2(n10956), .ZN(n10959) );
  INV_X1 U13974 ( .A(n15390), .ZN(n10957) );
  NAND2_X1 U13975 ( .A1(n10957), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10958) );
  NAND2_X1 U13976 ( .A1(n16455), .A2(n16456), .ZN(n10964) );
  AND2_X1 U13977 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16495) );
  NAND2_X1 U13978 ( .A1(n16495), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16493) );
  AND2_X1 U13979 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15518) );
  AND2_X1 U13980 ( .A1(n15518), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11339) );
  INV_X1 U13981 ( .A(n11339), .ZN(n10965) );
  OR2_X1 U13982 ( .A1(n10965), .A2(n15555), .ZN(n10966) );
  AND2_X1 U13983 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11335) );
  NAND2_X1 U13984 ( .A1(n10967), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15288) );
  INV_X1 U13985 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12341) );
  INV_X1 U13986 ( .A(n16527), .ZN(n10972) );
  NAND2_X1 U13987 ( .A1(n13319), .A2(n10972), .ZN(n11349) );
  INV_X1 U13988 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19392) );
  INV_X2 U13989 ( .A(n9736), .ZN(n11150) );
  AOI22_X1 U13990 ( .A1(n11150), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n9669), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10978) );
  NAND2_X1 U13991 ( .A1(n11147), .A2(n10976), .ZN(n10977) );
  OAI211_X1 U13992 ( .C1(n11175), .C2(n19392), .A(n10978), .B(n10977), .ZN(
        n14214) );
  NAND2_X1 U13993 ( .A1(n10979), .A2(n9668), .ZN(n10994) );
  MUX2_X1 U13994 ( .A(n13279), .B(n20106), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10980) );
  AND2_X1 U13995 ( .A1(n10994), .A2(n10980), .ZN(n10981) );
  INV_X1 U13996 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19091) );
  AOI21_X1 U13997 ( .B1(n10983), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10985) );
  NAND2_X1 U13998 ( .A1(n9658), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n10984) );
  INV_X1 U13999 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19354) );
  INV_X1 U14000 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20013) );
  XNOR2_X1 U14001 ( .A(n13607), .B(n10990), .ZN(n13616) );
  NAND2_X1 U14002 ( .A1(n10358), .A2(n13279), .ZN(n10986) );
  MUX2_X1 U14003 ( .A(n20098), .B(n10986), .S(n13484), .Z(n10987) );
  OAI21_X1 U14004 ( .B1(n10989), .B2(n10988), .A(n10987), .ZN(n13617) );
  NOR2_X1 U14005 ( .A1(n13616), .A2(n13617), .ZN(n10992) );
  NOR2_X1 U14006 ( .A1(n13607), .A2(n10990), .ZN(n10991) );
  NAND2_X1 U14007 ( .A1(n11147), .A2(n10993), .ZN(n10995) );
  OAI211_X1 U14008 ( .C1(n13484), .C2(n20088), .A(n10995), .B(n10994), .ZN(
        n10997) );
  XNOR2_X1 U14009 ( .A(n10998), .B(n10997), .ZN(n13804) );
  INV_X1 U14010 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20014) );
  AOI22_X1 U14011 ( .A1(n11150), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n9669), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10996) );
  OAI21_X1 U14012 ( .B1(n11175), .B2(n20014), .A(n10996), .ZN(n13803) );
  NOR2_X1 U14013 ( .A1(n13804), .A2(n13803), .ZN(n13805) );
  NOR2_X1 U14014 ( .A1(n10998), .A2(n10997), .ZN(n10999) );
  INV_X1 U14015 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n16471) );
  AOI22_X1 U14016 ( .A1(n9669), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11001) );
  NAND2_X1 U14017 ( .A1(n11150), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11000) );
  AND2_X1 U14018 ( .A1(n11001), .A2(n11000), .ZN(n11005) );
  INV_X1 U14019 ( .A(n11002), .ZN(n11003) );
  NAND2_X1 U14020 ( .A1(n11147), .A2(n11003), .ZN(n11004) );
  OAI211_X1 U14021 ( .C1(n11175), .C2(n16471), .A(n11005), .B(n11004), .ZN(
        n15109) );
  INV_X1 U14022 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n16460) );
  AOI22_X1 U14023 ( .A1(n11150), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n9669), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11008) );
  NAND2_X1 U14024 ( .A1(n11147), .A2(n11006), .ZN(n11007) );
  OAI211_X1 U14025 ( .C1(n11175), .C2(n16460), .A(n11008), .B(n11007), .ZN(
        n14301) );
  INV_X1 U14026 ( .A(n11009), .ZN(n11010) );
  NAND2_X1 U14027 ( .A1(n11147), .A2(n11010), .ZN(n11011) );
  INV_X1 U14028 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20019) );
  AOI22_X1 U14029 ( .A1(n11150), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n9669), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11013) );
  OAI21_X1 U14030 ( .B1(n11175), .B2(n20019), .A(n11013), .ZN(n15699) );
  NAND2_X1 U14031 ( .A1(n15698), .A2(n15699), .ZN(n11016) );
  NAND2_X1 U14032 ( .A1(n11147), .A2(n11014), .ZN(n11015) );
  INV_X1 U14033 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20021) );
  AOI22_X1 U14034 ( .A1(n11150), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n9669), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11017) );
  OAI21_X1 U14035 ( .B1(n11175), .B2(n20021), .A(n11017), .ZN(n14273) );
  INV_X1 U14036 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n11032) );
  AOI22_X1 U14037 ( .A1(n11150), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n9669), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11031) );
  AOI22_X1 U14038 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12555), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11021) );
  AOI22_X1 U14039 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11020) );
  AOI22_X1 U14040 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10612), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11019) );
  AOI22_X1 U14041 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n10542), .B1(
        n12557), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11018) );
  NAND4_X1 U14042 ( .A1(n11021), .A2(n11020), .A3(n11019), .A4(n11018), .ZN(
        n11029) );
  AOI22_X1 U14043 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n12569), .B1(
        n12563), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11027) );
  AOI22_X1 U14044 ( .A1(n12565), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__0__SCAN_IN), .B2(n12564), .ZN(n11023) );
  NAND2_X1 U14045 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11022) );
  AND2_X1 U14046 ( .A1(n11023), .A2(n11022), .ZN(n11026) );
  AOI22_X1 U14047 ( .A1(n12562), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12568), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11025) );
  NAND2_X1 U14048 ( .A1(n10534), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11024) );
  NAND4_X1 U14049 ( .A1(n11027), .A2(n11026), .A3(n11025), .A4(n11024), .ZN(
        n11028) );
  NAND2_X1 U14050 ( .A1(n11147), .A2(n19253), .ZN(n11030) );
  OAI211_X1 U14051 ( .C1(n11175), .C2(n11032), .A(n11031), .B(n11030), .ZN(
        n11033) );
  INV_X1 U14052 ( .A(n11033), .ZN(n15079) );
  INV_X1 U14053 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n16436) );
  AOI22_X1 U14054 ( .A1(n11150), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n9669), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11050) );
  AOI22_X1 U14055 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11038) );
  AOI22_X1 U14056 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10612), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11037) );
  AOI22_X1 U14057 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10534), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11036) );
  AOI22_X1 U14058 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n10542), .B1(
        n12557), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11035) );
  NAND4_X1 U14059 ( .A1(n11038), .A2(n11037), .A3(n11036), .A4(n11035), .ZN(
        n11048) );
  AOI22_X1 U14060 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12568), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11046) );
  AOI22_X1 U14061 ( .A1(n12565), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n12564), .ZN(n11040) );
  NAND2_X1 U14062 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11039) );
  OAI211_X1 U14063 ( .C1(n13749), .C2(n11041), .A(n11040), .B(n11039), .ZN(
        n11042) );
  INV_X1 U14064 ( .A(n11042), .ZN(n11045) );
  NAND2_X1 U14065 ( .A1(n12563), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11044) );
  NAND2_X1 U14066 ( .A1(n12562), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11043) );
  NAND4_X1 U14067 ( .A1(n11046), .A2(n11045), .A3(n11044), .A4(n11043), .ZN(
        n11047) );
  NAND2_X1 U14068 ( .A1(n11147), .A2(n13831), .ZN(n11049) );
  OAI211_X1 U14069 ( .C1(n11175), .C2(n16436), .A(n11050), .B(n11049), .ZN(
        n15065) );
  INV_X1 U14070 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n15053) );
  AOI22_X1 U14071 ( .A1(n11150), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n9669), .B2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11066) );
  AOI22_X1 U14072 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12556), .B1(
        n9659), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11054) );
  AOI22_X1 U14073 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n10542), .B1(
        n12557), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11053) );
  AOI22_X1 U14074 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10612), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11052) );
  AOI22_X1 U14075 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10534), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11051) );
  NAND4_X1 U14076 ( .A1(n11054), .A2(n11053), .A3(n11052), .A4(n11051), .ZN(
        n11064) );
  AOI22_X1 U14077 ( .A1(n12562), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12568), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11062) );
  INV_X1 U14078 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11057) );
  AOI22_X1 U14079 ( .A1(n12565), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n12564), .ZN(n11056) );
  NAND2_X1 U14080 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11055) );
  OAI211_X1 U14081 ( .C1(n13749), .C2(n11057), .A(n11056), .B(n11055), .ZN(
        n11058) );
  INV_X1 U14082 ( .A(n11058), .ZN(n11061) );
  NAND2_X1 U14083 ( .A1(n12563), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11060) );
  NAND2_X1 U14084 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11059) );
  NAND4_X1 U14085 ( .A1(n11062), .A2(n11061), .A3(n11060), .A4(n11059), .ZN(
        n11063) );
  NAND2_X1 U14086 ( .A1(n11147), .A2(n13882), .ZN(n11065) );
  OAI211_X1 U14087 ( .C1(n11175), .C2(n15053), .A(n11066), .B(n11065), .ZN(
        n15043) );
  INV_X1 U14088 ( .A(n15043), .ZN(n11067) );
  AOI22_X1 U14089 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11071) );
  AOI22_X1 U14090 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10612), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11070) );
  AOI22_X1 U14091 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10534), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11069) );
  AOI22_X1 U14092 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n10542), .B1(
        n12557), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11068) );
  NAND4_X1 U14093 ( .A1(n11071), .A2(n11070), .A3(n11069), .A4(n11068), .ZN(
        n11081) );
  AOI22_X1 U14094 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12568), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11079) );
  INV_X1 U14095 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11074) );
  AOI22_X1 U14096 ( .A1(n12565), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n12564), .ZN(n11073) );
  NAND2_X1 U14097 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11072) );
  OAI211_X1 U14098 ( .C1(n13749), .C2(n11074), .A(n11073), .B(n11072), .ZN(
        n11075) );
  INV_X1 U14099 ( .A(n11075), .ZN(n11078) );
  NAND2_X1 U14100 ( .A1(n12563), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11077) );
  NAND2_X1 U14101 ( .A1(n12562), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n11076) );
  NAND4_X1 U14102 ( .A1(n11079), .A2(n11078), .A3(n11077), .A4(n11076), .ZN(
        n11080) );
  AOI22_X1 U14103 ( .A1(n11170), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n11147), 
        .B2(n19241), .ZN(n11083) );
  AOI22_X1 U14104 ( .A1(n11150), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n9669), .B2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11082) );
  NAND2_X1 U14105 ( .A1(n11083), .A2(n11082), .ZN(n15650) );
  INV_X1 U14106 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19170) );
  AOI22_X1 U14107 ( .A1(n11150), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n9669), .B2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11098) );
  AOI22_X1 U14108 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12556), .B1(
        n10519), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11087) );
  AOI22_X1 U14109 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10542), .B1(
        n12557), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11086) );
  AOI22_X1 U14110 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10612), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11085) );
  AOI22_X1 U14111 ( .A1(n12555), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11084) );
  NAND4_X1 U14112 ( .A1(n11087), .A2(n11086), .A3(n11085), .A4(n11084), .ZN(
        n11096) );
  AOI22_X1 U14113 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12569), .B1(
        n12563), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11094) );
  BUF_X1 U14114 ( .A(n11088), .Z(n12564) );
  AOI22_X1 U14115 ( .A1(n12565), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n12564), .ZN(n11090) );
  NAND2_X1 U14116 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11089) );
  AND2_X1 U14117 ( .A1(n11090), .A2(n11089), .ZN(n11093) );
  AOI22_X1 U14118 ( .A1(n12562), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12568), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11092) );
  NAND2_X1 U14119 ( .A1(n10534), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11091) );
  NAND4_X1 U14120 ( .A1(n11094), .A2(n11093), .A3(n11092), .A4(n11091), .ZN(
        n11095) );
  OR2_X1 U14121 ( .A1(n11096), .A2(n11095), .ZN(n19240) );
  NAND2_X1 U14122 ( .A1(n11147), .A2(n19240), .ZN(n11097) );
  OAI211_X1 U14123 ( .C1(n11175), .C2(n19170), .A(n11098), .B(n11097), .ZN(
        n11099) );
  INV_X1 U14124 ( .A(n11099), .ZN(n15631) );
  INV_X1 U14125 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n16401) );
  AOI22_X1 U14126 ( .A1(n11150), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n9669), .B2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11115) );
  AOI22_X1 U14127 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11103) );
  AOI22_X1 U14128 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10612), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11102) );
  AOI22_X1 U14129 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10534), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11101) );
  AOI22_X1 U14130 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n10542), .B1(
        n12557), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11100) );
  NAND4_X1 U14131 ( .A1(n11103), .A2(n11102), .A3(n11101), .A4(n11100), .ZN(
        n11113) );
  AOI22_X1 U14132 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12568), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11111) );
  INV_X1 U14133 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11106) );
  AOI22_X1 U14134 ( .A1(n12565), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__5__SCAN_IN), .B2(n12564), .ZN(n11105) );
  NAND2_X1 U14135 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11104) );
  OAI211_X1 U14136 ( .C1(n13749), .C2(n11106), .A(n11105), .B(n11104), .ZN(
        n11107) );
  INV_X1 U14137 ( .A(n11107), .ZN(n11110) );
  NAND2_X1 U14138 ( .A1(n12563), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11109) );
  NAND2_X1 U14139 ( .A1(n12562), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11108) );
  NAND4_X1 U14140 ( .A1(n11111), .A2(n11110), .A3(n11109), .A4(n11108), .ZN(
        n11112) );
  NAND2_X1 U14141 ( .A1(n11147), .A2(n13911), .ZN(n11114) );
  OAI211_X1 U14142 ( .C1(n11175), .C2(n16401), .A(n11115), .B(n11114), .ZN(
        n15612) );
  INV_X1 U14143 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n11131) );
  AOI22_X1 U14144 ( .A1(n11150), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n9669), .B2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11130) );
  AOI22_X1 U14145 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12556), .B1(
        n9659), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11119) );
  AOI22_X1 U14146 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n10542), .B1(
        n12557), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11118) );
  AOI22_X1 U14147 ( .A1(n12555), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11117) );
  AOI22_X1 U14148 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10612), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11116) );
  NAND4_X1 U14149 ( .A1(n11119), .A2(n11118), .A3(n11117), .A4(n11116), .ZN(
        n11127) );
  AOI22_X1 U14150 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n12562), .B1(
        n12563), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11125) );
  AOI22_X1 U14151 ( .A1(n12565), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n12564), .ZN(n11121) );
  NAND2_X1 U14152 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11120) );
  AND2_X1 U14153 ( .A1(n11121), .A2(n11120), .ZN(n11124) );
  AOI22_X1 U14154 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12568), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11123) );
  NAND2_X1 U14155 ( .A1(n10534), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11122) );
  NAND4_X1 U14156 ( .A1(n11125), .A2(n11124), .A3(n11123), .A4(n11122), .ZN(
        n11126) );
  NOR2_X1 U14157 ( .A1(n11127), .A2(n11126), .ZN(n19236) );
  INV_X1 U14158 ( .A(n19236), .ZN(n11128) );
  NAND2_X1 U14159 ( .A1(n11147), .A2(n11128), .ZN(n11129) );
  OAI211_X1 U14160 ( .C1(n11175), .C2(n11131), .A(n11130), .B(n11129), .ZN(
        n11132) );
  INV_X1 U14161 ( .A(n11132), .ZN(n15030) );
  AOI22_X1 U14162 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11136) );
  AOI22_X1 U14163 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10612), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11135) );
  AOI22_X1 U14164 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10534), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11134) );
  AOI22_X1 U14165 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n10542), .B1(
        n12557), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11133) );
  NAND4_X1 U14166 ( .A1(n11136), .A2(n11135), .A3(n11134), .A4(n11133), .ZN(
        n11146) );
  AOI22_X1 U14167 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12568), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11144) );
  INV_X1 U14168 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11139) );
  AOI22_X1 U14169 ( .A1(n12565), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n12564), .ZN(n11138) );
  NAND2_X1 U14170 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11137) );
  OAI211_X1 U14171 ( .C1(n13749), .C2(n11139), .A(n11138), .B(n11137), .ZN(
        n11140) );
  INV_X1 U14172 ( .A(n11140), .ZN(n11143) );
  NAND2_X1 U14173 ( .A1(n12563), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11142) );
  NAND2_X1 U14174 ( .A1(n12562), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11141) );
  NAND4_X1 U14175 ( .A1(n11144), .A2(n11143), .A3(n11142), .A4(n11141), .ZN(
        n11145) );
  AOI22_X1 U14176 ( .A1(n11170), .A2(P2_REIP_REG_15__SCAN_IN), .B1(n11147), 
        .B2(n14029), .ZN(n11149) );
  AOI22_X1 U14177 ( .A1(n11150), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n9669), .B2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11148) );
  NAND2_X1 U14178 ( .A1(n11149), .A2(n11148), .ZN(n13409) );
  NAND2_X1 U14179 ( .A1(n13408), .A2(n13409), .ZN(n15021) );
  AOI222_X1 U14180 ( .A1(n11170), .A2(P2_REIP_REG_16__SCAN_IN), .B1(n11150), 
        .B2(P2_EAX_REG_16__SCAN_IN), .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), 
        .C2(n9669), .ZN(n15020) );
  INV_X1 U14181 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20035) );
  AOI22_X1 U14182 ( .A1(n11150), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n9669), .B2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11151) );
  OAI21_X1 U14183 ( .B1(n11175), .B2(n20035), .A(n11151), .ZN(n14353) );
  INV_X1 U14184 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n15355) );
  AOI22_X1 U14185 ( .A1(n11150), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n9669), .B2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11152) );
  OAI21_X1 U14186 ( .B1(n11175), .B2(n15355), .A(n11152), .ZN(n11153) );
  INV_X1 U14187 ( .A(n11153), .ZN(n14995) );
  INV_X1 U14188 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20038) );
  AOI22_X1 U14189 ( .A1(n11150), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n9669), .B2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11154) );
  OAI21_X1 U14190 ( .B1(n11175), .B2(n20038), .A(n11154), .ZN(n11155) );
  INV_X1 U14191 ( .A(n11155), .ZN(n15244) );
  INV_X1 U14192 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n11256) );
  AOI22_X1 U14193 ( .A1(n11150), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n9669), .B2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11156) );
  OAI21_X1 U14194 ( .B1(n11175), .B2(n11256), .A(n11156), .ZN(n11157) );
  INV_X1 U14195 ( .A(n11157), .ZN(n15528) );
  NOR2_X2 U14196 ( .A1(n15529), .A2(n15528), .ZN(n15530) );
  INV_X1 U14197 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20041) );
  AOI22_X1 U14198 ( .A1(n11150), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n9668), .B2(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11158) );
  OAI21_X1 U14199 ( .B1(n11175), .B2(n20041), .A(n11158), .ZN(n15235) );
  AND2_X2 U14200 ( .A1(n15530), .A2(n15235), .ZN(n15504) );
  INV_X1 U14201 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n11263) );
  AOI22_X1 U14202 ( .A1(n11150), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n9669), .B2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11159) );
  OAI21_X1 U14203 ( .B1(n11175), .B2(n11263), .A(n11159), .ZN(n15505) );
  INV_X1 U14204 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20044) );
  AOI22_X1 U14205 ( .A1(n11150), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n9668), .B2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11160) );
  OAI21_X1 U14206 ( .B1(n11175), .B2(n20044), .A(n11160), .ZN(n14983) );
  NAND2_X1 U14207 ( .A1(n11170), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11162) );
  AOI22_X1 U14208 ( .A1(n11150), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n9669), .B2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11161) );
  AND2_X1 U14209 ( .A1(n11162), .A2(n11161), .ZN(n14964) );
  NAND2_X1 U14210 ( .A1(n11170), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11164) );
  AOI22_X1 U14211 ( .A1(n11150), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n9669), .B2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11163) );
  AND2_X1 U14212 ( .A1(n11164), .A2(n11163), .ZN(n14949) );
  INV_X1 U14213 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20050) );
  AOI22_X1 U14214 ( .A1(n11150), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n9668), .B2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11165) );
  OAI21_X1 U14215 ( .B1(n11175), .B2(n20050), .A(n11165), .ZN(n15208) );
  NAND2_X1 U14216 ( .A1(n15209), .A2(n15208), .ZN(n13449) );
  NAND2_X1 U14217 ( .A1(n11170), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11167) );
  AOI22_X1 U14218 ( .A1(n11150), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n9669), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11166) );
  AND2_X1 U14219 ( .A1(n11167), .A2(n11166), .ZN(n13450) );
  OR2_X2 U14220 ( .A1(n13449), .A2(n13450), .ZN(n13452) );
  NAND2_X1 U14221 ( .A1(n11170), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11169) );
  AOI22_X1 U14222 ( .A1(n11150), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n9669), .B2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11168) );
  AND2_X1 U14223 ( .A1(n11169), .A2(n11168), .ZN(n12363) );
  OR2_X2 U14224 ( .A1(n13452), .A2(n12363), .ZN(n14448) );
  NAND2_X1 U14225 ( .A1(n11170), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11172) );
  AOI22_X1 U14226 ( .A1(n11150), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n9668), .B2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11171) );
  AND2_X1 U14227 ( .A1(n11172), .A2(n11171), .ZN(n14447) );
  INV_X1 U14228 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n14925) );
  AOI22_X1 U14229 ( .A1(n11150), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n9669), .B2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11173) );
  OAI21_X1 U14230 ( .B1(n11175), .B2(n14925), .A(n11173), .ZN(n13264) );
  NAND2_X1 U14231 ( .A1(n14449), .A2(n13264), .ZN(n13265) );
  INV_X1 U14232 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n20060) );
  AOI22_X1 U14233 ( .A1(n11150), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n9668), .B2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11174) );
  OAI21_X1 U14234 ( .B1(n11175), .B2(n20060), .A(n11174), .ZN(n11176) );
  INV_X1 U14235 ( .A(n11176), .ZN(n11177) );
  INV_X1 U14236 ( .A(n11179), .ZN(n11181) );
  NAND2_X1 U14237 ( .A1(n11181), .A2(n11180), .ZN(n14052) );
  OAI21_X1 U14238 ( .B1(n9666), .B2(n11178), .A(n14052), .ZN(n11182) );
  OR2_X1 U14239 ( .A1(n11185), .A2(n11184), .ZN(n11186) );
  NAND2_X1 U14240 ( .A1(n11187), .A2(n11186), .ZN(n14219) );
  INV_X1 U14241 ( .A(n14219), .ZN(n11194) );
  OR2_X1 U14242 ( .A1(n11286), .A2(n14304), .ZN(n11192) );
  AOI22_X1 U14243 ( .A1(n11188), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11190) );
  NAND2_X1 U14244 ( .A1(n9657), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11189) );
  AND2_X1 U14245 ( .A1(n11190), .A2(n11189), .ZN(n11191) );
  INV_X1 U14246 ( .A(n14218), .ZN(n11193) );
  NAND2_X1 U14247 ( .A1(n11194), .A2(n11193), .ZN(n13772) );
  OR2_X1 U14248 ( .A1(n11286), .A2(n14305), .ZN(n11198) );
  AOI22_X1 U14249 ( .A1(n11188), .A2(P2_EBX_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11196) );
  NAND2_X1 U14250 ( .A1(n9657), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n11195) );
  AND2_X1 U14251 ( .A1(n11196), .A2(n11195), .ZN(n11197) );
  AOI22_X1 U14252 ( .A1(n11188), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11200) );
  NAND2_X1 U14253 ( .A1(n9657), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11199) );
  OAI211_X1 U14254 ( .C1(n11286), .C2(n15695), .A(n11200), .B(n11199), .ZN(
        n13780) );
  OR2_X1 U14255 ( .A1(n11286), .A2(n16514), .ZN(n11204) );
  AOI22_X1 U14256 ( .A1(n11188), .A2(P2_EBX_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11202) );
  NAND2_X1 U14257 ( .A1(n9657), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11201) );
  AND2_X1 U14258 ( .A1(n11202), .A2(n11201), .ZN(n11203) );
  OR2_X1 U14259 ( .A1(n11286), .A2(n11205), .ZN(n11209) );
  AOI22_X1 U14260 ( .A1(n11188), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11207) );
  NAND2_X1 U14261 ( .A1(n9657), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11206) );
  AND2_X1 U14262 ( .A1(n11207), .A2(n11206), .ZN(n11208) );
  NAND2_X1 U14263 ( .A1(n11209), .A2(n11208), .ZN(n15077) );
  INV_X1 U14264 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15691) );
  OR2_X1 U14265 ( .A1(n11286), .A2(n15691), .ZN(n11213) );
  AOI22_X1 U14266 ( .A1(n11188), .A2(P2_EBX_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11211) );
  NAND2_X1 U14267 ( .A1(n9657), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11210) );
  AND2_X1 U14268 ( .A1(n11211), .A2(n11210), .ZN(n11212) );
  OR2_X1 U14269 ( .A1(n11286), .A2(n15674), .ZN(n11217) );
  AOI22_X1 U14270 ( .A1(n11188), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11215) );
  NAND2_X1 U14271 ( .A1(n9657), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11214) );
  AND2_X1 U14272 ( .A1(n11215), .A2(n11214), .ZN(n11216) );
  NAND2_X1 U14273 ( .A1(n11217), .A2(n11216), .ZN(n15048) );
  NAND2_X1 U14274 ( .A1(n15047), .A2(n15048), .ZN(n15049) );
  INV_X1 U14275 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15656) );
  OR2_X1 U14276 ( .A1(n11286), .A2(n15656), .ZN(n11221) );
  AOI22_X1 U14277 ( .A1(n11188), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11219) );
  NAND2_X1 U14278 ( .A1(n9657), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11218) );
  AND2_X1 U14279 ( .A1(n11219), .A2(n11218), .ZN(n11220) );
  OR2_X1 U14280 ( .A1(n11286), .A2(n15635), .ZN(n11225) );
  AOI22_X1 U14281 ( .A1(n11188), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11223) );
  NAND2_X1 U14282 ( .A1(n9657), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n11222) );
  AND2_X1 U14283 ( .A1(n11223), .A2(n11222), .ZN(n11224) );
  NAND2_X1 U14284 ( .A1(n11225), .A2(n11224), .ZN(n15633) );
  OR2_X1 U14285 ( .A1(n11286), .A2(n16392), .ZN(n11229) );
  AOI22_X1 U14286 ( .A1(n11188), .A2(P2_EBX_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11227) );
  NAND2_X1 U14287 ( .A1(n9657), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11226) );
  AND2_X1 U14288 ( .A1(n11227), .A2(n11226), .ZN(n11228) );
  OR2_X1 U14289 ( .A1(n11286), .A2(n11230), .ZN(n11234) );
  AOI22_X1 U14290 ( .A1(n11188), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11232) );
  NAND2_X1 U14291 ( .A1(n9657), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11231) );
  AND2_X1 U14292 ( .A1(n11232), .A2(n11231), .ZN(n11233) );
  NAND2_X1 U14293 ( .A1(n11234), .A2(n11233), .ZN(n15026) );
  OR2_X1 U14294 ( .A1(n11286), .A2(n15589), .ZN(n11238) );
  AOI22_X1 U14295 ( .A1(n11188), .A2(P2_EBX_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11236) );
  NAND2_X1 U14296 ( .A1(n9657), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11235) );
  AND2_X1 U14297 ( .A1(n11236), .A2(n11235), .ZN(n11237) );
  OR2_X1 U14298 ( .A1(n11286), .A2(n11239), .ZN(n11243) );
  NAND2_X1 U14299 ( .A1(n11281), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11241) );
  AOI22_X1 U14300 ( .A1(n11188), .A2(P2_EBX_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11240) );
  AND2_X1 U14301 ( .A1(n11241), .A2(n11240), .ZN(n11242) );
  NAND2_X1 U14302 ( .A1(n11243), .A2(n11242), .ZN(n15008) );
  OR2_X1 U14303 ( .A1(n11286), .A2(n10774), .ZN(n11247) );
  NAND2_X1 U14304 ( .A1(n11281), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11245) );
  AOI22_X1 U14305 ( .A1(n11188), .A2(P2_EBX_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n11244) );
  AND2_X1 U14306 ( .A1(n11245), .A2(n11244), .ZN(n11246) );
  OR2_X1 U14307 ( .A1(n11286), .A2(n15555), .ZN(n11251) );
  NAND2_X1 U14308 ( .A1(n9657), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11249) );
  AOI22_X1 U14309 ( .A1(n11188), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11248) );
  AND2_X1 U14310 ( .A1(n11249), .A2(n11248), .ZN(n11250) );
  NAND2_X1 U14311 ( .A1(n11251), .A2(n11250), .ZN(n14999) );
  OR2_X1 U14312 ( .A1(n11286), .A2(n15549), .ZN(n11253) );
  AOI22_X1 U14313 ( .A1(n11188), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11252) );
  OAI211_X1 U14314 ( .C1(n11296), .C2(n20038), .A(n11253), .B(n11252), .ZN(
        n15182) );
  NAND2_X1 U14315 ( .A1(n11188), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11255) );
  NAND2_X1 U14316 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11254) );
  OAI211_X1 U14317 ( .C1(n11296), .C2(n11256), .A(n11255), .B(n11254), .ZN(
        n11257) );
  AOI21_X1 U14318 ( .B1(n11298), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11257), .ZN(n15334) );
  NAND2_X1 U14319 ( .A1(n11188), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11259) );
  NAND2_X1 U14320 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11258) );
  OAI211_X1 U14321 ( .C1(n11296), .C2(n20041), .A(n11259), .B(n11258), .ZN(
        n11260) );
  AOI21_X1 U14322 ( .B1(n11298), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n11260), .ZN(n15174) );
  NAND2_X1 U14323 ( .A1(n11188), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11262) );
  NAND2_X1 U14324 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11261) );
  OAI211_X1 U14325 ( .C1(n11296), .C2(n11263), .A(n11262), .B(n11261), .ZN(
        n11264) );
  AOI21_X1 U14326 ( .B1(n11298), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n11264), .ZN(n15500) );
  OR2_X1 U14327 ( .A1(n11286), .A2(n15485), .ZN(n11268) );
  NAND2_X1 U14328 ( .A1(n11281), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11266) );
  AOI22_X1 U14329 ( .A1(n11188), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11265) );
  AND2_X1 U14330 ( .A1(n11266), .A2(n11265), .ZN(n11267) );
  NAND2_X1 U14331 ( .A1(n11268), .A2(n11267), .ZN(n14979) );
  OR2_X1 U14332 ( .A1(n11286), .A2(n15474), .ZN(n11272) );
  NAND2_X1 U14333 ( .A1(n9657), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11270) );
  AOI22_X1 U14334 ( .A1(n11188), .A2(P2_EBX_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n11269) );
  AND2_X1 U14335 ( .A1(n11270), .A2(n11269), .ZN(n11271) );
  NAND2_X1 U14336 ( .A1(n11272), .A2(n11271), .ZN(n14968) );
  INV_X1 U14337 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20048) );
  OR2_X1 U14338 ( .A1(n11286), .A2(n15456), .ZN(n11274) );
  AOI22_X1 U14339 ( .A1(n11188), .A2(P2_EBX_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n11273) );
  OAI211_X1 U14340 ( .C1(n11296), .C2(n20048), .A(n11274), .B(n11273), .ZN(
        n14954) );
  NAND2_X1 U14341 ( .A1(n11188), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n11276) );
  NAND2_X1 U14342 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11275) );
  OAI211_X1 U14343 ( .C1(n11296), .C2(n20050), .A(n11276), .B(n11275), .ZN(
        n11277) );
  AOI21_X1 U14344 ( .B1(n11298), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11277), .ZN(n15151) );
  INV_X1 U14345 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20053) );
  NAND2_X1 U14346 ( .A1(n11188), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11279) );
  NAND2_X1 U14347 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11278) );
  OAI211_X1 U14348 ( .C1(n11296), .C2(n20053), .A(n11279), .B(n11278), .ZN(
        n11280) );
  AOI21_X1 U14349 ( .B1(n11298), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11280), .ZN(n13448) );
  OR2_X1 U14350 ( .A1(n11286), .A2(n12341), .ZN(n11285) );
  NAND2_X1 U14351 ( .A1(n9657), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11283) );
  AOI22_X1 U14352 ( .A1(n11188), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11282) );
  AND2_X1 U14353 ( .A1(n11283), .A2(n11282), .ZN(n11284) );
  NAND2_X1 U14354 ( .A1(n11285), .A2(n11284), .ZN(n12346) );
  INV_X1 U14355 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20056) );
  OR2_X1 U14356 ( .A1(n11286), .A2(n15422), .ZN(n11288) );
  AOI22_X1 U14357 ( .A1(n11188), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11287) );
  OAI211_X1 U14358 ( .C1(n11296), .C2(n20056), .A(n11288), .B(n11287), .ZN(
        n12702) );
  NAND2_X1 U14359 ( .A1(n12347), .A2(n12702), .ZN(n12704) );
  INV_X1 U14360 ( .A(n12704), .ZN(n11293) );
  NAND2_X1 U14361 ( .A1(n11188), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11290) );
  NAND2_X1 U14362 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11289) );
  OAI211_X1 U14363 ( .C1(n11296), .C2(n14925), .A(n11290), .B(n11289), .ZN(
        n11291) );
  AOI21_X1 U14364 ( .B1(n11298), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n11291), .ZN(n12379) );
  INV_X1 U14365 ( .A(n12379), .ZN(n11292) );
  NAND2_X1 U14366 ( .A1(n11188), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n11295) );
  NAND2_X1 U14367 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11294) );
  OAI211_X1 U14368 ( .C1(n11296), .C2(n20060), .A(n11295), .B(n11294), .ZN(
        n11297) );
  AOI21_X1 U14369 ( .B1(n11298), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n11297), .ZN(n11299) );
  AND2_X1 U14370 ( .A1(n11300), .A2(n13618), .ZN(n16525) );
  INV_X1 U14371 ( .A(n11301), .ZN(n11302) );
  NAND2_X1 U14372 ( .A1(n13618), .A2(n14054), .ZN(n15575) );
  MUX2_X1 U14373 ( .A(n10917), .B(n11304), .S(n10353), .Z(n11305) );
  INV_X1 U14374 ( .A(n11305), .ZN(n11317) );
  NAND2_X1 U14375 ( .A1(n11306), .A2(n9676), .ZN(n14061) );
  NAND2_X1 U14376 ( .A1(n14061), .A2(n11307), .ZN(n11308) );
  NAND2_X1 U14377 ( .A1(n11308), .A2(n9860), .ZN(n11316) );
  INV_X1 U14378 ( .A(n11318), .ZN(n12700) );
  OAI21_X1 U14379 ( .B1(n11310), .B2(n12700), .A(n11309), .ZN(n11313) );
  NAND2_X1 U14380 ( .A1(n11311), .A2(n12700), .ZN(n13262) );
  OAI21_X1 U14381 ( .B1(n19416), .B2(n11309), .A(n13262), .ZN(n11312) );
  AOI21_X1 U14382 ( .B1(n11314), .B2(n11313), .A(n11312), .ZN(n11315) );
  NAND2_X1 U14383 ( .A1(n14066), .A2(n11318), .ZN(n11319) );
  NAND2_X1 U14384 ( .A1(n13618), .A2(n11319), .ZN(n15581) );
  NAND2_X1 U14385 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14459) );
  NAND2_X1 U14386 ( .A1(n14458), .A2(n14459), .ZN(n14465) );
  INV_X1 U14387 ( .A(n14465), .ZN(n14211) );
  NOR3_X1 U14388 ( .A1(n16534), .A2(n14305), .A3(n14304), .ZN(n15697) );
  NAND2_X1 U14389 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15697), .ZN(
        n16506) );
  NOR4_X1 U14390 ( .A1(n14211), .A2(n16514), .A3(n11205), .A4(n16506), .ZN(
        n11337) );
  OR2_X1 U14391 ( .A1(n16501), .A2(n11337), .ZN(n11326) );
  INV_X1 U14392 ( .A(n13618), .ZN(n11322) );
  NAND2_X1 U14393 ( .A1(n11320), .A2(n13484), .ZN(n20072) );
  NOR2_X1 U14394 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20072), .ZN(n11321) );
  AND2_X2 U14395 ( .A1(n11321), .A2(n14091), .ZN(n19198) );
  NAND2_X1 U14396 ( .A1(n11322), .A2(n19214), .ZN(n15716) );
  NAND2_X1 U14397 ( .A1(n15716), .A2(n15581), .ZN(n11325) );
  INV_X1 U14398 ( .A(n14459), .ZN(n11323) );
  NAND2_X1 U14399 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11323), .ZN(
        n11324) );
  NAND2_X1 U14400 ( .A1(n11325), .A2(n11336), .ZN(n14460) );
  NAND2_X1 U14401 ( .A1(n11326), .A2(n14460), .ZN(n15683) );
  NAND2_X1 U14402 ( .A1(n15608), .A2(n16501), .ZN(n15610) );
  NOR2_X1 U14403 ( .A1(n15656), .A2(n15674), .ZN(n15651) );
  NAND2_X1 U14404 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15651), .ZN(
        n11327) );
  NOR2_X1 U14405 ( .A1(n16493), .A2(n11327), .ZN(n15578) );
  NAND2_X1 U14406 ( .A1(n15578), .A2(n10232), .ZN(n15556) );
  NOR2_X1 U14407 ( .A1(n15556), .A2(n15555), .ZN(n11338) );
  NAND2_X1 U14408 ( .A1(n15608), .A2(n11338), .ZN(n11328) );
  NAND2_X1 U14409 ( .A1(n15610), .A2(n11328), .ZN(n15554) );
  OR2_X1 U14410 ( .A1(n16501), .A2(n11339), .ZN(n11329) );
  AND2_X1 U14411 ( .A1(n15554), .A2(n11329), .ZN(n15520) );
  OAI211_X1 U14412 ( .C1(n11335), .C2(n16501), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n15520), .ZN(n15476) );
  NAND2_X1 U14413 ( .A1(n15476), .A2(n15610), .ZN(n15457) );
  AND2_X1 U14414 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11340) );
  INV_X1 U14415 ( .A(n11340), .ZN(n11330) );
  NAND2_X1 U14416 ( .A1(n15610), .A2(n11330), .ZN(n11331) );
  NAND2_X1 U14417 ( .A1(n15457), .A2(n11331), .ZN(n15442) );
  NAND3_X1 U14418 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15413) );
  AND2_X1 U14419 ( .A1(n15610), .A2(n15413), .ZN(n11332) );
  NOR2_X1 U14420 ( .A1(n15442), .A2(n11332), .ZN(n15414) );
  OAI21_X1 U14421 ( .B1(n16501), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n15414), .ZN(n11333) );
  INV_X1 U14422 ( .A(n11333), .ZN(n11334) );
  OR2_X1 U14423 ( .A1(n11334), .A2(n10970), .ZN(n11346) );
  INV_X1 U14424 ( .A(n11335), .ZN(n15487) );
  NAND2_X1 U14425 ( .A1(n11336), .A2(n15575), .ZN(n14209) );
  NAND2_X1 U14426 ( .A1(n11339), .A2(n15547), .ZN(n15507) );
  NOR2_X1 U14427 ( .A1(n15487), .A2(n15507), .ZN(n15477) );
  NAND2_X1 U14428 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15477), .ZN(
        n15463) );
  INV_X1 U14429 ( .A(n15463), .ZN(n11341) );
  NAND2_X1 U14430 ( .A1(n11341), .A2(n11340), .ZN(n15440) );
  INV_X1 U14431 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11342) );
  NOR4_X1 U14432 ( .A1(n15440), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15413), .A4(n11342), .ZN(n11343) );
  NAND2_X1 U14433 ( .A1(n19198), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n13316) );
  INV_X1 U14434 ( .A(n13316), .ZN(n11344) );
  NOR2_X1 U14435 ( .A1(n11343), .A2(n11344), .ZN(n11345) );
  INV_X1 U14436 ( .A(n11347), .ZN(n11348) );
  OAI211_X1 U14437 ( .C1(n13322), .C2(n16490), .A(n11349), .B(n11348), .ZN(
        P2_U3015) );
  INV_X2 U14438 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11350) );
  AND2_X4 U14439 ( .A1(n11350), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13707) );
  NAND2_X1 U14440 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11354) );
  NAND2_X1 U14441 ( .A1(n11414), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11353) );
  NAND2_X1 U14442 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11352) );
  AND2_X4 U14443 ( .A1(n11366), .A2(n11355), .ZN(n12081) );
  NAND2_X1 U14444 ( .A1(n12081), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11351) );
  AND2_X4 U14445 ( .A1(n13707), .A2(n11355), .ZN(n11570) );
  NAND2_X1 U14446 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11359) );
  AND2_X2 U14447 ( .A1(n11360), .A2(n13702), .ZN(n11408) );
  NAND2_X1 U14448 ( .A1(n11408), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11358) );
  NAND2_X1 U14449 ( .A1(n11569), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11357) );
  AND2_X2 U14450 ( .A1(n11355), .A2(n11365), .ZN(n11428) );
  NAND2_X1 U14451 ( .A1(n11428), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11356) );
  NAND2_X1 U14452 ( .A1(n11480), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11364) );
  NOR2_X4 U14453 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13681) );
  AND2_X2 U14454 ( .A1(n13702), .A2(n13681), .ZN(n11429) );
  NAND2_X1 U14455 ( .A1(n11429), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11363) );
  AND2_X4 U14456 ( .A1(n13707), .A2(n13704), .ZN(n11550) );
  NAND2_X1 U14457 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11362) );
  NAND2_X1 U14458 ( .A1(n12267), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11361) );
  AND2_X2 U14459 ( .A1(n13707), .A2(n13681), .ZN(n11407) );
  NAND2_X1 U14460 ( .A1(n11407), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11370) );
  NAND2_X1 U14461 ( .A1(n11422), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11369) );
  NAND2_X1 U14462 ( .A1(n11430), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11368) );
  NAND2_X1 U14463 ( .A1(n12265), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11367) );
  NAND4_X4 U14464 ( .A1(n11374), .A2(n11373), .A3(n11372), .A4(n11371), .ZN(
        n11494) );
  NAND2_X1 U14465 ( .A1(n12142), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11378) );
  NAND2_X1 U14466 ( .A1(n11569), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11377) );
  NAND2_X1 U14467 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11376) );
  NAND2_X1 U14468 ( .A1(n11428), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11375) );
  NAND2_X1 U14469 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11382) );
  NAND2_X1 U14470 ( .A1(n11399), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11381) );
  NAND2_X1 U14471 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11380) );
  NAND2_X1 U14472 ( .A1(n12265), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11379) );
  NAND2_X1 U14473 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11386) );
  NAND2_X1 U14474 ( .A1(n11414), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11385) );
  NAND2_X1 U14475 ( .A1(n12081), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11384) );
  NAND2_X1 U14476 ( .A1(n12267), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11383) );
  NAND2_X1 U14477 ( .A1(n11408), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11390) );
  NAND2_X1 U14478 ( .A1(n11429), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11389) );
  NAND2_X1 U14479 ( .A1(n11430), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11388) );
  NAND2_X1 U14480 ( .A1(n11422), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11387) );
  INV_X1 U14482 ( .A(n12849), .ZN(n11406) );
  AOI22_X1 U14483 ( .A1(n11569), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11407), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11398) );
  AOI22_X1 U14484 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11428), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U14485 ( .A1(n11408), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11429), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11396) );
  AOI22_X1 U14486 ( .A1(n11430), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11395) );
  NAND4_X1 U14487 ( .A1(n11398), .A2(n11397), .A3(n11396), .A4(n11395), .ZN(
        n11405) );
  BUF_X4 U14488 ( .A(n11399), .Z(n12302) );
  AOI22_X1 U14489 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11403) );
  AOI22_X1 U14490 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11402) );
  AOI22_X1 U14491 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U14492 ( .A1(n11414), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12267), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11400) );
  NAND4_X1 U14493 ( .A1(n11403), .A2(n11402), .A3(n11401), .A4(n11400), .ZN(
        n11404) );
  NAND2_X1 U14494 ( .A1(n11406), .A2(n13629), .ZN(n11421) );
  AOI22_X1 U14495 ( .A1(n11480), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11412) );
  AOI22_X1 U14496 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12267), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11411) );
  AOI22_X1 U14497 ( .A1(n11569), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11407), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11410) );
  AOI22_X1 U14498 ( .A1(n11408), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11430), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11409) );
  AOI22_X1 U14499 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11428), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11417) );
  AOI22_X1 U14500 ( .A1(n11414), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11416) );
  AOI22_X1 U14501 ( .A1(n11429), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11415) );
  AND2_X2 U14502 ( .A1(n10251), .A2(n9715), .ZN(n11504) );
  NAND2_X1 U14504 ( .A1(n11419), .A2(n11563), .ZN(n11420) );
  NAND2_X1 U14505 ( .A1(n11421), .A2(n11420), .ZN(n11451) );
  INV_X2 U14506 ( .A(n11504), .ZN(n13331) );
  AOI22_X1 U14507 ( .A1(n11569), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11570), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11426) );
  AOI22_X1 U14508 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11425) );
  AOI22_X1 U14509 ( .A1(n11408), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11424) );
  AOI22_X1 U14510 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11423) );
  NAND4_X1 U14511 ( .A1(n11426), .A2(n11425), .A3(n11424), .A4(n11423), .ZN(
        n11436) );
  AOI22_X1 U14512 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11413), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11434) );
  INV_X1 U14513 ( .A(n11427), .ZN(n12164) );
  AOI22_X1 U14514 ( .A1(n12164), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11428), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11433) );
  AOI22_X1 U14515 ( .A1(n11429), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11430), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11432) );
  AOI22_X1 U14516 ( .A1(n11414), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12267), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11431) );
  NAND4_X1 U14517 ( .A1(n11434), .A2(n11433), .A3(n11432), .A4(n11431), .ZN(
        n11435) );
  NAND2_X1 U14518 ( .A1(n11508), .A2(n11437), .ZN(n11497) );
  NAND2_X1 U14519 ( .A1(n13821), .A2(n11497), .ZN(n11449) );
  AOI22_X1 U14520 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11441) );
  AOI22_X1 U14521 ( .A1(n11414), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11440) );
  AOI22_X1 U14522 ( .A1(n11429), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11430), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11439) );
  AOI22_X1 U14523 ( .A1(n11407), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11438) );
  NAND4_X1 U14524 ( .A1(n11441), .A2(n11440), .A3(n11439), .A4(n11438), .ZN(
        n11448) );
  AOI22_X1 U14525 ( .A1(n11569), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11570), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11446) );
  AOI22_X1 U14526 ( .A1(n11408), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11428), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11445) );
  AOI22_X1 U14527 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11444) );
  NAND4_X1 U14528 ( .A1(n11446), .A2(n11445), .A3(n11444), .A4(n11443), .ZN(
        n11447) );
  AND2_X2 U14529 ( .A1(n11451), .A2(n11450), .ZN(n12731) );
  INV_X1 U14530 ( .A(n12731), .ZN(n11525) );
  NAND2_X1 U14531 ( .A1(n12142), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11455) );
  NAND2_X1 U14532 ( .A1(n11569), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11454) );
  NAND2_X1 U14533 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11453) );
  NAND2_X1 U14534 ( .A1(n11428), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11452) );
  NAND2_X1 U14535 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11459) );
  NAND2_X1 U14536 ( .A1(n11480), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11458) );
  NAND2_X1 U14537 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11457) );
  NAND2_X1 U14538 ( .A1(n12265), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11456) );
  NAND2_X1 U14539 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11463) );
  NAND2_X1 U14540 ( .A1(n11414), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11462) );
  NAND2_X1 U14541 ( .A1(n12081), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11461) );
  NAND2_X1 U14542 ( .A1(n12267), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11460) );
  NAND2_X1 U14543 ( .A1(n11408), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11467) );
  NAND2_X1 U14544 ( .A1(n11429), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11466) );
  NAND2_X1 U14545 ( .A1(n11430), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11465) );
  NAND2_X1 U14546 ( .A1(n11422), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11464) );
  NAND4_X4 U14547 ( .A1(n11471), .A2(n11470), .A3(n11469), .A4(n11468), .ZN(
        n13918) );
  NAND2_X1 U14548 ( .A1(n11408), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11475) );
  NAND2_X1 U14549 ( .A1(n11414), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11474) );
  NAND2_X1 U14550 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11473) );
  NAND2_X1 U14551 ( .A1(n12265), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11472) );
  INV_X2 U14552 ( .A(n11427), .ZN(n12142) );
  NAND2_X1 U14553 ( .A1(n12142), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11479) );
  NAND2_X1 U14554 ( .A1(n11569), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11478) );
  NAND2_X1 U14555 ( .A1(n11413), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11477) );
  NAND2_X1 U14556 ( .A1(n11429), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11476) );
  NAND2_X1 U14557 ( .A1(n12267), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11483) );
  NAND2_X1 U14558 ( .A1(n12081), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11482) );
  NAND2_X1 U14559 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11481) );
  NAND3_X1 U14560 ( .A1(n11483), .A2(n11482), .A3(n11481), .ZN(n11484) );
  NAND2_X1 U14561 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11488) );
  NAND2_X1 U14562 ( .A1(n11428), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11487) );
  NAND2_X1 U14563 ( .A1(n11430), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11486) );
  NAND2_X1 U14564 ( .A1(n11422), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11485) );
  NAND2_X1 U14565 ( .A1(n20326), .A2(n13918), .ZN(n14009) );
  OR2_X1 U14566 ( .A1(n14009), .A2(n20347), .ZN(n11493) );
  NAND2_X1 U14567 ( .A1(n20316), .A2(n13943), .ZN(n13959) );
  NAND2_X1 U14568 ( .A1(n11510), .A2(n13331), .ZN(n11495) );
  AND2_X1 U14569 ( .A1(n11495), .A2(n11508), .ZN(n11529) );
  INV_X1 U14571 ( .A(n11506), .ZN(n11500) );
  INV_X1 U14572 ( .A(n11588), .ZN(n20339) );
  NAND2_X1 U14573 ( .A1(n20339), .A2(n13918), .ZN(n12742) );
  NAND2_X1 U14574 ( .A1(n11500), .A2(n14486), .ZN(n12852) );
  NAND4_X1 U14575 ( .A1(n11501), .A2(n11528), .A3(n11523), .A4(n12852), .ZN(
        n11502) );
  NAND2_X1 U14576 ( .A1(n11502), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11515) );
  NAND2_X2 U14577 ( .A1(n20326), .A2(n20316), .ZN(n11526) );
  NOR2_X1 U14578 ( .A1(n11526), .A2(n12849), .ZN(n11503) );
  NAND2_X1 U14579 ( .A1(n12731), .A2(n11503), .ZN(n13325) );
  NAND2_X1 U14580 ( .A1(n11509), .A2(n13918), .ZN(n14471) );
  XNOR2_X1 U14581 ( .A(n20896), .B(P1_STATE_REG_2__SCAN_IN), .ZN(n12714) );
  NAND2_X1 U14582 ( .A1(n13501), .A2(n12714), .ZN(n11513) );
  NAND2_X1 U14583 ( .A1(n9793), .A2(n11512), .ZN(n13330) );
  OR2_X2 U14584 ( .A1(n13330), .A2(n13821), .ZN(n12846) );
  NAND3_X1 U14585 ( .A1(n12739), .A2(n11513), .A3(n12846), .ZN(n11514) );
  NAND2_X1 U14586 ( .A1(n11514), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11520) );
  INV_X1 U14587 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n11516) );
  NAND2_X1 U14588 ( .A1(n11516), .A2(n16292), .ZN(n20958) );
  INV_X1 U14589 ( .A(n12324), .ZN(n11517) );
  NAND2_X1 U14590 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11601) );
  OAI21_X1 U14591 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n11601), .ZN(n20635) );
  NAND2_X1 U14592 ( .A1(n15913), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11595) );
  OAI21_X1 U14593 ( .B1(n11517), .B2(n20635), .A(n11595), .ZN(n11518) );
  INV_X1 U14594 ( .A(n11518), .ZN(n11519) );
  MUX2_X1 U14595 ( .A(n15913), .B(n12324), .S(n20751), .Z(n11521) );
  INV_X1 U14596 ( .A(n11521), .ZN(n11522) );
  INV_X1 U14597 ( .A(n11523), .ZN(n11524) );
  NAND2_X1 U14598 ( .A1(n11524), .A2(n13943), .ZN(n11536) );
  AND2_X1 U14599 ( .A1(n13629), .A2(n13918), .ZN(n11527) );
  OAI21_X1 U14600 ( .B1(n11529), .B2(n14009), .A(n11528), .ZN(n11534) );
  AND2_X1 U14601 ( .A1(n11526), .A2(n12864), .ZN(n13507) );
  NAND2_X1 U14602 ( .A1(n13507), .A2(n11530), .ZN(n11532) );
  INV_X1 U14603 ( .A(n20958), .ZN(n13718) );
  NAND2_X1 U14604 ( .A1(n11511), .A2(n11531), .ZN(n12860) );
  NAND4_X1 U14605 ( .A1(n11532), .A2(n13718), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .A4(n12860), .ZN(n11533) );
  NOR2_X1 U14606 ( .A1(n11534), .A2(n11533), .ZN(n11535) );
  INV_X1 U14607 ( .A(n11568), .ZN(n11537) );
  NAND2_X1 U14608 ( .A1(n11539), .A2(n11538), .ZN(n20753) );
  AOI22_X1 U14609 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12303), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11543) );
  AOI22_X1 U14610 ( .A1(n11480), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12120), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11542) );
  INV_X1 U14611 ( .A(n11550), .ZN(n11672) );
  AOI22_X1 U14612 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11541) );
  AOI22_X1 U14613 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11540) );
  NAND4_X1 U14614 ( .A1(n11543), .A2(n11542), .A3(n11541), .A4(n11540), .ZN(
        n11549) );
  AOI22_X1 U14615 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12142), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11547) );
  AOI22_X1 U14616 ( .A1(n11429), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11546) );
  BUF_X1 U14617 ( .A(n11612), .Z(n11551) );
  AOI22_X1 U14618 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11545) );
  AOI22_X1 U14619 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12267), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11544) );
  NAND4_X1 U14620 ( .A1(n11547), .A2(n11546), .A3(n11545), .A4(n11544), .ZN(
        n11548) );
  INV_X1 U14621 ( .A(n11562), .ZN(n11625) );
  AOI22_X1 U14622 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12266), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11555) );
  AOI22_X1 U14623 ( .A1(n12120), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11554) );
  AOI22_X1 U14624 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11553) );
  AOI22_X1 U14625 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11552) );
  NAND4_X1 U14626 ( .A1(n11555), .A2(n11554), .A3(n11553), .A4(n11552), .ZN(
        n11561) );
  AOI22_X1 U14627 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12142), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11559) );
  AOI22_X1 U14628 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11558) );
  AOI22_X1 U14629 ( .A1(n11480), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U14630 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12267), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11556) );
  NAND4_X1 U14631 ( .A1(n11559), .A2(n11558), .A3(n11557), .A4(n11556), .ZN(
        n11560) );
  NAND2_X1 U14632 ( .A1(n11589), .A2(n11562), .ZN(n11665) );
  OAI21_X1 U14633 ( .B1(n11562), .B2(n11589), .A(n11665), .ZN(n11564) );
  OAI211_X1 U14634 ( .C1(n11564), .C2(n14009), .A(n11563), .B(n11494), .ZN(
        n11565) );
  INV_X1 U14635 ( .A(n11565), .ZN(n11566) );
  NAND2_X1 U14636 ( .A1(n11567), .A2(n11566), .ZN(n11592) );
  AOI22_X1 U14637 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11574) );
  AOI22_X1 U14638 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12295), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11573) );
  AOI22_X1 U14639 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12303), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11572) );
  AOI22_X1 U14640 ( .A1(n12206), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11571) );
  NAND4_X1 U14641 ( .A1(n11574), .A2(n11573), .A3(n11572), .A4(n11571), .ZN(
        n11580) );
  AOI22_X1 U14642 ( .A1(n12266), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12120), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U14643 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11577) );
  AOI22_X1 U14644 ( .A1(n11408), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11576) );
  AOI22_X1 U14645 ( .A1(n12081), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11575) );
  NAND4_X1 U14646 ( .A1(n11578), .A2(n11577), .A3(n11576), .A4(n11575), .ZN(
        n11579) );
  NOR2_X1 U14647 ( .A1(n11649), .A2(n11747), .ZN(n11624) );
  NAND2_X1 U14648 ( .A1(n11624), .A2(n11589), .ZN(n11581) );
  NAND2_X1 U14649 ( .A1(n11813), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11583) );
  AOI21_X1 U14650 ( .B1(n20316), .B2(n11589), .A(n20971), .ZN(n11582) );
  OAI211_X1 U14651 ( .C1(n11585), .C2(n12845), .A(n11583), .B(n11582), .ZN(
        n11623) );
  INV_X1 U14652 ( .A(n11623), .ZN(n11584) );
  INV_X1 U14653 ( .A(n11744), .ZN(n11587) );
  INV_X1 U14654 ( .A(n11589), .ZN(n11586) );
  INV_X1 U14655 ( .A(n11773), .ZN(n11743) );
  NAND2_X1 U14656 ( .A1(n20316), .A2(n11588), .ZN(n11637) );
  OAI21_X1 U14657 ( .B1(n14009), .B2(n11589), .A(n11637), .ZN(n11590) );
  INV_X1 U14658 ( .A(n11590), .ZN(n11591) );
  NAND2_X1 U14659 ( .A1(n13665), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13664) );
  NAND2_X1 U14660 ( .A1(n20246), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20245) );
  INV_X1 U14661 ( .A(n11592), .ZN(n11593) );
  OR2_X1 U14662 ( .A1(n13664), .A2(n11593), .ZN(n11594) );
  INV_X1 U14663 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20282) );
  XNOR2_X1 U14664 ( .A(n11642), .B(n20282), .ZN(n13790) );
  NAND2_X1 U14665 ( .A1(n11595), .A2(n10010), .ZN(n11596) );
  NAND2_X1 U14666 ( .A1(n11597), .A2(n11596), .ZN(n11605) );
  AND2_X1 U14667 ( .A1(n15913), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11599) );
  INV_X1 U14668 ( .A(n11601), .ZN(n11600) );
  NAND2_X1 U14669 ( .A1(n11600), .A2(n11776), .ZN(n20666) );
  NAND2_X1 U14670 ( .A1(n11601), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11602) );
  NAND2_X1 U14671 ( .A1(n20666), .A2(n11602), .ZN(n20318) );
  NAND2_X1 U14672 ( .A1(n12324), .A2(n20318), .ZN(n11604) );
  NAND2_X1 U14673 ( .A1(n11606), .A2(n11604), .ZN(n11603) );
  AOI22_X1 U14674 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11611) );
  AOI22_X1 U14675 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11428), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11610) );
  AOI22_X1 U14676 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12266), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11609) );
  AOI22_X1 U14677 ( .A1(n12206), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11608) );
  NAND4_X1 U14678 ( .A1(n11611), .A2(n11610), .A3(n11609), .A4(n11608), .ZN(
        n11618) );
  AOI22_X1 U14679 ( .A1(n11480), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11616) );
  AOI22_X1 U14680 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11615) );
  AOI22_X1 U14681 ( .A1(n12120), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11614) );
  AOI22_X1 U14682 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12267), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11613) );
  NAND4_X1 U14683 ( .A1(n11616), .A2(n11615), .A3(n11614), .A4(n11613), .ZN(
        n11617) );
  INV_X1 U14684 ( .A(n11648), .ZN(n11620) );
  AOI22_X1 U14685 ( .A1(n11620), .A2(n11619), .B1(n11813), .B2(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11621) );
  XNOR2_X1 U14686 ( .A(n11622), .B(n11621), .ZN(n11633) );
  INV_X1 U14687 ( .A(n11624), .ZN(n11628) );
  NAND2_X1 U14688 ( .A1(n11813), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11627) );
  OR2_X1 U14689 ( .A1(n11648), .A2(n11625), .ZN(n11626) );
  XNOR2_X2 U14690 ( .A(n11629), .B(n11630), .ZN(n11832) );
  INV_X1 U14691 ( .A(n11630), .ZN(n11631) );
  AND2_X2 U14692 ( .A1(n11633), .A2(n11634), .ZN(n11662) );
  OR2_X1 U14693 ( .A1(n11830), .A2(n11743), .ZN(n11641) );
  XNOR2_X1 U14694 ( .A(n11665), .B(n11664), .ZN(n11639) );
  INV_X1 U14695 ( .A(n14009), .ZN(n20969) );
  INV_X1 U14696 ( .A(n11637), .ZN(n11638) );
  AOI21_X1 U14697 ( .B1(n11639), .B2(n20969), .A(n11638), .ZN(n11640) );
  NAND2_X1 U14698 ( .A1(n11641), .A2(n11640), .ZN(n13789) );
  NAND2_X1 U14699 ( .A1(n11642), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11643) );
  INV_X1 U14700 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n11644) );
  NAND2_X1 U14701 ( .A1(n11598), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11647) );
  NAND3_X1 U14702 ( .A1(n20710), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20551) );
  INV_X1 U14703 ( .A(n20571), .ZN(n11645) );
  NAND3_X1 U14704 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20825) );
  AOI21_X1 U14705 ( .B1(n20710), .B2(n11645), .A(n20873), .ZN(n20579) );
  AOI22_X1 U14706 ( .A1(n12324), .A2(n20579), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15913), .ZN(n11646) );
  XNOR2_X1 U14707 ( .A(n13638), .B(n20469), .ZN(n20578) );
  NAND2_X1 U14708 ( .A1(n20578), .A2(n20971), .ZN(n11661) );
  AOI22_X1 U14709 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11653) );
  AOI22_X1 U14710 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11428), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11652) );
  AOI22_X1 U14711 ( .A1(n11408), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12266), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11651) );
  AOI22_X1 U14712 ( .A1(n12206), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11650) );
  NAND4_X1 U14713 ( .A1(n11653), .A2(n11652), .A3(n11651), .A4(n11650), .ZN(
        n11659) );
  AOI22_X1 U14714 ( .A1(n11480), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U14715 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11656) );
  AOI22_X1 U14716 ( .A1(n12120), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11655) );
  INV_X1 U14717 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n20344) );
  AOI22_X1 U14718 ( .A1(n11414), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12267), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11654) );
  NAND4_X1 U14719 ( .A1(n11657), .A2(n11656), .A3(n11655), .A4(n11654), .ZN(
        n11658) );
  AOI22_X1 U14720 ( .A1(n11792), .A2(n11702), .B1(n11813), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11660) );
  NAND2_X1 U14721 ( .A1(n11665), .A2(n11664), .ZN(n11704) );
  INV_X1 U14722 ( .A(n11702), .ZN(n11666) );
  XNOR2_X1 U14723 ( .A(n11704), .B(n11666), .ZN(n11667) );
  NAND2_X1 U14724 ( .A1(n11667), .A2(n20969), .ZN(n11668) );
  NAND2_X1 U14725 ( .A1(n11669), .A2(n11668), .ZN(n13894) );
  NAND2_X1 U14726 ( .A1(n11670), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11671) );
  AOI22_X1 U14727 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11428), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U14728 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12302), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11675) );
  AOI22_X1 U14729 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12295), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11674) );
  AOI22_X1 U14730 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11673) );
  NAND4_X1 U14731 ( .A1(n11676), .A2(n11675), .A3(n11674), .A4(n11673), .ZN(
        n11682) );
  AOI22_X1 U14732 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11680) );
  AOI22_X1 U14733 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11429), .B1(
        n12120), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U14734 ( .A1(n12206), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U14735 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12267), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11677) );
  NAND4_X1 U14736 ( .A1(n11680), .A2(n11679), .A3(n11678), .A4(n11677), .ZN(
        n11681) );
  AOI22_X1 U14737 ( .A1(n11792), .A2(n11701), .B1(
        P1_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n11813), .ZN(n11683) );
  NAND2_X1 U14738 ( .A1(n11711), .A2(n11684), .ZN(n11859) );
  OR2_X1 U14739 ( .A1(n11859), .A2(n11743), .ZN(n11688) );
  NAND2_X1 U14740 ( .A1(n11704), .A2(n11702), .ZN(n11685) );
  XNOR2_X1 U14741 ( .A(n11685), .B(n11701), .ZN(n11686) );
  NAND2_X1 U14742 ( .A1(n11686), .A2(n20969), .ZN(n11687) );
  NAND2_X1 U14743 ( .A1(n11688), .A2(n11687), .ZN(n11689) );
  INV_X1 U14744 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12761) );
  XNOR2_X1 U14745 ( .A(n11689), .B(n12761), .ZN(n20236) );
  NAND2_X1 U14746 ( .A1(n20237), .A2(n20236), .ZN(n20235) );
  NAND2_X1 U14747 ( .A1(n11689), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11690) );
  NAND2_X1 U14748 ( .A1(n20235), .A2(n11690), .ZN(n16134) );
  AOI22_X1 U14749 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12142), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U14750 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11428), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U14751 ( .A1(n11408), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12266), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11692) );
  AOI22_X1 U14752 ( .A1(n12206), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11691) );
  NAND4_X1 U14753 ( .A1(n11694), .A2(n11693), .A3(n11692), .A4(n11691), .ZN(
        n11700) );
  AOI22_X1 U14754 ( .A1(n11480), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U14755 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11697) );
  AOI22_X1 U14756 ( .A1(n12120), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11696) );
  INV_X1 U14757 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20358) );
  AOI22_X1 U14758 ( .A1(n11414), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12267), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11695) );
  NAND4_X1 U14759 ( .A1(n11698), .A2(n11697), .A3(n11696), .A4(n11695), .ZN(
        n11699) );
  AOI22_X1 U14760 ( .A1(n11792), .A2(n11726), .B1(n11813), .B2(
        P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11712) );
  XNOR2_X1 U14761 ( .A(n11711), .B(n9986), .ZN(n11875) );
  NAND2_X1 U14762 ( .A1(n11875), .A2(n11773), .ZN(n11708) );
  AND2_X1 U14763 ( .A1(n11702), .A2(n11701), .ZN(n11703) );
  AND2_X1 U14764 ( .A1(n11704), .A2(n11703), .ZN(n11727) );
  INV_X1 U14765 ( .A(n11726), .ZN(n11705) );
  XNOR2_X1 U14766 ( .A(n11727), .B(n11705), .ZN(n11706) );
  NAND2_X1 U14767 ( .A1(n11706), .A2(n20969), .ZN(n11707) );
  NAND2_X1 U14768 ( .A1(n11708), .A2(n11707), .ZN(n11709) );
  INV_X1 U14769 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12872) );
  NAND2_X1 U14770 ( .A1(n11709), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11710) );
  AOI22_X1 U14771 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12142), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11716) );
  AOI22_X1 U14772 ( .A1(n12120), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U14773 ( .A1(n11414), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11714) );
  AOI22_X1 U14774 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11713) );
  NAND4_X1 U14775 ( .A1(n11716), .A2(n11715), .A3(n11714), .A4(n11713), .ZN(
        n11722) );
  AOI22_X1 U14776 ( .A1(n11408), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12266), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11720) );
  AOI22_X1 U14777 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11719) );
  AOI22_X1 U14778 ( .A1(n11480), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11718) );
  AOI22_X1 U14779 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12267), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11717) );
  NAND4_X1 U14780 ( .A1(n11720), .A2(n11719), .A3(n11718), .A4(n11717), .ZN(
        n11721) );
  AOI22_X1 U14781 ( .A1(n11792), .A2(n11735), .B1(n11813), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11724) );
  NAND2_X1 U14782 ( .A1(n11725), .A2(n11724), .ZN(n11884) );
  NAND2_X1 U14783 ( .A1(n11727), .A2(n11726), .ZN(n11736) );
  XNOR2_X1 U14784 ( .A(n11735), .B(n11736), .ZN(n11728) );
  NAND2_X1 U14785 ( .A1(n20969), .A2(n11728), .ZN(n11729) );
  INV_X1 U14786 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16126) );
  NAND2_X1 U14787 ( .A1(n11792), .A2(n11747), .ZN(n11732) );
  NAND2_X1 U14788 ( .A1(n11813), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11731) );
  NAND2_X1 U14789 ( .A1(n11732), .A2(n11731), .ZN(n11733) );
  INV_X1 U14790 ( .A(n11735), .ZN(n11737) );
  NOR2_X1 U14791 ( .A1(n11737), .A2(n11736), .ZN(n11746) );
  XNOR2_X1 U14792 ( .A(n11747), .B(n11746), .ZN(n11738) );
  NOR2_X1 U14793 ( .A1(n11738), .A2(n14009), .ZN(n11739) );
  AOI21_X1 U14794 ( .B1(n11885), .B2(n11773), .A(n11739), .ZN(n11741) );
  INV_X1 U14795 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11740) );
  NAND2_X1 U14796 ( .A1(n11741), .A2(n11740), .ZN(n16120) );
  INV_X1 U14797 ( .A(n11741), .ZN(n11742) );
  NAND2_X1 U14798 ( .A1(n11742), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16119) );
  NOR2_X1 U14799 ( .A1(n11744), .A2(n11743), .ZN(n11745) );
  NAND2_X1 U14800 ( .A1(n11747), .A2(n11746), .ZN(n11748) );
  INV_X1 U14801 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n14332) );
  NAND2_X1 U14802 ( .A1(n14333), .A2(n14332), .ZN(n11749) );
  NAND2_X1 U14803 ( .A1(n11750), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11751) );
  NAND2_X1 U14804 ( .A1(n16110), .A2(n16241), .ZN(n11753) );
  AND2_X1 U14805 ( .A1(n16086), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11754) );
  NOR2_X1 U14806 ( .A1(n14792), .A2(n11754), .ZN(n16092) );
  NAND2_X1 U14807 ( .A1(n16086), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11755) );
  NAND2_X1 U14808 ( .A1(n16092), .A2(n11755), .ZN(n16082) );
  NOR2_X1 U14809 ( .A1(n16086), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16102) );
  AND2_X1 U14810 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11756) );
  NOR2_X1 U14811 ( .A1(n16086), .A2(n11756), .ZN(n14801) );
  INV_X1 U14812 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16213) );
  XNOR2_X1 U14813 ( .A(n16086), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14784) );
  INV_X1 U14814 ( .A(n14784), .ZN(n11758) );
  INV_X1 U14815 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16202) );
  NAND2_X1 U14816 ( .A1(n16110), .A2(n16202), .ZN(n16095) );
  NAND2_X1 U14817 ( .A1(n16086), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14804) );
  INV_X1 U14818 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16240) );
  INV_X1 U14819 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16113) );
  NAND2_X1 U14820 ( .A1(n16240), .A2(n16113), .ZN(n11760) );
  NAND2_X1 U14821 ( .A1(n16086), .A2(n11760), .ZN(n14802) );
  OAI21_X1 U14822 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n16086), .ZN(n11761) );
  NAND2_X1 U14823 ( .A1(n14791), .A2(n11761), .ZN(n11762) );
  INV_X1 U14824 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16174) );
  XNOR2_X1 U14825 ( .A(n16086), .B(n16174), .ZN(n14777) );
  INV_X1 U14826 ( .A(n14768), .ZN(n11764) );
  NAND2_X1 U14827 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15931) );
  INV_X1 U14828 ( .A(n15931), .ZN(n11763) );
  NAND2_X1 U14829 ( .A1(n11764), .A2(n10230), .ZN(n11765) );
  INV_X1 U14830 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11766) );
  INV_X1 U14831 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14893) );
  NAND3_X1 U14832 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14735) );
  INV_X1 U14833 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14870) );
  INV_X1 U14834 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14882) );
  NAND2_X1 U14835 ( .A1(n14870), .A2(n14882), .ZN(n12708) );
  NAND2_X1 U14836 ( .A1(n11767), .A2(n16086), .ZN(n14738) );
  AND2_X1 U14837 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14846) );
  NAND2_X1 U14838 ( .A1(n16110), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11768) );
  INV_X1 U14839 ( .A(n12387), .ZN(n11769) );
  NOR2_X1 U14840 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12887) );
  INV_X1 U14841 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14845) );
  NAND2_X1 U14842 ( .A1(n14717), .A2(n14845), .ZN(n12389) );
  NAND2_X1 U14843 ( .A1(n11769), .A2(n12389), .ZN(n11770) );
  NAND2_X1 U14844 ( .A1(n15877), .A2(n20316), .ZN(n11772) );
  NAND3_X1 U14845 ( .A1(n11771), .A2(n11506), .A3(n11772), .ZN(n12728) );
  NOR2_X1 U14846 ( .A1(n12728), .A2(n12849), .ZN(n12736) );
  XNOR2_X1 U14847 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11786) );
  NAND2_X1 U14848 ( .A1(n20751), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11790) );
  NAND2_X1 U14849 ( .A1(n11786), .A2(n11787), .ZN(n11775) );
  NAND2_X1 U14850 ( .A1(n20638), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11774) );
  NAND2_X1 U14851 ( .A1(n11775), .A2(n11774), .ZN(n11800) );
  MUX2_X1 U14852 ( .A(n11776), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n11799) );
  NAND2_X1 U14853 ( .A1(n11800), .A2(n11799), .ZN(n11778) );
  NAND2_X1 U14854 ( .A1(n11776), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11777) );
  XNOR2_X1 U14855 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11784) );
  NOR2_X1 U14856 ( .A1(n13845), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11779) );
  NAND2_X1 U14857 ( .A1(n20303), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11780) );
  NOR2_X1 U14858 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20303), .ZN(
        n11782) );
  INV_X1 U14859 ( .A(n12723), .ZN(n11781) );
  NAND2_X1 U14860 ( .A1(n12723), .A2(n11792), .ZN(n11821) );
  NAND2_X1 U14861 ( .A1(n11798), .A2(n13943), .ZN(n11818) );
  NAND2_X1 U14862 ( .A1(n11813), .A2(n12721), .ZN(n11817) );
  INV_X1 U14863 ( .A(n11813), .ZN(n11809) );
  XNOR2_X1 U14864 ( .A(n11785), .B(n11784), .ZN(n12720) );
  XNOR2_X1 U14865 ( .A(n11787), .B(n11786), .ZN(n12719) );
  INV_X1 U14866 ( .A(n11798), .ZN(n11788) );
  NOR2_X1 U14867 ( .A1(n12719), .A2(n11788), .ZN(n11796) );
  NAND2_X1 U14868 ( .A1(n11510), .A2(n13918), .ZN(n11789) );
  NAND2_X1 U14869 ( .A1(n11789), .A2(n20326), .ZN(n11805) );
  OAI21_X1 U14870 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20751), .A(
        n11790), .ZN(n11793) );
  INV_X1 U14871 ( .A(n11793), .ZN(n11791) );
  OAI211_X1 U14872 ( .C1(n20316), .C2(n12849), .A(n11805), .B(n11791), .ZN(
        n11795) );
  OAI21_X1 U14873 ( .B1(n11806), .B2(n11793), .A(n11810), .ZN(n11794) );
  NAND2_X1 U14874 ( .A1(n11795), .A2(n11794), .ZN(n11797) );
  NAND2_X1 U14875 ( .A1(n11796), .A2(n11797), .ZN(n11804) );
  OAI211_X1 U14876 ( .C1(n11798), .C2(n11797), .A(n12719), .B(n11818), .ZN(
        n11803) );
  XNOR2_X1 U14877 ( .A(n11800), .B(n11799), .ZN(n12718) );
  NAND2_X1 U14878 ( .A1(n11813), .A2(n12718), .ZN(n11801) );
  OAI211_X1 U14879 ( .C1(n11806), .C2(n12718), .A(n11801), .B(n11805), .ZN(
        n11802) );
  NAND3_X1 U14880 ( .A1(n11804), .A2(n11803), .A3(n11802), .ZN(n11808) );
  AOI22_X1 U14881 ( .A1(n11809), .A2(n12720), .B1(n11808), .B2(n11807), .ZN(
        n11815) );
  INV_X1 U14882 ( .A(n12720), .ZN(n11811) );
  NOR2_X1 U14883 ( .A1(n11811), .A2(n11810), .ZN(n11814) );
  INV_X1 U14884 ( .A(n12721), .ZN(n11812) );
  OAI22_X1 U14885 ( .A1(n11815), .A2(n11814), .B1(n11813), .B2(n11812), .ZN(
        n11816) );
  OAI21_X1 U14886 ( .B1(n11818), .B2(n11817), .A(n11816), .ZN(n11819) );
  AOI21_X1 U14887 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20971), .A(
        n11819), .ZN(n11820) );
  NAND2_X1 U14888 ( .A1(n11821), .A2(n11820), .ZN(n11822) );
  INV_X2 U14889 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20968) );
  NOR2_X2 U14890 ( .A1(n14479), .A2(n20968), .ZN(n11843) );
  INV_X1 U14891 ( .A(n11893), .ZN(n12282) );
  XNOR2_X1 U14892 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13785) );
  NOR2_X1 U14893 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11824) );
  INV_X1 U14894 ( .A(n12315), .ZN(n12289) );
  NAND2_X1 U14895 ( .A1(n13785), .A2(n12289), .ZN(n11825) );
  NAND2_X1 U14896 ( .A1(n20968), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12321) );
  NAND2_X1 U14897 ( .A1(n11825), .A2(n12321), .ZN(n11826) );
  AOI21_X1 U14898 ( .B1(n12282), .B2(P1_EAX_REG_2__SCAN_IN), .A(n11826), .ZN(
        n11827) );
  INV_X1 U14899 ( .A(n11827), .ZN(n11828) );
  NOR2_X1 U14900 ( .A1(n13821), .A2(n20968), .ZN(n11842) );
  INV_X1 U14901 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13787) );
  OR2_X1 U14902 ( .A1(n12321), .A2(n13787), .ZN(n11848) );
  NAND2_X1 U14903 ( .A1(n13866), .A2(n11967), .ZN(n11837) );
  NAND2_X1 U14904 ( .A1(n11842), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11835) );
  AOI22_X1 U14905 ( .A1(n12282), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20968), .ZN(n11834) );
  AND2_X1 U14906 ( .A1(n11835), .A2(n11834), .ZN(n11836) );
  NAND2_X1 U14907 ( .A1(n11837), .A2(n11836), .ZN(n13828) );
  NAND2_X1 U14908 ( .A1(n11838), .A2(n11531), .ZN(n11839) );
  NAND2_X1 U14909 ( .A1(n11839), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13658) );
  INV_X1 U14911 ( .A(n11842), .ZN(n11864) );
  AOI22_X1 U14912 ( .A1(n11843), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20968), .ZN(n11844) );
  OAI21_X1 U14913 ( .B1(n9963), .B2(n11864), .A(n11844), .ZN(n11845) );
  AOI21_X1 U14914 ( .B1(n11841), .B2(n11967), .A(n11845), .ZN(n13659) );
  OR2_X1 U14915 ( .A1(n13658), .A2(n13659), .ZN(n13660) );
  NAND2_X1 U14916 ( .A1(n13659), .A2(n12289), .ZN(n11846) );
  NAND2_X1 U14917 ( .A1(n13660), .A2(n11846), .ZN(n13827) );
  NAND2_X1 U14918 ( .A1(n13828), .A2(n13827), .ZN(n13826) );
  INV_X1 U14919 ( .A(n13826), .ZN(n11847) );
  NAND2_X1 U14920 ( .A1(n10216), .A2(n11847), .ZN(n13784) );
  NAND2_X2 U14921 ( .A1(n13784), .A2(n11848), .ZN(n13841) );
  INV_X1 U14922 ( .A(n20305), .ZN(n11849) );
  NAND2_X1 U14923 ( .A1(n11849), .A2(n11967), .ZN(n11858) );
  INV_X1 U14924 ( .A(n11851), .ZN(n11853) );
  INV_X1 U14925 ( .A(n11861), .ZN(n11852) );
  OAI21_X1 U14926 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11853), .A(
        n11852), .ZN(n13973) );
  AOI22_X1 U14927 ( .A1(n12392), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n12289), .B2(n13973), .ZN(n11855) );
  NAND2_X1 U14928 ( .A1(n12282), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11854) );
  OAI211_X1 U14929 ( .C1(n11864), .C2(n13845), .A(n11855), .B(n11854), .ZN(
        n11856) );
  INV_X1 U14930 ( .A(n11856), .ZN(n11857) );
  NAND2_X1 U14931 ( .A1(n11858), .A2(n11857), .ZN(n13840) );
  INV_X1 U14932 ( .A(n11859), .ZN(n11860) );
  OAI21_X1 U14933 ( .B1(n11861), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n11869), .ZN(n20242) );
  INV_X1 U14934 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13642) );
  INV_X1 U14935 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21106) );
  OAI21_X1 U14936 ( .B1(n21106), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20968), .ZN(n11863) );
  NAND2_X1 U14937 ( .A1(n12282), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11862) );
  OAI211_X1 U14938 ( .C1(n11864), .C2(n13642), .A(n11863), .B(n11862), .ZN(
        n11865) );
  OAI21_X1 U14939 ( .B1(n20242), .B2(n12315), .A(n11865), .ZN(n11866) );
  INV_X1 U14940 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n11873) );
  INV_X1 U14941 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11868) );
  NAND2_X1 U14942 ( .A1(n11869), .A2(n11868), .ZN(n11871) );
  NAND2_X1 U14943 ( .A1(n11871), .A2(n11879), .ZN(n20170) );
  AOI22_X1 U14944 ( .A1(n20170), .A2(n12289), .B1(n12392), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11872) );
  OAI21_X1 U14945 ( .B1(n11893), .B2(n11873), .A(n11872), .ZN(n11874) );
  NAND2_X1 U14946 ( .A1(n11877), .A2(n11876), .ZN(n13930) );
  INV_X1 U14947 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n20220) );
  INV_X1 U14948 ( .A(n11886), .ZN(n11887) );
  INV_X1 U14949 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11880) );
  NAND2_X1 U14950 ( .A1(n11880), .A2(n11879), .ZN(n11881) );
  NAND2_X1 U14951 ( .A1(n11887), .A2(n11881), .ZN(n20158) );
  AOI22_X1 U14952 ( .A1(n20158), .A2(n11824), .B1(n12392), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11882) );
  OAI21_X1 U14953 ( .B1(n11893), .B2(n20220), .A(n11882), .ZN(n11883) );
  NOR2_X2 U14954 ( .A1(n13930), .A2(n13996), .ZN(n13994) );
  INV_X1 U14955 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11892) );
  NAND2_X1 U14956 ( .A1(n11885), .A2(n11967), .ZN(n11891) );
  INV_X1 U14957 ( .A(n11907), .ZN(n11889) );
  INV_X1 U14958 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20142) );
  NAND2_X1 U14959 ( .A1(n11887), .A2(n20142), .ZN(n11888) );
  NAND2_X1 U14960 ( .A1(n11889), .A2(n11888), .ZN(n20156) );
  AOI22_X1 U14961 ( .A1(n20156), .A2(n11824), .B1(n12392), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11890) );
  NAND2_X1 U14962 ( .A1(n13994), .A2(n14005), .ZN(n14003) );
  AOI22_X1 U14963 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11897) );
  BUF_X1 U14964 ( .A(n11408), .Z(n12301) );
  AOI22_X1 U14965 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11570), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11896) );
  AOI22_X1 U14966 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11895) );
  AOI22_X1 U14967 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11894) );
  NAND4_X1 U14968 ( .A1(n11897), .A2(n11896), .A3(n11895), .A4(n11894), .ZN(
        n11903) );
  AOI22_X1 U14969 ( .A1(n12120), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11901) );
  AOI22_X1 U14970 ( .A1(n12266), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11900) );
  AOI22_X1 U14971 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11899) );
  AOI22_X1 U14972 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11898) );
  NAND4_X1 U14973 ( .A1(n11901), .A2(n11900), .A3(n11899), .A4(n11898), .ZN(
        n11902) );
  OAI21_X1 U14974 ( .B1(n11903), .B2(n11902), .A(n11967), .ZN(n11906) );
  XNOR2_X1 U14975 ( .A(n11907), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14336) );
  AOI22_X1 U14976 ( .A1(n14336), .A2(n11824), .B1(n12392), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11905) );
  NAND2_X1 U14977 ( .A1(n12282), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11904) );
  XOR2_X1 U14978 ( .A(n11934), .B(n11935), .Z(n20131) );
  INV_X1 U14979 ( .A(n20131), .ZN(n11922) );
  AOI22_X1 U14980 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11911) );
  AOI22_X1 U14981 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11910) );
  AOI22_X1 U14982 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U14983 ( .A1(n12120), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11908) );
  NAND4_X1 U14984 ( .A1(n11911), .A2(n11910), .A3(n11909), .A4(n11908), .ZN(
        n11917) );
  AOI22_X1 U14985 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12142), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11915) );
  AOI22_X1 U14986 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11429), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11914) );
  AOI22_X1 U14987 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11913) );
  AOI22_X1 U14988 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11912) );
  NAND4_X1 U14989 ( .A1(n11915), .A2(n11914), .A3(n11913), .A4(n11912), .ZN(
        n11916) );
  NOR2_X1 U14990 ( .A1(n11917), .A2(n11916), .ZN(n11920) );
  NAND2_X1 U14991 ( .A1(n11843), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11919) );
  NAND2_X1 U14992 ( .A1(n12392), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11918) );
  OAI211_X1 U14993 ( .C1(n12016), .C2(n11920), .A(n11919), .B(n11918), .ZN(
        n11921) );
  AOI21_X1 U14994 ( .B1(n11922), .B2(n11824), .A(n11921), .ZN(n14265) );
  NAND2_X1 U14995 ( .A1(n14119), .A2(n11923), .ZN(n14264) );
  AOI22_X1 U14996 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11428), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11927) );
  AOI22_X1 U14997 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12295), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11926) );
  AOI22_X1 U14998 ( .A1(n12266), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12120), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11925) );
  AOI22_X1 U14999 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11924) );
  NAND4_X1 U15000 ( .A1(n11927), .A2(n11926), .A3(n11925), .A4(n11924), .ZN(
        n11933) );
  AOI22_X1 U15001 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12142), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11931) );
  AOI22_X1 U15002 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11930) );
  AOI22_X1 U15003 ( .A1(n11422), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11929) );
  AOI22_X1 U15004 ( .A1(n12081), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11928) );
  NAND4_X1 U15005 ( .A1(n11931), .A2(n11930), .A3(n11929), .A4(n11928), .ZN(
        n11932) );
  NOR2_X1 U15006 ( .A1(n11933), .A2(n11932), .ZN(n11938) );
  XNOR2_X1 U15007 ( .A(n11940), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14821) );
  NAND2_X1 U15008 ( .A1(n14821), .A2(n12289), .ZN(n11937) );
  AOI22_X1 U15009 ( .A1(n11843), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n12392), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11936) );
  OAI211_X1 U15010 ( .C1(n11938), .C2(n12016), .A(n11937), .B(n11936), .ZN(
        n14318) );
  NAND2_X1 U15011 ( .A1(n11843), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n11943) );
  OAI21_X1 U15012 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11941), .A(
        n11955), .ZN(n16118) );
  AOI22_X1 U15013 ( .A1(n12392), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n16118), .B2(n12289), .ZN(n11942) );
  NAND2_X1 U15014 ( .A1(n11943), .A2(n11942), .ZN(n14362) );
  AOI22_X1 U15015 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11947) );
  AOI22_X1 U15016 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12303), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11946) );
  AOI22_X1 U15017 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11945) );
  AOI22_X1 U15018 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11944) );
  NAND4_X1 U15019 ( .A1(n11947), .A2(n11946), .A3(n11945), .A4(n11944), .ZN(
        n11953) );
  AOI22_X1 U15020 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11951) );
  AOI22_X1 U15021 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11950) );
  AOI22_X1 U15022 ( .A1(n12266), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11949) );
  AOI22_X1 U15023 ( .A1(n12120), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11948) );
  NAND4_X1 U15024 ( .A1(n11951), .A2(n11950), .A3(n11949), .A4(n11948), .ZN(
        n11952) );
  OR2_X1 U15025 ( .A1(n11953), .A2(n11952), .ZN(n11954) );
  AND2_X1 U15026 ( .A1(n11967), .A2(n11954), .ZN(n14380) );
  XOR2_X1 U15027 ( .A(n14809), .B(n11987), .Z(n14811) );
  AOI22_X1 U15028 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11959) );
  AOI22_X1 U15029 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12266), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11958) );
  AOI22_X1 U15030 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12120), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U15031 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11956) );
  NAND4_X1 U15032 ( .A1(n11959), .A2(n11958), .A3(n11957), .A4(n11956), .ZN(
        n11965) );
  AOI22_X1 U15033 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11963) );
  AOI22_X1 U15034 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U15035 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11961) );
  AOI22_X1 U15036 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11960) );
  NAND4_X1 U15037 ( .A1(n11963), .A2(n11962), .A3(n11961), .A4(n11960), .ZN(
        n11964) );
  OR2_X1 U15038 ( .A1(n11965), .A2(n11964), .ZN(n11966) );
  AOI22_X1 U15039 ( .A1(n11967), .A2(n11966), .B1(n12392), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11969) );
  NAND2_X1 U15040 ( .A1(n11843), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11968) );
  OAI211_X1 U15041 ( .C1(n14811), .C2(n12315), .A(n11969), .B(n11968), .ZN(
        n14383) );
  XOR2_X1 U15042 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11970), .Z(
        n16107) );
  AOI22_X1 U15043 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11974) );
  AOI22_X1 U15044 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12302), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11973) );
  AOI22_X1 U15045 ( .A1(n11429), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11972) );
  AOI22_X1 U15046 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11971) );
  NAND4_X1 U15047 ( .A1(n11974), .A2(n11973), .A3(n11972), .A4(n11971), .ZN(
        n11980) );
  AOI22_X1 U15048 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12301), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11978) );
  AOI22_X1 U15049 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11551), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11977) );
  AOI22_X1 U15050 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12120), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U15051 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11975) );
  NAND4_X1 U15052 ( .A1(n11978), .A2(n11977), .A3(n11976), .A4(n11975), .ZN(
        n11979) );
  NOR2_X1 U15053 ( .A1(n11980), .A2(n11979), .ZN(n11983) );
  NAND2_X1 U15054 ( .A1(n11843), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11982) );
  NAND2_X1 U15055 ( .A1(n12392), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11981) );
  OAI211_X1 U15056 ( .C1(n12016), .C2(n11983), .A(n11982), .B(n11981), .ZN(
        n11984) );
  INV_X1 U15057 ( .A(n11984), .ZN(n11985) );
  OAI21_X1 U15058 ( .B1(n16107), .B2(n12315), .A(n11985), .ZN(n14382) );
  XNOR2_X1 U15059 ( .A(n12002), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16031) );
  AOI22_X1 U15060 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11991) );
  AOI22_X1 U15061 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11990) );
  AOI22_X1 U15062 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U15063 ( .A1(n12266), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11988) );
  NAND4_X1 U15064 ( .A1(n11991), .A2(n11990), .A3(n11989), .A4(n11988), .ZN(
        n11997) );
  AOI22_X1 U15065 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11995) );
  AOI22_X1 U15066 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11428), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11994) );
  AOI22_X1 U15067 ( .A1(n12120), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U15068 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11992) );
  NAND4_X1 U15069 ( .A1(n11995), .A2(n11994), .A3(n11993), .A4(n11992), .ZN(
        n11996) );
  NOR2_X1 U15070 ( .A1(n11997), .A2(n11996), .ZN(n12000) );
  NAND2_X1 U15071 ( .A1(n11843), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11999) );
  NAND2_X1 U15072 ( .A1(n12392), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11998) );
  OAI211_X1 U15073 ( .C1(n12016), .C2(n12000), .A(n11999), .B(n11998), .ZN(
        n12001) );
  AOI21_X1 U15074 ( .B1(n16031), .B2(n11824), .A(n12001), .ZN(n14374) );
  XOR2_X1 U15075 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n12020), .Z(
        n16098) );
  INV_X1 U15076 ( .A(n16098), .ZN(n12018) );
  AOI22_X1 U15077 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12006) );
  AOI22_X1 U15078 ( .A1(n12120), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12005) );
  AOI22_X1 U15079 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12004) );
  AOI22_X1 U15080 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12003) );
  NAND4_X1 U15081 ( .A1(n12006), .A2(n12005), .A3(n12004), .A4(n12003), .ZN(
        n12012) );
  AOI22_X1 U15082 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11428), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12010) );
  AOI22_X1 U15083 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12266), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12009) );
  AOI22_X1 U15084 ( .A1(n12206), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12008) );
  AOI22_X1 U15085 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12007) );
  NAND4_X1 U15086 ( .A1(n12010), .A2(n12009), .A3(n12008), .A4(n12007), .ZN(
        n12011) );
  NOR2_X1 U15087 ( .A1(n12012), .A2(n12011), .ZN(n12015) );
  NAND2_X1 U15088 ( .A1(n11843), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12014) );
  NAND2_X1 U15089 ( .A1(n12392), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12013) );
  OAI211_X1 U15090 ( .C1(n12016), .C2(n12015), .A(n12014), .B(n12013), .ZN(
        n12017) );
  AOI21_X1 U15091 ( .B1(n12018), .B2(n11824), .A(n12017), .ZN(n14645) );
  XNOR2_X1 U15092 ( .A(n12034), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14575) );
  AOI22_X1 U15093 ( .A1(n12266), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12024) );
  AOI22_X1 U15094 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12023) );
  AOI22_X1 U15095 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12022) );
  AOI22_X1 U15096 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12021) );
  NAND4_X1 U15097 ( .A1(n12024), .A2(n12023), .A3(n12022), .A4(n12021), .ZN(
        n12030) );
  AOI22_X1 U15098 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12142), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12028) );
  AOI22_X1 U15099 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12120), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12027) );
  AOI22_X1 U15100 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12026) );
  AOI22_X1 U15101 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12025) );
  NAND4_X1 U15102 ( .A1(n12028), .A2(n12027), .A3(n12026), .A4(n12025), .ZN(
        n12029) );
  OAI21_X1 U15103 ( .B1(n12030), .B2(n12029), .A(n12312), .ZN(n12032) );
  AOI22_X1 U15104 ( .A1(n11843), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20968), .ZN(n12031) );
  AOI21_X1 U15105 ( .B1(n12032), .B2(n12031), .A(n11824), .ZN(n12033) );
  AOI21_X1 U15106 ( .B1(n14575), .B2(n11824), .A(n12033), .ZN(n14566) );
  XOR2_X1 U15107 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12047), .Z(
        n16088) );
  AOI22_X1 U15108 ( .A1(n11843), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n12392), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12046) );
  AOI22_X1 U15109 ( .A1(n12142), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11428), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12038) );
  AOI22_X1 U15110 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12266), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12037) );
  AOI22_X1 U15111 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12036) );
  AOI22_X1 U15112 ( .A1(n12206), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12035) );
  NAND4_X1 U15113 ( .A1(n12038), .A2(n12037), .A3(n12036), .A4(n12035), .ZN(
        n12044) );
  AOI22_X1 U15114 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11570), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12042) );
  AOI22_X1 U15115 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12041) );
  AOI22_X1 U15116 ( .A1(n12120), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12040) );
  AOI22_X1 U15117 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12039) );
  NAND4_X1 U15118 ( .A1(n12042), .A2(n12041), .A3(n12040), .A4(n12039), .ZN(
        n12043) );
  OAI21_X1 U15119 ( .B1(n12044), .B2(n12043), .A(n12312), .ZN(n12045) );
  OAI211_X1 U15120 ( .C1(n16088), .C2(n12315), .A(n12046), .B(n12045), .ZN(
        n14638) );
  XNOR2_X1 U15121 ( .A(n12077), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16009) );
  NAND2_X1 U15122 ( .A1(n16009), .A2(n12289), .ZN(n12062) );
  AOI22_X1 U15123 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12142), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12051) );
  AOI22_X1 U15124 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11429), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U15125 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12049) );
  AOI22_X1 U15126 ( .A1(n12120), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12048) );
  NAND4_X1 U15127 ( .A1(n12051), .A2(n12050), .A3(n12049), .A4(n12048), .ZN(
        n12057) );
  AOI22_X1 U15128 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12303), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12055) );
  AOI22_X1 U15129 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12054) );
  AOI22_X1 U15130 ( .A1(n12206), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12053) );
  AOI22_X1 U15131 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12052) );
  NAND4_X1 U15132 ( .A1(n12055), .A2(n12054), .A3(n12053), .A4(n12052), .ZN(
        n12056) );
  NOR2_X1 U15133 ( .A1(n12057), .A2(n12056), .ZN(n12060) );
  AOI21_X1 U15134 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n16011), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12058) );
  AOI21_X1 U15135 ( .B1(n11843), .B2(P1_EAX_REG_18__SCAN_IN), .A(n12058), .ZN(
        n12059) );
  OAI21_X1 U15136 ( .B1(n12284), .B2(n12060), .A(n12059), .ZN(n12061) );
  NAND2_X1 U15137 ( .A1(n12062), .A2(n12061), .ZN(n14630) );
  AOI22_X1 U15138 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12142), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12066) );
  AOI22_X1 U15139 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12266), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12065) );
  AOI22_X1 U15140 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12064) );
  AOI22_X1 U15141 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12063) );
  NAND4_X1 U15142 ( .A1(n12066), .A2(n12065), .A3(n12064), .A4(n12063), .ZN(
        n12072) );
  AOI22_X1 U15143 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12070) );
  AOI22_X1 U15144 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U15145 ( .A1(n12120), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12068) );
  AOI22_X1 U15146 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12067) );
  NAND4_X1 U15147 ( .A1(n12070), .A2(n12069), .A3(n12068), .A4(n12067), .ZN(
        n12071) );
  NOR2_X1 U15148 ( .A1(n12072), .A2(n12071), .ZN(n12076) );
  NAND2_X1 U15149 ( .A1(n20968), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12073) );
  NAND2_X1 U15150 ( .A1(n12315), .A2(n12073), .ZN(n12074) );
  AOI21_X1 U15151 ( .B1(n11843), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12074), .ZN(
        n12075) );
  OAI21_X1 U15152 ( .B1(n12284), .B2(n12076), .A(n12075), .ZN(n12080) );
  OAI21_X1 U15153 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n12078), .A(
        n12111), .ZN(n16081) );
  OR2_X1 U15154 ( .A1(n12315), .A2(n16081), .ZN(n12079) );
  NAND2_X1 U15155 ( .A1(n12080), .A2(n12079), .ZN(n14620) );
  AOI22_X1 U15156 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12301), .B1(
        n12303), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12085) );
  AOI22_X1 U15157 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12302), .B1(
        n12120), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12084) );
  AOI22_X1 U15158 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12081), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12083) );
  AOI22_X1 U15159 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12082) );
  NAND4_X1 U15160 ( .A1(n12085), .A2(n12084), .A3(n12083), .A4(n12082), .ZN(
        n12091) );
  AOI22_X1 U15161 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12142), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12089) );
  AOI22_X1 U15162 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12088) );
  AOI22_X1 U15163 ( .A1(n11429), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12087) );
  AOI22_X1 U15164 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11551), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12086) );
  NAND4_X1 U15165 ( .A1(n12089), .A2(n12088), .A3(n12087), .A4(n12086), .ZN(
        n12090) );
  NOR2_X1 U15166 ( .A1(n12091), .A2(n12090), .ZN(n12094) );
  INV_X1 U15167 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16075) );
  AOI21_X1 U15168 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n16075), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12092) );
  AOI21_X1 U15169 ( .B1(n11843), .B2(P1_EAX_REG_20__SCAN_IN), .A(n12092), .ZN(
        n12093) );
  OAI21_X1 U15170 ( .B1(n12284), .B2(n12094), .A(n12093), .ZN(n12096) );
  XNOR2_X1 U15171 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n12111), .ZN(
        n16071) );
  NAND2_X1 U15172 ( .A1(n16071), .A2(n12289), .ZN(n12095) );
  AOI22_X1 U15173 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12100) );
  AOI22_X1 U15174 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12295), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12099) );
  AOI22_X1 U15175 ( .A1(n11480), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12098) );
  AOI22_X1 U15176 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12097) );
  NAND4_X1 U15177 ( .A1(n12100), .A2(n12099), .A3(n12098), .A4(n12097), .ZN(
        n12106) );
  AOI22_X1 U15178 ( .A1(n11429), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12120), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12104) );
  AOI22_X1 U15179 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12103) );
  AOI22_X1 U15180 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U15181 ( .A1(n12081), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12101) );
  NAND4_X1 U15182 ( .A1(n12104), .A2(n12103), .A3(n12102), .A4(n12101), .ZN(
        n12105) );
  NOR2_X1 U15183 ( .A1(n12106), .A2(n12105), .ZN(n12110) );
  NAND2_X1 U15184 ( .A1(n20968), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12107) );
  NAND2_X1 U15185 ( .A1(n12315), .A2(n12107), .ZN(n12108) );
  AOI21_X1 U15186 ( .B1(n11843), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12108), .ZN(
        n12109) );
  OAI21_X1 U15187 ( .B1(n12284), .B2(n12110), .A(n12109), .ZN(n12115) );
  OAI21_X1 U15188 ( .B1(n12113), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n12157), .ZN(n15981) );
  OR2_X1 U15189 ( .A1(n15981), .A2(n12315), .ZN(n12114) );
  AOI22_X1 U15190 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12119) );
  AOI22_X1 U15191 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12118) );
  AOI22_X1 U15192 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12117) );
  AOI22_X1 U15193 ( .A1(n11429), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12116) );
  NAND4_X1 U15194 ( .A1(n12119), .A2(n12118), .A3(n12117), .A4(n12116), .ZN(
        n12126) );
  AOI22_X1 U15195 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12120), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12124) );
  AOI22_X1 U15196 ( .A1(n11480), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12123) );
  AOI22_X1 U15197 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12122) );
  AOI22_X1 U15198 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12121) );
  NAND4_X1 U15199 ( .A1(n12124), .A2(n12123), .A3(n12122), .A4(n12121), .ZN(
        n12125) );
  NOR2_X1 U15200 ( .A1(n12126), .A2(n12125), .ZN(n12129) );
  INV_X1 U15201 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15974) );
  AOI21_X1 U15202 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15974), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12127) );
  AOI21_X1 U15203 ( .B1(n11843), .B2(P1_EAX_REG_22__SCAN_IN), .A(n12127), .ZN(
        n12128) );
  OAI21_X1 U15204 ( .B1(n12284), .B2(n12129), .A(n12128), .ZN(n12131) );
  XNOR2_X1 U15205 ( .A(n12157), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15979) );
  NAND2_X1 U15206 ( .A1(n15979), .A2(n12289), .ZN(n12130) );
  AOI22_X1 U15207 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12135) );
  AOI22_X1 U15208 ( .A1(n11408), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U15209 ( .A1(n12120), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U15210 ( .A1(n11414), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12132) );
  NAND4_X1 U15211 ( .A1(n12135), .A2(n12134), .A3(n12133), .A4(n12132), .ZN(
        n12141) );
  AOI22_X1 U15212 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12142), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12139) );
  AOI22_X1 U15213 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12266), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12138) );
  AOI22_X1 U15214 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12137) );
  AOI22_X1 U15215 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12136) );
  NAND4_X1 U15216 ( .A1(n12139), .A2(n12138), .A3(n12137), .A4(n12136), .ZN(
        n12140) );
  NOR2_X1 U15217 ( .A1(n12141), .A2(n12140), .ZN(n12162) );
  AOI22_X1 U15218 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12142), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12146) );
  AOI22_X1 U15219 ( .A1(n11408), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11428), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12145) );
  AOI22_X1 U15220 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12266), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12144) );
  AOI22_X1 U15221 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12143) );
  NAND4_X1 U15222 ( .A1(n12146), .A2(n12145), .A3(n12144), .A4(n12143), .ZN(
        n12152) );
  AOI22_X1 U15223 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12120), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12150) );
  AOI22_X1 U15224 ( .A1(n11414), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12149) );
  AOI22_X1 U15225 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U15226 ( .A1(n12206), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12147) );
  NAND4_X1 U15227 ( .A1(n12150), .A2(n12149), .A3(n12148), .A4(n12147), .ZN(
        n12151) );
  NOR2_X1 U15228 ( .A1(n12152), .A2(n12151), .ZN(n12163) );
  XNOR2_X1 U15229 ( .A(n12162), .B(n12163), .ZN(n12156) );
  NAND2_X1 U15230 ( .A1(n20968), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12153) );
  NAND2_X1 U15231 ( .A1(n12315), .A2(n12153), .ZN(n12154) );
  AOI21_X1 U15232 ( .B1(n11843), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12154), .ZN(
        n12155) );
  OAI21_X1 U15233 ( .B1(n12284), .B2(n12156), .A(n12155), .ZN(n12161) );
  OR2_X1 U15234 ( .A1(n12158), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12159) );
  NAND2_X1 U15235 ( .A1(n12196), .A2(n12159), .ZN(n16067) );
  NAND2_X1 U15236 ( .A1(n12161), .A2(n12160), .ZN(n14550) );
  NOR2_X1 U15237 ( .A1(n12163), .A2(n12162), .ZN(n12182) );
  AOI22_X1 U15238 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12168) );
  AOI22_X1 U15239 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12303), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12167) );
  AOI22_X1 U15240 ( .A1(n11408), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12266), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12166) );
  INV_X1 U15241 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n20330) );
  AOI22_X1 U15242 ( .A1(n12206), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12165) );
  NAND4_X1 U15243 ( .A1(n12168), .A2(n12167), .A3(n12166), .A4(n12165), .ZN(
        n12174) );
  AOI22_X1 U15244 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12172) );
  AOI22_X1 U15245 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12171) );
  AOI22_X1 U15246 ( .A1(n12120), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12170) );
  AOI22_X1 U15247 ( .A1(n11414), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12169) );
  NAND4_X1 U15248 ( .A1(n12172), .A2(n12171), .A3(n12170), .A4(n12169), .ZN(
        n12173) );
  OR2_X1 U15249 ( .A1(n12174), .A2(n12173), .ZN(n12181) );
  INV_X1 U15250 ( .A(n12181), .ZN(n12175) );
  XNOR2_X1 U15251 ( .A(n12182), .B(n12175), .ZN(n12176) );
  NAND2_X1 U15252 ( .A1(n12176), .A2(n12312), .ZN(n12180) );
  INV_X1 U15253 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15966) );
  AOI21_X1 U15254 ( .B1(n15966), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12177) );
  AOI21_X1 U15255 ( .B1(n11843), .B2(P1_EAX_REG_24__SCAN_IN), .A(n12177), .ZN(
        n12179) );
  XNOR2_X1 U15256 ( .A(n12196), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15963) );
  AOI21_X1 U15257 ( .B1(n12180), .B2(n12179), .A(n12178), .ZN(n14594) );
  NAND2_X1 U15258 ( .A1(n12182), .A2(n12181), .ZN(n12204) );
  AOI22_X1 U15259 ( .A1(n11480), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12266), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12186) );
  AOI22_X1 U15260 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12185) );
  AOI22_X1 U15261 ( .A1(n12206), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12184) );
  AOI22_X1 U15262 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12183) );
  NAND4_X1 U15263 ( .A1(n12186), .A2(n12185), .A3(n12184), .A4(n12183), .ZN(
        n12192) );
  AOI22_X1 U15264 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12142), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12190) );
  AOI22_X1 U15265 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12303), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U15266 ( .A1(n12120), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12188) );
  AOI22_X1 U15267 ( .A1(n11408), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12187) );
  NAND4_X1 U15268 ( .A1(n12190), .A2(n12189), .A3(n12188), .A4(n12187), .ZN(
        n12191) );
  NOR2_X1 U15269 ( .A1(n12192), .A2(n12191), .ZN(n12205) );
  XNOR2_X1 U15270 ( .A(n12204), .B(n12205), .ZN(n12195) );
  INV_X1 U15271 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12199) );
  AOI21_X1 U15272 ( .B1(n12199), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12193) );
  AOI21_X1 U15273 ( .B1(n11843), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12193), .ZN(
        n12194) );
  OAI21_X1 U15274 ( .B1(n12195), .B2(n12284), .A(n12194), .ZN(n12203) );
  INV_X1 U15275 ( .A(n12198), .ZN(n12200) );
  NAND2_X1 U15276 ( .A1(n12200), .A2(n12199), .ZN(n12201) );
  NAND2_X1 U15277 ( .A1(n12239), .A2(n12201), .ZN(n15946) );
  NAND2_X1 U15278 ( .A1(n14584), .A2(n14585), .ZN(n14537) );
  NOR2_X1 U15279 ( .A1(n12205), .A2(n12204), .ZN(n12234) );
  AOI22_X1 U15280 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12142), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U15281 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12303), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12209) );
  AOI22_X1 U15282 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12266), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12208) );
  AOI22_X1 U15283 ( .A1(n12206), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12207) );
  NAND4_X1 U15284 ( .A1(n12210), .A2(n12209), .A3(n12208), .A4(n12207), .ZN(
        n12216) );
  AOI22_X1 U15285 ( .A1(n11480), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12214) );
  AOI22_X1 U15286 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12213) );
  AOI22_X1 U15287 ( .A1(n12120), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12212) );
  AOI22_X1 U15288 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12211) );
  NAND4_X1 U15289 ( .A1(n12214), .A2(n12213), .A3(n12212), .A4(n12211), .ZN(
        n12215) );
  OR2_X1 U15290 ( .A1(n12216), .A2(n12215), .ZN(n12233) );
  XNOR2_X1 U15291 ( .A(n12234), .B(n12233), .ZN(n12220) );
  NAND2_X1 U15292 ( .A1(n20968), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12217) );
  NAND2_X1 U15293 ( .A1(n12315), .A2(n12217), .ZN(n12218) );
  AOI21_X1 U15294 ( .B1(n12282), .B2(P1_EAX_REG_26__SCAN_IN), .A(n12218), .ZN(
        n12219) );
  OAI21_X1 U15295 ( .B1(n12220), .B2(n12284), .A(n12219), .ZN(n12222) );
  XNOR2_X1 U15296 ( .A(n12239), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14740) );
  NAND2_X1 U15297 ( .A1(n14740), .A2(n12289), .ZN(n12221) );
  NAND2_X1 U15298 ( .A1(n12222), .A2(n12221), .ZN(n14538) );
  AOI22_X1 U15299 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12164), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U15300 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12266), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12225) );
  AOI22_X1 U15301 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12224) );
  AOI22_X1 U15302 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12223) );
  NAND4_X1 U15303 ( .A1(n12226), .A2(n12225), .A3(n12224), .A4(n12223), .ZN(
        n12232) );
  AOI22_X1 U15304 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n11551), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12230) );
  AOI22_X1 U15305 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12295), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12229) );
  AOI22_X1 U15306 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11570), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U15307 ( .A1(n12120), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12227) );
  NAND4_X1 U15308 ( .A1(n12230), .A2(n12229), .A3(n12228), .A4(n12227), .ZN(
        n12231) );
  NOR2_X1 U15309 ( .A1(n12232), .A2(n12231), .ZN(n12248) );
  NAND2_X1 U15310 ( .A1(n12234), .A2(n12233), .ZN(n12247) );
  XNOR2_X1 U15311 ( .A(n12248), .B(n12247), .ZN(n12238) );
  NAND2_X1 U15312 ( .A1(n20968), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12235) );
  NAND2_X1 U15313 ( .A1(n12315), .A2(n12235), .ZN(n12236) );
  AOI21_X1 U15314 ( .B1(n12282), .B2(P1_EAX_REG_27__SCAN_IN), .A(n12236), .ZN(
        n12237) );
  OAI21_X1 U15315 ( .B1(n12238), .B2(n12284), .A(n12237), .ZN(n12245) );
  INV_X1 U15316 ( .A(n12239), .ZN(n12240) );
  INV_X1 U15317 ( .A(n12241), .ZN(n12242) );
  INV_X1 U15318 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14526) );
  NAND2_X1 U15319 ( .A1(n12242), .A2(n14526), .ZN(n12243) );
  NAND2_X1 U15320 ( .A1(n12286), .A2(n12243), .ZN(n14731) );
  NAND2_X1 U15321 ( .A1(n12245), .A2(n12244), .ZN(n14521) );
  INV_X1 U15322 ( .A(n14521), .ZN(n12246) );
  NOR2_X1 U15323 ( .A1(n12248), .A2(n12247), .ZN(n12279) );
  AOI22_X1 U15324 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12142), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U15325 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11428), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12251) );
  AOI22_X1 U15326 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12266), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12250) );
  AOI22_X1 U15327 ( .A1(n12206), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12249) );
  NAND4_X1 U15328 ( .A1(n12252), .A2(n12251), .A3(n12250), .A4(n12249), .ZN(
        n12258) );
  AOI22_X1 U15329 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12256) );
  AOI22_X1 U15330 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12255) );
  AOI22_X1 U15331 ( .A1(n12120), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12254) );
  AOI22_X1 U15332 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12253) );
  NAND4_X1 U15333 ( .A1(n12256), .A2(n12255), .A3(n12254), .A4(n12253), .ZN(
        n12257) );
  OR2_X1 U15334 ( .A1(n12258), .A2(n12257), .ZN(n12278) );
  INV_X1 U15335 ( .A(n12278), .ZN(n12259) );
  XNOR2_X1 U15336 ( .A(n12279), .B(n12259), .ZN(n12260) );
  NAND2_X1 U15337 ( .A1(n12260), .A2(n12312), .ZN(n12264) );
  INV_X1 U15338 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13311) );
  AOI21_X1 U15339 ( .B1(n13311), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12261) );
  AOI21_X1 U15340 ( .B1(n12282), .B2(P1_EAX_REG_28__SCAN_IN), .A(n12261), .ZN(
        n12263) );
  XNOR2_X1 U15341 ( .A(n12286), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14435) );
  AOI22_X1 U15342 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12120), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12271) );
  AOI22_X1 U15343 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12270) );
  AOI22_X1 U15344 ( .A1(n12266), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12269) );
  AOI22_X1 U15345 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12267), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12268) );
  NAND4_X1 U15346 ( .A1(n12271), .A2(n12270), .A3(n12269), .A4(n12268), .ZN(
        n12277) );
  AOI22_X1 U15347 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12142), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12275) );
  AOI22_X1 U15348 ( .A1(n11570), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12303), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U15349 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12273) );
  AOI22_X1 U15350 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12272) );
  NAND4_X1 U15351 ( .A1(n12275), .A2(n12274), .A3(n12273), .A4(n12272), .ZN(
        n12276) );
  NOR2_X1 U15352 ( .A1(n12277), .A2(n12276), .ZN(n12293) );
  NAND2_X1 U15353 ( .A1(n12279), .A2(n12278), .ZN(n12292) );
  XNOR2_X1 U15354 ( .A(n12293), .B(n12292), .ZN(n12285) );
  NAND2_X1 U15355 ( .A1(n20968), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12280) );
  NAND2_X1 U15356 ( .A1(n12315), .A2(n12280), .ZN(n12281) );
  AOI21_X1 U15357 ( .B1(n12282), .B2(P1_EAX_REG_29__SCAN_IN), .A(n12281), .ZN(
        n12283) );
  OAI21_X1 U15358 ( .B1(n12285), .B2(n12284), .A(n12283), .ZN(n12291) );
  INV_X1 U15359 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14721) );
  NAND2_X1 U15360 ( .A1(n12287), .A2(n14721), .ZN(n12288) );
  NAND2_X1 U15361 ( .A1(n14719), .A2(n12289), .ZN(n12290) );
  NAND2_X1 U15362 ( .A1(n12291), .A2(n12290), .ZN(n14507) );
  NOR2_X1 U15363 ( .A1(n12293), .A2(n12292), .ZN(n12311) );
  AOI22_X1 U15364 ( .A1(n11612), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11550), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12299) );
  AOI22_X1 U15365 ( .A1(n12142), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11422), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U15366 ( .A1(n12120), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12265), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12297) );
  AOI22_X1 U15367 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12296) );
  NAND4_X1 U15368 ( .A1(n12299), .A2(n12298), .A3(n12297), .A4(n12296), .ZN(
        n12309) );
  AOI22_X1 U15369 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11570), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12307) );
  AOI22_X1 U15370 ( .A1(n12301), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12266), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12306) );
  AOI22_X1 U15371 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12305) );
  AOI22_X1 U15372 ( .A1(n12303), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12206), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12304) );
  NAND4_X1 U15373 ( .A1(n12307), .A2(n12306), .A3(n12305), .A4(n12304), .ZN(
        n12308) );
  NOR2_X1 U15374 ( .A1(n12309), .A2(n12308), .ZN(n12310) );
  XNOR2_X1 U15375 ( .A(n12311), .B(n12310), .ZN(n12313) );
  NAND2_X1 U15376 ( .A1(n12313), .A2(n12312), .ZN(n12319) );
  NAND2_X1 U15377 ( .A1(n20968), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12314) );
  NAND2_X1 U15378 ( .A1(n12315), .A2(n12314), .ZN(n12316) );
  AOI21_X1 U15379 ( .B1(n11843), .B2(P1_EAX_REG_30__SCAN_IN), .A(n12316), .ZN(
        n12318) );
  XNOR2_X1 U15380 ( .A(n12397), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14500) );
  AOI21_X1 U15381 ( .B1(n12319), .B2(n12318), .A(n12317), .ZN(n12391) );
  XNOR2_X1 U15382 ( .A(n14506), .B(n12320), .ZN(n14496) );
  NOR2_X1 U15383 ( .A1(n12321), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13878) );
  AND2_X1 U15384 ( .A1(n20971), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n16289) );
  INV_X1 U15385 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12396) );
  NOR2_X2 U15386 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20823) );
  OR2_X1 U15387 ( .A1(n12324), .A2(n20823), .ZN(n20974) );
  AND2_X1 U15388 ( .A1(n20974), .A2(n20971), .ZN(n12322) );
  NOR2_X1 U15389 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20968), .ZN(n20976) );
  AOI21_X1 U15390 ( .B1(n21106), .B2(P1_STATE2_REG_1__SCAN_IN), .A(n20976), 
        .ZN(n13663) );
  INV_X1 U15391 ( .A(n13663), .ZN(n12323) );
  NAND2_X1 U15392 ( .A1(n20249), .A2(n14500), .ZN(n12325) );
  INV_X2 U15393 ( .A(n10234), .ZN(n20290) );
  NAND2_X1 U15394 ( .A1(n20290), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14835) );
  OAI211_X1 U15395 ( .C1(n12396), .C2(n16074), .A(n12325), .B(n14835), .ZN(
        n12326) );
  AOI21_X1 U15396 ( .B1(n14496), .B2(n20313), .A(n12326), .ZN(n12327) );
  XNOR2_X1 U15397 ( .A(n12331), .B(n12330), .ZN(n15268) );
  INV_X1 U15398 ( .A(n12330), .ZN(n12332) );
  AOI22_X1 U15399 ( .A1(n15268), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n12332), .B2(n12331), .ZN(n12335) );
  XNOR2_X1 U15400 ( .A(n12333), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12334) );
  XNOR2_X1 U15401 ( .A(n12335), .B(n12334), .ZN(n12362) );
  AND2_X1 U15402 ( .A1(n12336), .A2(n13539), .ZN(n12337) );
  NAND2_X1 U15403 ( .A1(n12338), .A2(n12337), .ZN(n13473) );
  INV_X1 U15404 ( .A(n13473), .ZN(n12343) );
  NAND2_X1 U15405 ( .A1(n12362), .A2(n19397), .ZN(n12361) );
  NAND2_X1 U15406 ( .A1(n12340), .A2(n12341), .ZN(n12342) );
  NAND2_X1 U15407 ( .A1(n12339), .A2(n12342), .ZN(n12369) );
  NAND2_X1 U15408 ( .A1(n19860), .A2(n20072), .ZN(n20089) );
  NAND2_X1 U15409 ( .A1(n20089), .A2(n14091), .ZN(n12344) );
  NAND2_X1 U15410 ( .A1(n14091), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12426) );
  INV_X1 U15411 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19541) );
  NAND2_X1 U15412 ( .A1(n19541), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13390) );
  NAND2_X1 U15413 ( .A1(n12426), .A2(n13390), .ZN(n13498) );
  NAND2_X1 U15414 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n13379), .ZN(
        n13378) );
  INV_X1 U15415 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15383) );
  INV_X1 U15416 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n19141) );
  INV_X1 U15417 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15322) );
  INV_X1 U15418 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15297) );
  INV_X1 U15419 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n13436) );
  INV_X1 U15420 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15269) );
  INV_X1 U15421 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12356) );
  AND2_X1 U15422 ( .A1(n13442), .A2(n12356), .ZN(n12345) );
  NOR2_X1 U15423 ( .A1(n14920), .A2(n12345), .ZN(n14937) );
  INV_X1 U15424 ( .A(n12346), .ZN(n12349) );
  INV_X1 U15425 ( .A(n13447), .ZN(n12348) );
  AOI21_X1 U15426 ( .B1(n12349), .B2(n12348), .A(n12347), .ZN(n14936) );
  NOR2_X1 U15427 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16542) );
  INV_X1 U15428 ( .A(n16542), .ZN(n12350) );
  NAND2_X1 U15429 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n13543) );
  NAND2_X1 U15430 ( .A1(n12350), .A2(n13543), .ZN(n12351) );
  OR2_X1 U15431 ( .A1(n19860), .A2(n19541), .ZN(n20093) );
  INV_X1 U15432 ( .A(n20093), .ZN(n12354) );
  NAND2_X1 U15433 ( .A1(n14936), .A2(n19399), .ZN(n12355) );
  NAND2_X1 U15434 ( .A1(n19198), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12365) );
  OAI211_X1 U15435 ( .C1(n12356), .C2(n19394), .A(n12355), .B(n12365), .ZN(
        n12357) );
  AOI21_X1 U15436 ( .B1(n16473), .B2(n14937), .A(n12357), .ZN(n12358) );
  NAND2_X1 U15437 ( .A1(n12361), .A2(n12360), .ZN(P2_U2986) );
  NAND2_X1 U15438 ( .A1(n12362), .A2(n16530), .ZN(n12372) );
  NAND2_X1 U15439 ( .A1(n13452), .A2(n12363), .ZN(n12364) );
  INV_X1 U15440 ( .A(n15440), .ZN(n12366) );
  NAND2_X1 U15441 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15424) );
  AOI21_X1 U15442 ( .B1(n12366), .B2(n15424), .A(n15442), .ZN(n15423) );
  AOI21_X1 U15443 ( .B1(n12366), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12367) );
  NOR2_X1 U15444 ( .A1(n15423), .A2(n12367), .ZN(n12368) );
  NAND2_X1 U15445 ( .A1(n12372), .A2(n12371), .ZN(P2_U3018) );
  NAND2_X1 U15446 ( .A1(n12373), .A2(n15257), .ZN(n12378) );
  INV_X1 U15447 ( .A(n12374), .ZN(n12375) );
  NOR2_X1 U15448 ( .A1(n12376), .A2(n12375), .ZN(n12377) );
  XNOR2_X1 U15449 ( .A(n12378), .B(n12377), .ZN(n15419) );
  NAND2_X1 U15450 ( .A1(n12704), .A2(n12379), .ZN(n12380) );
  NAND2_X1 U15451 ( .A1(n19198), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15409) );
  NAND2_X1 U15452 ( .A1(n16447), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12382) );
  OAI211_X1 U15453 ( .C1(n15408), .C2(n16414), .A(n15409), .B(n12382), .ZN(
        n12383) );
  INV_X1 U15454 ( .A(n12383), .ZN(n12385) );
  INV_X1 U15455 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14926) );
  XNOR2_X1 U15456 ( .A(n13317), .B(n14926), .ZN(n14923) );
  INV_X1 U15457 ( .A(n14923), .ZN(n12384) );
  OAI211_X1 U15458 ( .C1(n15419), .C2(n16465), .A(n12386), .B(n10238), .ZN(
        P2_U2984) );
  OAI21_X1 U15459 ( .B1(n12389), .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n12388), .ZN(n12390) );
  XNOR2_X1 U15460 ( .A(n12390), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14834) );
  AOI22_X1 U15461 ( .A1(n11843), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12392), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12393) );
  NAND2_X1 U15462 ( .A1(n14489), .A2(n20313), .ZN(n12402) );
  XNOR2_X1 U15463 ( .A(n12398), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13948) );
  INV_X1 U15464 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21082) );
  NOR2_X1 U15465 ( .A1(n10234), .A2(n21082), .ZN(n14829) );
  AOI21_X1 U15466 ( .B1(n20244), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14829), .ZN(n12399) );
  OAI21_X1 U15467 ( .B1(n20243), .B2(n13948), .A(n12399), .ZN(n12400) );
  INV_X1 U15468 ( .A(n12400), .ZN(n12401) );
  OAI211_X1 U15469 ( .C1(n14834), .C2(n20115), .A(n12402), .B(n12401), .ZN(
        P1_U2968) );
  NAND2_X1 U15470 ( .A1(n13764), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12403) );
  NAND2_X1 U15471 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19765) );
  NAND2_X1 U15472 ( .A1(n19765), .A2(n20088), .ZN(n12405) );
  NAND2_X1 U15473 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19925) );
  INV_X1 U15474 ( .A(n19925), .ZN(n12404) );
  NAND2_X1 U15475 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12404), .ZN(
        n12422) );
  NAND2_X1 U15476 ( .A1(n12405), .A2(n12422), .ZN(n19537) );
  NOR2_X1 U15477 ( .A1(n19537), .A2(n19860), .ZN(n12406) );
  AOI21_X1 U15478 ( .B1(n12424), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12406), .ZN(n12407) );
  OAI21_X1 U15479 ( .B1(n12408), .B2(n12426), .A(n12407), .ZN(n12412) );
  INV_X1 U15480 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12410) );
  NAND2_X1 U15481 ( .A1(n12413), .A2(n12420), .ZN(n13669) );
  INV_X1 U15482 ( .A(n12426), .ZN(n12414) );
  NAND2_X1 U15483 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20098), .ZN(
        n19699) );
  NAND2_X1 U15484 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20106), .ZN(
        n19734) );
  AND2_X1 U15485 ( .A1(n19699), .A2(n19734), .ZN(n19535) );
  NOR2_X1 U15486 ( .A1(n19860), .A2(n19535), .ZN(n19598) );
  AOI21_X1 U15487 ( .B1(n12424), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n19598), .ZN(n12415) );
  NOR2_X1 U15488 ( .A1(n19860), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12417) );
  AOI21_X1 U15489 ( .B1(n12424), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n12417), .ZN(n12418) );
  OAI21_X2 U15490 ( .B1(n15709), .B2(n12426), .A(n12418), .ZN(n13608) );
  OAI22_X1 U15491 ( .A1(n13601), .A2(n13602), .B1(n12419), .B2(n13608), .ZN(
        n13670) );
  INV_X1 U15492 ( .A(n19860), .ZN(n20069) );
  INV_X1 U15493 ( .A(n12422), .ZN(n12421) );
  NAND2_X1 U15494 ( .A1(n12421), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19933) );
  NAND2_X1 U15495 ( .A1(n20081), .A2(n12422), .ZN(n12423) );
  AND3_X1 U15496 ( .A1(n20069), .A2(n19933), .A3(n12423), .ZN(n19799) );
  AOI21_X1 U15497 ( .B1(n12424), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19799), .ZN(n12425) );
  NOR2_X1 U15498 ( .A1(n12594), .A2(n14118), .ZN(n13736) );
  INV_X1 U15499 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12429) );
  NAND4_X1 U15500 ( .A1(n13882), .A2(n19240), .A3(n19241), .A4(n13831), .ZN(
        n12430) );
  NAND2_X1 U15501 ( .A1(n14028), .A2(n14029), .ZN(n19232) );
  INV_X1 U15502 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12432) );
  INV_X1 U15503 ( .A(n12563), .ZN(n12522) );
  INV_X1 U15504 ( .A(n12562), .ZN(n12521) );
  INV_X1 U15505 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12431) );
  OAI22_X1 U15506 ( .A1(n12432), .A2(n12522), .B1(n12521), .B2(n12431), .ZN(
        n12444) );
  AOI22_X1 U15507 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12436) );
  AOI22_X1 U15508 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10612), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12435) );
  AOI22_X1 U15509 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10534), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12434) );
  AOI22_X1 U15510 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n10542), .B1(
        n12557), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12433) );
  NAND4_X1 U15511 ( .A1(n12436), .A2(n12435), .A3(n12434), .A4(n12433), .ZN(
        n12443) );
  INV_X1 U15512 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12438) );
  INV_X1 U15513 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12437) );
  OAI22_X1 U15514 ( .A1(n12531), .A2(n12438), .B1(n12529), .B2(n12437), .ZN(
        n12442) );
  INV_X1 U15515 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n19744) );
  AOI22_X1 U15516 ( .A1(n12565), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__0__SCAN_IN), .B2(n12564), .ZN(n12440) );
  NAND2_X1 U15517 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12439) );
  OAI211_X1 U15518 ( .C1(n13749), .C2(n19744), .A(n12440), .B(n12439), .ZN(
        n12441) );
  NOR4_X1 U15519 ( .A1(n12444), .A2(n12443), .A3(n12442), .A4(n12441), .ZN(
        n19233) );
  NOR2_X2 U15520 ( .A1(n19232), .A2(n19233), .ZN(n14346) );
  AOI22_X1 U15521 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12448) );
  AOI22_X1 U15522 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10612), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12447) );
  AOI22_X1 U15523 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10534), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12446) );
  AOI22_X1 U15524 ( .A1(n10542), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n12557), .ZN(n12445) );
  NAND4_X1 U15525 ( .A1(n12448), .A2(n12447), .A3(n12446), .A4(n12445), .ZN(
        n12459) );
  AOI22_X1 U15526 ( .A1(n12565), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n12564), .ZN(n12450) );
  NAND2_X1 U15527 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12449) );
  OAI211_X1 U15528 ( .C1(n13749), .C2(n12451), .A(n12450), .B(n12449), .ZN(
        n12458) );
  INV_X1 U15529 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12452) );
  OAI22_X1 U15530 ( .A1(n12529), .A2(n12453), .B1(n12531), .B2(n12452), .ZN(
        n12457) );
  OAI22_X1 U15531 ( .A1(n12522), .A2(n12455), .B1(n12521), .B2(n12454), .ZN(
        n12456) );
  NAND2_X1 U15532 ( .A1(n14346), .A2(n14350), .ZN(n14348) );
  INV_X1 U15533 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12461) );
  INV_X1 U15534 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12460) );
  OAI22_X1 U15535 ( .A1(n12461), .A2(n12522), .B1(n12521), .B2(n12460), .ZN(
        n12474) );
  AOI22_X1 U15536 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12465) );
  AOI22_X1 U15537 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10612), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12464) );
  AOI22_X1 U15538 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10534), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12463) );
  AOI22_X1 U15539 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n10542), .B1(
        n12557), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12462) );
  NAND4_X1 U15540 ( .A1(n12465), .A2(n12464), .A3(n12463), .A4(n12462), .ZN(
        n12473) );
  INV_X1 U15541 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12467) );
  INV_X1 U15542 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12466) );
  OAI22_X1 U15543 ( .A1(n12531), .A2(n12467), .B1(n12529), .B2(n12466), .ZN(
        n12472) );
  INV_X1 U15544 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12470) );
  AOI22_X1 U15545 ( .A1(n12565), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__2__SCAN_IN), .B2(n12564), .ZN(n12469) );
  NAND2_X1 U15546 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n12468) );
  OAI211_X1 U15547 ( .C1(n13749), .C2(n12470), .A(n12469), .B(n12468), .ZN(
        n12471) );
  NOR4_X1 U15548 ( .A1(n12474), .A2(n12473), .A3(n12472), .A4(n12471), .ZN(
        n16344) );
  AOI22_X1 U15549 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12478) );
  AOI22_X1 U15550 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10612), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12477) );
  AOI22_X1 U15551 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10534), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12476) );
  AOI22_X1 U15552 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n10542), .B1(
        n12557), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12475) );
  NAND4_X1 U15553 ( .A1(n12478), .A2(n12477), .A3(n12476), .A4(n12475), .ZN(
        n12489) );
  AOI22_X1 U15554 ( .A1(n12565), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__3__SCAN_IN), .B2(n12564), .ZN(n12480) );
  NAND2_X1 U15555 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n12479) );
  OAI211_X1 U15556 ( .C1(n13749), .C2(n12481), .A(n12480), .B(n12479), .ZN(
        n12488) );
  INV_X1 U15557 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12483) );
  OAI22_X1 U15558 ( .A1(n12531), .A2(n12483), .B1(n12529), .B2(n12482), .ZN(
        n12487) );
  INV_X1 U15559 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12484) );
  OAI22_X1 U15560 ( .A1(n12485), .A2(n12522), .B1(n12521), .B2(n12484), .ZN(
        n12486) );
  INV_X1 U15561 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12491) );
  INV_X1 U15562 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12490) );
  OAI22_X1 U15563 ( .A1(n12491), .A2(n12522), .B1(n12521), .B2(n12490), .ZN(
        n12504) );
  AOI22_X1 U15564 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12495) );
  AOI22_X1 U15565 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10612), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12494) );
  AOI22_X1 U15566 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10534), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12493) );
  AOI22_X1 U15567 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n10542), .B1(
        n12557), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12492) );
  NAND4_X1 U15568 ( .A1(n12495), .A2(n12494), .A3(n12493), .A4(n12492), .ZN(
        n12503) );
  INV_X1 U15569 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12497) );
  INV_X1 U15570 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12496) );
  OAI22_X1 U15571 ( .A1(n12531), .A2(n12497), .B1(n12529), .B2(n12496), .ZN(
        n12502) );
  INV_X1 U15572 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12500) );
  AOI22_X1 U15573 ( .A1(n12565), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__4__SCAN_IN), .B2(n12564), .ZN(n12499) );
  NAND2_X1 U15574 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12498) );
  OAI211_X1 U15575 ( .C1(n13749), .C2(n12500), .A(n12499), .B(n12498), .ZN(
        n12501) );
  NOR4_X1 U15576 ( .A1(n12504), .A2(n12503), .A3(n12502), .A4(n12501), .ZN(
        n16342) );
  AOI22_X1 U15577 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12508) );
  AOI22_X1 U15578 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10612), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12507) );
  AOI22_X1 U15579 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10534), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12506) );
  AOI22_X1 U15580 ( .A1(n10542), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_7__5__SCAN_IN), .B2(n12557), .ZN(n12505) );
  NAND4_X1 U15581 ( .A1(n12508), .A2(n12507), .A3(n12506), .A4(n12505), .ZN(
        n12519) );
  INV_X1 U15582 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12511) );
  AOI22_X1 U15583 ( .A1(n12565), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__5__SCAN_IN), .B2(n12564), .ZN(n12510) );
  NAND2_X1 U15584 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n12509) );
  OAI211_X1 U15585 ( .C1(n13749), .C2(n12511), .A(n12510), .B(n12509), .ZN(
        n12518) );
  INV_X1 U15586 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12513) );
  INV_X1 U15587 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12512) );
  OAI22_X1 U15588 ( .A1(n12531), .A2(n12513), .B1(n12529), .B2(n12512), .ZN(
        n12517) );
  INV_X1 U15589 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12515) );
  INV_X1 U15590 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12514) );
  OAI22_X1 U15591 ( .A1(n12515), .A2(n12522), .B1(n12521), .B2(n12514), .ZN(
        n12516) );
  INV_X1 U15592 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12523) );
  INV_X1 U15593 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12520) );
  OAI22_X1 U15594 ( .A1(n12523), .A2(n12522), .B1(n12521), .B2(n12520), .ZN(
        n12538) );
  AOI22_X1 U15595 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12527) );
  AOI22_X1 U15596 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10612), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12526) );
  AOI22_X1 U15597 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10534), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12525) );
  AOI22_X1 U15598 ( .A1(n10542), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_7__6__SCAN_IN), .B2(n12557), .ZN(n12524) );
  NAND4_X1 U15599 ( .A1(n12527), .A2(n12526), .A3(n12525), .A4(n12524), .ZN(
        n12537) );
  INV_X1 U15600 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12530) );
  INV_X1 U15601 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12528) );
  OAI22_X1 U15602 ( .A1(n12531), .A2(n12530), .B1(n12529), .B2(n12528), .ZN(
        n12536) );
  AOI22_X1 U15603 ( .A1(n12565), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__6__SCAN_IN), .B2(n12564), .ZN(n12533) );
  NAND2_X1 U15604 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12532) );
  OAI211_X1 U15605 ( .C1(n13749), .C2(n12534), .A(n12533), .B(n12532), .ZN(
        n12535) );
  NOR4_X1 U15606 ( .A1(n12538), .A2(n12537), .A3(n12536), .A4(n12535), .ZN(
        n16339) );
  AOI22_X1 U15607 ( .A1(n9684), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(n9652), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12546) );
  AOI22_X1 U15608 ( .A1(n10481), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12545) );
  AOI22_X1 U15609 ( .A1(n9685), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12544) );
  NAND2_X1 U15610 ( .A1(n9649), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12542) );
  NAND2_X1 U15611 ( .A1(n12686), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12541) );
  NAND2_X1 U15612 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12540) );
  NAND2_X1 U15613 ( .A1(n12540), .A2(n12539), .ZN(n13248) );
  AND3_X1 U15614 ( .A1(n12542), .A2(n12541), .A3(n13248), .ZN(n12543) );
  NAND4_X1 U15615 ( .A1(n12546), .A2(n12545), .A3(n12544), .A4(n12543), .ZN(
        n12554) );
  AOI22_X1 U15616 ( .A1(n9680), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9652), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12552) );
  AOI22_X1 U15617 ( .A1(n9685), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12551) );
  AOI22_X1 U15618 ( .A1(n10481), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12550) );
  NAND2_X1 U15619 ( .A1(n12587), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12548) );
  NAND2_X1 U15620 ( .A1(n12686), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12547) );
  INV_X1 U15621 ( .A(n13248), .ZN(n13239) );
  AND3_X1 U15622 ( .A1(n12548), .A2(n12547), .A3(n13239), .ZN(n12549) );
  NAND4_X1 U15623 ( .A1(n12552), .A2(n12551), .A3(n12550), .A4(n12549), .ZN(
        n12553) );
  NAND2_X1 U15624 ( .A1(n9676), .A2(n12597), .ZN(n12576) );
  AOI22_X1 U15625 ( .A1(n9659), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12555), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12561) );
  AOI22_X1 U15626 ( .A1(n10519), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10612), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12560) );
  AOI22_X1 U15627 ( .A1(n12556), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10562), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12559) );
  AOI22_X1 U15628 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n10542), .B1(
        n12557), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12558) );
  NAND4_X1 U15629 ( .A1(n12561), .A2(n12560), .A3(n12559), .A4(n12558), .ZN(
        n12575) );
  AOI22_X1 U15630 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n12563), .B1(
        n12562), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12573) );
  AOI22_X1 U15631 ( .A1(n12565), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n12564), .ZN(n12567) );
  NAND2_X1 U15632 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12566) );
  AND2_X1 U15633 ( .A1(n12567), .A2(n12566), .ZN(n12572) );
  AOI22_X1 U15634 ( .A1(n12569), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12568), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12571) );
  NAND2_X1 U15635 ( .A1(n10534), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12570) );
  NAND4_X1 U15636 ( .A1(n12573), .A2(n12572), .A3(n12571), .A4(n12570), .ZN(
        n12574) );
  OR2_X1 U15637 ( .A1(n12575), .A2(n12574), .ZN(n12578) );
  XNOR2_X1 U15638 ( .A(n12576), .B(n12578), .ZN(n12600) );
  NAND2_X1 U15639 ( .A1(n9666), .A2(n12597), .ZN(n15229) );
  NAND2_X1 U15640 ( .A1(n12578), .A2(n12597), .ZN(n12603) );
  NAND2_X1 U15641 ( .A1(n10481), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12580) );
  AOI21_X1 U15642 ( .B1(n12686), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A(
        n13239), .ZN(n12579) );
  AND2_X1 U15643 ( .A1(n12580), .A2(n12579), .ZN(n12584) );
  AOI22_X1 U15644 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n9683), .B1(n9652), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12583) );
  AOI22_X1 U15645 ( .A1(n9685), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(n9649), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12582) );
  AOI22_X1 U15646 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12587), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12581) );
  NAND4_X1 U15647 ( .A1(n12584), .A2(n12583), .A3(n12582), .A4(n12581), .ZN(
        n12593) );
  NAND2_X1 U15648 ( .A1(n10481), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12586) );
  AOI21_X1 U15649 ( .B1(n12686), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n13248), .ZN(n12585) );
  AND2_X1 U15650 ( .A1(n12586), .A2(n12585), .ZN(n12591) );
  AOI22_X1 U15651 ( .A1(n9681), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9652), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12590) );
  AOI22_X1 U15652 ( .A1(n9685), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12589) );
  AOI22_X1 U15653 ( .A1(n12587), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12588) );
  NAND4_X1 U15654 ( .A1(n12591), .A2(n12590), .A3(n12589), .A4(n12588), .ZN(
        n12592) );
  NAND2_X1 U15655 ( .A1(n12593), .A2(n12592), .ZN(n12602) );
  XOR2_X1 U15656 ( .A(n12603), .B(n12602), .Z(n12595) );
  INV_X1 U15657 ( .A(n12594), .ZN(n13769) );
  NAND2_X1 U15658 ( .A1(n12595), .A2(n13769), .ZN(n15166) );
  INV_X1 U15659 ( .A(n12602), .ZN(n12596) );
  NAND2_X1 U15660 ( .A1(n9666), .A2(n12596), .ZN(n15167) );
  INV_X1 U15661 ( .A(n12597), .ZN(n12598) );
  NOR2_X1 U15662 ( .A1(n15167), .A2(n12598), .ZN(n12599) );
  NOR2_X1 U15663 ( .A1(n12603), .A2(n12602), .ZN(n12618) );
  AOI22_X1 U15664 ( .A1(n9685), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10481), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12609) );
  INV_X1 U15665 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n19888) );
  AOI22_X1 U15666 ( .A1(n9681), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9652), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12608) );
  AOI22_X1 U15667 ( .A1(n12587), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12607) );
  NAND2_X1 U15668 ( .A1(n9649), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12605) );
  NAND2_X1 U15669 ( .A1(n12686), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12604) );
  AND3_X1 U15670 ( .A1(n12605), .A2(n12604), .A3(n13239), .ZN(n12606) );
  NAND4_X1 U15671 ( .A1(n12609), .A2(n12608), .A3(n12607), .A4(n12606), .ZN(
        n12617) );
  NAND2_X1 U15672 ( .A1(n9685), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12611) );
  AOI21_X1 U15673 ( .B1(n12686), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n13239), .ZN(n12610) );
  AND2_X1 U15674 ( .A1(n12611), .A2(n12610), .ZN(n12615) );
  AOI22_X1 U15675 ( .A1(n9682), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(n9652), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12614) );
  AOI22_X1 U15676 ( .A1(n10481), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12613) );
  AOI22_X1 U15677 ( .A1(n12587), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12612) );
  NAND4_X1 U15678 ( .A1(n12615), .A2(n12614), .A3(n12613), .A4(n12612), .ZN(
        n12616) );
  AND2_X1 U15679 ( .A1(n12617), .A2(n12616), .ZN(n12619) );
  NAND2_X1 U15680 ( .A1(n12618), .A2(n12619), .ZN(n12659) );
  OAI211_X1 U15681 ( .C1(n12618), .C2(n12619), .A(n13769), .B(n12659), .ZN(
        n12622) );
  XNOR2_X1 U15682 ( .A(n12621), .B(n12623), .ZN(n15159) );
  INV_X1 U15683 ( .A(n12619), .ZN(n12620) );
  NOR2_X1 U15684 ( .A1(n9676), .A2(n12620), .ZN(n15162) );
  NAND2_X1 U15685 ( .A1(n15159), .A2(n15162), .ZN(n15161) );
  INV_X1 U15686 ( .A(n12621), .ZN(n12624) );
  NAND2_X1 U15687 ( .A1(n15161), .A2(n12625), .ZN(n12641) );
  NAND2_X1 U15688 ( .A1(n10481), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12627) );
  AOI21_X1 U15689 ( .B1(n12686), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A(
        n13239), .ZN(n12626) );
  AND2_X1 U15690 ( .A1(n12627), .A2(n12626), .ZN(n12631) );
  AOI22_X1 U15691 ( .A1(n9683), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n9652), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12630) );
  AOI22_X1 U15692 ( .A1(n9685), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(n9649), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12629) );
  AOI22_X1 U15693 ( .A1(n12587), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12628) );
  NAND4_X1 U15694 ( .A1(n12631), .A2(n12630), .A3(n12629), .A4(n12628), .ZN(
        n12639) );
  NAND2_X1 U15695 ( .A1(n10481), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12633) );
  AOI21_X1 U15696 ( .B1(n12686), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A(
        n13248), .ZN(n12632) );
  AND2_X1 U15697 ( .A1(n12633), .A2(n12632), .ZN(n12637) );
  AOI22_X1 U15698 ( .A1(n9683), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9652), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12636) );
  AOI22_X1 U15699 ( .A1(n9685), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12635) );
  AOI22_X1 U15700 ( .A1(n12587), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12634) );
  NAND4_X1 U15701 ( .A1(n12637), .A2(n12636), .A3(n12635), .A4(n12634), .ZN(
        n12638) );
  AND2_X1 U15702 ( .A1(n12639), .A2(n12638), .ZN(n12657) );
  XNOR2_X1 U15703 ( .A(n12659), .B(n12657), .ZN(n12640) );
  XNOR2_X1 U15704 ( .A(n12641), .B(n10233), .ZN(n15156) );
  NAND2_X1 U15705 ( .A1(n9666), .A2(n12657), .ZN(n15155) );
  NAND2_X1 U15706 ( .A1(n10481), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12644) );
  AOI21_X1 U15707 ( .B1(n12686), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A(
        n13239), .ZN(n12643) );
  AND2_X1 U15708 ( .A1(n12644), .A2(n12643), .ZN(n12648) );
  AOI22_X1 U15709 ( .A1(n9684), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(n9652), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12647) );
  AOI22_X1 U15710 ( .A1(n9685), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n9649), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12646) );
  AOI22_X1 U15711 ( .A1(n12587), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12645) );
  NAND4_X1 U15712 ( .A1(n12648), .A2(n12647), .A3(n12646), .A4(n12645), .ZN(
        n12656) );
  NAND2_X1 U15713 ( .A1(n10481), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12650) );
  AOI21_X1 U15714 ( .B1(n12686), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n13248), .ZN(n12649) );
  AND2_X1 U15715 ( .A1(n12650), .A2(n12649), .ZN(n12654) );
  AOI22_X1 U15716 ( .A1(n9683), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9652), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12653) );
  AOI22_X1 U15717 ( .A1(n9685), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12652) );
  AOI22_X1 U15718 ( .A1(n12587), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12651) );
  NAND4_X1 U15719 ( .A1(n12654), .A2(n12653), .A3(n12652), .A4(n12651), .ZN(
        n12655) );
  NAND2_X1 U15720 ( .A1(n12656), .A2(n12655), .ZN(n12660) );
  INV_X1 U15721 ( .A(n12660), .ZN(n12665) );
  INV_X1 U15722 ( .A(n12657), .ZN(n12658) );
  OR2_X1 U15723 ( .A1(n12659), .A2(n12658), .ZN(n12661) );
  INV_X1 U15724 ( .A(n12661), .ZN(n12662) );
  OR2_X1 U15725 ( .A1(n12661), .A2(n12660), .ZN(n15139) );
  OAI211_X1 U15726 ( .C1(n12665), .C2(n12662), .A(n15139), .B(n13769), .ZN(
        n12663) );
  NAND2_X1 U15727 ( .A1(n9666), .A2(n12665), .ZN(n15146) );
  NAND2_X1 U15728 ( .A1(n10481), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12667) );
  AOI21_X1 U15729 ( .B1(n12686), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n13239), .ZN(n12666) );
  AND2_X1 U15730 ( .A1(n12667), .A2(n12666), .ZN(n12671) );
  AOI22_X1 U15731 ( .A1(n9681), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(n9652), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12670) );
  AOI22_X1 U15732 ( .A1(n9685), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n9649), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12669) );
  AOI22_X1 U15733 ( .A1(n12587), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12668) );
  NAND4_X1 U15734 ( .A1(n12671), .A2(n12670), .A3(n12669), .A4(n12668), .ZN(
        n12679) );
  NAND2_X1 U15735 ( .A1(n10481), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12673) );
  AOI21_X1 U15736 ( .B1(n12686), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n13248), .ZN(n12672) );
  AND2_X1 U15737 ( .A1(n12673), .A2(n12672), .ZN(n12677) );
  AOI22_X1 U15738 ( .A1(n9680), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9652), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12676) );
  AOI22_X1 U15739 ( .A1(n9685), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12675) );
  AOI22_X1 U15740 ( .A1(n12587), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12674) );
  NAND4_X1 U15741 ( .A1(n12677), .A2(n12676), .A3(n12675), .A4(n12674), .ZN(
        n12678) );
  AND2_X1 U15742 ( .A1(n12679), .A2(n12678), .ZN(n15141) );
  NAND2_X1 U15743 ( .A1(n10481), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n12681) );
  AOI21_X1 U15744 ( .B1(n12686), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n13239), .ZN(n12680) );
  AND2_X1 U15745 ( .A1(n12681), .A2(n12680), .ZN(n12685) );
  AOI22_X1 U15746 ( .A1(n9682), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(n9652), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12684) );
  AOI22_X1 U15747 ( .A1(n9685), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12683) );
  AOI22_X1 U15748 ( .A1(n12587), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12682) );
  NAND4_X1 U15749 ( .A1(n12685), .A2(n12684), .A3(n12683), .A4(n12682), .ZN(
        n12694) );
  NAND2_X1 U15750 ( .A1(n10481), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12688) );
  AOI21_X1 U15751 ( .B1(n12686), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n13248), .ZN(n12687) );
  AND2_X1 U15752 ( .A1(n12688), .A2(n12687), .ZN(n12692) );
  AOI22_X1 U15753 ( .A1(n9681), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9652), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12691) );
  AOI22_X1 U15754 ( .A1(n9685), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12690) );
  AOI22_X1 U15755 ( .A1(n12587), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12689) );
  NAND4_X1 U15756 ( .A1(n12692), .A2(n12691), .A3(n12690), .A4(n12689), .ZN(
        n12693) );
  AND2_X1 U15757 ( .A1(n12694), .A2(n12693), .ZN(n12697) );
  NAND2_X1 U15758 ( .A1(n9676), .A2(n15141), .ZN(n12695) );
  NOR2_X1 U15759 ( .A1(n15139), .A2(n12695), .ZN(n12696) );
  NAND2_X1 U15760 ( .A1(n12696), .A2(n12697), .ZN(n13236) );
  OAI21_X1 U15761 ( .B1(n12697), .B2(n12696), .A(n13236), .ZN(n12698) );
  NAND2_X1 U15762 ( .A1(n12699), .A2(n12698), .ZN(n14446) );
  INV_X1 U15763 ( .A(n13261), .ZN(n14055) );
  INV_X1 U15764 ( .A(n14052), .ZN(n13746) );
  NAND2_X1 U15765 ( .A1(n14055), .A2(n13746), .ZN(n13480) );
  NAND2_X1 U15766 ( .A1(n14066), .A2(n12700), .ZN(n13753) );
  NAND2_X1 U15767 ( .A1(n13480), .A2(n13753), .ZN(n12701) );
  NAND2_X1 U15768 ( .A1(n19252), .A2(n13279), .ZN(n19254) );
  OR2_X1 U15769 ( .A1(n12347), .A2(n12702), .ZN(n12703) );
  NAND2_X1 U15770 ( .A1(n12704), .A2(n12703), .ZN(n16309) );
  NAND2_X1 U15771 ( .A1(n19259), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12705) );
  INV_X1 U15772 ( .A(n16063), .ZN(n14755) );
  INV_X1 U15773 ( .A(n12711), .ZN(n12710) );
  NOR4_X1 U15774 ( .A1(n12708), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12709) );
  NAND2_X1 U15775 ( .A1(n12710), .A2(n12709), .ZN(n12712) );
  INV_X1 U15776 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n12713) );
  NAND2_X1 U15777 ( .A1(n12714), .A2(n12713), .ZN(n15925) );
  INV_X1 U15778 ( .A(n15925), .ZN(n13916) );
  NAND2_X1 U15779 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20892) );
  OAI21_X1 U15780 ( .B1(n13943), .B2(n13916), .A(n20892), .ZN(n13942) );
  INV_X1 U15781 ( .A(n13942), .ZN(n12715) );
  NAND2_X1 U15782 ( .A1(n13676), .A2(n12715), .ZN(n12716) );
  NAND3_X1 U15783 ( .A1(n12716), .A2(n13918), .A3(n13821), .ZN(n12717) );
  NAND2_X1 U15784 ( .A1(n12717), .A2(n14477), .ZN(n12727) );
  NOR4_X1 U15785 ( .A1(n12721), .A2(n12720), .A3(n12719), .A4(n12718), .ZN(
        n12722) );
  OR2_X1 U15786 ( .A1(n12723), .A2(n12722), .ZN(n14473) );
  NAND2_X1 U15787 ( .A1(n13943), .A2(n15925), .ZN(n12724) );
  NAND2_X1 U15788 ( .A1(n12724), .A2(n20892), .ZN(n12725) );
  OR2_X1 U15789 ( .A1(n14473), .A2(n12725), .ZN(n12726) );
  MUX2_X1 U15790 ( .A(n12727), .B(n12726), .S(n13629), .Z(n12734) );
  INV_X1 U15791 ( .A(n12728), .ZN(n12737) );
  OAI21_X1 U15792 ( .B1(n20969), .B2(n12856), .A(n12859), .ZN(n12729) );
  NAND2_X1 U15793 ( .A1(n12737), .A2(n12729), .ZN(n12732) );
  NOR2_X1 U15794 ( .A1(n12849), .A2(n13918), .ZN(n12730) );
  NAND2_X1 U15795 ( .A1(n12731), .A2(n12730), .ZN(n14472) );
  NAND2_X1 U15796 ( .A1(n12732), .A2(n14472), .ZN(n13628) );
  INV_X1 U15797 ( .A(n14477), .ZN(n15911) );
  NOR2_X1 U15798 ( .A1(n15877), .A2(n20326), .ZN(n12853) );
  NAND2_X1 U15799 ( .A1(n15911), .A2(n12853), .ZN(n12733) );
  NAND3_X1 U15800 ( .A1(n12734), .A2(n13628), .A3(n12733), .ZN(n12735) );
  INV_X1 U15801 ( .A(n12736), .ZN(n12738) );
  NAND2_X1 U15802 ( .A1(n12737), .A2(n11512), .ZN(n13691) );
  AND2_X1 U15803 ( .A1(n12738), .A2(n13691), .ZN(n14478) );
  OAI211_X1 U15804 ( .C1(n20347), .C2(n12846), .A(n14478), .B(n12739), .ZN(
        n12740) );
  INV_X1 U15805 ( .A(n12864), .ZN(n13361) );
  NAND2_X1 U15806 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14485), .ZN(
        n12743) );
  AND2_X1 U15807 ( .A1(n12820), .A2(n12743), .ZN(n12744) );
  NAND2_X1 U15808 ( .A1(n12745), .A2(n12744), .ZN(n12749) );
  NAND2_X1 U15809 ( .A1(n9674), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12748) );
  INV_X1 U15810 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n12746) );
  NAND2_X1 U15811 ( .A1(n12864), .A2(n12746), .ZN(n12747) );
  NAND2_X1 U15812 ( .A1(n12748), .A2(n12747), .ZN(n13797) );
  XNOR2_X1 U15813 ( .A(n12749), .B(n13797), .ZN(n13984) );
  INV_X1 U15814 ( .A(n12749), .ZN(n12750) );
  AOI21_X1 U15815 ( .B1(n13984), .B2(n13357), .A(n12750), .ZN(n13901) );
  OR2_X1 U15816 ( .A1(n12840), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n12754) );
  NAND2_X1 U15817 ( .A1(n9674), .A2(n20282), .ZN(n12752) );
  INV_X1 U15818 ( .A(n13361), .ZN(n12780) );
  INV_X1 U15819 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13953) );
  NAND2_X1 U15820 ( .A1(n13357), .A2(n13953), .ZN(n12751) );
  NAND3_X1 U15821 ( .A1(n12752), .A2(n12780), .A3(n12751), .ZN(n12753) );
  NAND2_X1 U15822 ( .A1(n12754), .A2(n12753), .ZN(n13900) );
  NAND2_X1 U15823 ( .A1(n13901), .A2(n13900), .ZN(n13927) );
  NAND2_X1 U15824 ( .A1(n13357), .A2(n12864), .ZN(n12832) );
  INV_X1 U15825 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n12755) );
  NAND2_X1 U15826 ( .A1(n13357), .A2(n12755), .ZN(n12757) );
  NAND2_X1 U15827 ( .A1(n12864), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12756) );
  NAND3_X1 U15828 ( .A1(n12757), .A2(n9674), .A3(n12756), .ZN(n12758) );
  OAI21_X1 U15829 ( .B1(n12832), .B2(P1_EBX_REG_3__SCAN_IN), .A(n12758), .ZN(
        n13926) );
  MUX2_X1 U15830 ( .A(n12832), .B(n12780), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n12759) );
  OAI21_X1 U15831 ( .B1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n14486), .A(
        n12759), .ZN(n12760) );
  INV_X1 U15832 ( .A(n12760), .ZN(n13965) );
  OR2_X1 U15833 ( .A1(n12840), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n12765) );
  NAND2_X1 U15834 ( .A1(n9674), .A2(n12761), .ZN(n12763) );
  INV_X1 U15835 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n20191) );
  NAND2_X1 U15836 ( .A1(n13357), .A2(n20191), .ZN(n12762) );
  NAND3_X1 U15837 ( .A1(n12763), .A2(n12780), .A3(n12762), .ZN(n12764) );
  NAND2_X1 U15838 ( .A1(n12765), .A2(n12764), .ZN(n13966) );
  NAND2_X1 U15839 ( .A1(n13965), .A2(n13966), .ZN(n12766) );
  OR2_X1 U15840 ( .A1(n12840), .A2(P1_EBX_REG_6__SCAN_IN), .ZN(n12770) );
  NAND2_X1 U15841 ( .A1(n9674), .A2(n16126), .ZN(n12768) );
  INV_X1 U15842 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n13999) );
  NAND2_X1 U15843 ( .A1(n13357), .A2(n13999), .ZN(n12767) );
  NAND3_X1 U15844 ( .A1(n12768), .A2(n12780), .A3(n12767), .ZN(n12769) );
  NAND2_X1 U15845 ( .A1(n12770), .A2(n12769), .ZN(n13997) );
  INV_X1 U15846 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n20143) );
  NAND2_X1 U15847 ( .A1(n12835), .A2(n20143), .ZN(n12774) );
  NAND2_X1 U15848 ( .A1(n13357), .A2(n20143), .ZN(n12772) );
  NAND2_X1 U15849 ( .A1(n12780), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12771) );
  NAND3_X1 U15850 ( .A1(n12772), .A2(n9674), .A3(n12771), .ZN(n12773) );
  AND2_X1 U15851 ( .A1(n12774), .A2(n12773), .ZN(n14095) );
  OR2_X1 U15852 ( .A1(n12840), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n12779) );
  NAND2_X1 U15853 ( .A1(n9674), .A2(n14332), .ZN(n12777) );
  INV_X1 U15854 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n12775) );
  NAND2_X1 U15855 ( .A1(n13357), .A2(n12775), .ZN(n12776) );
  NAND3_X1 U15856 ( .A1(n12777), .A2(n12864), .A3(n12776), .ZN(n12778) );
  MUX2_X1 U15857 ( .A(n12832), .B(n12780), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n12781) );
  OAI21_X1 U15858 ( .B1(n14486), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n12781), .ZN(n14269) );
  MUX2_X1 U15859 ( .A(n12840), .B(n9674), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n12784) );
  NAND2_X1 U15860 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n14485), .ZN(
        n12782) );
  AND2_X1 U15861 ( .A1(n12820), .A2(n12782), .ZN(n12783) );
  NAND2_X1 U15862 ( .A1(n12784), .A2(n12783), .ZN(n14366) );
  INV_X1 U15863 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14369) );
  NAND2_X1 U15864 ( .A1(n12835), .A2(n14369), .ZN(n12788) );
  NAND2_X1 U15865 ( .A1(n13357), .A2(n14369), .ZN(n12786) );
  NAND2_X1 U15866 ( .A1(n12780), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12785) );
  NAND3_X1 U15867 ( .A1(n12786), .A2(n9674), .A3(n12785), .ZN(n12787) );
  AND2_X1 U15868 ( .A1(n12788), .A2(n12787), .ZN(n14365) );
  NAND2_X1 U15869 ( .A1(n14366), .A2(n14365), .ZN(n12789) );
  MUX2_X1 U15870 ( .A(n12840), .B(n9674), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n12792) );
  NAND2_X1 U15871 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14485), .ZN(
        n12790) );
  AND2_X1 U15872 ( .A1(n12820), .A2(n12790), .ZN(n12791) );
  NAND2_X1 U15873 ( .A1(n12792), .A2(n12791), .ZN(n14402) );
  INV_X1 U15874 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14392) );
  NAND2_X1 U15875 ( .A1(n12835), .A2(n14392), .ZN(n12796) );
  NAND2_X1 U15876 ( .A1(n13357), .A2(n14392), .ZN(n12794) );
  NAND2_X1 U15877 ( .A1(n12780), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12793) );
  NAND3_X1 U15878 ( .A1(n12794), .A2(n9674), .A3(n12793), .ZN(n12795) );
  AND2_X1 U15879 ( .A1(n12796), .A2(n12795), .ZN(n14384) );
  MUX2_X1 U15880 ( .A(n12832), .B(n12780), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12798) );
  OAI21_X1 U15881 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n14486), .A(
        n12798), .ZN(n12799) );
  INV_X1 U15882 ( .A(n12799), .ZN(n14647) );
  MUX2_X1 U15883 ( .A(n12840), .B(n9674), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n12802) );
  NAND2_X1 U15884 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n14485), .ZN(
        n12800) );
  AND2_X1 U15885 ( .A1(n12820), .A2(n12800), .ZN(n12801) );
  NAND2_X1 U15886 ( .A1(n12802), .A2(n12801), .ZN(n14648) );
  MUX2_X1 U15887 ( .A(n12840), .B(n9674), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n12804) );
  NAND2_X1 U15888 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n14485), .ZN(
        n12803) );
  MUX2_X1 U15889 ( .A(n12832), .B(n12780), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n12805) );
  OAI21_X1 U15890 ( .B1(n14486), .B2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n12805), .ZN(n12806) );
  INV_X1 U15891 ( .A(n12806), .ZN(n14634) );
  MUX2_X1 U15892 ( .A(n12840), .B(n12742), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n12809) );
  NAND2_X1 U15893 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n14485), .ZN(
        n12807) );
  AND2_X1 U15894 ( .A1(n12820), .A2(n12807), .ZN(n12808) );
  NAND2_X1 U15895 ( .A1(n12809), .A2(n12808), .ZN(n14626) );
  INV_X1 U15896 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n16002) );
  NAND2_X1 U15897 ( .A1(n13357), .A2(n16002), .ZN(n12811) );
  NAND2_X1 U15898 ( .A1(n12780), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12810) );
  NAND3_X1 U15899 ( .A1(n12811), .A2(n12742), .A3(n12810), .ZN(n12812) );
  OAI21_X1 U15900 ( .B1(n12832), .B2(P1_EBX_REG_19__SCAN_IN), .A(n12812), .ZN(
        n14622) );
  MUX2_X1 U15901 ( .A(n12840), .B(n9674), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n12814) );
  NAND2_X1 U15902 ( .A1(n14485), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12813) );
  AND3_X1 U15903 ( .A1(n12814), .A2(n12820), .A3(n12813), .ZN(n14614) );
  INV_X1 U15904 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15984) );
  NAND2_X1 U15905 ( .A1(n12835), .A2(n15984), .ZN(n12818) );
  NAND2_X1 U15906 ( .A1(n13357), .A2(n15984), .ZN(n12816) );
  NAND2_X1 U15907 ( .A1(n12864), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12815) );
  NAND3_X1 U15908 ( .A1(n12816), .A2(n9674), .A3(n12815), .ZN(n12817) );
  AND2_X1 U15909 ( .A1(n12818), .A2(n12817), .ZN(n14609) );
  MUX2_X1 U15910 ( .A(n12840), .B(n9674), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n12822) );
  NAND2_X1 U15911 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n14485), .ZN(
        n12819) );
  AND2_X1 U15912 ( .A1(n12820), .A2(n12819), .ZN(n12821) );
  NAND2_X1 U15913 ( .A1(n12822), .A2(n12821), .ZN(n14601) );
  INV_X1 U15914 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n12823) );
  NAND2_X1 U15915 ( .A1(n13357), .A2(n12823), .ZN(n12825) );
  NAND2_X1 U15916 ( .A1(n12780), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12824) );
  NAND3_X1 U15917 ( .A1(n12825), .A2(n12742), .A3(n12824), .ZN(n12826) );
  OAI21_X1 U15918 ( .B1(n12832), .B2(P1_EBX_REG_23__SCAN_IN), .A(n12826), .ZN(
        n14556) );
  MUX2_X1 U15919 ( .A(n12840), .B(n9674), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n12828) );
  NAND2_X1 U15920 ( .A1(n14485), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12827) );
  AND2_X1 U15921 ( .A1(n12828), .A2(n12827), .ZN(n14595) );
  INV_X1 U15922 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14590) );
  NAND2_X1 U15923 ( .A1(n13357), .A2(n14590), .ZN(n12830) );
  NAND2_X1 U15924 ( .A1(n12780), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12829) );
  NAND3_X1 U15925 ( .A1(n12830), .A2(n12742), .A3(n12829), .ZN(n12831) );
  OAI21_X1 U15926 ( .B1(n12832), .B2(P1_EBX_REG_25__SCAN_IN), .A(n12831), .ZN(
        n14587) );
  MUX2_X1 U15927 ( .A(n12840), .B(n9674), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n12834) );
  NAND2_X1 U15928 ( .A1(n14485), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12833) );
  NAND2_X1 U15929 ( .A1(n12834), .A2(n12833), .ZN(n14534) );
  INV_X1 U15930 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14582) );
  NAND2_X1 U15931 ( .A1(n12835), .A2(n14582), .ZN(n12839) );
  NAND2_X1 U15932 ( .A1(n13357), .A2(n14582), .ZN(n12837) );
  NAND2_X1 U15933 ( .A1(n12780), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12836) );
  NAND3_X1 U15934 ( .A1(n12837), .A2(n12742), .A3(n12836), .ZN(n12838) );
  AND2_X1 U15935 ( .A1(n12839), .A2(n12838), .ZN(n14522) );
  MUX2_X1 U15936 ( .A(n12840), .B(n9674), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n12842) );
  NAND2_X1 U15937 ( .A1(n14485), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12841) );
  NAND2_X1 U15938 ( .A1(n12842), .A2(n12841), .ZN(n12843) );
  OR2_X1 U15939 ( .A1(n14524), .A2(n12843), .ZN(n12844) );
  NAND2_X1 U15940 ( .A1(n13676), .A2(n20969), .ZN(n15904) );
  OAI21_X1 U15941 ( .B1(n12846), .B2(n12845), .A(n15904), .ZN(n12847) );
  NAND2_X1 U15942 ( .A1(n20290), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n13310) );
  INV_X1 U15943 ( .A(n13310), .ZN(n12848) );
  AOI21_X1 U15944 ( .B1(n14440), .B2(n20292), .A(n12848), .ZN(n12892) );
  NAND2_X1 U15945 ( .A1(n12874), .A2(n15880), .ZN(n16165) );
  INV_X1 U15946 ( .A(n13959), .ZN(n12850) );
  NAND2_X1 U15947 ( .A1(n12850), .A2(n12849), .ZN(n12851) );
  AND2_X1 U15948 ( .A1(n12852), .A2(n12851), .ZN(n12863) );
  NAND2_X1 U15949 ( .A1(n12863), .A2(n12853), .ZN(n14470) );
  INV_X1 U15950 ( .A(n14470), .ZN(n12854) );
  INV_X1 U15951 ( .A(n20276), .ZN(n20261) );
  INV_X1 U15952 ( .A(n12855), .ZN(n13674) );
  INV_X1 U15953 ( .A(n12856), .ZN(n12857) );
  AOI21_X1 U15954 ( .B1(n12857), .B2(n13943), .A(n20316), .ZN(n12858) );
  NAND2_X1 U15955 ( .A1(n12859), .A2(n12858), .ZN(n13677) );
  OAI211_X1 U15956 ( .C1(n13674), .C2(n13918), .A(n13677), .B(n12860), .ZN(
        n12868) );
  OAI21_X1 U15957 ( .B1(n11563), .B2(n13331), .A(n14479), .ZN(n12861) );
  OAI21_X1 U15958 ( .B1(n12861), .B2(n11511), .A(n13943), .ZN(n12862) );
  OAI211_X1 U15959 ( .C1(n11771), .C2(n12864), .A(n12863), .B(n12862), .ZN(
        n12865) );
  INV_X1 U15960 ( .A(n12865), .ZN(n12866) );
  NAND2_X1 U15961 ( .A1(n12867), .A2(n12866), .ZN(n13680) );
  OR2_X1 U15962 ( .A1(n12868), .A2(n13680), .ZN(n12869) );
  NAND2_X1 U15963 ( .A1(n12874), .A2(n12869), .ZN(n16172) );
  NAND2_X1 U15964 ( .A1(n20261), .A2(n16172), .ZN(n13794) );
  INV_X1 U15965 ( .A(n13794), .ZN(n12870) );
  NAND2_X1 U15966 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16150) );
  NAND4_X1 U15967 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16173) );
  NOR2_X1 U15968 ( .A1(n16174), .A2(n16173), .ZN(n12884) );
  AND2_X1 U15969 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n12884), .ZN(
        n12873) );
  NAND2_X1 U15970 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16243) );
  INV_X1 U15971 ( .A(n16243), .ZN(n16264) );
  NAND4_X1 U15972 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A4(n16264), .ZN(n16220) );
  NOR2_X1 U15973 ( .A1(n16113), .A2(n16220), .ZN(n16228) );
  NAND2_X1 U15974 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16228), .ZN(
        n12883) );
  NAND2_X1 U15975 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20256) );
  INV_X1 U15976 ( .A(n20256), .ZN(n12871) );
  INV_X1 U15977 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n16168) );
  INV_X1 U15978 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20300) );
  OAI21_X1 U15979 ( .B1(n16168), .B2(n20300), .A(n20282), .ZN(n20273) );
  NAND2_X1 U15980 ( .A1(n12871), .A2(n20273), .ZN(n16282) );
  NOR2_X1 U15981 ( .A1(n12872), .A2(n16282), .ZN(n12882) );
  INV_X1 U15982 ( .A(n12882), .ZN(n16280) );
  NOR2_X1 U15983 ( .A1(n12883), .A2(n16280), .ZN(n16169) );
  NAND2_X1 U15984 ( .A1(n12873), .A2(n16169), .ZN(n16155) );
  NAND2_X1 U15985 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20259) );
  NOR2_X1 U15986 ( .A1(n20259), .A2(n20256), .ZN(n16257) );
  NAND2_X1 U15987 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n16257), .ZN(
        n16244) );
  NOR2_X1 U15988 ( .A1(n16244), .A2(n12883), .ZN(n16211) );
  NAND2_X1 U15989 ( .A1(n16165), .A2(n16172), .ZN(n20260) );
  INV_X1 U15990 ( .A(n20260), .ZN(n16258) );
  AOI21_X1 U15991 ( .B1(n16211), .B2(n12873), .A(n16258), .ZN(n12875) );
  OAI22_X1 U15992 ( .A1(n20290), .A2(n12874), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n16172), .ZN(n20258) );
  AOI211_X1 U15993 ( .C1(n20276), .C2(n16155), .A(n12875), .B(n20258), .ZN(
        n16156) );
  NOR2_X1 U15994 ( .A1(n15931), .A2(n16155), .ZN(n14889) );
  NOR2_X1 U15995 ( .A1(n16188), .A2(n20258), .ZN(n16259) );
  AOI21_X1 U15996 ( .B1(n16156), .B2(n14889), .A(n16259), .ZN(n16145) );
  AOI21_X1 U15997 ( .B1(n16188), .B2(n16150), .A(n16145), .ZN(n16144) );
  INV_X1 U15998 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16143) );
  NAND2_X1 U15999 ( .A1(n20276), .A2(n16143), .ZN(n12876) );
  AND2_X1 U16000 ( .A1(n16144), .A2(n12876), .ZN(n14881) );
  NOR2_X1 U16001 ( .A1(n14882), .A2(n16143), .ZN(n14871) );
  INV_X1 U16002 ( .A(n16165), .ZN(n13795) );
  NAND2_X1 U16003 ( .A1(n13795), .A2(n14735), .ZN(n12878) );
  NAND2_X1 U16004 ( .A1(n20276), .A2(n14882), .ZN(n12877) );
  OAI211_X1 U16005 ( .C1(n14871), .C2(n16172), .A(n12878), .B(n12877), .ZN(
        n12879) );
  INV_X1 U16006 ( .A(n12879), .ZN(n12880) );
  NAND2_X1 U16007 ( .A1(n14869), .A2(n20293), .ZN(n14860) );
  AND2_X1 U16008 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12881) );
  NAND2_X1 U16009 ( .A1(n14869), .A2(n12881), .ZN(n14859) );
  NAND3_X1 U16010 ( .A1(n14860), .A2(n14859), .A3(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12890) );
  NAND2_X1 U16011 ( .A1(n16165), .A2(n16168), .ZN(n20294) );
  AND4_X1 U16012 ( .A1(n12884), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n11763), .A4(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12885) );
  INV_X1 U16013 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14864) );
  NOR2_X1 U16014 ( .A1(n14735), .A2(n14864), .ZN(n12886) );
  NOR2_X1 U16015 ( .A1(n12887), .A2(n14846), .ZN(n12888) );
  NAND2_X1 U16016 ( .A1(n14858), .A2(n12888), .ZN(n12889) );
  INV_X1 U16017 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17184) );
  NAND3_X1 U16018 ( .A1(n19025), .A2(n19014), .A3(n10055), .ZN(n12912) );
  INV_X1 U16019 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12895) );
  INV_X2 U16020 ( .A(n12990), .ZN(n12928) );
  AOI22_X1 U16021 ( .A1(n12945), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17352), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12894) );
  OAI21_X1 U16022 ( .B1(n12918), .B2(n17184), .A(n12894), .ZN(n12911) );
  INV_X1 U16023 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17179) );
  AOI22_X1 U16024 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17320), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12909) );
  INV_X1 U16025 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17106) );
  INV_X1 U16026 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17107) );
  OAI22_X1 U16027 ( .A1(n17367), .A2(n17106), .B1(n17249), .B2(n17107), .ZN(
        n12907) );
  NOR2_X2 U16028 ( .A1(n12899), .A2(n17060), .ZN(n13080) );
  AOI22_X1 U16029 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12905) );
  AOI22_X1 U16030 ( .A1(n17384), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12904) );
  NAND2_X4 U16031 ( .A1(n18850), .A2(n12902), .ZN(n17380) );
  AOI22_X1 U16032 ( .A1(n17321), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17392), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12903) );
  NAND3_X1 U16033 ( .A1(n12905), .A2(n12904), .A3(n12903), .ZN(n12906) );
  AOI211_X1 U16034 ( .C1(n17336), .C2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n12907), .B(n12906), .ZN(n12908) );
  OAI211_X1 U16035 ( .C1(n17268), .C2(n17179), .A(n12909), .B(n12908), .ZN(
        n12910) );
  INV_X2 U16036 ( .A(n17249), .ZN(n13039) );
  INV_X1 U16037 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17205) );
  AOI22_X1 U16038 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17320), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12913) );
  OAI21_X1 U16039 ( .B1(n15784), .B2(n17205), .A(n12913), .ZN(n12917) );
  INV_X1 U16040 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17313) );
  AOI22_X1 U16041 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12915) );
  INV_X2 U16042 ( .A(n17396), .ZN(n17217) );
  AOI22_X1 U16043 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17352), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12914) );
  OAI211_X1 U16044 ( .C1(n17358), .C2(n17313), .A(n12915), .B(n12914), .ZN(
        n12916) );
  AOI211_X1 U16045 ( .C1(n17374), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n12917), .B(n12916), .ZN(n12925) );
  AOI22_X1 U16046 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12919) );
  OAI21_X1 U16047 ( .B1(n12918), .B2(n17302), .A(n12919), .ZN(n12923) );
  AOI22_X1 U16048 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17321), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12921) );
  INV_X1 U16049 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17305) );
  NAND3_X1 U16050 ( .A1(n12921), .A2(n10222), .A3(n12920), .ZN(n12922) );
  INV_X1 U16051 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17319) );
  INV_X2 U16052 ( .A(n15833), .ZN(n17356) );
  AOI22_X1 U16053 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17356), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12936) );
  INV_X1 U16054 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17218) );
  INV_X2 U16055 ( .A(n12918), .ZN(n17339) );
  AOI22_X1 U16056 ( .A1(n12945), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12927) );
  INV_X1 U16057 ( .A(n17303), .ZN(n17375) );
  AOI22_X1 U16058 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12926) );
  OAI211_X1 U16059 ( .C1(n17249), .C2(n17218), .A(n12927), .B(n12926), .ZN(
        n12934) );
  INV_X2 U16060 ( .A(n12928), .ZN(n17381) );
  AOI22_X1 U16061 ( .A1(n17381), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12932) );
  AOI22_X1 U16062 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17336), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12931) );
  INV_X2 U16063 ( .A(n17120), .ZN(n17384) );
  AOI22_X1 U16064 ( .A1(n17384), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17320), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12930) );
  NAND2_X1 U16065 ( .A1(n17392), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12929) );
  NAND4_X1 U16066 ( .A1(n12932), .A2(n12931), .A3(n12930), .A4(n12929), .ZN(
        n12933) );
  AOI211_X1 U16067 ( .C1(n17321), .C2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n12934), .B(n12933), .ZN(n12935) );
  INV_X1 U16068 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17424) );
  AOI22_X1 U16069 ( .A1(n17352), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12937) );
  OAI21_X1 U16070 ( .B1(n17268), .B2(n17424), .A(n12937), .ZN(n12943) );
  AOI22_X1 U16071 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17320), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12941) );
  INV_X1 U16072 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17348) );
  AOI22_X1 U16073 ( .A1(n17321), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17392), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12944) );
  INV_X1 U16074 ( .A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15754) );
  OAI22_X1 U16075 ( .A1(n17249), .A2(n15754), .B1(n12918), .B2(n17232), .ZN(
        n12950) );
  AOI22_X1 U16076 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17356), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12948) );
  AOI22_X1 U16077 ( .A1(n9665), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12945), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12947) );
  NAND3_X1 U16078 ( .A1(n12948), .A2(n12947), .A3(n12946), .ZN(n12949) );
  NOR3_X1 U16079 ( .A1(n12951), .A2(n12950), .A3(n12949), .ZN(n12952) );
  AOI22_X1 U16080 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17320), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12956) );
  INV_X1 U16081 ( .A(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17359) );
  INV_X1 U16082 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17366) );
  AOI22_X1 U16083 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n13117), .ZN(n12958) );
  AOI22_X1 U16084 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n12990), .B1(
        n9665), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12957) );
  OAI211_X1 U16085 ( .C1(n17380), .C2(n17366), .A(n12958), .B(n12957), .ZN(
        n12959) );
  AOI22_X1 U16086 ( .A1(n12938), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n14415), .ZN(n12964) );
  AOI22_X1 U16087 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n17382), .B1(
        n12945), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12963) );
  AOI22_X1 U16088 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17356), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12962) );
  NAND2_X1 U16089 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n13039), .ZN(
        n12961) );
  NAND2_X2 U16090 ( .A1(n12965), .A2(n10235), .ZN(n17585) );
  AOI22_X1 U16091 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17320), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12976) );
  INV_X1 U16092 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15807) );
  AOI22_X1 U16093 ( .A1(n17384), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17381), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12967) );
  AOI22_X1 U16094 ( .A1(n13117), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12966) );
  OAI211_X1 U16095 ( .C1(n17249), .C2(n15807), .A(n12967), .B(n12966), .ZN(
        n12974) );
  AOI22_X1 U16096 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12972) );
  AOI22_X1 U16097 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12971) );
  AOI22_X1 U16098 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12945), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12970) );
  NAND2_X1 U16099 ( .A1(n17392), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12969) );
  NAND4_X1 U16100 ( .A1(n12972), .A2(n12971), .A3(n12970), .A4(n12969), .ZN(
        n12973) );
  AOI211_X1 U16101 ( .C1(n17321), .C2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n12974), .B(n12973), .ZN(n12975) );
  OAI211_X1 U16102 ( .C1(n14414), .C2(n15825), .A(n12976), .B(n12975), .ZN(
        n17566) );
  INV_X1 U16103 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17406) );
  AOI22_X1 U16104 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17321), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12986) );
  INV_X1 U16105 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17119) );
  AOI22_X1 U16106 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17381), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12978) );
  AOI22_X1 U16107 ( .A1(n17384), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17306), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12977) );
  OAI211_X1 U16108 ( .C1(n17358), .C2(n17119), .A(n12978), .B(n12977), .ZN(
        n12984) );
  AOI22_X1 U16109 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12982) );
  AOI22_X1 U16110 ( .A1(n12945), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12981) );
  AOI22_X1 U16111 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17336), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12980) );
  NAND2_X1 U16112 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12979) );
  NAND4_X1 U16113 ( .A1(n12982), .A2(n12981), .A3(n12980), .A4(n12979), .ZN(
        n12983) );
  AOI211_X1 U16114 ( .C1(n17374), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n12984), .B(n12983), .ZN(n12985) );
  XOR2_X1 U16115 ( .A(n17563), .B(n12987), .Z(n13016) );
  INV_X1 U16116 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19020) );
  NOR2_X1 U16117 ( .A1(n17585), .A2(n19020), .ZN(n13000) );
  INV_X1 U16118 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15762) );
  AOI22_X1 U16119 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12989) );
  AOI22_X1 U16120 ( .A1(n17382), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12988) );
  OAI211_X1 U16121 ( .C1(n17358), .C2(n15762), .A(n12989), .B(n12988), .ZN(
        n12999) );
  AOI22_X1 U16122 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12938), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12994) );
  AOI22_X1 U16123 ( .A1(n12945), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12990), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12993) );
  AOI22_X1 U16124 ( .A1(n17384), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12968), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12992) );
  NAND2_X1 U16125 ( .A1(n17321), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12991) );
  NAND4_X1 U16126 ( .A1(n12994), .A2(n12993), .A3(n12992), .A4(n12991), .ZN(
        n12998) );
  AOI22_X1 U16127 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12996) );
  INV_X1 U16128 ( .A(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17395) );
  NAND3_X1 U16129 ( .A1(n12996), .A2(n12995), .A3(n10223), .ZN(n12997) );
  NOR2_X1 U16130 ( .A1(n18072), .A2(n18079), .ZN(n18071) );
  NOR2_X1 U16131 ( .A1(n13000), .A2(n18071), .ZN(n18062) );
  NOR2_X1 U16132 ( .A1(n18062), .A2(n18063), .ZN(n13004) );
  NOR2_X1 U16133 ( .A1(n13001), .A2(n13002), .ZN(n13003) );
  XNOR2_X1 U16134 ( .A(n13155), .B(n13005), .ZN(n13006) );
  NOR2_X1 U16135 ( .A1(n13007), .A2(n13006), .ZN(n13008) );
  XNOR2_X1 U16136 ( .A(n13007), .B(n13006), .ZN(n18049) );
  INV_X1 U16137 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18050) );
  NOR2_X1 U16138 ( .A1(n18049), .A2(n18050), .ZN(n18048) );
  INV_X1 U16139 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18338) );
  XOR2_X1 U16140 ( .A(n18338), .B(n13011), .Z(n18034) );
  XNOR2_X1 U16141 ( .A(n17566), .B(n13012), .ZN(n13013) );
  NOR2_X1 U16142 ( .A1(n13014), .A2(n13013), .ZN(n13015) );
  INV_X1 U16143 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18344) );
  NOR2_X1 U16144 ( .A1(n18344), .A2(n18026), .ZN(n18025) );
  NOR2_X2 U16145 ( .A1(n13015), .A2(n18025), .ZN(n18017) );
  INV_X1 U16146 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18336) );
  XOR2_X1 U16147 ( .A(n18336), .B(n13016), .Z(n18016) );
  INV_X1 U16148 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18324) );
  NOR2_X1 U16149 ( .A1(n13019), .A2(n13018), .ZN(n13020) );
  NOR2_X2 U16150 ( .A1(n18006), .A2(n13020), .ZN(n13022) );
  INV_X1 U16151 ( .A(n13022), .ZN(n13021) );
  INV_X1 U16152 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18312) );
  NAND2_X2 U16153 ( .A1(n13021), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18272) );
  NAND2_X1 U16154 ( .A1(n13022), .A2(n18312), .ZN(n17959) );
  INV_X1 U16155 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17981) );
  INV_X1 U16156 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18286) );
  NOR2_X1 U16157 ( .A1(n17981), .A2(n18286), .ZN(n17963) );
  NAND2_X1 U16158 ( .A1(n17963), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18262) );
  INV_X1 U16159 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18261) );
  NOR2_X1 U16160 ( .A1(n18262), .A2(n18261), .ZN(n18231) );
  INV_X1 U16161 ( .A(n18231), .ZN(n18258) );
  NAND2_X1 U16162 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17910) );
  NOR2_X1 U16163 ( .A1(n18258), .A2(n17910), .ZN(n18208) );
  NAND2_X1 U16164 ( .A1(n18208), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13221) );
  OR2_X2 U16165 ( .A1(n17931), .A2(n13221), .ZN(n13026) );
  NAND2_X1 U16166 ( .A1(n13026), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13024) );
  INV_X1 U16167 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18213) );
  NAND2_X1 U16168 ( .A1(n13024), .A2(n13023), .ZN(n13025) );
  INV_X1 U16169 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17933) );
  NOR2_X1 U16170 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18222) );
  AOI21_X1 U16171 ( .B1(n17907), .B2(n18222), .A(n10059), .ZN(n17873) );
  INV_X1 U16172 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18200) );
  NAND2_X1 U16173 ( .A1(n17869), .A2(n18200), .ZN(n17868) );
  NAND2_X2 U16174 ( .A1(n17868), .A2(n17819), .ZN(n17781) );
  NOR2_X1 U16175 ( .A1(n18213), .A2(n18200), .ZN(n18193) );
  NAND2_X1 U16176 ( .A1(n18193), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18162) );
  INV_X1 U16177 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18183) );
  INV_X1 U16178 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18150) );
  NOR2_X1 U16179 ( .A1(n18183), .A2(n18150), .ZN(n18164) );
  NAND2_X1 U16180 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18164), .ZN(
        n18144) );
  NOR2_X1 U16181 ( .A1(n18162), .A2(n18144), .ZN(n18148) );
  NAND2_X1 U16182 ( .A1(n18148), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18152) );
  INV_X1 U16183 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18129) );
  NOR2_X1 U16184 ( .A1(n18152), .A2(n18129), .ZN(n17774) );
  NAND2_X1 U16185 ( .A1(n17858), .A2(n18183), .ZN(n13027) );
  INV_X1 U16186 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17823) );
  NAND2_X1 U16187 ( .A1(n17821), .A2(n17823), .ZN(n17797) );
  NAND2_X1 U16188 ( .A1(n18193), .A2(n17798), .ZN(n17818) );
  INV_X1 U16189 ( .A(n18144), .ZN(n18155) );
  AND2_X1 U16190 ( .A1(n18155), .A2(n10239), .ZN(n13030) );
  INV_X1 U16191 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18115) );
  NAND2_X1 U16192 ( .A1(n17819), .A2(n10068), .ZN(n13031) );
  OAI211_X1 U16193 ( .C1(n13032), .C2(n18115), .A(n13031), .B(n10212), .ZN(
        n17746) );
  NAND2_X1 U16194 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18087) );
  INV_X1 U16195 ( .A(n18087), .ZN(n13033) );
  NOR2_X1 U16196 ( .A1(n17819), .A2(n13033), .ZN(n13034) );
  NOR2_X2 U16197 ( .A1(n17745), .A2(n13035), .ZN(n13036) );
  AOI21_X1 U16198 ( .B1(n10059), .B2(n17735), .A(n17733), .ZN(n17709) );
  INV_X1 U16199 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15858) );
  OAI22_X1 U16200 ( .A1(n15858), .A2(n17819), .B1(n10059), .B2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17708) );
  NOR2_X1 U16201 ( .A1(n17709), .A2(n17708), .ZN(n17710) );
  INV_X1 U16202 ( .A(n17735), .ZN(n13227) );
  INV_X1 U16203 ( .A(n16559), .ZN(n17559) );
  NAND2_X1 U16204 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18112) );
  INV_X1 U16205 ( .A(n18112), .ZN(n18108) );
  NAND3_X1 U16206 ( .A1(n18108), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13292) );
  NOR2_X1 U16207 ( .A1(n18152), .A2(n13292), .ZN(n13231) );
  INV_X1 U16208 ( .A(n13231), .ZN(n16568) );
  NAND3_X1 U16209 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(n18090), .ZN(n16584) );
  INV_X1 U16210 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17418) );
  AOI22_X1 U16211 ( .A1(n17384), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13038) );
  OAI21_X1 U16212 ( .B1(n15784), .B2(n17418), .A(n13038), .ZN(n13044) );
  AOI22_X1 U16213 ( .A1(n17381), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13042) );
  AOI22_X1 U16214 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13041) );
  AOI22_X1 U16215 ( .A1(n13039), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17392), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13040) );
  NAND3_X1 U16216 ( .A1(n13042), .A2(n13041), .A3(n13040), .ZN(n13043) );
  AOI211_X1 U16217 ( .C1(n13080), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n13044), .B(n13043), .ZN(n13049) );
  INV_X1 U16218 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15747) );
  OAI22_X1 U16219 ( .A1(n17367), .A2(n17302), .B1(n17268), .B2(n15747), .ZN(
        n13048) );
  AOI22_X1 U16220 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17320), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13046) );
  NAND3_X1 U16221 ( .A1(n13046), .A2(n10224), .A3(n13045), .ZN(n13047) );
  INV_X1 U16222 ( .A(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17172) );
  AOI22_X1 U16223 ( .A1(n17382), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13059) );
  INV_X1 U16224 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17175) );
  AOI22_X1 U16225 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17356), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13051) );
  AOI22_X1 U16226 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17352), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13050) );
  OAI211_X1 U16227 ( .C1(n17249), .C2(n17175), .A(n13051), .B(n13050), .ZN(
        n13057) );
  AOI22_X1 U16228 ( .A1(n12945), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13055) );
  AOI22_X1 U16229 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13054) );
  AOI22_X1 U16230 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13053) );
  NAND2_X1 U16231 ( .A1(n17392), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n13052) );
  NAND4_X1 U16232 ( .A1(n13055), .A2(n13054), .A3(n13053), .A4(n13052), .ZN(
        n13056) );
  AOI22_X1 U16233 ( .A1(n17356), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13061) );
  AOI22_X1 U16234 ( .A1(n12945), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17352), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13060) );
  OAI211_X1 U16235 ( .C1(n17358), .C2(n15825), .A(n13061), .B(n13060), .ZN(
        n13067) );
  AOI22_X1 U16236 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13065) );
  AOI22_X1 U16237 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13080), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13064) );
  AOI22_X1 U16238 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17321), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13063) );
  NAND2_X1 U16239 ( .A1(n14415), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n13062) );
  NAND4_X1 U16240 ( .A1(n13065), .A2(n13064), .A3(n13063), .A4(n13062), .ZN(
        n13066) );
  INV_X2 U16241 ( .A(n18439), .ZN(n17446) );
  AOI22_X1 U16242 ( .A1(n17381), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13079) );
  AOI22_X1 U16243 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13080), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13071) );
  AOI22_X1 U16244 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13070) );
  OAI211_X1 U16245 ( .C1(n17358), .C2(n17348), .A(n13071), .B(n13070), .ZN(
        n13077) );
  AOI22_X1 U16246 ( .A1(n12945), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13075) );
  AOI22_X1 U16247 ( .A1(n9665), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13074) );
  AOI22_X1 U16248 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17320), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13073) );
  NAND2_X1 U16249 ( .A1(n17374), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n13072) );
  NAND4_X1 U16250 ( .A1(n13075), .A2(n13074), .A3(n13073), .A4(n13072), .ZN(
        n13076) );
  AOI22_X1 U16251 ( .A1(n17382), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13091) );
  INV_X1 U16252 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13090) );
  INV_X1 U16253 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17284) );
  AOI22_X1 U16254 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13080), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13082) );
  AOI22_X1 U16255 ( .A1(n12945), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17352), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13081) );
  OAI211_X1 U16256 ( .C1(n17358), .C2(n17284), .A(n13082), .B(n13081), .ZN(
        n13083) );
  INV_X1 U16257 ( .A(n13083), .ZN(n13089) );
  AOI22_X1 U16258 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17306), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13087) );
  AOI22_X1 U16259 ( .A1(n9665), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13086) );
  AOI22_X1 U16260 ( .A1(n17356), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17320), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13085) );
  NAND2_X1 U16261 ( .A1(n17374), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n13084) );
  NAND4_X1 U16262 ( .A1(n13087), .A2(n13086), .A3(n13085), .A4(n13084), .ZN(
        n13088) );
  INV_X1 U16263 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17420) );
  AOI22_X1 U16264 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17320), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13101) );
  INV_X1 U16265 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17330) );
  AOI22_X1 U16266 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13080), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13093) );
  AOI22_X1 U16267 ( .A1(n17382), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13092) );
  OAI211_X1 U16268 ( .C1(n17358), .C2(n17330), .A(n13093), .B(n13092), .ZN(
        n13099) );
  AOI22_X1 U16269 ( .A1(n9665), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13097) );
  AOI22_X1 U16270 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17352), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13096) );
  AOI22_X1 U16271 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13095) );
  NAND2_X1 U16272 ( .A1(n17321), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n13094) );
  NAND4_X1 U16273 ( .A1(n13097), .A2(n13096), .A3(n13095), .A4(n13094), .ZN(
        n13098) );
  NAND2_X1 U16274 ( .A1(n18449), .A2(n18429), .ZN(n13150) );
  INV_X1 U16275 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17379) );
  AOI22_X1 U16276 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13109) );
  INV_X1 U16277 ( .A(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13103) );
  AOI22_X1 U16278 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13039), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13102) );
  OAI21_X1 U16279 ( .B1(n15833), .B2(n13103), .A(n13102), .ZN(n13107) );
  INV_X1 U16280 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15770) );
  AOI22_X1 U16281 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13105) );
  AOI22_X1 U16282 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13104) );
  OAI211_X1 U16283 ( .C1(n17358), .C2(n15770), .A(n13105), .B(n13104), .ZN(
        n13106) );
  AOI211_X1 U16284 ( .C1(n17321), .C2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n13107), .B(n13106), .ZN(n13108) );
  OAI211_X1 U16285 ( .C1(n15784), .C2(n17379), .A(n13109), .B(n13108), .ZN(
        n13110) );
  INV_X1 U16286 ( .A(n13110), .ZN(n13115) );
  AOI22_X1 U16287 ( .A1(n9665), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17352), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13111) );
  OAI21_X1 U16288 ( .B1(n17355), .B2(n17267), .A(n13111), .ZN(n13113) );
  INV_X1 U16289 ( .A(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17248) );
  AOI22_X1 U16290 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13116) );
  OAI21_X1 U16291 ( .B1(n14414), .B2(n17248), .A(n13116), .ZN(n13128) );
  AOI22_X1 U16292 ( .A1(n17382), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17352), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13120) );
  AOI22_X1 U16293 ( .A1(n13117), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13119) );
  AOI22_X1 U16294 ( .A1(n17374), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17392), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13118) );
  NAND3_X1 U16295 ( .A1(n13120), .A2(n13119), .A3(n13118), .ZN(n13126) );
  AOI22_X1 U16296 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17306), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13124) );
  INV_X1 U16297 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17247) );
  OAI22_X1 U16298 ( .A1(n17380), .A2(n17247), .B1(n15833), .B2(n17354), .ZN(
        n13121) );
  NAND3_X1 U16299 ( .A1(n13124), .A2(n13123), .A3(n13122), .ZN(n13125) );
  AOI211_X4 U16300 ( .C1(n9662), .C2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n13128), .B(n13127), .ZN(n17658) );
  NAND2_X1 U16301 ( .A1(n18444), .A2(n17446), .ZN(n14409) );
  NAND3_X1 U16302 ( .A1(n13134), .A2(n13136), .A3(n14409), .ZN(n13129) );
  INV_X1 U16303 ( .A(n16551), .ZN(n13130) );
  NOR2_X1 U16304 ( .A1(n17658), .A2(n18424), .ZN(n13216) );
  NAND2_X1 U16305 ( .A1(n13216), .A2(n18444), .ZN(n13209) );
  OAI21_X1 U16306 ( .B1(n16584), .B2(n16559), .A(n18839), .ZN(n13131) );
  INV_X1 U16307 ( .A(n13131), .ZN(n13132) );
  NAND2_X1 U16308 ( .A1(n17658), .A2(n18411), .ZN(n13137) );
  NAND2_X1 U16309 ( .A1(n13136), .A2(n13137), .ZN(n19068) );
  NAND2_X1 U16310 ( .A1(n13199), .A2(n17436), .ZN(n13138) );
  NOR2_X1 U16311 ( .A1(n17446), .A2(n18434), .ZN(n13141) );
  NAND4_X1 U16312 ( .A1(n13149), .A2(n13139), .A3(n13141), .A4(n18444), .ZN(
        n13153) );
  NOR2_X1 U16313 ( .A1(n13140), .A2(n13153), .ZN(n13213) );
  NOR2_X1 U16314 ( .A1(n16695), .A2(n13136), .ZN(n16713) );
  NAND2_X1 U16315 ( .A1(n13140), .A2(n18439), .ZN(n13218) );
  AOI21_X1 U16316 ( .B1(n18449), .B2(n15943), .A(n13137), .ZN(n13210) );
  AOI21_X1 U16317 ( .B1(n13138), .B2(n13218), .A(n13210), .ZN(n13148) );
  INV_X1 U16318 ( .A(n13139), .ZN(n13147) );
  AND4_X1 U16319 ( .A1(n13151), .A2(n14409), .A3(n13140), .A4(n14411), .ZN(
        n13146) );
  NOR2_X1 U16320 ( .A1(n17446), .A2(n17436), .ZN(n13198) );
  NOR3_X1 U16321 ( .A1(n13142), .A2(n13141), .A3(n18424), .ZN(n13144) );
  OAI21_X1 U16322 ( .B1(n13198), .B2(n17527), .A(n18434), .ZN(n13143) );
  OAI21_X1 U16323 ( .B1(n13198), .B2(n13144), .A(n13143), .ZN(n13145) );
  AOI211_X1 U16324 ( .C1(n13149), .C2(n13147), .A(n13146), .B(n13145), .ZN(
        n13212) );
  NAND2_X1 U16325 ( .A1(n17578), .A2(n13157), .ZN(n13156) );
  NAND2_X1 U16326 ( .A1(n13156), .A2(n13155), .ZN(n13167) );
  NAND2_X1 U16327 ( .A1(n13169), .A2(n17566), .ZN(n13173) );
  NOR2_X1 U16328 ( .A1(n17563), .A2(n13173), .ZN(n13177) );
  NAND2_X1 U16329 ( .A1(n13177), .A2(n16559), .ZN(n13178) );
  INV_X1 U16330 ( .A(n13155), .ZN(n17574) );
  XOR2_X1 U16331 ( .A(n13156), .B(n17574), .Z(n13164) );
  NOR2_X1 U16332 ( .A1(n18050), .A2(n13164), .ZN(n13165) );
  XOR2_X1 U16333 ( .A(n17578), .B(n13157), .Z(n13158) );
  NOR2_X1 U16334 ( .A1(n13158), .A2(n13001), .ZN(n13163) );
  XOR2_X1 U16335 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n13158), .Z(
        n18061) );
  INV_X1 U16336 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19035) );
  NOR2_X1 U16337 ( .A1(n13160), .A2(n19035), .ZN(n13162) );
  NAND3_X1 U16338 ( .A1(n13161), .A2(n13160), .A3(n19035), .ZN(n13159) );
  OAI221_X1 U16339 ( .B1(n13162), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n13161), .C2(n13160), .A(n13159), .ZN(n18060) );
  NOR2_X1 U16340 ( .A1(n18061), .A2(n18060), .ZN(n18059) );
  NOR2_X1 U16341 ( .A1(n13166), .A2(n18338), .ZN(n13168) );
  XNOR2_X1 U16342 ( .A(n13167), .B(n17571), .ZN(n18037) );
  XNOR2_X1 U16343 ( .A(n13169), .B(n17566), .ZN(n13171) );
  NOR2_X1 U16344 ( .A1(n13170), .A2(n13171), .ZN(n13172) );
  XNOR2_X1 U16345 ( .A(n13173), .B(n17563), .ZN(n13175) );
  NOR2_X1 U16346 ( .A1(n13174), .A2(n13175), .ZN(n13176) );
  XNOR2_X1 U16347 ( .A(n13175), .B(n13174), .ZN(n18012) );
  XNOR2_X1 U16348 ( .A(n13177), .B(n16559), .ZN(n13180) );
  INV_X1 U16349 ( .A(n13178), .ZN(n13183) );
  OR2_X1 U16350 ( .A1(n13180), .A2(n13179), .ZN(n18001) );
  OAI21_X1 U16351 ( .B1(n13183), .B2(n13182), .A(n18001), .ZN(n13181) );
  INV_X1 U16352 ( .A(n13221), .ZN(n18187) );
  INV_X1 U16353 ( .A(n17726), .ZN(n18092) );
  NAND2_X1 U16354 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13185) );
  INV_X1 U16355 ( .A(n13298), .ZN(n16587) );
  NAND2_X1 U16356 ( .A1(n19018), .A2(n19008), .ZN(n19009) );
  NOR2_X1 U16357 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19009), .ZN(n19070) );
  OAI22_X1 U16358 ( .A1(n19031), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n18864), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13202) );
  NAND2_X1 U16359 ( .A1(n18414), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13201) );
  NOR2_X1 U16360 ( .A1(n13202), .A2(n13201), .ZN(n13186) );
  AOI21_X1 U16361 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18864), .A(
        n13186), .ZN(n13192) );
  AOI22_X1 U16362 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n18884), .B2(n19025), .ZN(
        n13191) );
  NOR2_X1 U16363 ( .A1(n13192), .A2(n13191), .ZN(n13187) );
  AOI21_X1 U16364 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n18884), .A(
        n13187), .ZN(n13188) );
  AOI22_X1 U16365 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18849), .B1(
        n13188), .B2(n19014), .ZN(n13193) );
  NOR2_X1 U16366 ( .A1(n13188), .A2(n19014), .ZN(n13194) );
  NAND2_X1 U16367 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18849), .ZN(
        n13189) );
  OAI22_X1 U16368 ( .A1(n13193), .A2(n18887), .B1(n13194), .B2(n13189), .ZN(
        n13190) );
  INV_X1 U16369 ( .A(n13190), .ZN(n13197) );
  OAI211_X1 U16370 ( .C1(n18414), .C2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n13201), .B(n13197), .ZN(n13208) );
  XNOR2_X1 U16371 ( .A(n13192), .B(n13191), .ZN(n13207) );
  INV_X1 U16372 ( .A(n13207), .ZN(n13196) );
  OAI21_X1 U16373 ( .B1(n18887), .B2(n13194), .A(n13193), .ZN(n13195) );
  AOI21_X1 U16374 ( .B1(n13197), .B2(n13196), .A(n13205), .ZN(n13203) );
  OAI21_X1 U16375 ( .B1(n13202), .B2(n13208), .A(n13203), .ZN(n14407) );
  INV_X1 U16376 ( .A(n14407), .ZN(n18845) );
  INV_X1 U16377 ( .A(n13198), .ZN(n13200) );
  OAI21_X1 U16378 ( .B1(n18424), .B2(n13200), .A(n13199), .ZN(n13214) );
  XOR2_X1 U16379 ( .A(n13202), .B(n13201), .Z(n13206) );
  INV_X1 U16380 ( .A(n13203), .ZN(n13204) );
  OAI21_X1 U16381 ( .B1(n13208), .B2(n13207), .A(n16690), .ZN(n18838) );
  INV_X1 U16382 ( .A(n13210), .ZN(n13211) );
  OAI211_X1 U16383 ( .C1(n13213), .C2(n16551), .A(n13212), .B(n13211), .ZN(
        n15847) );
  NAND2_X1 U16384 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n19050) );
  INV_X1 U16385 ( .A(n19050), .ZN(n19057) );
  NAND2_X1 U16386 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18931), .ZN(n19066) );
  INV_X2 U16387 ( .A(n19066), .ZN(n19000) );
  NAND2_X1 U16388 ( .A1(n19000), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18996) );
  NOR2_X1 U16389 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18919) );
  INV_X1 U16390 ( .A(n18919), .ZN(n13215) );
  NAND3_X1 U16391 ( .A1(n18931), .A2(n18990), .A3(n13215), .ZN(n18924) );
  INV_X1 U16392 ( .A(n18924), .ZN(n19055) );
  AOI211_X1 U16393 ( .C1(n17658), .C2(n18424), .A(n13216), .B(n19055), .ZN(
        n13217) );
  NOR2_X1 U16394 ( .A1(n19057), .A2(n13217), .ZN(n16694) );
  NAND3_X1 U16395 ( .A1(n16694), .A2(n13218), .A3(n16690), .ZN(n13219) );
  NAND2_X1 U16396 ( .A1(n19018), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18909) );
  NAND2_X1 U16397 ( .A1(n18380), .A2(n18386), .ZN(n18378) );
  INV_X1 U16398 ( .A(n18859), .ZN(n18851) );
  NOR2_X1 U16399 ( .A1(n18880), .A2(n18851), .ZN(n18287) );
  INV_X1 U16400 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17727) );
  INV_X1 U16401 ( .A(n18857), .ZN(n18871) );
  NAND2_X1 U16402 ( .A1(n18871), .A2(n18859), .ZN(n18306) );
  NAND2_X1 U16403 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18185) );
  INV_X1 U16404 ( .A(n18185), .ZN(n18346) );
  NOR3_X1 U16405 ( .A1(n18050), .A2(n18338), .A3(n18344), .ZN(n18186) );
  NAND2_X1 U16406 ( .A1(n18346), .A2(n18186), .ZN(n18305) );
  NAND3_X1 U16407 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18243) );
  NOR2_X1 U16408 ( .A1(n18305), .A2(n18243), .ZN(n18151) );
  INV_X1 U16409 ( .A(n18151), .ZN(n18274) );
  NOR2_X1 U16410 ( .A1(n13221), .A2(n18274), .ZN(n18086) );
  AOI21_X1 U16411 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18348) );
  INV_X1 U16412 ( .A(n18348), .ZN(n18365) );
  NAND2_X1 U16413 ( .A1(n18186), .A2(n18365), .ZN(n18307) );
  NOR2_X1 U16414 ( .A1(n18243), .A2(n18307), .ZN(n18205) );
  NAND2_X1 U16415 ( .A1(n18187), .A2(n18205), .ZN(n18190) );
  OAI21_X1 U16416 ( .B1(n16568), .B2(n18190), .A(n18880), .ZN(n18089) );
  OAI221_X1 U16417 ( .B1(n18367), .B2(n13231), .C1(n18367), .C2(n18086), .A(
        n18089), .ZN(n13222) );
  AOI221_X1 U16418 ( .B1(n19035), .B2(n18857), .C1(n17727), .C2(n18857), .A(
        n13222), .ZN(n13293) );
  OAI21_X1 U16419 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18287), .A(
        n13293), .ZN(n15857) );
  AOI211_X1 U16420 ( .C1(n18252), .C2(n16587), .A(n18388), .B(n15857), .ZN(
        n13223) );
  INV_X2 U16421 ( .A(n18380), .ZN(n18393) );
  NOR2_X1 U16422 ( .A1(n18393), .A2(n15858), .ZN(n13225) );
  AND3_X1 U16423 ( .A1(n15858), .A2(n13228), .A3(n13227), .ZN(n13230) );
  AND2_X1 U16424 ( .A1(n17708), .A2(n17733), .ZN(n13229) );
  NAND2_X1 U16425 ( .A1(n18394), .A2(n18839), .ZN(n18401) );
  AOI21_X1 U16426 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18857), .A(
        n18851), .ZN(n18366) );
  INV_X1 U16427 ( .A(n18086), .ZN(n18147) );
  OAI22_X1 U16428 ( .A1(n18844), .A2(n18190), .B1(n18366), .B2(n18147), .ZN(
        n13290) );
  NAND2_X1 U16429 ( .A1(n17559), .A2(n18839), .ZN(n18248) );
  OAI22_X1 U16430 ( .A1(n18843), .A2(n18227), .B1(n18218), .B2(n18248), .ZN(
        n18188) );
  NOR2_X1 U16431 ( .A1(n13290), .A2(n18188), .ZN(n18136) );
  NAND2_X1 U16432 ( .A1(n13231), .A2(n18142), .ZN(n18093) );
  NAND2_X1 U16433 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n15858), .ZN(
        n17732) );
  NAND2_X1 U16434 ( .A1(n18393), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17716) );
  INV_X1 U16435 ( .A(n13236), .ZN(n13237) );
  NOR2_X1 U16436 ( .A1(n13238), .A2(n13237), .ZN(n13258) );
  INV_X1 U16437 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13242) );
  AOI22_X1 U16438 ( .A1(n9685), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12587), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13241) );
  AOI21_X1 U16439 ( .B1(n9652), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A(n13239), .ZN(n13240) );
  OAI211_X1 U16440 ( .C1(n9654), .C2(n13242), .A(n13241), .B(n13240), .ZN(
        n13256) );
  AOI22_X1 U16441 ( .A1(n10481), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13244) );
  AOI22_X1 U16442 ( .A1(n9680), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12686), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13243) );
  NAND2_X1 U16443 ( .A1(n13244), .A2(n13243), .ZN(n13255) );
  INV_X1 U16444 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13245) );
  NOR2_X1 U16445 ( .A1(n13246), .A2(n13245), .ZN(n13247) );
  AOI211_X1 U16446 ( .C1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .C2(n10481), .A(
        n13248), .B(n13247), .ZN(n13253) );
  AOI22_X1 U16447 ( .A1(n9681), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9652), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13252) );
  AOI22_X1 U16448 ( .A1(n12587), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10485), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13251) );
  AOI22_X1 U16449 ( .A1(n9685), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9649), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13250) );
  NAND4_X1 U16450 ( .A1(n13253), .A2(n13252), .A3(n13251), .A4(n13250), .ZN(
        n13254) );
  OAI21_X1 U16451 ( .B1(n13256), .B2(n13255), .A(n13254), .ZN(n13257) );
  XNOR2_X1 U16452 ( .A(n13258), .B(n13257), .ZN(n14445) );
  INV_X1 U16453 ( .A(n11178), .ZN(n13470) );
  AND2_X1 U16454 ( .A1(n11309), .A2(n14909), .ZN(n13468) );
  NAND2_X1 U16455 ( .A1(n13470), .A2(n13468), .ZN(n13259) );
  NOR2_X1 U16456 ( .A1(n13472), .A2(n13259), .ZN(n13260) );
  AOI21_X1 U16457 ( .B1(n13261), .B2(n14054), .A(n13260), .ZN(n13481) );
  NAND2_X1 U16458 ( .A1(n13481), .A2(n13262), .ZN(n13263) );
  NAND2_X1 U16459 ( .A1(n19293), .A2(n10979), .ZN(n19325) );
  OR2_X1 U16460 ( .A1(n14449), .A2(n13264), .ZN(n13266) );
  NAND2_X1 U16461 ( .A1(n19293), .A2(n13267), .ZN(n15247) );
  NOR4_X1 U16462 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13271) );
  NOR4_X1 U16463 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n13270) );
  NOR4_X1 U16464 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13269) );
  NOR4_X1 U16465 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n13268) );
  NAND4_X1 U16466 ( .A1(n13271), .A2(n13270), .A3(n13269), .A4(n13268), .ZN(
        n13276) );
  NOR4_X1 U16467 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n13274) );
  NOR4_X1 U16468 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13273) );
  NOR4_X1 U16469 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13272) );
  INV_X1 U16470 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20016) );
  NAND4_X1 U16471 ( .A1(n13274), .A2(n13273), .A3(n13272), .A4(n20016), .ZN(
        n13275) );
  MUX2_X1 U16472 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n15220), .Z(n19275) );
  INV_X1 U16473 ( .A(n19275), .ZN(n19375) );
  INV_X1 U16474 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13277) );
  OAI22_X1 U16475 ( .A1(n15247), .A2(n19375), .B1(n19293), .B2(n13277), .ZN(
        n13278) );
  AOI21_X1 U16476 ( .B1(n15407), .B2(n19321), .A(n13278), .ZN(n13282) );
  AND2_X1 U16477 ( .A1(n13279), .A2(n13764), .ZN(n13280) );
  NAND2_X1 U16478 ( .A1(n19293), .A2(n13280), .ZN(n13612) );
  NOR2_X2 U16479 ( .A1(n13612), .A2(n14108), .ZN(n19266) );
  NOR2_X2 U16480 ( .A1(n13612), .A2(n14107), .ZN(n19265) );
  AOI22_X1 U16481 ( .A1(n19266), .A2(BUF2_REG_30__SCAN_IN), .B1(n19265), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n13281) );
  AND2_X1 U16482 ( .A1(n13282), .A2(n13281), .ZN(n13283) );
  OAI21_X1 U16483 ( .B1(n14445), .B2(n19325), .A(n13283), .ZN(P2_U2889) );
  INV_X1 U16484 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16579) );
  NOR2_X1 U16485 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16579), .ZN(
        n13289) );
  INV_X1 U16486 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19019) );
  INV_X1 U16487 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16586) );
  AOI22_X1 U16488 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17819), .B1(
        n10059), .B2(n19019), .ZN(n13286) );
  NAND2_X1 U16489 ( .A1(n13284), .A2(n13286), .ZN(n13288) );
  AOI22_X1 U16490 ( .A1(n13285), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n15917), .B2(n17819), .ZN(n13287) );
  OAI22_X1 U16491 ( .A1(n13289), .A2(n13288), .B1(n13287), .B2(n13286), .ZN(
        n16562) );
  NAND2_X1 U16492 ( .A1(n16562), .A2(n18315), .ZN(n13305) );
  NAND3_X1 U16493 ( .A1(n19019), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13300) );
  INV_X1 U16494 ( .A(n13300), .ZN(n13297) );
  INV_X1 U16495 ( .A(n18152), .ZN(n13291) );
  NAND2_X1 U16496 ( .A1(n13291), .A2(n13290), .ZN(n18111) );
  NAND2_X1 U16497 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18394), .ZN(
        n18094) );
  NOR4_X1 U16498 ( .A1(n13292), .A2(n15858), .A3(n18111), .A4(n18094), .ZN(
        n15856) );
  INV_X1 U16499 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18993) );
  NOR2_X1 U16500 ( .A1(n18993), .A2(n18380), .ZN(n16558) );
  NOR3_X1 U16501 ( .A1(n17727), .A2(n15858), .A3(n16586), .ZN(n16569) );
  OAI211_X1 U16502 ( .C1(n18233), .C2(n16569), .A(n18394), .B(n13293), .ZN(
        n13294) );
  NAND2_X1 U16503 ( .A1(n18380), .A2(n13294), .ZN(n15922) );
  NAND2_X1 U16504 ( .A1(n18394), .A2(n18309), .ZN(n18381) );
  AOI221_X1 U16505 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15922), 
        .C1(n18381), .C2(n15922), .A(n19019), .ZN(n13295) );
  AOI211_X1 U16506 ( .C1(n13297), .C2(n15856), .A(n16558), .B(n13295), .ZN(
        n13303) );
  NAND2_X1 U16507 ( .A1(n17726), .A2(n16569), .ZN(n16567) );
  OR2_X1 U16508 ( .A1(n16579), .A2(n16567), .ZN(n13296) );
  AOI22_X1 U16509 ( .A1(n13298), .A2(n13297), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n13296), .ZN(n16565) );
  OR2_X1 U16510 ( .A1(n16565), .A2(n18391), .ZN(n13302) );
  NAND2_X1 U16511 ( .A1(n16569), .A2(n18090), .ZN(n16566) );
  OAI21_X1 U16512 ( .B1(n16579), .B2(n16566), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13299) );
  OAI21_X1 U16513 ( .B1(n13300), .B2(n16584), .A(n13299), .ZN(n16560) );
  NAND2_X1 U16514 ( .A1(n17559), .A2(n18384), .ZN(n18319) );
  INV_X1 U16515 ( .A(n18319), .ZN(n15859) );
  NAND2_X1 U16516 ( .A1(n13305), .A2(n13304), .ZN(P3_U2831) );
  NAND2_X1 U16517 ( .A1(n13309), .A2(n13308), .ZN(n14442) );
  INV_X1 U16518 ( .A(n20313), .ZN(n20254) );
  OAI21_X1 U16519 ( .B1(n16074), .B2(n13311), .A(n13310), .ZN(n13312) );
  NAND2_X1 U16520 ( .A1(n16447), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13315) );
  OAI211_X1 U16521 ( .C1(n16334), .C2(n16414), .A(n13316), .B(n13315), .ZN(
        n13318) );
  NOR2_X1 U16522 ( .A1(n13318), .A2(n10220), .ZN(n13321) );
  NAND2_X1 U16523 ( .A1(n13319), .A2(n19400), .ZN(n13320) );
  INV_X1 U16524 ( .A(n20892), .ZN(n15924) );
  OAI21_X1 U16525 ( .B1(n15924), .B2(n13323), .A(n13691), .ZN(n13324) );
  NAND2_X1 U16526 ( .A1(n13324), .A2(n14477), .ZN(n13329) );
  INV_X1 U16527 ( .A(n13326), .ZN(n13851) );
  INV_X1 U16528 ( .A(n14473), .ZN(n13327) );
  NAND3_X1 U16529 ( .A1(n13851), .A2(n13327), .A3(n20892), .ZN(n13328) );
  NAND4_X1 U16530 ( .A1(n20372), .A2(n20347), .A3(n14483), .A4(n13331), .ZN(
        n13352) );
  OR2_X1 U16531 ( .A1(n13330), .A2(n13352), .ZN(n13332) );
  NOR4_X1 U16532 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13337) );
  NOR4_X1 U16533 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n13336) );
  NOR4_X1 U16534 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13335) );
  NOR4_X1 U16535 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n13334) );
  AND4_X1 U16536 ( .A1(n13337), .A2(n13336), .A3(n13335), .A4(n13334), .ZN(
        n13342) );
  NOR4_X1 U16537 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n13340) );
  NOR4_X1 U16538 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n13339) );
  NOR4_X1 U16539 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13338) );
  INV_X1 U16540 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20904) );
  AND4_X1 U16541 ( .A1(n13340), .A2(n13339), .A3(n13338), .A4(n20904), .ZN(
        n13341) );
  NAND2_X1 U16542 ( .A1(n13342), .A2(n13341), .ZN(n13343) );
  NOR3_X1 U16543 ( .A1(n16057), .A2(n20311), .A3(n13821), .ZN(n13344) );
  AOI22_X1 U16544 ( .A1(n14708), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n16057), .ZN(n13345) );
  INV_X1 U16545 ( .A(n13345), .ZN(n13348) );
  INV_X1 U16546 ( .A(n20311), .ZN(n20312) );
  NOR2_X1 U16547 ( .A1(n13821), .A2(n20312), .ZN(n13346) );
  NAND2_X1 U16548 ( .A1(n14711), .A2(n13346), .ZN(n14691) );
  INV_X1 U16549 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20371) );
  NOR2_X1 U16550 ( .A1(n14691), .A2(n20371), .ZN(n13347) );
  NOR2_X1 U16551 ( .A1(n13348), .A2(n13347), .ZN(n13351) );
  AND2_X1 U16552 ( .A1(n14711), .A2(n20372), .ZN(n13349) );
  NAND2_X1 U16553 ( .A1(n14489), .A2(n13349), .ZN(n13350) );
  NAND2_X1 U16554 ( .A1(n13351), .A2(n13350), .ZN(P1_U2873) );
  NOR2_X1 U16555 ( .A1(n13352), .A2(n14485), .ZN(n13353) );
  NAND2_X1 U16556 ( .A1(n9793), .A2(n13353), .ZN(n13354) );
  OR2_X1 U16557 ( .A1(n14486), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13358) );
  INV_X1 U16558 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n13356) );
  NAND2_X1 U16559 ( .A1(n13357), .A2(n13356), .ZN(n13359) );
  NAND2_X1 U16560 ( .A1(n13358), .A2(n13359), .ZN(n13362) );
  MUX2_X1 U16561 ( .A(n13362), .B(n13359), .S(n13361), .Z(n14508) );
  NAND2_X1 U16562 ( .A1(n14510), .A2(n13361), .ZN(n13364) );
  OR2_X1 U16563 ( .A1(n13360), .A2(n13362), .ZN(n13363) );
  NAND2_X1 U16564 ( .A1(n13364), .A2(n13363), .ZN(n13366) );
  AOI22_X1 U16565 ( .A1(n14486), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n14485), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14484) );
  INV_X1 U16566 ( .A(n14484), .ZN(n13365) );
  INV_X1 U16567 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14503) );
  NOR2_X1 U16568 ( .A1(n14642), .A2(n14503), .ZN(n13367) );
  AOI21_X1 U16569 ( .B1(n10231), .B2(n13368), .A(n13367), .ZN(n13369) );
  NOR2_X1 U16570 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13372) );
  NOR4_X1 U16571 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13371) );
  NAND4_X1 U16572 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13372), .A4(n13371), .ZN(n13375) );
  NOR2_X1 U16573 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13375), .ZN(n16676)
         );
  INV_X1 U16574 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n21118) );
  NOR3_X1 U16575 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        n21118), .ZN(n13374) );
  NOR4_X1 U16576 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(P1_BE_N_REG_2__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n13373)
         );
  NAND4_X1 U16577 ( .A1(n20311), .A2(P1_W_R_N_REG_SCAN_IN), .A3(n13374), .A4(
        n13373), .ZN(U214) );
  NOR2_X1 U16578 ( .A1(n15220), .A2(n13375), .ZN(n16600) );
  NAND2_X1 U16579 ( .A1(n16600), .A2(U214), .ZN(U212) );
  AOI21_X1 U16580 ( .B1(n15383), .B2(n13386), .A(n13420), .ZN(n13404) );
  AOI21_X1 U16581 ( .B1(n16409), .B2(n13384), .A(n9773), .ZN(n19166) );
  AOI21_X1 U16582 ( .B1(n19187), .B2(n13382), .A(n13385), .ZN(n19192) );
  AOI21_X1 U16583 ( .B1(n16445), .B2(n9746), .A(n13383), .ZN(n15063) );
  AOI21_X1 U16584 ( .B1(n15394), .B2(n13380), .A(n13376), .ZN(n15392) );
  AOI21_X1 U16585 ( .B1(n16470), .B2(n13378), .A(n13381), .ZN(n19223) );
  AOI21_X1 U16586 ( .B1(n16484), .B2(n13377), .A(n13379), .ZN(n16472) );
  MUX2_X1 U16587 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n15720) );
  INV_X1 U16588 ( .A(n15720), .ZN(n14296) );
  MUX2_X1 U16589 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B(n13550), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n14251) );
  NAND2_X1 U16590 ( .A1(n14296), .A2(n14251), .ZN(n15132) );
  INV_X1 U16591 ( .A(n15132), .ZN(n15122) );
  OAI21_X1 U16592 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n13377), .ZN(n15136) );
  NAND2_X1 U16593 ( .A1(n15122), .A2(n15136), .ZN(n15117) );
  NOR2_X1 U16594 ( .A1(n16472), .A2(n15117), .ZN(n15102) );
  OAI21_X1 U16595 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13379), .A(
        n13378), .ZN(n19404) );
  NAND2_X1 U16596 ( .A1(n15102), .A2(n19404), .ZN(n19222) );
  NOR2_X1 U16597 ( .A1(n19223), .A2(n19222), .ZN(n19204) );
  OAI21_X1 U16598 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13381), .A(
        n13380), .ZN(n19205) );
  NAND2_X1 U16599 ( .A1(n19204), .A2(n19205), .ZN(n14272) );
  NOR2_X1 U16600 ( .A1(n15392), .A2(n14272), .ZN(n15085) );
  OAI21_X1 U16601 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n13376), .A(
        n9746), .ZN(n16459) );
  NAND2_X1 U16602 ( .A1(n15085), .A2(n16459), .ZN(n15073) );
  NOR2_X1 U16603 ( .A1(n15063), .A2(n15073), .ZN(n15057) );
  OAI21_X1 U16604 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n13383), .A(
        n13382), .ZN(n16435) );
  NAND2_X1 U16605 ( .A1(n15057), .A2(n16435), .ZN(n19191) );
  NOR2_X1 U16606 ( .A1(n19192), .A2(n19191), .ZN(n19176) );
  OAI21_X1 U16607 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n13385), .A(
        n13384), .ZN(n19177) );
  NAND2_X1 U16608 ( .A1(n19176), .A2(n19177), .ZN(n19161) );
  NOR2_X1 U16609 ( .A1(n19166), .A2(n19161), .ZN(n15036) );
  OAI21_X1 U16610 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n9773), .A(
        n13386), .ZN(n16400) );
  NAND2_X1 U16611 ( .A1(n15036), .A2(n16400), .ZN(n13391) );
  NOR2_X1 U16612 ( .A1(n13404), .A2(n13391), .ZN(n15016) );
  NAND2_X1 U16613 ( .A1(n14091), .A2(n19926), .ZN(n13389) );
  OR2_X1 U16614 ( .A1(n13390), .A2(n13389), .ZN(n16312) );
  INV_X1 U16615 ( .A(n16312), .ZN(n19227) );
  AOI211_X1 U16616 ( .C1(n13404), .C2(n13391), .A(n15016), .B(n15103), .ZN(
        n13419) );
  INV_X1 U16617 ( .A(n13392), .ZN(n13393) );
  NAND2_X1 U16618 ( .A1(n13393), .A2(n13539), .ZN(n13394) );
  NOR2_X1 U16619 ( .A1(n13395), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n13410) );
  OR2_X1 U16620 ( .A1(n19390), .A2(n13410), .ZN(n16297) );
  NAND2_X1 U16621 ( .A1(n19541), .A2(n14909), .ZN(n13405) );
  INV_X1 U16622 ( .A(n13405), .ZN(n13413) );
  NOR2_X1 U16623 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n13413), .ZN(n13396) );
  NAND2_X1 U16624 ( .A1(n13508), .A2(n13396), .ZN(n13397) );
  INV_X1 U16625 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n13403) );
  NAND2_X1 U16626 ( .A1(n13470), .A2(n13539), .ZN(n13398) );
  NOR2_X1 U16627 ( .A1(n13484), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19632) );
  INV_X1 U16628 ( .A(n19632), .ZN(n14198) );
  NOR2_X1 U16629 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n14198), .ZN(n13399) );
  NAND2_X1 U16630 ( .A1(n13399), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n16536) );
  AND3_X1 U16631 ( .A1(n19214), .A2(n16312), .A3(n16536), .ZN(n13400) );
  AND2_X2 U16632 ( .A1(n19215), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19221) );
  INV_X1 U16633 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20031) );
  OAI21_X1 U16634 ( .B1(n19215), .B2(n20031), .A(n19214), .ZN(n13401) );
  AOI21_X1 U16635 ( .B1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n19221), .A(
        n13401), .ZN(n13402) );
  OAI21_X1 U16636 ( .B1(n19218), .B2(n13403), .A(n13402), .ZN(n13418) );
  INV_X1 U16637 ( .A(n13404), .ZN(n15384) );
  NAND3_X1 U16638 ( .A1(n13414), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n13405), 
        .ZN(n13406) );
  NOR2_X2 U16639 ( .A1(n13464), .A2(n13406), .ZN(n19189) );
  OAI22_X1 U16640 ( .A1(n19151), .A2(n15384), .B1(n13407), .B2(n19216), .ZN(
        n13417) );
  OAI21_X1 U16641 ( .B1(n13408), .B2(n13409), .A(n15021), .ZN(n19273) );
  INV_X1 U16642 ( .A(n13410), .ZN(n14092) );
  AOI21_X1 U16643 ( .B1(n13412), .B2(n15027), .A(n13411), .ZN(n15598) );
  INV_X1 U16644 ( .A(n15598), .ZN(n14030) );
  INV_X1 U16645 ( .A(n13464), .ZN(n14907) );
  AND2_X1 U16646 ( .A1(n13414), .A2(n13413), .ZN(n13415) );
  NAND2_X1 U16647 ( .A1(n14907), .A2(n13415), .ZN(n19129) );
  OAI22_X1 U16648 ( .A1(n19273), .A2(n19231), .B1(n14030), .B2(n19129), .ZN(
        n13416) );
  OR4_X1 U16649 ( .A1(n13419), .A2(n13418), .A3(n13417), .A4(n13416), .ZN(
        P2_U2840) );
  OAI21_X1 U16650 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n13420), .A(
        n13421), .ZN(n15371) );
  AND2_X1 U16651 ( .A1(n15016), .A2(n15371), .ZN(n19147) );
  AND2_X1 U16652 ( .A1(n13421), .A2(n19141), .ZN(n13422) );
  OR2_X1 U16653 ( .A1(n13422), .A2(n13424), .ZN(n19146) );
  OAI21_X1 U16654 ( .B1(n10105), .B2(n19147), .A(n19146), .ZN(n19148) );
  NOR2_X1 U16655 ( .A1(n13424), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13425) );
  NOR2_X1 U16656 ( .A1(n13427), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13428) );
  OR2_X1 U16657 ( .A1(n13429), .A2(n13428), .ZN(n19131) );
  OAI21_X1 U16658 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n13429), .A(
        n13431), .ZN(n19113) );
  AOI21_X1 U16659 ( .B1(n15322), .B2(n13431), .A(n13430), .ZN(n19099) );
  INV_X1 U16660 ( .A(n19099), .ZN(n13432) );
  OAI21_X1 U16661 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n13430), .A(
        n13434), .ZN(n16386) );
  INV_X1 U16662 ( .A(n16386), .ZN(n15871) );
  AOI21_X1 U16663 ( .B1(n15297), .B2(n13434), .A(n13433), .ZN(n15300) );
  INV_X1 U16664 ( .A(n15300), .ZN(n13435) );
  OAI21_X1 U16665 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n13433), .A(
        n13437), .ZN(n16375) );
  INV_X1 U16666 ( .A(n16375), .ZN(n14961) );
  AND2_X1 U16667 ( .A1(n13437), .A2(n13436), .ZN(n13438) );
  NOR2_X1 U16668 ( .A1(n9776), .A2(n13438), .ZN(n15290) );
  OR2_X1 U16669 ( .A1(n9776), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13439) );
  NAND2_X1 U16670 ( .A1(n13440), .A2(n13439), .ZN(n15281) );
  INV_X1 U16671 ( .A(n15281), .ZN(n16325) );
  NAND2_X1 U16672 ( .A1(n13440), .A2(n15269), .ZN(n13441) );
  NAND2_X1 U16673 ( .A1(n13442), .A2(n13441), .ZN(n15270) );
  OAI21_X1 U16674 ( .B1(n16324), .B2(n15270), .A(n19227), .ZN(n13444) );
  OAI21_X1 U16675 ( .B1(n16324), .B2(n10085), .A(n15270), .ZN(n14938) );
  INV_X1 U16676 ( .A(n14938), .ZN(n13443) );
  AOI21_X1 U16677 ( .B1(n19151), .B2(n13444), .A(n13443), .ZN(n13457) );
  OAI22_X1 U16678 ( .A1(n13445), .A2(n19216), .B1(n20053), .B2(n19215), .ZN(
        n13456) );
  AOI22_X1 U16679 ( .A1(n19183), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n19221), .ZN(n13446) );
  INV_X1 U16680 ( .A(n13446), .ZN(n13455) );
  AOI21_X1 U16681 ( .B1(n13448), .B2(n15153), .A(n13447), .ZN(n15438) );
  INV_X1 U16682 ( .A(n15438), .ZN(n13453) );
  NAND2_X1 U16683 ( .A1(n13449), .A2(n13450), .ZN(n13451) );
  NAND2_X1 U16684 ( .A1(n13452), .A2(n13451), .ZN(n15436) );
  OAI22_X1 U16685 ( .A1(n13453), .A2(n19129), .B1(n15436), .B2(n19231), .ZN(
        n13454) );
  OR4_X1 U16686 ( .A1(n13457), .A2(n13456), .A3(n13455), .A4(n13454), .ZN(
        P2_U2828) );
  NOR3_X1 U16687 ( .A1(n14909), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n14091), 
        .ZN(n16538) );
  INV_X1 U16688 ( .A(n13543), .ZN(n13458) );
  NAND2_X1 U16689 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13458), .ZN(n15935) );
  INV_X1 U16690 ( .A(n15935), .ZN(n16539) );
  NOR3_X1 U16691 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n13459) );
  NOR4_X1 U16692 ( .A1(n16538), .A2(n16539), .A3(n16542), .A4(n13459), .ZN(
        P2_U3178) );
  OR2_X1 U16693 ( .A1(n10888), .A2(n16548), .ZN(n13460) );
  NOR2_X1 U16694 ( .A1(n13472), .A2(n13460), .ZN(n15131) );
  INV_X1 U16695 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13461) );
  OR2_X1 U16696 ( .A1(n19860), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13466) );
  OAI211_X1 U16697 ( .C1(n15131), .C2(n13461), .A(n13509), .B(n13466), .ZN(
        P2_U2814) );
  INV_X1 U16698 ( .A(n11309), .ZN(n13465) );
  INV_X1 U16699 ( .A(n13466), .ZN(n13462) );
  OAI21_X1 U16700 ( .B1(n13462), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n13464), 
        .ZN(n13463) );
  OAI21_X1 U16701 ( .B1(n13465), .B2(n13464), .A(n13463), .ZN(P2_U3612) );
  INV_X1 U16702 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n13467) );
  OAI22_X1 U16703 ( .A1(n14907), .A2(n13467), .B1(n14091), .B2(n13466), .ZN(
        P2_U2816) );
  NOR2_X1 U16704 ( .A1(n13468), .A2(n13477), .ZN(n13469) );
  NAND2_X1 U16705 ( .A1(n13470), .A2(n13469), .ZN(n13471) );
  NOR2_X1 U16706 ( .A1(n13472), .A2(n13471), .ZN(n14059) );
  OR2_X1 U16707 ( .A1(n14059), .A2(n16548), .ZN(n14918) );
  INV_X1 U16708 ( .A(n14918), .ZN(n13474) );
  OAI21_X1 U16709 ( .B1(n13474), .B2(n15936), .A(n13473), .ZN(P2_U2819) );
  INV_X1 U16710 ( .A(n10888), .ZN(n13475) );
  NAND2_X1 U16711 ( .A1(n13540), .A2(n13477), .ZN(n13483) );
  INV_X1 U16712 ( .A(n13478), .ZN(n13479) );
  AND3_X1 U16713 ( .A1(n13481), .A2(n13480), .A3(n13479), .ZN(n13482) );
  NAND2_X1 U16714 ( .A1(n13483), .A2(n13482), .ZN(n14077) );
  OAI22_X1 U16715 ( .A1(n15935), .A2(n15936), .B1(n13484), .B2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n13485) );
  AOI21_X1 U16716 ( .B1(n14077), .B2(n13539), .A(n13485), .ZN(n15737) );
  INV_X1 U16717 ( .A(n15737), .ZN(n13491) );
  NOR3_X1 U16718 ( .A1(n13488), .A2(n13487), .A3(n13486), .ZN(n14056) );
  INV_X1 U16719 ( .A(n20072), .ZN(n15733) );
  NAND3_X1 U16720 ( .A1(n13491), .A2(n14056), .A3(n15733), .ZN(n13489) );
  OAI21_X1 U16721 ( .B1(n13491), .B2(n13490), .A(n13489), .ZN(P2_U3595) );
  INV_X1 U16722 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13494) );
  INV_X1 U16723 ( .A(n14289), .ZN(n13493) );
  INV_X1 U16724 ( .A(n13546), .ZN(n13492) );
  AOI21_X1 U16725 ( .B1(n13494), .B2(n13493), .A(n13492), .ZN(n15714) );
  OAI21_X1 U16726 ( .B1(n13496), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13495), .ZN(n15713) );
  NAND2_X1 U16727 ( .A1(n19198), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n15708) );
  OAI21_X1 U16728 ( .B1(n16463), .B2(n15713), .A(n15708), .ZN(n13497) );
  AOI21_X1 U16729 ( .B1(n19397), .B2(n15714), .A(n13497), .ZN(n13500) );
  OAI21_X1 U16730 ( .B1(n16447), .B2(n13498), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13499) );
  OAI211_X1 U16731 ( .C1(n16414), .C2(n15709), .A(n13500), .B(n13499), .ZN(
        P2_U3014) );
  NOR2_X1 U16732 ( .A1(n14472), .A2(n14473), .ZN(n13533) );
  NAND2_X1 U16733 ( .A1(n13533), .A2(n14483), .ZN(n13504) );
  NOR2_X1 U16734 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20817), .ZN(n14130) );
  INV_X1 U16735 ( .A(n14011), .ZN(n13502) );
  AOI211_X1 U16736 ( .C1(P1_MEMORYFETCH_REG_SCAN_IN), .C2(n13504), .A(n14130), 
        .B(n13502), .ZN(n13503) );
  INV_X1 U16737 ( .A(n13503), .ZN(P1_U2801) );
  INV_X1 U16738 ( .A(n20973), .ZN(n13506) );
  OAI21_X1 U16739 ( .B1(n14130), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n13506), 
        .ZN(n13505) );
  OAI21_X1 U16740 ( .B1(n13507), .B2(n13506), .A(n13505), .ZN(P1_U3487) );
  INV_X1 U16741 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n15201) );
  AOI21_X2 U16742 ( .B1(n13508), .B2(n14909), .A(n13593), .ZN(n19388) );
  NAND2_X1 U16743 ( .A1(n19388), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13514) );
  NOR3_X1 U16744 ( .A1(n13509), .A2(n9666), .A3(n20003), .ZN(n19359) );
  INV_X1 U16745 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13510) );
  OR2_X1 U16746 ( .A1(n15220), .A2(n13510), .ZN(n13512) );
  NAND2_X1 U16747 ( .A1(n14107), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13511) );
  AND2_X1 U16748 ( .A1(n13512), .A2(n13511), .ZN(n19282) );
  INV_X1 U16749 ( .A(n19282), .ZN(n13513) );
  NAND2_X1 U16750 ( .A1(n19359), .A2(n13513), .ZN(n13528) );
  OAI211_X1 U16751 ( .C1(n19390), .C2(n15201), .A(n13514), .B(n13528), .ZN(
        P2_U2963) );
  INV_X1 U16752 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n13519) );
  NAND2_X1 U16753 ( .A1(n19388), .A2(P2_LWORD_REG_13__SCAN_IN), .ZN(n13518) );
  INV_X1 U16754 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16621) );
  OR2_X1 U16755 ( .A1(n15220), .A2(n16621), .ZN(n13516) );
  NAND2_X1 U16756 ( .A1(n14107), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13515) );
  AND2_X1 U16757 ( .A1(n13516), .A2(n13515), .ZN(n19278) );
  INV_X1 U16758 ( .A(n19278), .ZN(n13517) );
  NAND2_X1 U16759 ( .A1(n19359), .A2(n13517), .ZN(n13520) );
  OAI211_X1 U16760 ( .C1(n13519), .C2(n19390), .A(n13518), .B(n13520), .ZN(
        P2_U2980) );
  INV_X1 U16761 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14451) );
  NAND2_X1 U16762 ( .A1(n19388), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13521) );
  OAI211_X1 U16763 ( .C1(n19390), .C2(n14451), .A(n13521), .B(n13520), .ZN(
        P2_U2965) );
  INV_X1 U16764 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n13527) );
  NAND2_X1 U16765 ( .A1(n19388), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n13526) );
  INV_X1 U16766 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n13522) );
  OR2_X1 U16767 ( .A1(n15220), .A2(n13522), .ZN(n13524) );
  NAND2_X1 U16768 ( .A1(n14107), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13523) );
  AND2_X1 U16769 ( .A1(n13524), .A2(n13523), .ZN(n19287) );
  INV_X1 U16770 ( .A(n19287), .ZN(n13525) );
  NAND2_X1 U16771 ( .A1(n19359), .A2(n13525), .ZN(n13531) );
  OAI211_X1 U16772 ( .C1(n13527), .C2(n19390), .A(n13526), .B(n13531), .ZN(
        P2_U2976) );
  INV_X1 U16773 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n13530) );
  NAND2_X1 U16774 ( .A1(n19388), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13529) );
  OAI211_X1 U16775 ( .C1(n19390), .C2(n13530), .A(n13529), .B(n13528), .ZN(
        P2_U2978) );
  INV_X1 U16776 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n15215) );
  NAND2_X1 U16777 ( .A1(n19388), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13532) );
  OAI211_X1 U16778 ( .C1(n19390), .C2(n15215), .A(n13532), .B(n13531), .ZN(
        P2_U2961) );
  INV_X1 U16779 ( .A(n13533), .ZN(n13535) );
  INV_X1 U16780 ( .A(n13501), .ZN(n13534) );
  AOI22_X1 U16781 ( .A1(n13535), .A2(n13534), .B1(n15911), .B2(n11526), .ZN(
        n14482) );
  INV_X1 U16782 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n13536) );
  AOI21_X1 U16783 ( .B1(n14482), .B2(n14483), .A(n13536), .ZN(n13538) );
  NOR3_X1 U16784 ( .A1(n20958), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(n20971), 
        .ZN(n13537) );
  OR2_X1 U16785 ( .A1(n13538), .A2(n13537), .ZN(P1_U2803) );
  NAND2_X1 U16786 ( .A1(n13540), .A2(n13539), .ZN(n13541) );
  NAND2_X1 U16787 ( .A1(n13541), .A2(n19390), .ZN(n13542) );
  NAND2_X1 U16788 ( .A1(n19331), .A2(n14899), .ZN(n13734) );
  NOR2_X1 U16789 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13543), .ZN(n13728) );
  AOI22_X1 U16790 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n19339), .B1(n19356), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13544) );
  OAI21_X1 U16791 ( .B1(n13277), .B2(n13734), .A(n13544), .ZN(P2_U2921) );
  OAI21_X1 U16792 ( .B1(n14255), .B2(n13546), .A(n13545), .ZN(n13547) );
  XOR2_X1 U16793 ( .A(n13547), .B(n13550), .Z(n13622) );
  AOI21_X1 U16794 ( .B1(n13550), .B2(n13549), .A(n13548), .ZN(n13623) );
  INV_X1 U16795 ( .A(n13623), .ZN(n13551) );
  OAI22_X1 U16796 ( .A1(n16463), .A2(n13551), .B1(n20013), .B2(n19214), .ZN(
        n13552) );
  AOI21_X1 U16797 ( .B1(n19397), .B2(n13622), .A(n13552), .ZN(n13554) );
  MUX2_X1 U16798 ( .A(n19405), .B(n19394), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n13553) );
  OAI211_X1 U16799 ( .C1(n16414), .C2(n10460), .A(n13554), .B(n13553), .ZN(
        P2_U3013) );
  INV_X1 U16800 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n15230) );
  AOI22_X1 U16801 ( .A1(n13728), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13555) );
  OAI21_X1 U16802 ( .B1(n15230), .B2(n13734), .A(n13555), .ZN(P2_U2928) );
  INV_X1 U16803 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n19366) );
  AOI22_X1 U16804 ( .A1(n13728), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13556) );
  OAI21_X1 U16805 ( .B1(n19366), .B2(n13734), .A(n13556), .ZN(P2_U2927) );
  AOI22_X1 U16806 ( .A1(n13728), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13557) );
  OAI21_X1 U16807 ( .B1(n15215), .B2(n13734), .A(n13557), .ZN(P2_U2926) );
  AOI22_X1 U16808 ( .A1(n13728), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13558) );
  OAI21_X1 U16809 ( .B1(n15201), .B2(n13734), .A(n13558), .ZN(P2_U2924) );
  INV_X1 U16810 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n19374) );
  AOI22_X1 U16811 ( .A1(n19356), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13559) );
  OAI21_X1 U16812 ( .B1(n19374), .B2(n13734), .A(n13559), .ZN(P2_U2923) );
  INV_X1 U16813 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n13561) );
  OAI22_X1 U16814 ( .A1(n15220), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n14108), .ZN(n19413) );
  NOR2_X1 U16815 ( .A1(n19376), .A2(n19413), .ZN(n13578) );
  AOI21_X1 U16816 ( .B1(n13593), .B2(P2_EAX_REG_18__SCAN_IN), .A(n13578), .ZN(
        n13560) );
  OAI21_X1 U16817 ( .B1(n13599), .B2(n13561), .A(n13560), .ZN(P2_U2954) );
  INV_X1 U16818 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n13563) );
  INV_X1 U16819 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16638) );
  INV_X1 U16820 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18436) );
  AOI22_X1 U16821 ( .A1(n14108), .A2(n16638), .B1(n18436), .B2(n14107), .ZN(
        n16353) );
  INV_X1 U16822 ( .A(n16353), .ZN(n19418) );
  NOR2_X1 U16823 ( .A1(n19376), .A2(n19418), .ZN(n13586) );
  AOI21_X1 U16824 ( .B1(n13593), .B2(P2_EAX_REG_20__SCAN_IN), .A(n13586), .ZN(
        n13562) );
  OAI21_X1 U16825 ( .B1(n13599), .B2(n13563), .A(n13562), .ZN(P2_U2956) );
  INV_X1 U16826 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n13565) );
  AOI22_X1 U16827 ( .A1(n14108), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n14107), .ZN(n19319) );
  NOR2_X1 U16828 ( .A1(n19376), .A2(n19319), .ZN(n13589) );
  AOI21_X1 U16829 ( .B1(n13593), .B2(P2_EAX_REG_19__SCAN_IN), .A(n13589), .ZN(
        n13564) );
  OAI21_X1 U16830 ( .B1(n13599), .B2(n13565), .A(n13564), .ZN(P2_U2955) );
  INV_X1 U16831 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n13567) );
  AOI22_X1 U16832 ( .A1(n14108), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n14107), .ZN(n19441) );
  NOR2_X1 U16833 ( .A1(n19376), .A2(n19441), .ZN(n13570) );
  AOI21_X1 U16834 ( .B1(n13593), .B2(P2_EAX_REG_7__SCAN_IN), .A(n13570), .ZN(
        n13566) );
  OAI21_X1 U16835 ( .B1(n13599), .B2(n13567), .A(n13566), .ZN(P2_U2974) );
  INV_X1 U16836 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n13569) );
  INV_X1 U16837 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16634) );
  INV_X1 U16838 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18446) );
  AOI22_X1 U16839 ( .A1(n14108), .A2(n16634), .B1(n18446), .B2(n14107), .ZN(
        n16347) );
  INV_X1 U16840 ( .A(n16347), .ZN(n19431) );
  NOR2_X1 U16841 ( .A1(n19376), .A2(n19431), .ZN(n13573) );
  AOI21_X1 U16842 ( .B1(n13593), .B2(P2_EAX_REG_6__SCAN_IN), .A(n13573), .ZN(
        n13568) );
  OAI21_X1 U16843 ( .B1(n13599), .B2(n13569), .A(n13568), .ZN(P2_U2973) );
  INV_X1 U16844 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n13572) );
  AOI21_X1 U16845 ( .B1(n13593), .B2(P2_EAX_REG_23__SCAN_IN), .A(n13570), .ZN(
        n13571) );
  OAI21_X1 U16846 ( .B1(n13599), .B2(n13572), .A(n13571), .ZN(P2_U2959) );
  INV_X1 U16847 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n13575) );
  AOI21_X1 U16848 ( .B1(n13593), .B2(P2_EAX_REG_22__SCAN_IN), .A(n13573), .ZN(
        n13574) );
  OAI21_X1 U16849 ( .B1(n13599), .B2(n13575), .A(n13574), .ZN(P2_U2958) );
  INV_X1 U16850 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n13577) );
  AOI22_X1 U16851 ( .A1(n14108), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n14107), .ZN(n19424) );
  NOR2_X1 U16852 ( .A1(n19376), .A2(n19424), .ZN(n13583) );
  AOI21_X1 U16853 ( .B1(n13593), .B2(P2_EAX_REG_21__SCAN_IN), .A(n13583), .ZN(
        n13576) );
  OAI21_X1 U16854 ( .B1(n13599), .B2(n13577), .A(n13576), .ZN(P2_U2957) );
  INV_X1 U16855 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n13580) );
  AOI21_X1 U16856 ( .B1(P2_EAX_REG_2__SCAN_IN), .B2(n13593), .A(n13578), .ZN(
        n13579) );
  OAI21_X1 U16857 ( .B1(n13599), .B2(n13580), .A(n13579), .ZN(P2_U2969) );
  INV_X1 U16858 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n13582) );
  AOI22_X1 U16859 ( .A1(n14108), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n14107), .ZN(n19330) );
  NOR2_X1 U16860 ( .A1(n19376), .A2(n19330), .ZN(n13592) );
  AOI21_X1 U16861 ( .B1(P2_EAX_REG_1__SCAN_IN), .B2(n13593), .A(n13592), .ZN(
        n13581) );
  OAI21_X1 U16862 ( .B1(n13599), .B2(n13582), .A(n13581), .ZN(P2_U2968) );
  INV_X1 U16863 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n13585) );
  AOI21_X1 U16864 ( .B1(P2_EAX_REG_5__SCAN_IN), .B2(n13593), .A(n13583), .ZN(
        n13584) );
  OAI21_X1 U16865 ( .B1(n13599), .B2(n13585), .A(n13584), .ZN(P2_U2972) );
  INV_X1 U16866 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n13588) );
  AOI21_X1 U16867 ( .B1(P2_EAX_REG_4__SCAN_IN), .B2(n13593), .A(n13586), .ZN(
        n13587) );
  OAI21_X1 U16868 ( .B1(n13599), .B2(n13588), .A(n13587), .ZN(P2_U2971) );
  INV_X1 U16869 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n13591) );
  AOI21_X1 U16870 ( .B1(P2_EAX_REG_3__SCAN_IN), .B2(n13593), .A(n13589), .ZN(
        n13590) );
  OAI21_X1 U16871 ( .B1(n13599), .B2(n13591), .A(n13590), .ZN(P2_U2970) );
  INV_X1 U16872 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n13595) );
  AOI21_X1 U16873 ( .B1(n13593), .B2(P2_EAX_REG_17__SCAN_IN), .A(n13592), .ZN(
        n13594) );
  OAI21_X1 U16874 ( .B1(n13599), .B2(n13595), .A(n13594), .ZN(P2_U2953) );
  INV_X1 U16875 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n13597) );
  OAI22_X1 U16876 ( .A1(n14107), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n14108), .ZN(n19407) );
  INV_X1 U16877 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13596) );
  OAI222_X1 U16878 ( .A1(n13597), .A2(n13599), .B1(n19376), .B2(n19407), .C1(
        n19390), .C2(n13596), .ZN(P2_U2967) );
  INV_X1 U16879 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13600) );
  AOI22_X1 U16880 ( .A1(n14108), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n14107), .ZN(n19272) );
  INV_X1 U16881 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13598) );
  OAI222_X1 U16882 ( .A1(n13600), .A2(n13599), .B1(n19376), .B2(n19272), .C1(
        n19390), .C2(n13598), .ZN(P2_U2982) );
  MUX2_X1 U16883 ( .A(n14258), .B(n10460), .S(n19252), .Z(n13603) );
  OAI21_X1 U16884 ( .B1(n20091), .B2(n19254), .A(n13603), .ZN(P2_U2886) );
  NOR2_X1 U16885 ( .A1(n13605), .A2(n13604), .ZN(n13606) );
  NOR2_X1 U16886 ( .A1(n13607), .A2(n13606), .ZN(n15712) );
  INV_X1 U16887 ( .A(n15712), .ZN(n13615) );
  INV_X1 U16888 ( .A(n19321), .ZN(n15223) );
  INV_X1 U16889 ( .A(n13608), .ZN(n15722) );
  INV_X1 U16890 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19410) );
  NAND2_X1 U16891 ( .A1(n9676), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13609) );
  NAND4_X1 U16892 ( .A1(n10357), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13609), 
        .A4(n13484), .ZN(n13610) );
  NOR2_X1 U16893 ( .A1(n20101), .A2(n13615), .ZN(n19324) );
  AOI211_X1 U16894 ( .C1(n20101), .C2(n13615), .A(n19325), .B(n19324), .ZN(
        n13611) );
  AOI21_X1 U16895 ( .B1(P2_EAX_REG_0__SCAN_IN), .B2(n19320), .A(n13611), .ZN(
        n13614) );
  NAND2_X1 U16896 ( .A1(n15247), .A2(n13612), .ZN(n19295) );
  INV_X1 U16897 ( .A(n19407), .ZN(n19360) );
  NAND2_X1 U16898 ( .A1(n19295), .A2(n19360), .ZN(n13613) );
  OAI211_X1 U16899 ( .C1(n13615), .C2(n15223), .A(n13614), .B(n13613), .ZN(
        P2_U2919) );
  OAI21_X1 U16900 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n14459), .ZN(n13626) );
  XNOR2_X1 U16901 ( .A(n13616), .B(n13617), .ZN(n20096) );
  NOR3_X1 U16902 ( .A1(n13618), .A2(n19198), .A3(n13550), .ZN(n13619) );
  AOI21_X1 U16903 ( .B1(n19198), .B2(P2_REIP_REG_1__SCAN_IN), .A(n13619), .ZN(
        n13620) );
  OAI21_X1 U16904 ( .B1(n10460), .B2(n15710), .A(n13620), .ZN(n13621) );
  AOI21_X1 U16905 ( .B1(n16502), .B2(n20096), .A(n13621), .ZN(n13625) );
  AOI22_X1 U16906 ( .A1(n10972), .A2(n13623), .B1(n16530), .B2(n13622), .ZN(
        n13624) );
  OAI211_X1 U16907 ( .C1(n16501), .C2(n13626), .A(n13625), .B(n13624), .ZN(
        P2_U3045) );
  OAI211_X1 U16908 ( .C1(n13959), .C2(n13629), .A(n13628), .B(n13627), .ZN(
        n13630) );
  NOR2_X1 U16909 ( .A1(n13631), .A2(n13630), .ZN(n13634) );
  NOR2_X1 U16910 ( .A1(n15925), .A2(n15924), .ZN(n13632) );
  OAI211_X1 U16911 ( .C1(n15880), .C2(n13676), .A(n13632), .B(n14477), .ZN(
        n13633) );
  NAND2_X1 U16912 ( .A1(n13634), .A2(n13633), .ZN(n15889) );
  NAND2_X1 U16913 ( .A1(n15889), .A2(n14483), .ZN(n13636) );
  NAND2_X1 U16914 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16295) );
  NOR2_X1 U16915 ( .A1(n20971), .A2(n16295), .ZN(n13860) );
  NAND2_X1 U16916 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13860), .ZN(n13635) );
  NAND2_X1 U16917 ( .A1(n13636), .A2(n13635), .ZN(n13640) );
  AND2_X1 U16918 ( .A1(n20971), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13637) );
  OR2_X1 U16919 ( .A1(n13640), .A2(n13637), .ZN(n20953) );
  INV_X1 U16920 ( .A(n20469), .ZN(n20707) );
  OR2_X1 U16921 ( .A1(n13638), .A2(n20707), .ZN(n13639) );
  XNOR2_X1 U16922 ( .A(n13639), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20185) );
  NAND4_X1 U16923 ( .A1(n20185), .A2(n13718), .A3(n13851), .A4(n13640), .ZN(
        n13641) );
  OAI21_X1 U16924 ( .B1(n13642), .B2(n20953), .A(n13641), .ZN(P1_U3468) );
  OAI21_X1 U16925 ( .B1(n13645), .B2(n13644), .A(n13643), .ZN(n13646) );
  INV_X1 U16926 ( .A(n13646), .ZN(n14467) );
  AND2_X1 U16927 ( .A1(n19198), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n14461) );
  NAND2_X1 U16928 ( .A1(n13648), .A2(n13647), .ZN(n13649) );
  NAND2_X1 U16929 ( .A1(n13650), .A2(n13649), .ZN(n14457) );
  INV_X1 U16930 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13651) );
  OAI22_X1 U16931 ( .A1(n16465), .A2(n14457), .B1(n19394), .B2(n13651), .ZN(
        n13652) );
  AOI211_X1 U16932 ( .C1(n14467), .C2(n19400), .A(n14461), .B(n13652), .ZN(
        n13655) );
  NAND2_X1 U16933 ( .A1(n13653), .A2(n19399), .ZN(n13654) );
  OAI211_X1 U16934 ( .C1(n15136), .C2(n19405), .A(n13655), .B(n13654), .ZN(
        P2_U3012) );
  NOR2_X1 U16935 ( .A1(n19259), .A2(n15709), .ZN(n13656) );
  AOI21_X1 U16936 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n19259), .A(n13656), .ZN(
        n13657) );
  OAI21_X1 U16937 ( .B1(n19254), .B2(n20101), .A(n13657), .ZN(P2_U2887) );
  INV_X1 U16938 ( .A(n13658), .ZN(n13662) );
  INV_X1 U16939 ( .A(n13659), .ZN(n13661) );
  OAI21_X1 U16940 ( .B1(n13662), .B2(n13661), .A(n13660), .ZN(n13990) );
  NAND2_X1 U16941 ( .A1(n13663), .A2(n16074), .ZN(n13667) );
  AND2_X1 U16942 ( .A1(n20290), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13799) );
  OAI21_X1 U16943 ( .B1(n13665), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13664), .ZN(n13802) );
  NOR2_X1 U16944 ( .A1(n13802), .A2(n20115), .ZN(n13666) );
  AOI211_X1 U16945 ( .C1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n13667), .A(
        n13799), .B(n13666), .ZN(n13668) );
  OAI21_X1 U16946 ( .B1(n20254), .B2(n13990), .A(n13668), .ZN(P1_U2999) );
  INV_X1 U16947 ( .A(n13670), .ZN(n13671) );
  MUX2_X1 U16948 ( .A(n15123), .B(n15129), .S(n19252), .Z(n13672) );
  OAI21_X1 U16949 ( .B1(n20084), .B2(n19254), .A(n13672), .ZN(P2_U2885) );
  NAND2_X1 U16950 ( .A1(n13674), .A2(n13330), .ZN(n13675) );
  NOR2_X1 U16951 ( .A1(n13676), .A2(n13675), .ZN(n13678) );
  NAND3_X1 U16952 ( .A1(n13678), .A2(n13326), .A3(n13677), .ZN(n13679) );
  NOR2_X1 U16953 ( .A1(n13680), .A2(n13679), .ZN(n15878) );
  NAND2_X1 U16954 ( .A1(n15880), .A2(n10010), .ZN(n13703) );
  INV_X1 U16955 ( .A(n15877), .ZN(n13683) );
  INV_X1 U16956 ( .A(n13859), .ZN(n13682) );
  INV_X1 U16957 ( .A(n13704), .ZN(n13713) );
  NAND3_X1 U16958 ( .A1(n13683), .A2(n13682), .A3(n13713), .ZN(n13684) );
  OAI211_X1 U16959 ( .C1(n13673), .C2(n15878), .A(n13703), .B(n13684), .ZN(
        n15882) );
  INV_X1 U16960 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13685) );
  AOI22_X1 U16961 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n20300), .B2(n13685), .ZN(
        n13699) );
  NAND2_X1 U16962 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13697) );
  NOR2_X1 U16963 ( .A1(n13699), .A2(n13697), .ZN(n13687) );
  NOR3_X1 U16964 ( .A1(n13859), .A2(n13704), .A3(n20950), .ZN(n13686) );
  AOI211_X1 U16965 ( .C1(n15882), .C2(n13718), .A(n13687), .B(n13686), .ZN(
        n13689) );
  NAND2_X1 U16966 ( .A1(n20955), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13688) );
  OAI21_X1 U16967 ( .B1(n13689), .B2(n20955), .A(n13688), .ZN(P1_U3473) );
  XNOR2_X1 U16968 ( .A(n9985), .B(n13704), .ZN(n13698) );
  AND2_X1 U16969 ( .A1(n11511), .A2(n13698), .ZN(n13693) );
  NAND2_X1 U16970 ( .A1(n13691), .A2(n14470), .ZN(n13705) );
  INV_X1 U16971 ( .A(n13698), .ZN(n13692) );
  AOI22_X1 U16972 ( .A1(n15878), .A2(n13693), .B1(n13705), .B2(n13692), .ZN(
        n13696) );
  NAND2_X1 U16973 ( .A1(n15880), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13694) );
  MUX2_X1 U16974 ( .A(n13694), .B(n13703), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n13695) );
  OAI211_X1 U16975 ( .C1(n13690), .C2(n15878), .A(n13696), .B(n13695), .ZN(
        n13847) );
  INV_X1 U16976 ( .A(n13697), .ZN(n20952) );
  AOI222_X1 U16977 ( .A1(n13847), .A2(n13718), .B1(n20952), .B2(n13699), .C1(
        n13861), .C2(n13698), .ZN(n13701) );
  NAND2_X1 U16978 ( .A1(n20955), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13700) );
  OAI21_X1 U16979 ( .B1(n13701), .B2(n20955), .A(n13700), .ZN(P1_U3472) );
  INV_X1 U16980 ( .A(n20578), .ZN(n13873) );
  INV_X1 U16981 ( .A(n15880), .ZN(n13711) );
  AOI21_X1 U16982 ( .B1(n13707), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n13702), .ZN(n13710) );
  OR2_X1 U16983 ( .A1(n13703), .A2(n13845), .ZN(n13709) );
  MUX2_X1 U16984 ( .A(n13702), .B(n13845), .S(n13704), .Z(n13706) );
  OAI21_X1 U16985 ( .B1(n13707), .B2(n13706), .A(n13705), .ZN(n13708) );
  OAI211_X1 U16986 ( .C1(n13711), .C2(n13710), .A(n13709), .B(n13708), .ZN(
        n13712) );
  INV_X1 U16987 ( .A(n13712), .ZN(n13716) );
  AOI21_X1 U16988 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13713), .A(
        n13702), .ZN(n13714) );
  NAND2_X1 U16989 ( .A1(n11672), .A2(n13714), .ZN(n13717) );
  NAND3_X1 U16990 ( .A1(n15878), .A2(n11511), .A3(n13717), .ZN(n13715) );
  OAI211_X1 U16991 ( .C1(n13873), .C2(n15878), .A(n13716), .B(n13715), .ZN(
        n13844) );
  AOI22_X1 U16992 ( .A1(n13844), .A2(n13718), .B1(n13717), .B2(n13861), .ZN(
        n13720) );
  NAND2_X1 U16993 ( .A1(n20955), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13719) );
  OAI21_X1 U16994 ( .B1(n13720), .B2(n20955), .A(n13719), .ZN(P1_U3469) );
  INV_X1 U16995 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13722) );
  AOI22_X1 U16996 ( .A1(n13728), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19355), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13721) );
  OAI21_X1 U16997 ( .B1(n13722), .B2(n13734), .A(n13721), .ZN(P2_U2933) );
  INV_X1 U16998 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n19370) );
  AOI22_X1 U16999 ( .A1(n13728), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19355), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13723) );
  OAI21_X1 U17000 ( .B1(n19370), .B2(n13734), .A(n13723), .ZN(P2_U2925) );
  INV_X1 U17001 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15238) );
  AOI22_X1 U17002 ( .A1(n13728), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19355), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13724) );
  OAI21_X1 U17003 ( .B1(n15238), .B2(n13734), .A(n13724), .ZN(P2_U2930) );
  INV_X1 U17004 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13726) );
  AOI22_X1 U17005 ( .A1(n13728), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19355), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13725) );
  OAI21_X1 U17006 ( .B1(n13726), .B2(n13734), .A(n13725), .ZN(P2_U2931) );
  INV_X1 U17007 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n15246) );
  AOI22_X1 U17008 ( .A1(n13728), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19355), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13727) );
  OAI21_X1 U17009 ( .B1(n15246), .B2(n13734), .A(n13727), .ZN(P2_U2932) );
  INV_X1 U17010 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13730) );
  AOI22_X1 U17011 ( .A1(n13728), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19355), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13729) );
  OAI21_X1 U17012 ( .B1(n13730), .B2(n13734), .A(n13729), .ZN(P2_U2929) );
  INV_X1 U17013 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14355) );
  AOI22_X1 U17014 ( .A1(n19356), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19355), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13731) );
  OAI21_X1 U17015 ( .B1(n14355), .B2(n13734), .A(n13731), .ZN(P2_U2934) );
  INV_X1 U17016 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n19362) );
  AOI22_X1 U17017 ( .A1(n19356), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19355), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13732) );
  OAI21_X1 U17018 ( .B1(n19362), .B2(n13734), .A(n13732), .ZN(P2_U2935) );
  AOI22_X1 U17019 ( .A1(n19356), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19355), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13733) );
  OAI21_X1 U17020 ( .B1(n14451), .B2(n13734), .A(n13733), .ZN(P2_U2922) );
  INV_X1 U17021 ( .A(n13735), .ZN(n13739) );
  NAND2_X1 U17022 ( .A1(n13737), .A2(n13736), .ZN(n13766) );
  NAND2_X1 U17023 ( .A1(n13738), .A2(n13766), .ZN(n13740) );
  NAND2_X1 U17024 ( .A1(n13739), .A2(n13740), .ZN(n13742) );
  INV_X1 U17025 ( .A(n13740), .ZN(n13741) );
  NAND2_X1 U17026 ( .A1(n13741), .A2(n13735), .ZN(n13768) );
  INV_X1 U17027 ( .A(n20074), .ZN(n19299) );
  NOR2_X1 U17028 ( .A1(n13743), .A2(n19259), .ZN(n13744) );
  AOI21_X1 U17029 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n19259), .A(n13744), .ZN(
        n13745) );
  OAI21_X1 U17030 ( .B1(n19299), .B2(n19254), .A(n13745), .ZN(P2_U2884) );
  OR2_X1 U17031 ( .A1(n14054), .A2(n13746), .ZN(n14035) );
  INV_X1 U17032 ( .A(n13747), .ZN(n13748) );
  NAND2_X1 U17033 ( .A1(n13748), .A2(n10588), .ZN(n14033) );
  AOI22_X1 U17034 ( .A1(n14035), .A2(n14033), .B1(n10872), .B2(n10393), .ZN(
        n13751) );
  OR2_X1 U17035 ( .A1(n13743), .A2(n14066), .ZN(n13750) );
  OAI211_X1 U17036 ( .C1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(n13751), .A(
        n13750), .B(n13749), .ZN(n14048) );
  AOI22_X1 U17037 ( .A1(n20074), .A2(n16543), .B1(n15733), .B2(n14048), .ZN(
        n13758) );
  NAND2_X1 U17038 ( .A1(n13753), .A2(n13752), .ZN(n14040) );
  INV_X1 U17039 ( .A(n10872), .ZN(n13754) );
  NAND2_X1 U17040 ( .A1(n10393), .A2(n13754), .ZN(n14037) );
  NAND2_X1 U17041 ( .A1(n14037), .A2(n14033), .ZN(n13755) );
  AOI21_X1 U17042 ( .B1(n14040), .B2(n9654), .A(n13755), .ZN(n14046) );
  INV_X1 U17043 ( .A(n14046), .ZN(n13756) );
  AOI21_X1 U17044 ( .B1(n15733), .B2(n13756), .A(n15737), .ZN(n13757) );
  OAI22_X1 U17045 ( .A1(n13758), .A2(n15737), .B1(n13757), .B2(n14045), .ZN(
        P2_U3596) );
  XOR2_X1 U17046 ( .A(n13759), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13763)
         );
  AOI21_X1 U17047 ( .B1(n13760), .B2(n13779), .A(n9783), .ZN(n16517) );
  NOR2_X1 U17048 ( .A1(n19252), .A2(n10720), .ZN(n13761) );
  AOI21_X1 U17049 ( .B1(n16517), .B2(n19252), .A(n13761), .ZN(n13762) );
  OAI21_X1 U17050 ( .B1(n13763), .B2(n19254), .A(n13762), .ZN(P2_U2880) );
  NAND2_X1 U17051 ( .A1(n13764), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13765) );
  AND2_X1 U17052 ( .A1(n13766), .A2(n13765), .ZN(n13767) );
  AND2_X1 U17053 ( .A1(n13768), .A2(n13767), .ZN(n15095) );
  INV_X1 U17054 ( .A(n15095), .ZN(n13771) );
  NAND2_X1 U17055 ( .A1(n13769), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n15094) );
  INV_X1 U17056 ( .A(n15094), .ZN(n13770) );
  NAND2_X1 U17057 ( .A1(n13771), .A2(n13770), .ZN(n15096) );
  XOR2_X1 U17058 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n15096), .Z(n13776)
         );
  AND2_X1 U17059 ( .A1(n13772), .A2(n13773), .ZN(n13774) );
  OR2_X1 U17060 ( .A1(n13781), .A2(n13774), .ZN(n14299) );
  MUX2_X1 U17061 ( .A(n14299), .B(n10673), .S(n19259), .Z(n13775) );
  OAI21_X1 U17062 ( .B1(n13776), .B2(n19254), .A(n13775), .ZN(P2_U2882) );
  INV_X1 U17063 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n19213) );
  INV_X1 U17064 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13777) );
  NOR2_X1 U17065 ( .A1(n15096), .A2(n13777), .ZN(n13778) );
  OAI211_X1 U17066 ( .C1(n13778), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n19260), .B(n13759), .ZN(n13783) );
  OAI21_X1 U17067 ( .B1(n13781), .B2(n13780), .A(n13779), .ZN(n15702) );
  INV_X1 U17068 ( .A(n15702), .ZN(n19207) );
  NAND2_X1 U17069 ( .A1(n19207), .A2(n19252), .ZN(n13782) );
  OAI211_X1 U17070 ( .C1(n19252), .C2(n19213), .A(n13783), .B(n13782), .ZN(
        P2_U2881) );
  OAI21_X1 U17071 ( .B1(n10216), .B2(n11847), .A(n13784), .ZN(n13963) );
  INV_X1 U17072 ( .A(n13785), .ZN(n13950) );
  INV_X1 U17073 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n13786) );
  OAI22_X1 U17074 ( .A1(n16074), .A2(n13787), .B1(n10234), .B2(n13786), .ZN(
        n13788) );
  AOI21_X1 U17075 ( .B1(n13950), .B2(n20249), .A(n13788), .ZN(n13793) );
  OR2_X1 U17076 ( .A1(n13790), .A2(n13789), .ZN(n20277) );
  NAND3_X1 U17077 ( .A1(n20277), .A2(n13791), .A3(n20250), .ZN(n13792) );
  OAI211_X1 U17078 ( .C1(n13963), .C2(n20254), .A(n13793), .B(n13792), .ZN(
        P1_U2997) );
  AOI21_X1 U17079 ( .B1(n20276), .B2(n16168), .A(n20258), .ZN(n20301) );
  INV_X1 U17080 ( .A(n20301), .ZN(n13796) );
  OAI22_X1 U17081 ( .A1(n13796), .A2(n13795), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n13794), .ZN(n13801) );
  OR2_X1 U17082 ( .A1(n14486), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13798) );
  AND2_X1 U17083 ( .A1(n13798), .A2(n13797), .ZN(n13985) );
  AOI21_X1 U17084 ( .B1(n20292), .B2(n13985), .A(n13799), .ZN(n13800) );
  OAI211_X1 U17085 ( .C1(n16225), .C2(n13802), .A(n13801), .B(n13800), .ZN(
        P1_U3031) );
  NAND2_X1 U17086 ( .A1(n13804), .A2(n13803), .ZN(n13807) );
  INV_X1 U17087 ( .A(n13805), .ZN(n13806) );
  AND2_X1 U17088 ( .A1(n13807), .A2(n13806), .ZN(n19298) );
  XNOR2_X1 U17089 ( .A(n20084), .B(n19298), .ZN(n13812) );
  INV_X1 U17090 ( .A(n20096), .ZN(n13808) );
  NAND2_X1 U17091 ( .A1(n20091), .A2(n13808), .ZN(n13809) );
  OAI21_X1 U17092 ( .B1(n20091), .B2(n13808), .A(n13809), .ZN(n19323) );
  NOR2_X1 U17093 ( .A1(n19323), .A2(n19324), .ZN(n19322) );
  INV_X1 U17094 ( .A(n13809), .ZN(n13810) );
  NOR2_X1 U17095 ( .A1(n19322), .A2(n13810), .ZN(n13811) );
  NOR2_X1 U17096 ( .A1(n13811), .A2(n13812), .ZN(n19297) );
  AOI21_X1 U17097 ( .B1(n13812), .B2(n13811), .A(n19297), .ZN(n13815) );
  INV_X1 U17098 ( .A(n19413), .ZN(n16359) );
  AOI22_X1 U17099 ( .A1(n19295), .A2(n16359), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19320), .ZN(n13814) );
  INV_X1 U17100 ( .A(n19298), .ZN(n20086) );
  NAND2_X1 U17101 ( .A1(n20086), .A2(n19321), .ZN(n13813) );
  OAI211_X1 U17102 ( .C1(n13815), .C2(n19325), .A(n13814), .B(n13813), .ZN(
        P2_U2917) );
  NAND2_X1 U17103 ( .A1(n11510), .A2(n14479), .ZN(n13819) );
  AND2_X1 U17104 ( .A1(n13819), .A2(n13821), .ZN(n13816) );
  NAND2_X1 U17105 ( .A1(n20312), .A2(DATAI_2_), .ZN(n13818) );
  NAND2_X1 U17106 ( .A1(n20311), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13817) );
  AND2_X1 U17107 ( .A1(n13818), .A2(n13817), .ZN(n20332) );
  INV_X1 U17108 ( .A(n13819), .ZN(n13820) );
  INV_X1 U17109 ( .A(n13821), .ZN(n13822) );
  AND2_X1 U17110 ( .A1(n14711), .A2(n13822), .ZN(n13823) );
  INV_X1 U17111 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20227) );
  OAI222_X1 U17112 ( .A1(n13963), .A2(n14715), .B1(n20332), .B2(n14713), .C1(
        n14711), .C2(n20227), .ZN(P1_U2902) );
  NAND2_X1 U17113 ( .A1(n20312), .A2(DATAI_0_), .ZN(n13825) );
  NAND2_X1 U17114 ( .A1(n20311), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13824) );
  AND2_X1 U17115 ( .A1(n13825), .A2(n13824), .ZN(n20317) );
  INV_X1 U17116 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20234) );
  OAI222_X1 U17117 ( .A1(n13990), .A2(n14715), .B1(n20317), .B2(n14713), .C1(
        n14711), .C2(n20234), .ZN(P1_U2904) );
  OAI21_X1 U17118 ( .B1(n13828), .B2(n13827), .A(n13826), .ZN(n20253) );
  NAND2_X1 U17119 ( .A1(n20312), .A2(DATAI_1_), .ZN(n13830) );
  NAND2_X1 U17120 ( .A1(n20311), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13829) );
  AND2_X1 U17121 ( .A1(n13830), .A2(n13829), .ZN(n20327) );
  INV_X1 U17122 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20229) );
  OAI222_X1 U17123 ( .A1(n20253), .A2(n14715), .B1(n20327), .B2(n14713), .C1(
        n14711), .C2(n20229), .ZN(P1_U2903) );
  INV_X1 U17124 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n13838) );
  NAND2_X1 U17125 ( .A1(n9697), .A2(n13831), .ZN(n19247) );
  OAI211_X1 U17126 ( .C1(n9697), .C2(n13831), .A(n19247), .B(n19260), .ZN(
        n13837) );
  NAND2_X1 U17127 ( .A1(n13833), .A2(n13832), .ZN(n13835) );
  INV_X1 U17128 ( .A(n15047), .ZN(n13834) );
  NAND2_X1 U17129 ( .A1(n19252), .A2(n16442), .ZN(n13836) );
  OAI211_X1 U17130 ( .C1(n19252), .C2(n13838), .A(n13837), .B(n13836), .ZN(
        P2_U2878) );
  OAI21_X1 U17131 ( .B1(n13841), .B2(n13840), .A(n13839), .ZN(n13980) );
  NAND2_X1 U17132 ( .A1(n20312), .A2(DATAI_3_), .ZN(n13843) );
  NAND2_X1 U17133 ( .A1(n20311), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13842) );
  AND2_X1 U17134 ( .A1(n13843), .A2(n13842), .ZN(n20340) );
  INV_X1 U17135 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20225) );
  OAI222_X1 U17136 ( .A1(n13980), .A2(n14715), .B1(n20340), .B2(n14713), .C1(
        n14711), .C2(n20225), .ZN(P1_U2901) );
  INV_X1 U17137 ( .A(n15889), .ZN(n15884) );
  NOR2_X1 U17138 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n15884), .ZN(n13850) );
  MUX2_X1 U17139 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n13844), .S(
        n15889), .Z(n15894) );
  INV_X1 U17140 ( .A(n15894), .ZN(n13846) );
  INV_X1 U17141 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21100) );
  NAND2_X1 U17142 ( .A1(n21100), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13854) );
  OAI22_X1 U17143 ( .A1(n13846), .A2(P1_STATE2_REG_1__SCAN_IN), .B1(n13845), 
        .B2(n13854), .ZN(n13849) );
  NOR2_X1 U17144 ( .A1(n13847), .A2(n15884), .ZN(n15888) );
  NAND2_X1 U17145 ( .A1(n13854), .A2(n15888), .ZN(n13848) );
  OAI211_X1 U17146 ( .C1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(n13850), .A(
        n13849), .B(n13848), .ZN(n15900) );
  AOI21_X1 U17147 ( .B1(n20185), .B2(n13851), .A(n15884), .ZN(n13853) );
  OAI21_X1 U17148 ( .B1(n15889), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n16292), .ZN(n13852) );
  OR2_X1 U17149 ( .A1(n13853), .A2(n13852), .ZN(n13857) );
  INV_X1 U17150 ( .A(n13854), .ZN(n13855) );
  NAND2_X1 U17151 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n13855), .ZN(
        n13856) );
  NAND2_X1 U17152 ( .A1(n13857), .A2(n13856), .ZN(n15899) );
  INV_X1 U17153 ( .A(n15899), .ZN(n13858) );
  OAI21_X1 U17154 ( .B1(n15900), .B2(n13859), .A(n13858), .ZN(n13863) );
  OAI21_X1 U17155 ( .B1(n13863), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13860), .ZN(
        n13862) );
  NAND2_X1 U17156 ( .A1(n20968), .A2(n16292), .ZN(n20970) );
  NAND2_X1 U17157 ( .A1(n13862), .A2(n20475), .ZN(n20302) );
  NOR2_X1 U17158 ( .A1(n13863), .A2(n16295), .ZN(n15908) );
  INV_X1 U17159 ( .A(n11841), .ZN(n15879) );
  AND2_X1 U17160 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n11516), .ZN(n14896) );
  OAI22_X1 U17161 ( .A1(n11838), .A2(n20817), .B1(n15879), .B2(n14896), .ZN(
        n13864) );
  OAI21_X1 U17162 ( .B1(n15908), .B2(n13864), .A(n20302), .ZN(n13865) );
  OAI21_X1 U17163 ( .B1(n20302), .B2(n20751), .A(n13865), .ZN(P1_U3478) );
  INV_X1 U17164 ( .A(n13878), .ZN(n13867) );
  OR2_X1 U17165 ( .A1(n9675), .A2(n13867), .ZN(n20386) );
  INV_X1 U17166 ( .A(n20386), .ZN(n13869) );
  INV_X1 U17167 ( .A(n9675), .ZN(n13872) );
  NOR2_X1 U17168 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20817), .ZN(n20410) );
  INV_X1 U17169 ( .A(n20410), .ZN(n20705) );
  OAI22_X1 U17170 ( .A1(n13872), .A2(n20705), .B1(n13673), .B2(n14896), .ZN(
        n13868) );
  OAI21_X1 U17171 ( .B1(n13869), .B2(n13868), .A(n20302), .ZN(n13870) );
  OAI21_X1 U17172 ( .B1(n20302), .B2(n20638), .A(n13870), .ZN(P1_U3477) );
  INV_X1 U17173 ( .A(n20302), .ZN(n13881) );
  INV_X1 U17174 ( .A(n11830), .ZN(n13871) );
  OAI21_X1 U17175 ( .B1(n13872), .B2(n20553), .A(n20675), .ZN(n13877) );
  OAI22_X1 U17176 ( .A1(n20305), .A2(n20705), .B1(n13873), .B2(n14896), .ZN(
        n13876) );
  INV_X1 U17177 ( .A(n13874), .ZN(n13875) );
  NOR2_X1 U17178 ( .A1(n20702), .A2(n20386), .ZN(n20757) );
  AOI211_X1 U17179 ( .C1(n13878), .C2(n13877), .A(n13876), .B(n20757), .ZN(
        n13880) );
  NAND2_X1 U17180 ( .A1(n13881), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13879) );
  OAI21_X1 U17181 ( .B1(n13881), .B2(n13880), .A(n13879), .ZN(P1_U3475) );
  INV_X1 U17182 ( .A(n13882), .ZN(n19248) );
  NOR2_X1 U17183 ( .A1(n19247), .A2(n19248), .ZN(n19246) );
  XNOR2_X1 U17184 ( .A(n19246), .B(n19241), .ZN(n13889) );
  NAND2_X1 U17185 ( .A1(n13883), .A2(n15049), .ZN(n13885) );
  INV_X1 U17186 ( .A(n15632), .ZN(n13884) );
  AND2_X1 U17187 ( .A1(n13885), .A2(n13884), .ZN(n19194) );
  NOR2_X1 U17188 ( .A1(n19252), .A2(n13886), .ZN(n13887) );
  AOI21_X1 U17189 ( .B1(n19194), .B2(n19252), .A(n13887), .ZN(n13888) );
  OAI21_X1 U17190 ( .B1(n13889), .B2(n19254), .A(n13888), .ZN(P2_U2876) );
  XOR2_X1 U17191 ( .A(n13839), .B(n13890), .Z(n20239) );
  INV_X1 U17192 ( .A(n20239), .ZN(n13925) );
  NOR2_X1 U17193 ( .A1(n20311), .A2(DATAI_4_), .ZN(n13891) );
  AOI21_X1 U17194 ( .B1(n20311), .B2(n16638), .A(n13891), .ZN(n20348) );
  AOI22_X1 U17195 ( .A1(n16059), .A2(n20348), .B1(n16057), .B2(
        P1_EAX_REG_4__SCAN_IN), .ZN(n13892) );
  OAI21_X1 U17196 ( .B1(n13925), .B2(n14715), .A(n13892), .ZN(P1_U2900) );
  OAI21_X1 U17197 ( .B1(n13895), .B2(n13894), .A(n13893), .ZN(n20267) );
  INV_X1 U17198 ( .A(n13980), .ZN(n13898) );
  AOI22_X1 U17199 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20290), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n13896) );
  OAI21_X1 U17200 ( .B1(n20243), .B2(n13973), .A(n13896), .ZN(n13897) );
  AOI21_X1 U17201 ( .B1(n13898), .B2(n20313), .A(n13897), .ZN(n13899) );
  OAI21_X1 U17202 ( .B1(n20267), .B2(n20115), .A(n13899), .ZN(P1_U2996) );
  OR2_X1 U17203 ( .A1(n13901), .A2(n13900), .ZN(n13902) );
  NAND2_X1 U17204 ( .A1(n13927), .A2(n13902), .ZN(n20287) );
  OAI22_X1 U17205 ( .A1(n20287), .A2(n14643), .B1(n13953), .B2(n14642), .ZN(
        n13903) );
  INV_X1 U17206 ( .A(n13903), .ZN(n13904) );
  OAI21_X1 U17207 ( .B1(n13963), .B2(n14655), .A(n13904), .ZN(P1_U2870) );
  NAND2_X1 U17208 ( .A1(n13906), .A2(n13905), .ZN(n13908) );
  INV_X1 U17209 ( .A(n15025), .ZN(n13907) );
  AND2_X1 U17210 ( .A1(n13908), .A2(n13907), .ZN(n19165) );
  INV_X1 U17211 ( .A(n19165), .ZN(n13914) );
  OAI211_X1 U17212 ( .C1(n9771), .C2(n13911), .A(n13910), .B(n19260), .ZN(
        n13913) );
  NAND2_X1 U17213 ( .A1(n19259), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13912) );
  OAI211_X1 U17214 ( .C1(n13914), .C2(n19259), .A(n13913), .B(n13912), .ZN(
        P2_U2874) );
  INV_X1 U17215 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14176) );
  NAND3_X1 U17216 ( .A1(n15880), .A2(n14483), .A3(n14477), .ZN(n13915) );
  NAND2_X1 U17217 ( .A1(n13915), .A2(n14193), .ZN(n13917) );
  NAND2_X1 U17218 ( .A1(n20201), .A2(n13918), .ZN(n14249) );
  NOR2_X1 U17219 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16295), .ZN(n14243) );
  AOI22_X1 U17220 ( .A1(n14243), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20218), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13919) );
  OAI21_X1 U17221 ( .B1(n14176), .B2(n14249), .A(n13919), .ZN(P1_U2913) );
  INV_X1 U17222 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n14671) );
  AOI22_X1 U17223 ( .A1(n14243), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20218), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13920) );
  OAI21_X1 U17224 ( .B1(n14671), .B2(n14249), .A(n13920), .ZN(P1_U2911) );
  INV_X1 U17225 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14167) );
  AOI22_X1 U17226 ( .A1(n20231), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20218), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13921) );
  OAI21_X1 U17227 ( .B1(n14167), .B2(n14249), .A(n13921), .ZN(P1_U2909) );
  INV_X1 U17228 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14140) );
  AOI22_X1 U17229 ( .A1(n20231), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20218), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13922) );
  OAI21_X1 U17230 ( .B1(n14140), .B2(n14249), .A(n13922), .ZN(P1_U2907) );
  INV_X1 U17231 ( .A(n14642), .ZN(n14653) );
  AOI22_X1 U17232 ( .A1(n13368), .A2(n13985), .B1(P1_EBX_REG_0__SCAN_IN), .B2(
        n14653), .ZN(n13923) );
  OAI21_X1 U17233 ( .B1(n13990), .B2(n14655), .A(n13923), .ZN(P1_U2872) );
  XNOR2_X1 U17234 ( .A(n13964), .B(n13966), .ZN(n20257) );
  AOI22_X1 U17235 ( .A1(n20257), .A2(n13368), .B1(n14653), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n13924) );
  OAI21_X1 U17236 ( .B1(n13925), .B2(n14655), .A(n13924), .ZN(P1_U2868) );
  NAND2_X1 U17237 ( .A1(n13927), .A2(n13926), .ZN(n13928) );
  AND2_X1 U17238 ( .A1(n13964), .A2(n13928), .ZN(n20266) );
  AOI22_X1 U17239 ( .A1(n20266), .A2(n13368), .B1(n14653), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n13929) );
  OAI21_X1 U17240 ( .B1(n13980), .B2(n14655), .A(n13929), .ZN(P1_U2869) );
  NAND2_X1 U17241 ( .A1(n13932), .A2(n13931), .ZN(n13933) );
  AND2_X1 U17242 ( .A1(n13930), .A2(n13933), .ZN(n20179) );
  INV_X1 U17243 ( .A(n20179), .ZN(n13970) );
  INV_X1 U17244 ( .A(DATAI_5_), .ZN(n21041) );
  NAND2_X1 U17245 ( .A1(n20312), .A2(n21041), .ZN(n13935) );
  INV_X1 U17246 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16636) );
  NAND2_X1 U17247 ( .A1(n20311), .A2(n16636), .ZN(n13934) );
  AND2_X1 U17248 ( .A1(n13935), .A2(n13934), .ZN(n20354) );
  INV_X1 U17249 ( .A(n20354), .ZN(n13936) );
  OAI222_X1 U17250 ( .A1(n13970), .A2(n14715), .B1(n13936), .B2(n14713), .C1(
        n14711), .C2(n11873), .ZN(P1_U2899) );
  OR2_X1 U17251 ( .A1(n11516), .A2(n20970), .ZN(n15909) );
  NAND2_X1 U17252 ( .A1(n11824), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13937) );
  MUX2_X1 U17253 ( .A(n15909), .B(n13937), .S(n20971), .Z(n13938) );
  NAND2_X1 U17254 ( .A1(n13938), .A2(n10234), .ZN(n13939) );
  NOR2_X1 U17255 ( .A1(n13948), .A2(n16292), .ZN(n13940) );
  NOR2_X1 U17256 ( .A1(n13960), .A2(n11526), .ZN(n13941) );
  OR2_X1 U17257 ( .A1(n20165), .A2(n13941), .ZN(n20198) );
  OR2_X1 U17258 ( .A1(n13942), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13945) );
  INV_X1 U17259 ( .A(n13945), .ZN(n15906) );
  OR2_X1 U17260 ( .A1(n20175), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n14022) );
  NAND2_X1 U17261 ( .A1(n14022), .A2(n20144), .ZN(n13972) );
  AND2_X1 U17262 ( .A1(n13943), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13954) );
  INV_X1 U17263 ( .A(n13954), .ZN(n13944) );
  AND2_X1 U17264 ( .A1(n13945), .A2(n13944), .ZN(n13946) );
  NOR2_X1 U17265 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n20175), .ZN(n13971) );
  AOI22_X1 U17266 ( .A1(n20186), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n13971), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n13952) );
  AND2_X1 U17267 ( .A1(n13948), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13949) );
  NAND2_X1 U17268 ( .A1(n20171), .A2(n13950), .ZN(n13951) );
  OAI211_X1 U17269 ( .C1(n20190), .C2(n13953), .A(n13952), .B(n13951), .ZN(
        n13958) );
  OAI21_X1 U17270 ( .B1(n15924), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n13954), 
        .ZN(n13955) );
  NOR2_X1 U17271 ( .A1(n20162), .A2(n20287), .ZN(n13957) );
  AOI211_X1 U17272 ( .C1(n13972), .C2(P1_REIP_REG_2__SCAN_IN), .A(n13958), .B(
        n13957), .ZN(n13962) );
  INV_X1 U17273 ( .A(n13690), .ZN(n20308) );
  NOR2_X1 U17274 ( .A1(n13960), .A2(n13959), .ZN(n20184) );
  NAND2_X1 U17275 ( .A1(n20308), .A2(n20184), .ZN(n13961) );
  OAI211_X1 U17276 ( .C1(n13963), .C2(n14024), .A(n13962), .B(n13961), .ZN(
        P1_U2838) );
  INV_X1 U17277 ( .A(n13964), .ZN(n13967) );
  AOI21_X1 U17278 ( .B1(n13967), .B2(n13966), .A(n13965), .ZN(n13968) );
  NOR2_X1 U17279 ( .A1(n13968), .A2(n9772), .ZN(n20178) );
  AOI22_X1 U17280 ( .A1(n20178), .A2(n13368), .B1(n14653), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n13969) );
  OAI21_X1 U17281 ( .B1(n13970), .B2(n14640), .A(n13969), .ZN(P1_U2867) );
  OAI21_X1 U17282 ( .B1(n13972), .B2(n13971), .A(P1_REIP_REG_3__SCAN_IN), .ZN(
        n13979) );
  INV_X1 U17283 ( .A(n13973), .ZN(n13974) );
  AOI22_X1 U17284 ( .A1(n13974), .A2(n20171), .B1(n20186), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13978) );
  INV_X1 U17285 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20905) );
  AND3_X1 U17286 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(n20905), .ZN(n13975) );
  AOI22_X1 U17287 ( .A1(n20146), .A2(n13975), .B1(n20196), .B2(n20266), .ZN(
        n13977) );
  NAND2_X1 U17288 ( .A1(n20173), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n13976) );
  NAND4_X1 U17289 ( .A1(n13979), .A2(n13978), .A3(n13977), .A4(n13976), .ZN(
        n13982) );
  NOR2_X1 U17290 ( .A1(n13980), .A2(n14024), .ZN(n13981) );
  AOI211_X1 U17291 ( .C1(n20184), .C2(n20578), .A(n13982), .B(n13981), .ZN(
        n13983) );
  INV_X1 U17292 ( .A(n13983), .ZN(P1_U2837) );
  XNOR2_X1 U17293 ( .A(n13984), .B(n14485), .ZN(n20289) );
  INV_X1 U17294 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n14020) );
  OAI222_X1 U17295 ( .A1(n20289), .A2(n14643), .B1(n14020), .B2(n14633), .C1(
        n14640), .C2(n20253), .ZN(P1_U2871) );
  NAND2_X1 U17296 ( .A1(n20175), .A2(n20144), .ZN(n15970) );
  NAND2_X1 U17297 ( .A1(n15970), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13989) );
  NAND2_X1 U17298 ( .A1(n20196), .A2(n13985), .ZN(n13988) );
  NAND2_X1 U17299 ( .A1(n20173), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13987) );
  OAI21_X1 U17300 ( .B1(n20186), .B2(n20171), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13986) );
  NAND4_X1 U17301 ( .A1(n13989), .A2(n13988), .A3(n13987), .A4(n13986), .ZN(
        n13992) );
  NOR2_X1 U17302 ( .A1(n13990), .A2(n14024), .ZN(n13991) );
  AOI211_X1 U17303 ( .C1(n20184), .C2(n11841), .A(n13992), .B(n13991), .ZN(
        n13993) );
  INV_X1 U17304 ( .A(n13993), .ZN(P1_U2840) );
  AOI21_X1 U17305 ( .B1(n13996), .B2(n13930), .A(n13995), .ZN(n20166) );
  NOR2_X1 U17306 ( .A1(n9772), .A2(n13997), .ZN(n13998) );
  OR2_X1 U17307 ( .A1(n14096), .A2(n13998), .ZN(n20161) );
  OAI22_X1 U17308 ( .A1(n20161), .A2(n14643), .B1(n13999), .B2(n14642), .ZN(
        n14000) );
  AOI21_X1 U17309 ( .B1(n20166), .B2(n14001), .A(n14000), .ZN(n14002) );
  INV_X1 U17310 ( .A(n14002), .ZN(P1_U2866) );
  OAI21_X1 U17311 ( .B1(n13995), .B2(n14005), .A(n14004), .ZN(n20149) );
  INV_X1 U17312 ( .A(DATAI_7_), .ZN(n21035) );
  NAND2_X1 U17313 ( .A1(n20312), .A2(n21035), .ZN(n14007) );
  INV_X1 U17314 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16632) );
  NAND2_X1 U17315 ( .A1(n20311), .A2(n16632), .ZN(n14006) );
  AND2_X1 U17316 ( .A1(n14007), .A2(n14006), .ZN(n20376) );
  INV_X1 U17317 ( .A(n20376), .ZN(n14008) );
  OAI222_X1 U17318 ( .A1(n20149), .A2(n14715), .B1(n14008), .B2(n14713), .C1(
        n14711), .C2(n11892), .ZN(P1_U2897) );
  AND2_X1 U17319 ( .A1(n14009), .A2(n15924), .ZN(n14010) );
  NOR2_X2 U17320 ( .A1(n14190), .A2(n20326), .ZN(n14179) );
  INV_X1 U17321 ( .A(n14179), .ZN(n14014) );
  INV_X1 U17322 ( .A(DATAI_15_), .ZN(n21060) );
  INV_X1 U17323 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n16617) );
  MUX2_X1 U17324 ( .A(n21060), .B(n16617), .S(n20311), .Z(n14714) );
  INV_X1 U17325 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n14013) );
  INV_X1 U17326 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14712) );
  OAI222_X1 U17327 ( .A1(n14014), .A2(n14714), .B1(n14013), .B2(n14012), .C1(
        n14712), .C2(n14193), .ZN(P1_U2967) );
  INV_X1 U17328 ( .A(n20166), .ZN(n14017) );
  NOR2_X1 U17329 ( .A1(n20311), .A2(DATAI_6_), .ZN(n14015) );
  AOI21_X1 U17330 ( .B1(n20311), .B2(n16634), .A(n14015), .ZN(n20361) );
  INV_X1 U17331 ( .A(n20361), .ZN(n14016) );
  OAI222_X1 U17332 ( .A1(n14017), .A2(n14715), .B1(n14016), .B2(n14713), .C1(
        n20220), .C2(n14711), .ZN(P1_U2898) );
  INV_X1 U17333 ( .A(n13673), .ZN(n20783) );
  INV_X1 U17334 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20248) );
  INV_X1 U17335 ( .A(n20144), .ZN(n14128) );
  AOI22_X1 U17336 ( .A1(n20171), .A2(n20248), .B1(n14128), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n14019) );
  NAND2_X1 U17337 ( .A1(n20186), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14018) );
  OAI211_X1 U17338 ( .C1(n20190), .C2(n14020), .A(n14019), .B(n14018), .ZN(
        n14021) );
  INV_X1 U17339 ( .A(n14021), .ZN(n14023) );
  OAI211_X1 U17340 ( .C1(n20162), .C2(n20289), .A(n14023), .B(n14022), .ZN(
        n14026) );
  NOR2_X1 U17341 ( .A1(n20253), .A2(n14024), .ZN(n14025) );
  AOI211_X1 U17342 ( .C1(n20184), .C2(n20783), .A(n14026), .B(n14025), .ZN(
        n14027) );
  INV_X1 U17343 ( .A(n14027), .ZN(P1_U2839) );
  XNOR2_X1 U17344 ( .A(n14028), .B(n14029), .ZN(n14032) );
  MUX2_X1 U17345 ( .A(n13403), .B(n14030), .S(n19252), .Z(n14031) );
  OAI21_X1 U17346 ( .B1(n14032), .B2(n19254), .A(n14031), .ZN(P2_U2872) );
  OR2_X1 U17347 ( .A1(n15129), .A2(n14066), .ZN(n14043) );
  NAND2_X1 U17348 ( .A1(n9654), .A2(n14033), .ZN(n14034) );
  INV_X1 U17349 ( .A(n14034), .ZN(n14041) );
  NOR2_X1 U17350 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14038) );
  NAND2_X1 U17351 ( .A1(n14035), .A2(n14034), .ZN(n14036) );
  OAI21_X1 U17352 ( .B1(n14038), .B2(n14037), .A(n14036), .ZN(n14039) );
  AOI21_X1 U17353 ( .B1(n14041), .B2(n14040), .A(n14039), .ZN(n14042) );
  NAND2_X1 U17354 ( .A1(n14043), .A2(n14042), .ZN(n15732) );
  INV_X1 U17355 ( .A(n14077), .ZN(n14044) );
  MUX2_X1 U17356 ( .A(n15732), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n14044), .Z(n14090) );
  AOI21_X1 U17357 ( .B1(n14077), .B2(n14046), .A(n14045), .ZN(n14047) );
  OR2_X1 U17358 ( .A1(n14048), .A2(n14047), .ZN(n14050) );
  OR2_X1 U17359 ( .A1(n14077), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14049) );
  NAND2_X1 U17360 ( .A1(n14050), .A2(n14049), .ZN(n14078) );
  INV_X1 U17361 ( .A(n14078), .ZN(n14089) );
  OAI22_X1 U17362 ( .A1(n14055), .A2(n14052), .B1(n14051), .B2(n11178), .ZN(
        n14053) );
  AOI21_X1 U17363 ( .B1(n14055), .B2(n14054), .A(n14053), .ZN(n14915) );
  OR2_X1 U17364 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(P2_MORE_REG_SCAN_IN), .ZN(
        n14058) );
  AOI211_X1 U17365 ( .C1(n14059), .C2(n14058), .A(n14057), .B(n14056), .ZN(
        n14060) );
  OAI211_X1 U17366 ( .C1(n14077), .C2(n13490), .A(n14915), .B(n14060), .ZN(
        n14088) );
  NAND2_X1 U17367 ( .A1(n20081), .A2(n20088), .ZN(n19504) );
  INV_X1 U17368 ( .A(n19504), .ZN(n19474) );
  NOR2_X1 U17369 ( .A1(n14078), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14085) );
  OR2_X1 U17370 ( .A1(n15709), .A2(n14066), .ZN(n14065) );
  INV_X1 U17371 ( .A(n11180), .ZN(n14062) );
  NAND2_X1 U17372 ( .A1(n14062), .A2(n14061), .ZN(n14073) );
  MUX2_X1 U17373 ( .A(n14073), .B(n10393), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n14063) );
  INV_X1 U17374 ( .A(n14063), .ZN(n14064) );
  NAND2_X1 U17375 ( .A1(n14065), .A2(n14064), .ZN(n15721) );
  NOR2_X1 U17376 ( .A1(n15721), .A2(n20106), .ZN(n14083) );
  INV_X1 U17377 ( .A(n14066), .ZN(n14067) );
  NAND2_X1 U17378 ( .A1(n14068), .A2(n14067), .ZN(n14076) );
  INV_X1 U17379 ( .A(n9677), .ZN(n14071) );
  NAND2_X1 U17380 ( .A1(n14069), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14070) );
  NAND2_X1 U17381 ( .A1(n14071), .A2(n14070), .ZN(n14072) );
  AOI22_X1 U17382 ( .A1(n14074), .A2(n10393), .B1(n14073), .B2(n14072), .ZN(
        n14075) );
  NAND2_X1 U17383 ( .A1(n14076), .A2(n14075), .ZN(n15728) );
  NAND2_X1 U17384 ( .A1(n15728), .A2(n20098), .ZN(n14082) );
  OAI21_X1 U17385 ( .B1(n15728), .B2(n20098), .A(n14077), .ZN(n14081) );
  NOR2_X1 U17386 ( .A1(n14078), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14079) );
  AOI211_X1 U17387 ( .C1(n14090), .C2(n20081), .A(n19474), .B(n14079), .ZN(
        n14080) );
  AOI211_X1 U17388 ( .C1(n14083), .C2(n14082), .A(n14081), .B(n14080), .ZN(
        n14084) );
  AOI211_X1 U17389 ( .C1(n14090), .C2(n19474), .A(n14085), .B(n14084), .ZN(
        n14086) );
  NOR2_X1 U17390 ( .A1(n14086), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n14087) );
  AOI211_X1 U17391 ( .C1(n14090), .C2(n14089), .A(n14088), .B(n14087), .ZN(
        n16549) );
  AOI21_X1 U17392 ( .B1(n16549), .B2(n11320), .A(n14091), .ZN(n14194) );
  OR3_X1 U17393 ( .A1(n13392), .A2(n9676), .A3(n14092), .ZN(n14094) );
  NOR2_X1 U17394 ( .A1(n14093), .A2(n19926), .ZN(n14906) );
  NAND2_X1 U17395 ( .A1(n14094), .A2(n14906), .ZN(n14195) );
  OAI21_X1 U17396 ( .B1(n14194), .B2(n14195), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n16544) );
  INV_X1 U17397 ( .A(n16544), .ZN(n14199) );
  OAI21_X1 U17398 ( .B1(n14199), .B2(n13484), .A(n15935), .ZN(P2_U3593) );
  OAI21_X1 U17399 ( .B1(n14096), .B2(n14095), .A(n14123), .ZN(n16266) );
  OAI222_X1 U17400 ( .A1(n16266), .A2(n14643), .B1(n20143), .B2(n14633), .C1(
        n14640), .C2(n20149), .ZN(P1_U2865) );
  NAND2_X1 U17401 ( .A1(n19989), .A2(n19473), .ZN(n14098) );
  AOI21_X1 U17402 ( .B1(n14098), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19860), 
        .ZN(n14102) );
  NAND2_X1 U17403 ( .A1(n19474), .A2(n20098), .ZN(n19448) );
  NOR2_X1 U17404 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19448), .ZN(
        n19430) );
  INV_X1 U17405 ( .A(n19430), .ZN(n19439) );
  AND2_X1 U17406 ( .A1(n19933), .A2(n19439), .ZN(n14105) );
  NAND2_X1 U17407 ( .A1(n14102), .A2(n14105), .ZN(n14101) );
  OAI211_X1 U17408 ( .C1(n10641), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19860), 
        .B(n19439), .ZN(n14099) );
  AND2_X1 U17409 ( .A1(n14099), .A2(n19936), .ZN(n14100) );
  NAND2_X1 U17410 ( .A1(n14101), .A2(n14100), .ZN(n19443) );
  INV_X1 U17411 ( .A(n14102), .ZN(n14106) );
  OAI21_X1 U17412 ( .B1(n14103), .B2(n19430), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14104) );
  NOR2_X2 U17413 ( .A1(n19865), .A2(n19330), .ZN(n19943) );
  INV_X1 U17414 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20325) );
  INV_X1 U17415 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18421) );
  OAI22_X2 U17416 ( .A1(n20325), .A2(n19427), .B1(n18421), .B2(n19428), .ZN(
        n19944) );
  INV_X1 U17417 ( .A(n19944), .ZN(n14111) );
  AOI22_X2 U17418 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19437), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19436), .ZN(n19947) );
  INV_X1 U17419 ( .A(n19947), .ZN(n19878) );
  NOR2_X2 U17420 ( .A1(n19438), .A2(n9666), .ZN(n19942) );
  AOI22_X1 U17421 ( .A1(n19878), .A2(n19465), .B1(n19430), .B2(n19942), .ZN(
        n14110) );
  OAI21_X1 U17422 ( .B1(n19989), .B2(n14111), .A(n14110), .ZN(n14112) );
  AOI21_X1 U17423 ( .B1(n19442), .B2(n19943), .A(n14112), .ZN(n14113) );
  OAI21_X1 U17424 ( .B1(n19435), .B2(n14114), .A(n14113), .ZN(P2_U3049) );
  NOR2_X2 U17425 ( .A1(n19865), .A2(n19319), .ZN(n19955) );
  NAND2_X1 U17426 ( .A1(n19442), .A2(n19955), .ZN(n14117) );
  INV_X1 U17427 ( .A(n19989), .ZN(n19975) );
  INV_X1 U17428 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20338) );
  INV_X1 U17429 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n18430) );
  OR2_X1 U17430 ( .A1(n19438), .A2(n10356), .ZN(n19889) );
  AOI22_X1 U17431 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19437), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19436), .ZN(n19890) );
  OAI22_X1 U17432 ( .A1(n19889), .A2(n19439), .B1(n19890), .B2(n19473), .ZN(
        n14115) );
  AOI21_X1 U17433 ( .B1(n19975), .B2(n19892), .A(n14115), .ZN(n14116) );
  OAI211_X1 U17434 ( .C1(n19435), .C2(n14118), .A(n14117), .B(n14116), .ZN(
        P2_U3051) );
  AOI21_X1 U17435 ( .B1(n14120), .B2(n14004), .A(n14119), .ZN(n14338) );
  INV_X1 U17436 ( .A(n14338), .ZN(n14138) );
  MUX2_X1 U17437 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n20311), .Z(
        n14677) );
  AOI22_X1 U17438 ( .A1(n16059), .A2(n14677), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n16057), .ZN(n14121) );
  OAI21_X1 U17439 ( .B1(n14138), .B2(n14715), .A(n14121), .ZN(P1_U2896) );
  INV_X1 U17440 ( .A(n14268), .ZN(n14122) );
  AOI21_X1 U17441 ( .B1(n14124), .B2(n14123), .A(n14122), .ZN(n16255) );
  AOI22_X1 U17442 ( .A1(n16255), .A2(n13368), .B1(n14653), .B2(
        P1_EBX_REG_8__SCAN_IN), .ZN(n14125) );
  OAI21_X1 U17443 ( .B1(n14138), .B2(n14640), .A(n14125), .ZN(P1_U2864) );
  INV_X1 U17444 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n14126) );
  INV_X1 U17445 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20147) );
  NAND4_X1 U17446 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n20174)
         );
  NAND2_X1 U17447 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20145) );
  NOR3_X1 U17448 ( .A1(n20147), .A2(n20174), .A3(n20145), .ZN(n14127) );
  AND3_X1 U17449 ( .A1(n20146), .A2(n14126), .A3(n14127), .ZN(n14136) );
  NAND2_X1 U17450 ( .A1(n20173), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n14134) );
  NAND2_X1 U17451 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n14127), .ZN(n20134) );
  NOR2_X1 U17452 ( .A1(n14128), .A2(n20134), .ZN(n14554) );
  NOR2_X1 U17453 ( .A1(n15968), .A2(n14554), .ZN(n14129) );
  NAND2_X1 U17454 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n14129), .ZN(n14131) );
  NAND2_X1 U17455 ( .A1(n14130), .A2(n20144), .ZN(n20187) );
  NAND2_X1 U17456 ( .A1(n14131), .A2(n20187), .ZN(n14132) );
  AOI21_X1 U17457 ( .B1(n20186), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n14132), .ZN(n14133) );
  OAI211_X1 U17458 ( .C1(n20189), .C2(n14336), .A(n14134), .B(n14133), .ZN(
        n14135) );
  AOI211_X1 U17459 ( .C1(n16255), .C2(n20196), .A(n14136), .B(n14135), .ZN(
        n14137) );
  OAI21_X1 U17460 ( .B1(n14138), .B2(n20148), .A(n14137), .ZN(P1_U2832) );
  MUX2_X1 U17461 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n20311), .Z(
        n14660) );
  NAND2_X1 U17462 ( .A1(n14179), .A2(n14660), .ZN(n14184) );
  NAND2_X1 U17463 ( .A1(n14187), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n14139) );
  OAI211_X1 U17464 ( .C1(n14140), .C2(n14193), .A(n14184), .B(n14139), .ZN(
        P1_U2950) );
  INV_X1 U17465 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20208) );
  INV_X1 U17466 ( .A(DATAI_12_), .ZN(n21043) );
  NOR2_X1 U17467 ( .A1(n20312), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14141) );
  AOI21_X1 U17468 ( .B1(n21043), .B2(n20312), .A(n14141), .ZN(n16054) );
  NAND2_X1 U17469 ( .A1(n14179), .A2(n16054), .ZN(n14164) );
  NAND2_X1 U17470 ( .A1(n14187), .A2(P1_LWORD_REG_12__SCAN_IN), .ZN(n14142) );
  OAI211_X1 U17471 ( .C1(n20208), .C2(n14193), .A(n14164), .B(n14142), .ZN(
        P1_U2964) );
  INV_X1 U17472 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20212) );
  MUX2_X1 U17473 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n20311), .Z(
        n14667) );
  NAND2_X1 U17474 ( .A1(n14179), .A2(n14667), .ZN(n14169) );
  NAND2_X1 U17475 ( .A1(n14187), .A2(P1_LWORD_REG_10__SCAN_IN), .ZN(n14143) );
  OAI211_X1 U17476 ( .C1(n20212), .C2(n14193), .A(n14169), .B(n14143), .ZN(
        P1_U2962) );
  INV_X1 U17477 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20214) );
  INV_X1 U17478 ( .A(DATAI_9_), .ZN(n21103) );
  MUX2_X1 U17479 ( .A(n21103), .B(n13522), .S(n20311), .Z(n14672) );
  INV_X1 U17480 ( .A(n14672), .ZN(n14144) );
  NAND2_X1 U17481 ( .A1(n14179), .A2(n14144), .ZN(n14171) );
  NAND2_X1 U17482 ( .A1(n14187), .A2(P1_LWORD_REG_9__SCAN_IN), .ZN(n14145) );
  OAI211_X1 U17483 ( .C1(n20214), .C2(n14193), .A(n14171), .B(n14145), .ZN(
        P1_U2961) );
  INV_X1 U17484 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20210) );
  MUX2_X1 U17485 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n20311), .Z(
        n16058) );
  NAND2_X1 U17486 ( .A1(n14179), .A2(n16058), .ZN(n14166) );
  NAND2_X1 U17487 ( .A1(n14187), .A2(P1_LWORD_REG_11__SCAN_IN), .ZN(n14146) );
  OAI211_X1 U17488 ( .C1(n20210), .C2(n14193), .A(n14166), .B(n14146), .ZN(
        P1_U2963) );
  NAND2_X1 U17489 ( .A1(n14179), .A2(n20376), .ZN(n14175) );
  NAND2_X1 U17490 ( .A1(n14190), .A2(P1_LWORD_REG_7__SCAN_IN), .ZN(n14147) );
  OAI211_X1 U17491 ( .C1(n11892), .C2(n14193), .A(n14175), .B(n14147), .ZN(
        P1_U2959) );
  INV_X1 U17492 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20204) );
  MUX2_X1 U17493 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n20311), .Z(
        n14656) );
  NAND2_X1 U17494 ( .A1(n14179), .A2(n14656), .ZN(n14189) );
  NAND2_X1 U17495 ( .A1(n14187), .A2(P1_LWORD_REG_14__SCAN_IN), .ZN(n14148) );
  OAI211_X1 U17496 ( .C1(n20204), .C2(n14193), .A(n14189), .B(n14148), .ZN(
        P1_U2966) );
  NAND2_X1 U17497 ( .A1(n14179), .A2(n20354), .ZN(n14162) );
  NAND2_X1 U17498 ( .A1(n14190), .A2(P1_LWORD_REG_5__SCAN_IN), .ZN(n14149) );
  OAI211_X1 U17499 ( .C1(n11873), .C2(n14193), .A(n14162), .B(n14149), .ZN(
        P1_U2957) );
  INV_X1 U17500 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14232) );
  INV_X1 U17501 ( .A(n20340), .ZN(n14150) );
  NAND2_X1 U17502 ( .A1(n14179), .A2(n14150), .ZN(n14155) );
  NAND2_X1 U17503 ( .A1(n14190), .A2(P1_UWORD_REG_3__SCAN_IN), .ZN(n14151) );
  OAI211_X1 U17504 ( .C1(n14232), .C2(n14193), .A(n14155), .B(n14151), .ZN(
        P1_U2940) );
  INV_X1 U17505 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14238) );
  INV_X1 U17506 ( .A(n20332), .ZN(n14699) );
  NAND2_X1 U17507 ( .A1(n14179), .A2(n14699), .ZN(n14178) );
  NAND2_X1 U17508 ( .A1(n14190), .A2(P1_UWORD_REG_2__SCAN_IN), .ZN(n14152) );
  OAI211_X1 U17509 ( .C1(n14238), .C2(n14193), .A(n14178), .B(n14152), .ZN(
        P1_U2939) );
  INV_X1 U17510 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20223) );
  NAND2_X1 U17511 ( .A1(n14179), .A2(n20348), .ZN(n14182) );
  NAND2_X1 U17512 ( .A1(n14187), .A2(P1_LWORD_REG_4__SCAN_IN), .ZN(n14153) );
  OAI211_X1 U17513 ( .C1(n20223), .C2(n14193), .A(n14182), .B(n14153), .ZN(
        P1_U2956) );
  NAND2_X1 U17514 ( .A1(n14187), .A2(P1_LWORD_REG_3__SCAN_IN), .ZN(n14154) );
  OAI211_X1 U17515 ( .C1(n20225), .C2(n14193), .A(n14155), .B(n14154), .ZN(
        P1_U2955) );
  INV_X1 U17516 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20216) );
  NAND2_X1 U17517 ( .A1(n14179), .A2(n14677), .ZN(n14173) );
  NAND2_X1 U17518 ( .A1(n14187), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n14156) );
  OAI211_X1 U17519 ( .C1(n20216), .C2(n14193), .A(n14173), .B(n14156), .ZN(
        P1_U2960) );
  INV_X1 U17520 ( .A(n20327), .ZN(n14702) );
  NAND2_X1 U17521 ( .A1(n14179), .A2(n14702), .ZN(n14192) );
  NAND2_X1 U17522 ( .A1(n14187), .A2(P1_LWORD_REG_1__SCAN_IN), .ZN(n14157) );
  OAI211_X1 U17523 ( .C1(n20229), .C2(n14193), .A(n14192), .B(n14157), .ZN(
        P1_U2953) );
  NAND2_X1 U17524 ( .A1(n14179), .A2(n20361), .ZN(n14160) );
  NAND2_X1 U17525 ( .A1(n14190), .A2(P1_LWORD_REG_6__SCAN_IN), .ZN(n14158) );
  OAI211_X1 U17526 ( .C1(n14193), .C2(n20220), .A(n14160), .B(n14158), .ZN(
        P1_U2958) );
  INV_X1 U17527 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14236) );
  NAND2_X1 U17528 ( .A1(n14190), .A2(P1_UWORD_REG_6__SCAN_IN), .ZN(n14159) );
  OAI211_X1 U17529 ( .C1(n14236), .C2(n14193), .A(n14160), .B(n14159), .ZN(
        P1_U2943) );
  INV_X1 U17530 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n14230) );
  NAND2_X1 U17531 ( .A1(n14190), .A2(P1_UWORD_REG_5__SCAN_IN), .ZN(n14161) );
  OAI211_X1 U17532 ( .C1(n14230), .C2(n14193), .A(n14162), .B(n14161), .ZN(
        P1_U2942) );
  INV_X1 U17533 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n14250) );
  NAND2_X1 U17534 ( .A1(n14187), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n14163) );
  OAI211_X1 U17535 ( .C1(n14250), .C2(n14193), .A(n14164), .B(n14163), .ZN(
        P1_U2949) );
  NAND2_X1 U17536 ( .A1(n14187), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n14165) );
  OAI211_X1 U17537 ( .C1(n14167), .C2(n14193), .A(n14166), .B(n14165), .ZN(
        P1_U2948) );
  INV_X1 U17538 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14234) );
  NAND2_X1 U17539 ( .A1(n14190), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n14168) );
  OAI211_X1 U17540 ( .C1(n14234), .C2(n14193), .A(n14169), .B(n14168), .ZN(
        P1_U2947) );
  NAND2_X1 U17541 ( .A1(n14190), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n14170) );
  OAI211_X1 U17542 ( .C1(n14193), .C2(n14671), .A(n14171), .B(n14170), .ZN(
        P1_U2946) );
  INV_X1 U17543 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14240) );
  NAND2_X1 U17544 ( .A1(n14190), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n14172) );
  OAI211_X1 U17545 ( .C1(n14240), .C2(n14193), .A(n14173), .B(n14172), .ZN(
        P1_U2945) );
  NAND2_X1 U17546 ( .A1(n14190), .A2(P1_UWORD_REG_7__SCAN_IN), .ZN(n14174) );
  OAI211_X1 U17547 ( .C1(n14176), .C2(n14193), .A(n14175), .B(n14174), .ZN(
        P1_U2944) );
  NAND2_X1 U17548 ( .A1(n14187), .A2(P1_LWORD_REG_2__SCAN_IN), .ZN(n14177) );
  OAI211_X1 U17549 ( .C1(n20227), .C2(n14193), .A(n14178), .B(n14177), .ZN(
        P1_U2954) );
  INV_X1 U17550 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14247) );
  INV_X1 U17551 ( .A(n20317), .ZN(n14706) );
  NAND2_X1 U17552 ( .A1(n14179), .A2(n14706), .ZN(n14186) );
  NAND2_X1 U17553 ( .A1(n14190), .A2(P1_UWORD_REG_0__SCAN_IN), .ZN(n14180) );
  OAI211_X1 U17554 ( .C1(n14247), .C2(n14193), .A(n14186), .B(n14180), .ZN(
        P1_U2937) );
  INV_X1 U17555 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14245) );
  NAND2_X1 U17556 ( .A1(n14190), .A2(P1_UWORD_REG_4__SCAN_IN), .ZN(n14181) );
  OAI211_X1 U17557 ( .C1(n14245), .C2(n14193), .A(n14182), .B(n14181), .ZN(
        P1_U2941) );
  INV_X1 U17558 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20206) );
  NAND2_X1 U17559 ( .A1(n14187), .A2(P1_LWORD_REG_13__SCAN_IN), .ZN(n14183) );
  OAI211_X1 U17560 ( .C1(n20206), .C2(n14193), .A(n14184), .B(n14183), .ZN(
        P1_U2965) );
  NAND2_X1 U17561 ( .A1(n14187), .A2(P1_LWORD_REG_0__SCAN_IN), .ZN(n14185) );
  OAI211_X1 U17562 ( .C1(n20234), .C2(n14193), .A(n14186), .B(n14185), .ZN(
        P1_U2952) );
  INV_X1 U17563 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n14228) );
  NAND2_X1 U17564 ( .A1(n14187), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n14188) );
  OAI211_X1 U17565 ( .C1(n14228), .C2(n14193), .A(n14189), .B(n14188), .ZN(
        P1_U2951) );
  INV_X1 U17566 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14242) );
  NAND2_X1 U17567 ( .A1(n14190), .A2(P1_UWORD_REG_1__SCAN_IN), .ZN(n14191) );
  OAI211_X1 U17568 ( .C1(n14242), .C2(n14193), .A(n14192), .B(n14191), .ZN(
        P1_U2938) );
  INV_X1 U17569 ( .A(n14194), .ZN(n14196) );
  NOR2_X1 U17570 ( .A1(n14195), .A2(n14909), .ZN(n16541) );
  AOI21_X1 U17571 ( .B1(n14196), .B2(n16541), .A(n16538), .ZN(n14201) );
  NAND2_X1 U17572 ( .A1(n20003), .A2(n19926), .ZN(n14197) );
  NAND3_X1 U17573 ( .A1(n14199), .A2(n14198), .A3(n14197), .ZN(n14200) );
  MUX2_X1 U17574 ( .A(n14201), .B(n14200), .S(n11320), .Z(n14202) );
  NAND2_X1 U17575 ( .A1(n14202), .A2(n16312), .ZN(P2_U3177) );
  XOR2_X1 U17576 ( .A(n14204), .B(n14203), .Z(n19396) );
  INV_X1 U17577 ( .A(n19396), .ZN(n14226) );
  XNOR2_X1 U17578 ( .A(n14205), .B(n14304), .ZN(n14208) );
  NAND2_X1 U17579 ( .A1(n16478), .A2(n14206), .ZN(n14207) );
  XNOR2_X1 U17580 ( .A(n14208), .B(n14207), .ZN(n19401) );
  NAND2_X1 U17581 ( .A1(n14465), .A2(n14209), .ZN(n16535) );
  INV_X1 U17582 ( .A(n16535), .ZN(n15696) );
  NAND2_X1 U17583 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15696), .ZN(
        n14303) );
  OR2_X1 U17584 ( .A1(n16501), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14213) );
  INV_X1 U17585 ( .A(n15575), .ZN(n14212) );
  INV_X1 U17586 ( .A(n14460), .ZN(n14210) );
  AOI21_X1 U17587 ( .B1(n14212), .B2(n14211), .A(n14210), .ZN(n16533) );
  NAND2_X1 U17588 ( .A1(n14213), .A2(n16533), .ZN(n14302) );
  OR2_X1 U17589 ( .A1(n14214), .A2(n9784), .ZN(n14216) );
  INV_X1 U17590 ( .A(n14300), .ZN(n14215) );
  AND2_X1 U17591 ( .A1(n14216), .A2(n14215), .ZN(n19305) );
  INV_X1 U17592 ( .A(n19305), .ZN(n14217) );
  OAI22_X1 U17593 ( .A1(n16522), .A2(n14217), .B1(n19392), .B2(n19214), .ZN(
        n14222) );
  NAND2_X1 U17594 ( .A1(n14219), .A2(n14218), .ZN(n14220) );
  NAND2_X1 U17595 ( .A1(n13772), .A2(n14220), .ZN(n19263) );
  NOR2_X1 U17596 ( .A1(n19263), .A2(n15710), .ZN(n14221) );
  AOI211_X1 U17597 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n14302), .A(
        n14222), .B(n14221), .ZN(n14223) );
  OAI21_X1 U17598 ( .B1(n14303), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n14223), .ZN(n14224) );
  AOI21_X1 U17599 ( .B1(n19401), .B2(n10972), .A(n14224), .ZN(n14225) );
  OAI21_X1 U17600 ( .B1(n14226), .B2(n16490), .A(n14225), .ZN(P2_U3042) );
  AOI22_X1 U17601 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20231), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n20230), .ZN(n14227) );
  OAI21_X1 U17602 ( .B1(n14228), .B2(n14249), .A(n14227), .ZN(P1_U2906) );
  AOI22_X1 U17603 ( .A1(n14243), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20230), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n14229) );
  OAI21_X1 U17604 ( .B1(n14230), .B2(n14249), .A(n14229), .ZN(P1_U2915) );
  AOI22_X1 U17605 ( .A1(n14243), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20230), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n14231) );
  OAI21_X1 U17606 ( .B1(n14232), .B2(n14249), .A(n14231), .ZN(P1_U2917) );
  AOI22_X1 U17607 ( .A1(n14243), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20230), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n14233) );
  OAI21_X1 U17608 ( .B1(n14234), .B2(n14249), .A(n14233), .ZN(P1_U2910) );
  AOI22_X1 U17609 ( .A1(n14243), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20230), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n14235) );
  OAI21_X1 U17610 ( .B1(n14236), .B2(n14249), .A(n14235), .ZN(P1_U2914) );
  AOI22_X1 U17611 ( .A1(n14243), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20230), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n14237) );
  OAI21_X1 U17612 ( .B1(n14238), .B2(n14249), .A(n14237), .ZN(P1_U2918) );
  AOI22_X1 U17613 ( .A1(n14243), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20230), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n14239) );
  OAI21_X1 U17614 ( .B1(n14240), .B2(n14249), .A(n14239), .ZN(P1_U2912) );
  AOI22_X1 U17615 ( .A1(n14243), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20230), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n14241) );
  OAI21_X1 U17616 ( .B1(n14242), .B2(n14249), .A(n14241), .ZN(P1_U2919) );
  AOI22_X1 U17617 ( .A1(n14243), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20230), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n14244) );
  OAI21_X1 U17618 ( .B1(n14245), .B2(n14249), .A(n14244), .ZN(P1_U2916) );
  AOI22_X1 U17619 ( .A1(n20231), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(n20230), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n14246) );
  OAI21_X1 U17620 ( .B1(n14247), .B2(n14249), .A(n14246), .ZN(P1_U2920) );
  AOI22_X1 U17621 ( .A1(n20231), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20230), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n14248) );
  OAI21_X1 U17622 ( .B1(n14250), .B2(n14249), .A(n14248), .ZN(P1_U2908) );
  INV_X1 U17623 ( .A(n14251), .ZN(n14252) );
  NAND2_X1 U17624 ( .A1(n14252), .A2(n15720), .ZN(n14253) );
  AND2_X1 U17625 ( .A1(n15132), .A2(n14253), .ZN(n14254) );
  NAND2_X1 U17626 ( .A1(n13426), .A2(n14254), .ZN(n15727) );
  INV_X1 U17627 ( .A(n19221), .ZN(n19186) );
  MUX2_X1 U17628 ( .A(n19151), .B(n19186), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n14263) );
  INV_X1 U17629 ( .A(n14255), .ZN(n14256) );
  AOI22_X1 U17630 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19199), .B1(n19189), 
        .B2(n14256), .ZN(n14257) );
  OAI21_X1 U17631 ( .B1(n19218), .B2(n14258), .A(n14257), .ZN(n14259) );
  AOI21_X1 U17632 ( .B1(n19209), .B2(n20096), .A(n14259), .ZN(n14260) );
  OAI21_X1 U17633 ( .B1(n10460), .B2(n19129), .A(n14260), .ZN(n14261) );
  AOI21_X1 U17634 ( .B1(n20094), .B2(n15131), .A(n14261), .ZN(n14262) );
  OAI211_X1 U17635 ( .C1(n15727), .C2(n16312), .A(n14263), .B(n14262), .ZN(
        P2_U2854) );
  NAND2_X1 U17636 ( .A1(n14266), .A2(n14265), .ZN(n14267) );
  NAND2_X1 U17637 ( .A1(n14264), .A2(n14267), .ZN(n20132) );
  INV_X1 U17638 ( .A(n14321), .ZN(n14367) );
  AOI21_X1 U17639 ( .B1(n14269), .B2(n14268), .A(n14367), .ZN(n20130) );
  AOI22_X1 U17640 ( .A1(n20130), .A2(n13368), .B1(n14653), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n14270) );
  OAI21_X1 U17641 ( .B1(n20132), .B2(n14655), .A(n14270), .ZN(P1_U2863) );
  OAI222_X1 U17642 ( .A1(n20132), .A2(n14715), .B1(n14672), .B2(n14713), .C1(
        n20214), .C2(n14711), .ZN(P1_U2895) );
  OAI21_X1 U17643 ( .B1(n14272), .B2(n16312), .A(n19151), .ZN(n14287) );
  INV_X1 U17644 ( .A(n15392), .ZN(n14271) );
  NAND3_X1 U17645 ( .A1(n15133), .A2(n14272), .A3(n14271), .ZN(n14285) );
  OR2_X1 U17646 ( .A1(n14274), .A2(n14273), .ZN(n14276) );
  NAND2_X1 U17647 ( .A1(n14276), .A2(n14275), .ZN(n19292) );
  NAND2_X1 U17648 ( .A1(n19221), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14277) );
  OAI21_X1 U17649 ( .B1(n19231), .B2(n19292), .A(n14277), .ZN(n14280) );
  NAND2_X1 U17650 ( .A1(n16517), .A2(n19226), .ZN(n14278) );
  OAI211_X1 U17651 ( .C1(n20021), .C2(n19215), .A(n14278), .B(n19214), .ZN(
        n14279) );
  NOR2_X1 U17652 ( .A1(n14280), .A2(n14279), .ZN(n14284) );
  NAND2_X1 U17653 ( .A1(n14281), .A2(n19189), .ZN(n14283) );
  NAND2_X1 U17654 ( .A1(n19183), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n14282) );
  NAND4_X1 U17655 ( .A1(n14285), .A2(n14284), .A3(n14283), .A4(n14282), .ZN(
        n14286) );
  AOI21_X1 U17656 ( .B1(n15392), .B2(n14287), .A(n14286), .ZN(n14288) );
  INV_X1 U17657 ( .A(n14288), .ZN(P2_U2848) );
  OAI21_X1 U17658 ( .B1(n19167), .B2(n19221), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14295) );
  NAND2_X1 U17659 ( .A1(n19209), .A2(n15712), .ZN(n14291) );
  AOI22_X1 U17660 ( .A1(n19199), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n19189), 
        .B2(n14289), .ZN(n14290) );
  OAI211_X1 U17661 ( .C1(n19129), .C2(n15709), .A(n14291), .B(n14290), .ZN(
        n14293) );
  INV_X1 U17662 ( .A(n15131), .ZN(n15098) );
  NOR2_X1 U17663 ( .A1(n20101), .A2(n15098), .ZN(n14292) );
  AOI211_X1 U17664 ( .C1(P2_EBX_REG_0__SCAN_IN), .C2(n19183), .A(n14293), .B(
        n14292), .ZN(n14294) );
  OAI211_X1 U17665 ( .C1(n14296), .C2(n15103), .A(n14295), .B(n14294), .ZN(
        P2_U2855) );
  XNOR2_X1 U17666 ( .A(n14298), .B(n14297), .ZN(n16466) );
  INV_X1 U17667 ( .A(n14299), .ZN(n19225) );
  XNOR2_X1 U17668 ( .A(n14301), .B(n14300), .ZN(n19303) );
  NAND2_X1 U17669 ( .A1(n14302), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14308) );
  AOI221_X1 U17670 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n14305), .C2(n14304), .A(
        n14303), .ZN(n14306) );
  AOI21_X1 U17671 ( .B1(n19198), .B2(P2_REIP_REG_5__SCAN_IN), .A(n14306), .ZN(
        n14307) );
  OAI211_X1 U17672 ( .C1(n19303), .C2(n16522), .A(n14308), .B(n14307), .ZN(
        n14316) );
  AND2_X1 U17673 ( .A1(n14310), .A2(n14309), .ZN(n14311) );
  OAI22_X1 U17674 ( .A1(n14314), .A2(n14313), .B1(n14312), .B2(n14311), .ZN(
        n16464) );
  NOR2_X1 U17675 ( .A1(n16464), .A2(n16527), .ZN(n14315) );
  AOI211_X1 U17676 ( .C1(n16525), .C2(n19225), .A(n14316), .B(n14315), .ZN(
        n14317) );
  OAI21_X1 U17677 ( .B1(n16490), .B2(n16466), .A(n14317), .ZN(P2_U3041) );
  AOI21_X1 U17678 ( .B1(n11939), .B2(n14264), .A(n14320), .ZN(n14823) );
  INV_X1 U17679 ( .A(n14823), .ZN(n14330) );
  XNOR2_X1 U17680 ( .A(n14321), .B(n14366), .ZN(n16242) );
  NAND2_X1 U17681 ( .A1(n20173), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n14323) );
  AOI21_X1 U17682 ( .B1(n20186), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n20177), .ZN(n14322) );
  OAI211_X1 U17683 ( .C1(n20189), .C2(n14821), .A(n14323), .B(n14322), .ZN(
        n14326) );
  INV_X1 U17684 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n14324) );
  OAI21_X1 U17685 ( .B1(n15968), .B2(n14554), .A(P1_REIP_REG_9__SCAN_IN), .ZN(
        n20136) );
  NAND2_X1 U17686 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n14569) );
  INV_X1 U17687 ( .A(n14554), .ZN(n14568) );
  OAI21_X1 U17688 ( .B1(n14569), .B2(n14568), .A(n15970), .ZN(n16051) );
  AOI21_X1 U17689 ( .B1(n14324), .B2(n20136), .A(n16051), .ZN(n14325) );
  AOI211_X1 U17690 ( .C1(n20196), .C2(n16242), .A(n14326), .B(n14325), .ZN(
        n14327) );
  OAI21_X1 U17691 ( .B1(n14330), .B2(n20148), .A(n14327), .ZN(P1_U2830) );
  AOI22_X1 U17692 ( .A1(n16242), .A2(n13368), .B1(n14653), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n14328) );
  OAI21_X1 U17693 ( .B1(n14330), .B2(n14655), .A(n14328), .ZN(P1_U2862) );
  AOI22_X1 U17694 ( .A1(n16059), .A2(n14667), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n16057), .ZN(n14329) );
  OAI21_X1 U17695 ( .B1(n14330), .B2(n14715), .A(n14329), .ZN(P1_U2894) );
  XNOR2_X1 U17696 ( .A(n14333), .B(n14332), .ZN(n14334) );
  XNOR2_X1 U17697 ( .A(n14331), .B(n14334), .ZN(n16260) );
  INV_X1 U17698 ( .A(n16260), .ZN(n14340) );
  AOI22_X1 U17699 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n20290), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n14335) );
  OAI21_X1 U17700 ( .B1(n20243), .B2(n14336), .A(n14335), .ZN(n14337) );
  AOI21_X1 U17701 ( .B1(n14338), .B2(n20313), .A(n14337), .ZN(n14339) );
  OAI21_X1 U17702 ( .B1(n14340), .B2(n20115), .A(n14339), .ZN(P1_U2991) );
  INV_X1 U17703 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16241) );
  MUX2_X1 U17704 ( .A(n16241), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .S(
        n16086), .Z(n14341) );
  XNOR2_X1 U17705 ( .A(n14342), .B(n14341), .ZN(n16251) );
  NAND2_X1 U17706 ( .A1(n16251), .A2(n20250), .ZN(n14345) );
  OAI22_X1 U17707 ( .A1(n16074), .A2(n11934), .B1(n10234), .B2(n20133), .ZN(
        n14343) );
  AOI21_X1 U17708 ( .B1(n20131), .B2(n20249), .A(n14343), .ZN(n14344) );
  OAI211_X1 U17709 ( .C1(n20254), .C2(n20132), .A(n14345), .B(n14344), .ZN(
        P1_U2990) );
  OAI21_X1 U17710 ( .B1(n14347), .B2(n14350), .A(n14349), .ZN(n15187) );
  OR2_X1 U17711 ( .A1(n14353), .A2(n14352), .ZN(n14354) );
  NAND2_X1 U17712 ( .A1(n14351), .A2(n14354), .ZN(n19156) );
  INV_X1 U17713 ( .A(n19156), .ZN(n15574) );
  OAI22_X1 U17714 ( .A1(n15247), .A2(n19330), .B1(n19293), .B2(n14355), .ZN(
        n14359) );
  INV_X1 U17715 ( .A(n19266), .ZN(n15250) );
  INV_X1 U17716 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n14357) );
  INV_X1 U17717 ( .A(n19265), .ZN(n15248) );
  INV_X1 U17718 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n14356) );
  OAI22_X1 U17719 ( .A1(n15250), .A2(n14357), .B1(n15248), .B2(n14356), .ZN(
        n14358) );
  AOI211_X1 U17720 ( .C1(n19321), .C2(n15574), .A(n14359), .B(n14358), .ZN(
        n14360) );
  OAI21_X1 U17721 ( .B1(n15187), .B2(n19325), .A(n14360), .ZN(P2_U2902) );
  OR2_X1 U17722 ( .A1(n14320), .A2(n14362), .ZN(n14363) );
  AND2_X1 U17723 ( .A1(n14361), .A2(n14363), .ZN(n14381) );
  INV_X1 U17724 ( .A(n14380), .ZN(n14364) );
  XNOR2_X1 U17725 ( .A(n14381), .B(n14364), .ZN(n16115) );
  INV_X1 U17726 ( .A(n16115), .ZN(n16061) );
  AOI21_X1 U17727 ( .B1(n14367), .B2(n14366), .A(n14365), .ZN(n14368) );
  OR2_X1 U17728 ( .A1(n14368), .A2(n14404), .ZN(n16046) );
  OAI22_X1 U17729 ( .A1(n16046), .A2(n14643), .B1(n14369), .B2(n14633), .ZN(
        n14370) );
  INV_X1 U17730 ( .A(n14370), .ZN(n14371) );
  OAI21_X1 U17731 ( .B1(n16061), .B2(n14655), .A(n14371), .ZN(P1_U2861) );
  NAND2_X1 U17732 ( .A1(n14373), .A2(n14374), .ZN(n14375) );
  AND2_X1 U17733 ( .A1(n14644), .A2(n14375), .ZN(n16036) );
  INV_X1 U17734 ( .A(n16036), .ZN(n14378) );
  AOI22_X1 U17735 ( .A1(n16059), .A2(n14656), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n16057), .ZN(n14376) );
  OAI21_X1 U17736 ( .B1(n14378), .B2(n14715), .A(n14376), .ZN(P1_U2890) );
  XNOR2_X1 U17737 ( .A(n14646), .B(n14648), .ZN(n16204) );
  AOI22_X1 U17738 ( .A1(n16204), .A2(n13368), .B1(n14653), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n14377) );
  OAI21_X1 U17739 ( .B1(n14378), .B2(n14640), .A(n14377), .ZN(P1_U2858) );
  INV_X1 U17740 ( .A(n14361), .ZN(n14379) );
  AOI21_X1 U17741 ( .B1(n14381), .B2(n14380), .A(n14379), .ZN(n14401) );
  INV_X1 U17742 ( .A(n14382), .ZN(n14400) );
  NOR2_X1 U17743 ( .A1(n14401), .A2(n14400), .ZN(n14399) );
  OAI21_X1 U17744 ( .B1(n14399), .B2(n14383), .A(n14373), .ZN(n14814) );
  NAND2_X1 U17745 ( .A1(n14404), .A2(n14402), .ZN(n14386) );
  INV_X1 U17746 ( .A(n14384), .ZN(n14385) );
  NAND2_X1 U17747 ( .A1(n14386), .A2(n14385), .ZN(n14387) );
  NAND2_X1 U17748 ( .A1(n14387), .A2(n14646), .ZN(n16219) );
  OAI22_X1 U17749 ( .A1(n16219), .A2(n14643), .B1(n14392), .B2(n14633), .ZN(
        n14388) );
  INV_X1 U17750 ( .A(n14388), .ZN(n14389) );
  OAI21_X1 U17751 ( .B1(n14814), .B2(n14655), .A(n14389), .ZN(P1_U2859) );
  NAND2_X1 U17752 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14391) );
  INV_X1 U17753 ( .A(n14391), .ZN(n14390) );
  OAI21_X1 U17754 ( .B1(n14390), .B2(n15968), .A(n16051), .ZN(n16042) );
  NOR3_X1 U17755 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n14391), .A3(n16053), 
        .ZN(n14396) );
  OAI22_X1 U17756 ( .A1(n16219), .A2(n20162), .B1(n14392), .B2(n20190), .ZN(
        n14393) );
  AOI21_X1 U17757 ( .B1(n14811), .B2(n20171), .A(n14393), .ZN(n14394) );
  OAI211_X1 U17758 ( .C1(n20141), .C2(n14809), .A(n14394), .B(n20187), .ZN(
        n14395) );
  AOI211_X1 U17759 ( .C1(P1_REIP_REG_13__SCAN_IN), .C2(n16042), .A(n14396), 
        .B(n14395), .ZN(n14397) );
  OAI21_X1 U17760 ( .B1(n14814), .B2(n20148), .A(n14397), .ZN(P1_U2827) );
  AOI22_X1 U17761 ( .A1(n16059), .A2(n14660), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n16057), .ZN(n14398) );
  OAI21_X1 U17762 ( .B1(n14814), .B2(n14715), .A(n14398), .ZN(P1_U2891) );
  AOI21_X1 U17763 ( .B1(n14401), .B2(n14400), .A(n14399), .ZN(n16106) );
  INV_X1 U17764 ( .A(n16106), .ZN(n16056) );
  INV_X1 U17765 ( .A(n14402), .ZN(n14403) );
  XNOR2_X1 U17766 ( .A(n14404), .B(n14403), .ZN(n16040) );
  INV_X1 U17767 ( .A(n16040), .ZN(n16232) );
  INV_X1 U17768 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14405) );
  OAI222_X1 U17769 ( .A1(n16056), .A2(n14655), .B1(n14643), .B2(n16232), .C1(
        n14633), .C2(n14405), .ZN(P1_U2860) );
  INV_X1 U17770 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n14412) );
  INV_X1 U17771 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n16943) );
  INV_X1 U17772 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n16960) );
  INV_X1 U17773 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17397) );
  INV_X1 U17774 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17026) );
  NOR4_X1 U17775 ( .A1(n18449), .A2(n18434), .A3(n14409), .A4(n14408), .ZN(
        n14410) );
  NAND4_X1 U17776 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .A4(P3_EBX_REG_2__SCAN_IN), .ZN(n15820) );
  NAND3_X1 U17777 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(n17408), .ZN(n17373) );
  NAND2_X1 U17778 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17371), .ZN(n17370) );
  NAND2_X1 U17779 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n17351), .ZN(n17333) );
  NOR2_X1 U17780 ( .A1(n16943), .A2(n17333), .ZN(n17317) );
  NAND2_X1 U17781 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17317), .ZN(n15836) );
  AOI21_X1 U17782 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17317), .A(
        P3_EBX_REG_14__SCAN_IN), .ZN(n14413) );
  NOR2_X1 U17783 ( .A1(n17297), .A2(n14413), .ZN(n14426) );
  AOI22_X1 U17784 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14425) );
  AOI22_X1 U17785 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14424) );
  AOI22_X1 U17786 ( .A1(n13039), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17392), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14423) );
  OAI22_X1 U17787 ( .A1(n15784), .A2(n17107), .B1(n17380), .B2(n17179), .ZN(
        n14421) );
  AOI22_X1 U17788 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14419) );
  AOI22_X1 U17789 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17381), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14418) );
  AOI22_X1 U17790 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14417) );
  NAND2_X1 U17791 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n14416) );
  NAND4_X1 U17792 ( .A1(n14419), .A2(n14418), .A3(n14417), .A4(n14416), .ZN(
        n14420) );
  AOI211_X1 U17793 ( .C1(n17320), .C2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        n14421), .B(n14420), .ZN(n14422) );
  NAND4_X1 U17794 ( .A1(n14425), .A2(n14424), .A3(n14423), .A4(n14422), .ZN(
        n17531) );
  MUX2_X1 U17795 ( .A(n14426), .B(n17531), .S(n17432), .Z(P3_U2689) );
  AOI22_X1 U17796 ( .A1(n14705), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n16057), .ZN(n14428) );
  AOI22_X1 U17797 ( .A1(n14708), .A2(DATAI_28_), .B1(n14707), .B2(n16054), 
        .ZN(n14427) );
  OAI211_X1 U17798 ( .C1(n14442), .C2(n14715), .A(n14428), .B(n14427), .ZN(
        P1_U2876) );
  INV_X1 U17799 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14438) );
  INV_X1 U17800 ( .A(n14440), .ZN(n14429) );
  OAI222_X1 U17801 ( .A1(n14438), .A2(n14642), .B1(n14643), .B2(n14429), .C1(
        n14442), .C2(n14640), .ZN(P1_U2844) );
  INV_X1 U17802 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20919) );
  NAND3_X1 U17803 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .A3(P1_REIP_REG_11__SCAN_IN), .ZN(n16033) );
  NOR2_X1 U17804 ( .A1(n20919), .A2(n16033), .ZN(n14570) );
  NAND4_X1 U17805 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n14570), .A3(
        P1_REIP_REG_16__SCAN_IN), .A4(P1_REIP_REG_15__SCAN_IN), .ZN(n15967) );
  NAND3_X1 U17806 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .A3(P1_REIP_REG_18__SCAN_IN), .ZN(n15971) );
  INV_X1 U17807 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14551) );
  NOR4_X1 U17808 ( .A1(n15967), .A2(n15971), .A3(n14551), .A4(n14569), .ZN(
        n14430) );
  NAND3_X1 U17809 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .A3(n14430), .ZN(n14552) );
  NOR2_X1 U17810 ( .A1(n20134), .A2(n14552), .ZN(n15958) );
  NAND2_X1 U17811 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n15958), .ZN(n14540) );
  NAND2_X1 U17812 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14431) );
  NOR2_X1 U17813 ( .A1(n14540), .A2(n14431), .ZN(n14528) );
  NAND2_X1 U17814 ( .A1(n14528), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14432) );
  NOR2_X1 U17815 ( .A1(n20175), .A2(n14432), .ZN(n14513) );
  NAND2_X1 U17816 ( .A1(n20144), .A2(n14528), .ZN(n14525) );
  NAND2_X1 U17817 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n14433) );
  OAI21_X1 U17818 ( .B1(n14525), .B2(n14433), .A(n15970), .ZN(n14516) );
  INV_X1 U17819 ( .A(n14516), .ZN(n14434) );
  OAI21_X1 U17820 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(n14513), .A(n14434), 
        .ZN(n14437) );
  AOI22_X1 U17821 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n20186), .B1(
        n20171), .B2(n14435), .ZN(n14436) );
  OAI211_X1 U17822 ( .C1(n20190), .C2(n14438), .A(n14437), .B(n14436), .ZN(
        n14439) );
  AOI21_X1 U17823 ( .B1(n14440), .B2(n20196), .A(n14439), .ZN(n14441) );
  OAI21_X1 U17824 ( .B1(n14442), .B2(n20148), .A(n14441), .ZN(P1_U2812) );
  MUX2_X1 U17825 ( .A(n15408), .B(n14443), .S(n19259), .Z(n14444) );
  OAI21_X1 U17826 ( .B1(n14445), .B2(n19254), .A(n14444), .ZN(P2_U2857) );
  NAND2_X1 U17827 ( .A1(n14446), .A2(n19308), .ZN(n14456) );
  AND2_X1 U17828 ( .A1(n14448), .A2(n14447), .ZN(n14450) );
  INV_X1 U17829 ( .A(n16317), .ZN(n14453) );
  OAI22_X1 U17830 ( .A1(n15247), .A2(n19278), .B1(n19293), .B2(n14451), .ZN(
        n14452) );
  AOI21_X1 U17831 ( .B1(n19321), .B2(n14453), .A(n14452), .ZN(n14455) );
  AOI22_X1 U17832 ( .A1(n19266), .A2(BUF2_REG_29__SCAN_IN), .B1(n19265), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n14454) );
  OAI211_X1 U17833 ( .C1(n13238), .C2(n14456), .A(n14455), .B(n14454), .ZN(
        P2_U2890) );
  NOR2_X1 U17834 ( .A1(n16490), .A2(n14457), .ZN(n14464) );
  NOR3_X1 U17835 ( .A1(n15581), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A3(
        n14459), .ZN(n14463) );
  AOI221_X1 U17836 ( .B1(n15575), .B2(n14460), .C1(n14459), .C2(n14460), .A(
        n14458), .ZN(n14462) );
  NOR4_X1 U17837 ( .A1(n14464), .A2(n14463), .A3(n14462), .A4(n14461), .ZN(
        n14469) );
  OAI22_X1 U17838 ( .A1(n19298), .A2(n16522), .B1(n15575), .B2(n14465), .ZN(
        n14466) );
  AOI21_X1 U17839 ( .B1(n10972), .B2(n14467), .A(n14466), .ZN(n14468) );
  OAI211_X1 U17840 ( .C1(n15129), .C2(n15710), .A(n14469), .B(n14468), .ZN(
        P2_U3044) );
  MUX2_X1 U17841 ( .A(n14471), .B(n14470), .S(n14477), .Z(n14476) );
  INV_X1 U17842 ( .A(n14472), .ZN(n14474) );
  NAND2_X1 U17843 ( .A1(n14474), .A2(n14473), .ZN(n14475) );
  OAI211_X1 U17844 ( .C1(n14478), .C2(n14477), .A(n14476), .B(n14475), .ZN(
        n14480) );
  AND2_X1 U17845 ( .A1(n14480), .A2(n14479), .ZN(n15896) );
  NAND3_X1 U17846 ( .A1(n14485), .A2(n11526), .A3(n15925), .ZN(n14481) );
  NAND2_X1 U17847 ( .A1(n14481), .A2(n20892), .ZN(n20967) );
  NAND2_X1 U17848 ( .A1(n14482), .A2(n20967), .ZN(n15895) );
  AND2_X1 U17849 ( .A1(n15895), .A2(n14483), .ZN(n20116) );
  MUX2_X1 U17850 ( .A(P1_MORE_REG_SCAN_IN), .B(n15896), .S(n20116), .Z(
        P1_U3484) );
  MUX2_X1 U17851 ( .A(n14484), .B(n12780), .S(n14510), .Z(n14488) );
  AOI22_X1 U17852 ( .A1(n14486), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n14485), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14487) );
  NAND2_X1 U17853 ( .A1(n14489), .A2(n20165), .ZN(n14495) );
  INV_X1 U17854 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21046) );
  OAI21_X1 U17855 ( .B1(n21046), .B2(n21174), .A(n20146), .ZN(n14490) );
  NAND2_X1 U17856 ( .A1(n14516), .A2(n14490), .ZN(n14498) );
  INV_X1 U17857 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14580) );
  INV_X1 U17858 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14491) );
  OAI22_X1 U17859 ( .A1(n20190), .A2(n14580), .B1(n14491), .B2(n20141), .ZN(
        n14493) );
  NAND3_X1 U17860 ( .A1(n14513), .A2(P1_REIP_REG_29__SCAN_IN), .A3(
        P1_REIP_REG_28__SCAN_IN), .ZN(n14497) );
  NOR3_X1 U17861 ( .A1(n14497), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n21174), 
        .ZN(n14492) );
  AOI211_X1 U17862 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14498), .A(n14493), 
        .B(n14492), .ZN(n14494) );
  OAI211_X1 U17863 ( .C1(n14826), .C2(n20162), .A(n14495), .B(n14494), .ZN(
        P1_U2809) );
  INV_X1 U17864 ( .A(n14497), .ZN(n14499) );
  OAI21_X1 U17865 ( .B1(n14499), .B2(P1_REIP_REG_30__SCAN_IN), .A(n14498), 
        .ZN(n14502) );
  AOI22_X1 U17866 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n20186), .B1(
        n20171), .B2(n14500), .ZN(n14501) );
  OAI211_X1 U17867 ( .C1(n20190), .C2(n14503), .A(n14502), .B(n14501), .ZN(
        n14504) );
  AOI21_X1 U17868 ( .B1(n10231), .B2(n20196), .A(n14504), .ZN(n14505) );
  OAI21_X1 U17869 ( .B1(n14659), .B2(n20148), .A(n14505), .ZN(P1_U2810) );
  AOI21_X1 U17870 ( .B1(n14507), .B2(n13308), .A(n14506), .ZN(n14723) );
  INV_X1 U17871 ( .A(n14723), .ZN(n14663) );
  NAND2_X1 U17872 ( .A1(n13360), .A2(n14508), .ZN(n14509) );
  INV_X1 U17873 ( .A(n14719), .ZN(n14511) );
  OAI22_X1 U17874 ( .A1(n14721), .A2(n20141), .B1(n20189), .B2(n14511), .ZN(
        n14512) );
  AOI21_X1 U17875 ( .B1(n20173), .B2(P1_EBX_REG_29__SCAN_IN), .A(n14512), .ZN(
        n14515) );
  NAND3_X1 U17876 ( .A1(n14513), .A2(P1_REIP_REG_28__SCAN_IN), .A3(n21046), 
        .ZN(n14514) );
  OAI211_X1 U17877 ( .C1(n14516), .C2(n21046), .A(n14515), .B(n14514), .ZN(
        n14517) );
  AOI21_X1 U17878 ( .B1(n14844), .B2(n20196), .A(n14517), .ZN(n14518) );
  OAI21_X1 U17879 ( .B1(n14663), .B2(n20148), .A(n14518), .ZN(P1_U2811) );
  INV_X1 U17880 ( .A(n14519), .ZN(n14520) );
  AOI21_X1 U17881 ( .B1(n14521), .B2(n14520), .A(n13306), .ZN(n14733) );
  INV_X1 U17882 ( .A(n14733), .ZN(n14666) );
  NOR2_X1 U17883 ( .A1(n14536), .A2(n14522), .ZN(n14523) );
  OR2_X1 U17884 ( .A1(n14524), .A2(n14523), .ZN(n14854) );
  INV_X1 U17885 ( .A(n14854), .ZN(n14532) );
  NAND2_X1 U17886 ( .A1(n15970), .A2(n14525), .ZN(n14541) );
  INV_X1 U17887 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21053) );
  OAI22_X1 U17888 ( .A1(n14526), .A2(n20141), .B1(n20189), .B2(n14731), .ZN(
        n14527) );
  AOI21_X1 U17889 ( .B1(n20173), .B2(P1_EBX_REG_27__SCAN_IN), .A(n14527), .ZN(
        n14530) );
  NAND3_X1 U17890 ( .A1(n20146), .A2(n14528), .A3(n21053), .ZN(n14529) );
  OAI211_X1 U17891 ( .C1(n14541), .C2(n21053), .A(n14530), .B(n14529), .ZN(
        n14531) );
  AOI21_X1 U17892 ( .B1(n14532), .B2(n20196), .A(n14531), .ZN(n14533) );
  OAI21_X1 U17893 ( .B1(n14666), .B2(n20148), .A(n14533), .ZN(P1_U2813) );
  NOR2_X1 U17894 ( .A1(n14589), .A2(n14534), .ZN(n14535) );
  OR2_X1 U17895 ( .A1(n14536), .A2(n14535), .ZN(n14867) );
  AOI21_X1 U17896 ( .B1(n14538), .B2(n14537), .A(n14519), .ZN(n14744) );
  NAND2_X1 U17897 ( .A1(n14744), .A2(n20165), .ZN(n14547) );
  INV_X1 U17898 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14742) );
  INV_X1 U17899 ( .A(n14740), .ZN(n14539) );
  OAI22_X1 U17900 ( .A1(n14742), .A2(n20141), .B1(n20189), .B2(n14539), .ZN(
        n14545) );
  INV_X1 U17901 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n14543) );
  INV_X1 U17902 ( .A(n14540), .ZN(n15945) );
  NAND3_X1 U17903 ( .A1(n20146), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n15945), 
        .ZN(n14542) );
  AOI21_X1 U17904 ( .B1(n14543), .B2(n14542), .A(n14541), .ZN(n14544) );
  AOI211_X1 U17905 ( .C1(n20173), .C2(P1_EBX_REG_26__SCAN_IN), .A(n14545), .B(
        n14544), .ZN(n14546) );
  OAI211_X1 U17906 ( .C1(n20162), .C2(n14867), .A(n14547), .B(n14546), .ZN(
        P1_U2814) );
  AOI21_X1 U17907 ( .B1(n14550), .B2(n14548), .A(n14549), .ZN(n16064) );
  INV_X1 U17908 ( .A(n16064), .ZN(n14682) );
  INV_X1 U17909 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n16154) );
  INV_X1 U17910 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21073) );
  NOR2_X1 U17911 ( .A1(n15967), .A2(n16053), .ZN(n16013) );
  NAND3_X1 U17912 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .A3(n16013), .ZN(n15999) );
  NOR2_X1 U17913 ( .A1(n21073), .A2(n15999), .ZN(n15990) );
  NAND2_X1 U17914 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n15990), .ZN(n15975) );
  OAI21_X1 U17915 ( .B1(n16154), .B2(n15975), .A(n14551), .ZN(n14562) );
  INV_X1 U17916 ( .A(n14552), .ZN(n14553) );
  AOI21_X1 U17917 ( .B1(n14554), .B2(n14553), .A(n15968), .ZN(n15957) );
  INV_X1 U17918 ( .A(n14596), .ZN(n14555) );
  AOI21_X1 U17919 ( .B1(n14556), .B2(n14603), .A(n14555), .ZN(n16139) );
  INV_X1 U17920 ( .A(n16139), .ZN(n14560) );
  INV_X1 U17921 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14557) );
  OAI22_X1 U17922 ( .A1(n14557), .A2(n20141), .B1(n20189), .B2(n16067), .ZN(
        n14558) );
  AOI21_X1 U17923 ( .B1(n20173), .B2(P1_EBX_REG_23__SCAN_IN), .A(n14558), .ZN(
        n14559) );
  OAI21_X1 U17924 ( .B1(n14560), .B2(n20162), .A(n14559), .ZN(n14561) );
  AOI21_X1 U17925 ( .B1(n14562), .B2(n15957), .A(n14561), .ZN(n14563) );
  OAI21_X1 U17926 ( .B1(n14682), .B2(n20148), .A(n14563), .ZN(P1_U2817) );
  AOI21_X1 U17927 ( .B1(n14566), .B2(n14564), .A(n14565), .ZN(n14567) );
  INV_X1 U17928 ( .A(n14567), .ZN(n14790) );
  NOR2_X1 U17929 ( .A1(n14569), .A2(n14568), .ZN(n14571) );
  AOI21_X1 U17930 ( .B1(n14571), .B2(n14570), .A(n15968), .ZN(n16035) );
  NOR3_X1 U17931 ( .A1(n20919), .A2(n16033), .A3(n16053), .ZN(n16026) );
  INV_X1 U17932 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20923) );
  INV_X1 U17933 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n16195) );
  XOR2_X1 U17934 ( .A(n20923), .B(n16195), .Z(n14572) );
  AOI22_X1 U17935 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n16035), .B1(n16026), 
        .B2(n14572), .ZN(n14579) );
  AND2_X1 U17936 ( .A1(n14650), .A2(n14573), .ZN(n14574) );
  OR2_X1 U17937 ( .A1(n14574), .A2(n14635), .ZN(n16189) );
  INV_X1 U17938 ( .A(n14575), .ZN(n14788) );
  AOI22_X1 U17939 ( .A1(P1_EBX_REG_16__SCAN_IN), .A2(n20173), .B1(n14788), 
        .B2(n20171), .ZN(n14576) );
  OAI21_X1 U17940 ( .B1(n20162), .B2(n16189), .A(n14576), .ZN(n14577) );
  AOI211_X1 U17941 ( .C1(n20186), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n14577), .B(n20177), .ZN(n14578) );
  OAI211_X1 U17942 ( .C1(n14790), .C2(n20148), .A(n14579), .B(n14578), .ZN(
        P1_U2824) );
  OAI22_X1 U17943 ( .A1(n14826), .A2(n14643), .B1(n14580), .B2(n14642), .ZN(
        P1_U2841) );
  AOI22_X1 U17944 ( .A1(n14844), .A2(n13368), .B1(n14653), .B2(
        P1_EBX_REG_29__SCAN_IN), .ZN(n14581) );
  OAI21_X1 U17945 ( .B1(n14663), .B2(n14655), .A(n14581), .ZN(P1_U2843) );
  OAI222_X1 U17946 ( .A1(n14582), .A2(n14642), .B1(n14643), .B2(n14854), .C1(
        n14666), .C2(n14640), .ZN(P1_U2845) );
  INV_X1 U17947 ( .A(n14744), .ZN(n14670) );
  INV_X1 U17948 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14583) );
  OAI222_X1 U17949 ( .A1(n14640), .A2(n14670), .B1(n14633), .B2(n14583), .C1(
        n14867), .C2(n14643), .ZN(P1_U2846) );
  OR2_X1 U17950 ( .A1(n14584), .A2(n14585), .ZN(n14586) );
  AND2_X1 U17951 ( .A1(n14537), .A2(n14586), .ZN(n15953) );
  INV_X1 U17952 ( .A(n15953), .ZN(n14676) );
  AND2_X1 U17953 ( .A1(n14598), .A2(n14587), .ZN(n14588) );
  NOR2_X1 U17954 ( .A1(n14589), .A2(n14588), .ZN(n15952) );
  NOR2_X1 U17955 ( .A1(n14633), .A2(n14590), .ZN(n14591) );
  AOI21_X1 U17956 ( .B1(n15952), .B2(n13368), .A(n14591), .ZN(n14592) );
  OAI21_X1 U17957 ( .B1(n14676), .B2(n14655), .A(n14592), .ZN(P1_U2847) );
  INV_X1 U17958 ( .A(n14584), .ZN(n14593) );
  OAI21_X1 U17959 ( .B1(n14594), .B2(n14549), .A(n14593), .ZN(n15960) );
  INV_X1 U17960 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14599) );
  NAND2_X1 U17961 ( .A1(n14596), .A2(n14595), .ZN(n14597) );
  NAND2_X1 U17962 ( .A1(n14598), .A2(n14597), .ZN(n15959) );
  OAI222_X1 U17963 ( .A1(n14655), .A2(n15960), .B1(n14633), .B2(n14599), .C1(
        n15959), .C2(n14643), .ZN(P1_U2848) );
  AOI22_X1 U17964 ( .A1(n16139), .A2(n13368), .B1(n14653), .B2(
        P1_EBX_REG_23__SCAN_IN), .ZN(n14600) );
  OAI21_X1 U17965 ( .B1(n14682), .B2(n14655), .A(n14600), .ZN(P1_U2849) );
  OR2_X1 U17966 ( .A1(n14611), .A2(n14601), .ZN(n14602) );
  NAND2_X1 U17967 ( .A1(n14603), .A2(n14602), .ZN(n16146) );
  INV_X1 U17968 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14605) );
  OAI21_X1 U17969 ( .B1(n10152), .B2(n9781), .A(n14548), .ZN(n15976) );
  OAI222_X1 U17970 ( .A1(n16146), .A2(n14643), .B1(n14633), .B2(n14605), .C1(
        n14640), .C2(n15976), .ZN(P1_U2850) );
  OR2_X1 U17971 ( .A1(n14606), .A2(n14607), .ZN(n14608) );
  AND2_X1 U17972 ( .A1(n14604), .A2(n14608), .ZN(n15987) );
  INV_X1 U17973 ( .A(n15987), .ZN(n14688) );
  NOR2_X1 U17974 ( .A1(n14615), .A2(n14609), .ZN(n14610) );
  OR2_X1 U17975 ( .A1(n14611), .A2(n14610), .ZN(n15988) );
  OAI22_X1 U17976 ( .A1(n15988), .A2(n14643), .B1(n15984), .B2(n14642), .ZN(
        n14612) );
  INV_X1 U17977 ( .A(n14612), .ZN(n14613) );
  OAI21_X1 U17978 ( .B1(n14688), .B2(n14655), .A(n14613), .ZN(P1_U2851) );
  AND2_X1 U17979 ( .A1(n14624), .A2(n14614), .ZN(n14616) );
  OR2_X1 U17980 ( .A1(n14616), .A2(n14615), .ZN(n15995) );
  INV_X1 U17981 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15994) );
  INV_X1 U17982 ( .A(n14606), .ZN(n14618) );
  OAI21_X1 U17983 ( .B1(n14619), .B2(n14617), .A(n14618), .ZN(n16069) );
  OAI222_X1 U17984 ( .A1(n15995), .A2(n14643), .B1(n14633), .B2(n15994), .C1(
        n14640), .C2(n16069), .ZN(P1_U2852) );
  AND2_X1 U17985 ( .A1(n9730), .A2(n14620), .ZN(n14621) );
  NOR2_X1 U17986 ( .A1(n14617), .A2(n14621), .ZN(n16078) );
  INV_X1 U17987 ( .A(n16078), .ZN(n14698) );
  NAND2_X1 U17988 ( .A1(n14628), .A2(n14622), .ZN(n14623) );
  AND2_X1 U17989 ( .A1(n14624), .A2(n14623), .ZN(n16159) );
  AOI22_X1 U17990 ( .A1(n16159), .A2(n13368), .B1(n14653), .B2(
        P1_EBX_REG_19__SCAN_IN), .ZN(n14625) );
  OAI21_X1 U17991 ( .B1(n14698), .B2(n14655), .A(n14625), .ZN(P1_U2853) );
  OR2_X1 U17992 ( .A1(n14637), .A2(n14626), .ZN(n14627) );
  NAND2_X1 U17993 ( .A1(n14628), .A2(n14627), .ZN(n16179) );
  INV_X1 U17994 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14632) );
  NAND2_X1 U17995 ( .A1(n14629), .A2(n14630), .ZN(n14631) );
  NAND2_X1 U17996 ( .A1(n9730), .A2(n14631), .ZN(n16014) );
  OAI222_X1 U17997 ( .A1(n16179), .A2(n14643), .B1(n14633), .B2(n14632), .C1(
        n14640), .C2(n16014), .ZN(P1_U2854) );
  NOR2_X1 U17998 ( .A1(n14635), .A2(n14634), .ZN(n14636) );
  OR2_X1 U17999 ( .A1(n14637), .A2(n14636), .ZN(n16019) );
  INV_X1 U18000 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14639) );
  OAI21_X1 U18001 ( .B1(n14565), .B2(n14638), .A(n14629), .ZN(n16018) );
  OAI222_X1 U18002 ( .A1(n16019), .A2(n14643), .B1(n14639), .B2(n14642), .C1(
        n16018), .C2(n14640), .ZN(P1_U2855) );
  INV_X1 U18003 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14641) );
  OAI222_X1 U18004 ( .A1(n16189), .A2(n14643), .B1(n14642), .B2(n14641), .C1(
        n14640), .C2(n14790), .ZN(P1_U2856) );
  AOI21_X1 U18005 ( .B1(n14645), .B2(n14644), .A(n10162), .ZN(n16099) );
  INV_X1 U18006 ( .A(n16099), .ZN(n14716) );
  INV_X1 U18007 ( .A(n14646), .ZN(n14649) );
  AOI21_X1 U18008 ( .B1(n14649), .B2(n14648), .A(n14647), .ZN(n14652) );
  INV_X1 U18009 ( .A(n14650), .ZN(n14651) );
  NOR2_X1 U18010 ( .A1(n14652), .A2(n14651), .ZN(n16200) );
  AOI22_X1 U18011 ( .A1(n16200), .A2(n13368), .B1(n14653), .B2(
        P1_EBX_REG_15__SCAN_IN), .ZN(n14654) );
  OAI21_X1 U18012 ( .B1(n14716), .B2(n14655), .A(n14654), .ZN(P1_U2857) );
  AOI22_X1 U18013 ( .A1(n14705), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n16057), .ZN(n14658) );
  AOI22_X1 U18014 ( .A1(n14708), .A2(DATAI_30_), .B1(n14707), .B2(n14656), 
        .ZN(n14657) );
  OAI211_X1 U18015 ( .C1(n14659), .C2(n14715), .A(n14658), .B(n14657), .ZN(
        P1_U2874) );
  AOI22_X1 U18016 ( .A1(n14705), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n16057), .ZN(n14662) );
  AOI22_X1 U18017 ( .A1(n14708), .A2(DATAI_29_), .B1(n14707), .B2(n14660), 
        .ZN(n14661) );
  OAI211_X1 U18018 ( .C1(n14663), .C2(n14715), .A(n14662), .B(n14661), .ZN(
        P1_U2875) );
  AOI22_X1 U18019 ( .A1(n14705), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n16057), .ZN(n14665) );
  AOI22_X1 U18020 ( .A1(n14708), .A2(DATAI_27_), .B1(n14707), .B2(n16058), 
        .ZN(n14664) );
  OAI211_X1 U18021 ( .C1(n14666), .C2(n14715), .A(n14665), .B(n14664), .ZN(
        P1_U2877) );
  AOI22_X1 U18022 ( .A1(n14705), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n16057), .ZN(n14669) );
  AOI22_X1 U18023 ( .A1(n14708), .A2(DATAI_26_), .B1(n14707), .B2(n14667), 
        .ZN(n14668) );
  OAI211_X1 U18024 ( .C1(n14670), .C2(n14715), .A(n14669), .B(n14668), .ZN(
        P1_U2878) );
  OAI22_X1 U18025 ( .A1(n14691), .A2(n20325), .B1(n14671), .B2(n14711), .ZN(
        n14674) );
  INV_X1 U18026 ( .A(n14707), .ZN(n14692) );
  NOR2_X1 U18027 ( .A1(n14692), .A2(n14672), .ZN(n14673) );
  AOI211_X1 U18028 ( .C1(n14708), .C2(DATAI_25_), .A(n14674), .B(n14673), .ZN(
        n14675) );
  OAI21_X1 U18029 ( .B1(n14676), .B2(n14715), .A(n14675), .ZN(P1_U2879) );
  AOI22_X1 U18030 ( .A1(n14705), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n16057), .ZN(n14679) );
  AOI22_X1 U18031 ( .A1(n14708), .A2(DATAI_24_), .B1(n14707), .B2(n14677), 
        .ZN(n14678) );
  OAI211_X1 U18032 ( .C1(n15960), .C2(n14715), .A(n14679), .B(n14678), .ZN(
        P1_U2880) );
  AOI22_X1 U18033 ( .A1(n14705), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n16057), .ZN(n14681) );
  AOI22_X1 U18034 ( .A1(n14708), .A2(DATAI_23_), .B1(n14707), .B2(n20376), 
        .ZN(n14680) );
  OAI211_X1 U18035 ( .C1(n14682), .C2(n14715), .A(n14681), .B(n14680), .ZN(
        P1_U2881) );
  AOI22_X1 U18036 ( .A1(n14705), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n16057), .ZN(n14684) );
  AOI22_X1 U18037 ( .A1(n14708), .A2(DATAI_22_), .B1(n14707), .B2(n20361), 
        .ZN(n14683) );
  OAI211_X1 U18038 ( .C1(n15976), .C2(n14715), .A(n14684), .B(n14683), .ZN(
        P1_U2882) );
  INV_X1 U18039 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20355) );
  OAI22_X1 U18040 ( .A1(n14691), .A2(n20355), .B1(n14230), .B2(n14711), .ZN(
        n14685) );
  INV_X1 U18041 ( .A(n14685), .ZN(n14687) );
  AOI22_X1 U18042 ( .A1(n14708), .A2(DATAI_21_), .B1(n14707), .B2(n20354), 
        .ZN(n14686) );
  OAI211_X1 U18043 ( .C1(n14688), .C2(n14715), .A(n14687), .B(n14686), .ZN(
        P1_U2883) );
  AOI22_X1 U18044 ( .A1(n14705), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n16057), .ZN(n14690) );
  AOI22_X1 U18045 ( .A1(n14708), .A2(DATAI_20_), .B1(n14707), .B2(n20348), 
        .ZN(n14689) );
  OAI211_X1 U18046 ( .C1(n16069), .C2(n14715), .A(n14690), .B(n14689), .ZN(
        P1_U2884) );
  INV_X1 U18047 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20341) );
  NOR2_X1 U18048 ( .A1(n14691), .A2(n20341), .ZN(n14696) );
  INV_X1 U18049 ( .A(n14708), .ZN(n14694) );
  INV_X1 U18050 ( .A(DATAI_19_), .ZN(n14693) );
  OAI22_X1 U18051 ( .A1(n14694), .A2(n14693), .B1(n20340), .B2(n14692), .ZN(
        n14695) );
  AOI211_X1 U18052 ( .C1(n16057), .C2(P1_EAX_REG_19__SCAN_IN), .A(n14696), .B(
        n14695), .ZN(n14697) );
  OAI21_X1 U18053 ( .B1(n14698), .B2(n14715), .A(n14697), .ZN(P1_U2885) );
  AOI22_X1 U18054 ( .A1(n14705), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n16057), .ZN(n14701) );
  AOI22_X1 U18055 ( .A1(n14708), .A2(DATAI_18_), .B1(n14707), .B2(n14699), 
        .ZN(n14700) );
  OAI211_X1 U18056 ( .C1(n16014), .C2(n14715), .A(n14701), .B(n14700), .ZN(
        P1_U2886) );
  AOI22_X1 U18057 ( .A1(n14705), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n16057), .ZN(n14704) );
  AOI22_X1 U18058 ( .A1(n14708), .A2(DATAI_17_), .B1(n14707), .B2(n14702), 
        .ZN(n14703) );
  OAI211_X1 U18059 ( .C1(n16018), .C2(n14715), .A(n14704), .B(n14703), .ZN(
        P1_U2887) );
  AOI22_X1 U18060 ( .A1(n14705), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n16057), .ZN(n14710) );
  AOI22_X1 U18061 ( .A1(n14708), .A2(DATAI_16_), .B1(n14707), .B2(n14706), 
        .ZN(n14709) );
  OAI211_X1 U18062 ( .C1(n14790), .C2(n14715), .A(n14710), .B(n14709), .ZN(
        P1_U2888) );
  OAI222_X1 U18063 ( .A1(n14716), .A2(n14715), .B1(n14714), .B2(n14713), .C1(
        n14712), .C2(n14711), .ZN(P1_U2889) );
  XNOR2_X1 U18064 ( .A(n14718), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14853) );
  NAND2_X1 U18065 ( .A1(n20249), .A2(n14719), .ZN(n14720) );
  NAND2_X1 U18066 ( .A1(n20290), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14847) );
  OAI211_X1 U18067 ( .C1(n14721), .C2(n16074), .A(n14720), .B(n14847), .ZN(
        n14722) );
  AOI21_X1 U18068 ( .B1(n14723), .B2(n20313), .A(n14722), .ZN(n14724) );
  OAI21_X1 U18069 ( .B1(n14853), .B2(n20115), .A(n14724), .ZN(P1_U2970) );
  OR2_X1 U18070 ( .A1(n14726), .A2(n14725), .ZN(n14727) );
  MUX2_X1 U18071 ( .A(n14728), .B(n14727), .S(n16110), .Z(n14729) );
  INV_X1 U18072 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14857) );
  XNOR2_X1 U18073 ( .A(n14729), .B(n14857), .ZN(n14863) );
  NOR2_X1 U18074 ( .A1(n10234), .A2(n21053), .ZN(n14856) );
  AOI21_X1 U18075 ( .B1(n20244), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14856), .ZN(n14730) );
  OAI21_X1 U18076 ( .B1(n20243), .B2(n14731), .A(n14730), .ZN(n14732) );
  AOI21_X1 U18077 ( .B1(n14733), .B2(n20313), .A(n14732), .ZN(n14734) );
  OAI21_X1 U18078 ( .B1(n20115), .B2(n14863), .A(n14734), .ZN(P1_U2972) );
  NAND2_X1 U18079 ( .A1(n16063), .A2(n9814), .ZN(n14736) );
  NAND2_X1 U18080 ( .A1(n14736), .A2(n16110), .ZN(n14737) );
  NAND2_X1 U18081 ( .A1(n14738), .A2(n14737), .ZN(n14739) );
  XNOR2_X1 U18082 ( .A(n14739), .B(n14864), .ZN(n14874) );
  NAND2_X1 U18083 ( .A1(n20249), .A2(n14740), .ZN(n14741) );
  NAND2_X1 U18084 ( .A1(n20290), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14865) );
  OAI211_X1 U18085 ( .C1(n16074), .C2(n14742), .A(n14741), .B(n14865), .ZN(
        n14743) );
  AOI21_X1 U18086 ( .B1(n14744), .B2(n20313), .A(n14743), .ZN(n14745) );
  OAI21_X1 U18087 ( .B1(n20115), .B2(n14874), .A(n14745), .ZN(P1_U2973) );
  MUX2_X1 U18088 ( .A(n14882), .B(n14746), .S(n16086), .Z(n14747) );
  INV_X1 U18089 ( .A(n14747), .ZN(n14750) );
  NAND2_X1 U18090 ( .A1(n14756), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14749) );
  NAND2_X1 U18091 ( .A1(n14750), .A2(n14749), .ZN(n14751) );
  XNOR2_X1 U18092 ( .A(n14751), .B(n14870), .ZN(n14880) );
  INV_X1 U18093 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21116) );
  NOR2_X1 U18094 ( .A1(n10234), .A2(n21116), .ZN(n14876) );
  AOI21_X1 U18095 ( .B1(n20244), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n14876), .ZN(n14752) );
  OAI21_X1 U18096 ( .B1(n20243), .B2(n15946), .A(n14752), .ZN(n14753) );
  AOI21_X1 U18097 ( .B1(n15953), .B2(n20313), .A(n14753), .ZN(n14754) );
  OAI21_X1 U18098 ( .B1(n20115), .B2(n14880), .A(n14754), .ZN(P1_U2974) );
  NAND2_X1 U18099 ( .A1(n14756), .A2(n14755), .ZN(n14757) );
  MUX2_X1 U18100 ( .A(n14757), .B(n14756), .S(n16110), .Z(n14758) );
  XNOR2_X1 U18101 ( .A(n14758), .B(n14882), .ZN(n14888) );
  NAND2_X1 U18102 ( .A1(n20290), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14883) );
  OAI21_X1 U18103 ( .B1(n16074), .B2(n15966), .A(n14883), .ZN(n14760) );
  NOR2_X1 U18104 ( .A1(n15960), .A2(n20254), .ZN(n14759) );
  AOI211_X1 U18105 ( .C1(n20249), .C2(n15963), .A(n14760), .B(n14759), .ZN(
        n14761) );
  OAI21_X1 U18106 ( .B1(n20115), .B2(n14888), .A(n14761), .ZN(P1_U2975) );
  OAI22_X1 U18107 ( .A1(n16074), .A2(n15974), .B1(n10234), .B2(n16154), .ZN(
        n14762) );
  AOI21_X1 U18108 ( .B1(n15979), .B2(n20249), .A(n14762), .ZN(n14767) );
  NAND2_X1 U18109 ( .A1(n14764), .A2(n14763), .ZN(n14765) );
  XNOR2_X1 U18110 ( .A(n14765), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16149) );
  NAND2_X1 U18111 ( .A1(n16149), .A2(n20250), .ZN(n14766) );
  OAI211_X1 U18112 ( .C1(n15976), .C2(n20254), .A(n14767), .B(n14766), .ZN(
        P1_U2977) );
  OR3_X1 U18113 ( .A1(n16163), .A2(n16086), .A3(n11766), .ZN(n14770) );
  NAND2_X1 U18114 ( .A1(n16086), .A2(n16174), .ZN(n16076) );
  OR3_X1 U18115 ( .A1(n14778), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n16076), .ZN(n14769) );
  NAND2_X1 U18116 ( .A1(n14770), .A2(n14769), .ZN(n15927) );
  NAND2_X1 U18117 ( .A1(n15927), .A2(n15934), .ZN(n15929) );
  OAI22_X1 U18118 ( .A1(n15929), .A2(n16110), .B1(n15934), .B2(n14770), .ZN(
        n14771) );
  XNOR2_X1 U18119 ( .A(n14771), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14895) );
  NAND2_X1 U18120 ( .A1(n20290), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14890) );
  NAND2_X1 U18121 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14772) );
  OAI211_X1 U18122 ( .C1(n20243), .C2(n15981), .A(n14890), .B(n14772), .ZN(
        n14773) );
  AOI21_X1 U18123 ( .B1(n15987), .B2(n20313), .A(n14773), .ZN(n14774) );
  OAI21_X1 U18124 ( .B1(n14895), .B2(n20115), .A(n14774), .ZN(P1_U2978) );
  INV_X1 U18125 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n14775) );
  OAI22_X1 U18126 ( .A1(n16074), .A2(n16011), .B1(n10234), .B2(n14775), .ZN(
        n14776) );
  AOI21_X1 U18127 ( .B1(n16009), .B2(n20249), .A(n14776), .ZN(n14780) );
  OR2_X1 U18128 ( .A1(n14778), .A2(n14777), .ZN(n16164) );
  NAND3_X1 U18129 ( .A1(n16164), .A2(n16163), .A3(n20250), .ZN(n14779) );
  OAI211_X1 U18130 ( .C1(n16014), .C2(n20254), .A(n14780), .B(n14779), .ZN(
        P1_U2981) );
  INV_X1 U18131 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n14786) );
  OAI21_X1 U18132 ( .B1(n14781), .B2(n14782), .A(n14791), .ZN(n16094) );
  OAI21_X1 U18133 ( .B1(n16082), .B2(n16094), .A(n16095), .ZN(n14783) );
  XOR2_X1 U18134 ( .A(n14784), .B(n14783), .Z(n16192) );
  AOI22_X1 U18135 ( .A1(n20250), .A2(n16192), .B1(n20290), .B2(
        P1_REIP_REG_16__SCAN_IN), .ZN(n14785) );
  OAI21_X1 U18136 ( .B1(n16074), .B2(n14786), .A(n14785), .ZN(n14787) );
  AOI21_X1 U18137 ( .B1(n14788), .B2(n20249), .A(n14787), .ZN(n14789) );
  OAI21_X1 U18138 ( .B1(n14790), .B2(n20254), .A(n14789), .ZN(P1_U2983) );
  NAND2_X1 U18139 ( .A1(n14781), .A2(n14791), .ZN(n16083) );
  AOI21_X1 U18140 ( .B1(n16083), .B2(n14793), .A(n14792), .ZN(n14795) );
  AOI22_X1 U18141 ( .A1(n16086), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n10013), .B2(n16110), .ZN(n14794) );
  XNOR2_X1 U18142 ( .A(n14795), .B(n14794), .ZN(n16206) );
  INV_X1 U18143 ( .A(n16206), .ZN(n14799) );
  AOI22_X1 U18144 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20290), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n14796) );
  OAI21_X1 U18145 ( .B1(n20243), .B2(n16031), .A(n14796), .ZN(n14797) );
  AOI21_X1 U18146 ( .B1(n16036), .B2(n20313), .A(n14797), .ZN(n14798) );
  OAI21_X1 U18147 ( .B1(n14799), .B2(n20115), .A(n14798), .ZN(P1_U2985) );
  OR2_X1 U18148 ( .A1(n14781), .A2(n14801), .ZN(n14803) );
  NAND2_X1 U18149 ( .A1(n14803), .A2(n14802), .ZN(n16105) );
  INV_X1 U18150 ( .A(n14804), .ZN(n14805) );
  NOR2_X1 U18151 ( .A1(n10237), .A2(n16102), .ZN(n14806) );
  XOR2_X1 U18152 ( .A(n14807), .B(n14806), .Z(n16216) );
  NAND2_X1 U18153 ( .A1(n16216), .A2(n20250), .ZN(n14813) );
  INV_X1 U18154 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14809) );
  INV_X1 U18155 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n14808) );
  OAI22_X1 U18156 ( .A1(n16074), .A2(n14809), .B1(n10234), .B2(n14808), .ZN(
        n14810) );
  AOI21_X1 U18157 ( .B1(n14811), .B2(n20249), .A(n14810), .ZN(n14812) );
  OAI211_X1 U18158 ( .C1(n20254), .C2(n14814), .A(n14813), .B(n14812), .ZN(
        P1_U2986) );
  NAND2_X1 U18159 ( .A1(n14815), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14817) );
  XNOR2_X1 U18160 ( .A(n14781), .B(n16240), .ZN(n14816) );
  MUX2_X1 U18161 ( .A(n14817), .B(n14816), .S(n16110), .Z(n14819) );
  INV_X1 U18162 ( .A(n14815), .ZN(n14818) );
  NAND3_X1 U18163 ( .A1(n14818), .A2(n16086), .A3(n16240), .ZN(n16111) );
  NAND2_X1 U18164 ( .A1(n14819), .A2(n16111), .ZN(n16246) );
  INV_X1 U18165 ( .A(n16246), .ZN(n14825) );
  AOI22_X1 U18166 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n20290), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14820) );
  OAI21_X1 U18167 ( .B1(n20243), .B2(n14821), .A(n14820), .ZN(n14822) );
  AOI21_X1 U18168 ( .B1(n14823), .B2(n20313), .A(n14822), .ZN(n14824) );
  OAI21_X1 U18169 ( .B1(n14825), .B2(n20115), .A(n14824), .ZN(P1_U2989) );
  INV_X1 U18170 ( .A(n14826), .ZN(n14830) );
  NAND3_X1 U18171 ( .A1(n14858), .A2(n14846), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14837) );
  INV_X1 U18172 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14827) );
  NOR3_X1 U18173 ( .A1(n14837), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14827), .ZN(n14828) );
  AOI211_X1 U18174 ( .C1(n14830), .C2(n20292), .A(n14829), .B(n14828), .ZN(
        n14833) );
  OR2_X1 U18175 ( .A1(n14859), .A2(n10042), .ZN(n14831) );
  NAND2_X1 U18176 ( .A1(n14831), .A2(n14860), .ZN(n14843) );
  OAI211_X1 U18177 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n20293), .A(
        n14843), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14838) );
  NAND3_X1 U18178 ( .A1(n14838), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14860), .ZN(n14832) );
  OAI211_X1 U18179 ( .C1(n14834), .C2(n16225), .A(n14833), .B(n14832), .ZN(
        P1_U3000) );
  INV_X1 U18180 ( .A(n14835), .ZN(n14836) );
  AOI21_X1 U18181 ( .B1(n10231), .B2(n20292), .A(n14836), .ZN(n14841) );
  INV_X1 U18182 ( .A(n14837), .ZN(n14839) );
  OAI21_X1 U18183 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14839), .A(
        n14838), .ZN(n14840) );
  OAI211_X1 U18184 ( .C1(n14842), .C2(n16225), .A(n14841), .B(n14840), .ZN(
        P1_U3001) );
  INV_X1 U18185 ( .A(n14843), .ZN(n14851) );
  INV_X1 U18186 ( .A(n14844), .ZN(n14849) );
  NAND3_X1 U18187 ( .A1(n14858), .A2(n14846), .A3(n14845), .ZN(n14848) );
  OAI211_X1 U18188 ( .C1(n14849), .C2(n20288), .A(n14848), .B(n14847), .ZN(
        n14850) );
  AOI21_X1 U18189 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n14851), .A(
        n14850), .ZN(n14852) );
  OAI21_X1 U18190 ( .B1(n14853), .B2(n16225), .A(n14852), .ZN(P1_U3002) );
  NOR2_X1 U18191 ( .A1(n14854), .A2(n20288), .ZN(n14855) );
  AOI211_X1 U18192 ( .C1(n14858), .C2(n14857), .A(n14856), .B(n14855), .ZN(
        n14862) );
  NAND3_X1 U18193 ( .A1(n14860), .A2(n14859), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14861) );
  OAI211_X1 U18194 ( .C1(n14863), .C2(n16225), .A(n14862), .B(n14861), .ZN(
        P1_U3004) );
  NAND3_X1 U18195 ( .A1(n16138), .A2(n9814), .A3(n14864), .ZN(n14866) );
  OAI211_X1 U18196 ( .C1(n20288), .C2(n14867), .A(n14866), .B(n14865), .ZN(
        n14868) );
  INV_X1 U18197 ( .A(n14868), .ZN(n14873) );
  INV_X1 U18198 ( .A(n14869), .ZN(n14877) );
  AND3_X1 U18199 ( .A1(n16138), .A2(n14871), .A3(n14870), .ZN(n14875) );
  OAI21_X1 U18200 ( .B1(n14877), .B2(n14875), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14872) );
  OAI211_X1 U18201 ( .C1(n14874), .C2(n16225), .A(n14873), .B(n14872), .ZN(
        P1_U3005) );
  AOI211_X1 U18202 ( .C1(n20292), .C2(n15952), .A(n14876), .B(n14875), .ZN(
        n14879) );
  NAND2_X1 U18203 ( .A1(n14877), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14878) );
  OAI211_X1 U18204 ( .C1(n14880), .C2(n16225), .A(n14879), .B(n14878), .ZN(
        P1_U3006) );
  OAI21_X1 U18205 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n20279), .A(
        n14881), .ZN(n14886) );
  NAND3_X1 U18206 ( .A1(n16138), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n14882), .ZN(n14884) );
  OAI211_X1 U18207 ( .C1(n20288), .C2(n15959), .A(n14884), .B(n14883), .ZN(
        n14885) );
  AOI21_X1 U18208 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14886), .A(
        n14885), .ZN(n14887) );
  OAI21_X1 U18209 ( .B1(n14888), .B2(n16225), .A(n14887), .ZN(P1_U3007) );
  INV_X1 U18210 ( .A(n16273), .ZN(n16265) );
  AND2_X1 U18211 ( .A1(n16265), .A2(n14889), .ZN(n16151) );
  NAND2_X1 U18212 ( .A1(n16145), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14891) );
  OAI211_X1 U18213 ( .C1(n20288), .C2(n15988), .A(n14891), .B(n14890), .ZN(
        n14892) );
  AOI21_X1 U18214 ( .B1(n16151), .B2(n14893), .A(n14892), .ZN(n14894) );
  OAI21_X1 U18215 ( .B1(n14895), .B2(n16225), .A(n14894), .ZN(P1_U3010) );
  NAND2_X1 U18216 ( .A1(n9675), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20671) );
  XNOR2_X1 U18217 ( .A(n11830), .B(n20671), .ZN(n14897) );
  OAI22_X1 U18218 ( .A1(n14897), .A2(n20817), .B1(n13690), .B2(n14896), .ZN(
        n14898) );
  MUX2_X1 U18219 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n14898), .S(
        n20302), .Z(P1_U3476) );
  INV_X1 U18220 ( .A(n19996), .ZN(n14900) );
  OAI21_X1 U18221 ( .B1(n14900), .B2(n19541), .A(n14899), .ZN(n14903) );
  NAND2_X1 U18222 ( .A1(n14901), .A2(n14900), .ZN(n14902) );
  MUX2_X1 U18223 ( .A(n14903), .B(n14902), .S(n9676), .Z(n14905) );
  OAI22_X1 U18224 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16542), .B1(n20003), 
        .B2(n19926), .ZN(n14904) );
  NAND2_X1 U18225 ( .A1(n14905), .A2(n14904), .ZN(n14911) );
  NOR2_X1 U18226 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n14906), .ZN(n14908) );
  AOI211_X1 U18227 ( .C1(n14909), .C2(n19356), .A(n14908), .B(n14907), .ZN(
        n14910) );
  MUX2_X1 U18228 ( .A(n14911), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n14910), 
        .Z(P2_U3610) );
  INV_X1 U18229 ( .A(n14912), .ZN(n14914) );
  MUX2_X1 U18230 ( .A(n14914), .B(n16540), .S(n9676), .Z(n14917) );
  OAI21_X1 U18231 ( .B1(n14917), .B2(n14916), .A(n14915), .ZN(n14919) );
  MUX2_X1 U18232 ( .A(n14919), .B(P2_MORE_REG_SCAN_IN), .S(n14918), .Z(
        P2_U3609) );
  AOI21_X1 U18233 ( .B1(n14938), .B2(n13426), .A(n14937), .ZN(n16311) );
  NOR2_X1 U18234 ( .A1(n14920), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14921) );
  OR2_X1 U18235 ( .A1(n13317), .A2(n14921), .ZN(n16310) );
  OR2_X1 U18236 ( .A1(n15103), .A2(n14923), .ZN(n16303) );
  OAI21_X1 U18237 ( .B1(n14922), .B2(n16312), .A(n19151), .ZN(n14924) );
  NAND2_X1 U18238 ( .A1(n14924), .A2(n14923), .ZN(n14935) );
  OAI22_X1 U18239 ( .A1(n19186), .A2(n14926), .B1(n14925), .B2(n19215), .ZN(
        n14927) );
  OR2_X1 U18240 ( .A1(n14927), .A2(n10244), .ZN(n14928) );
  OAI211_X1 U18241 ( .C1(n16313), .C2(n16303), .A(n14935), .B(n14934), .ZN(
        P2_U2825) );
  INV_X1 U18242 ( .A(n14936), .ZN(n15144) );
  AOI21_X1 U18243 ( .B1(n14938), .B2(n14937), .A(n16312), .ZN(n14940) );
  INV_X1 U18244 ( .A(n16311), .ZN(n14939) );
  OAI21_X1 U18245 ( .B1(n19167), .B2(n14940), .A(n14939), .ZN(n14946) );
  NAND2_X1 U18246 ( .A1(n19183), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n14942) );
  AOI22_X1 U18247 ( .A1(n19221), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(
        n19199), .B2(P2_REIP_REG_28__SCAN_IN), .ZN(n14941) );
  OAI211_X1 U18248 ( .C1(n19231), .C2(n15197), .A(n14942), .B(n14941), .ZN(
        n14943) );
  AOI21_X1 U18249 ( .B1(n14944), .B2(n19189), .A(n14943), .ZN(n14945) );
  OAI211_X1 U18250 ( .C1(n19129), .C2(n15144), .A(n14946), .B(n14945), .ZN(
        P2_U2827) );
  INV_X1 U18251 ( .A(n14947), .ZN(n14960) );
  AOI21_X1 U18252 ( .B1(n9738), .B2(n15290), .A(n16312), .ZN(n14948) );
  OAI21_X1 U18253 ( .B1(n14948), .B2(n19167), .A(n16326), .ZN(n14959) );
  AND2_X1 U18254 ( .A1(n14966), .A2(n14949), .ZN(n14950) );
  NOR2_X1 U18255 ( .A1(n15209), .A2(n14950), .ZN(n15461) );
  AOI22_X1 U18256 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n19183), .B1(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n19221), .ZN(n14951) );
  OAI21_X1 U18257 ( .B1(n19215), .B2(n20048), .A(n14951), .ZN(n14957) );
  OR2_X1 U18258 ( .A1(n14953), .A2(n14954), .ZN(n14955) );
  NAND2_X1 U18259 ( .A1(n14952), .A2(n14955), .ZN(n15458) );
  NOR2_X1 U18260 ( .A1(n15458), .A2(n19129), .ZN(n14956) );
  AOI211_X1 U18261 ( .C1(n19209), .C2(n15461), .A(n14957), .B(n14956), .ZN(
        n14958) );
  OAI211_X1 U18262 ( .C1(n19216), .C2(n14960), .A(n14959), .B(n14958), .ZN(
        P2_U2830) );
  AOI21_X1 U18263 ( .B1(n14977), .B2(n14961), .A(n16312), .ZN(n14962) );
  OAI21_X1 U18264 ( .B1(n19167), .B2(n14962), .A(n9738), .ZN(n14973) );
  NAND2_X1 U18265 ( .A1(n14963), .A2(n14964), .ZN(n14965) );
  NAND2_X1 U18266 ( .A1(n14966), .A2(n14965), .ZN(n15479) );
  AOI22_X1 U18267 ( .A1(n19221), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n19199), .B2(P2_REIP_REG_24__SCAN_IN), .ZN(n14967) );
  OAI21_X1 U18268 ( .B1(n15479), .B2(n19231), .A(n14967), .ZN(n14971) );
  NOR2_X1 U18269 ( .A1(n14981), .A2(n14968), .ZN(n14969) );
  OR2_X1 U18270 ( .A1(n14953), .A2(n14969), .ZN(n15478) );
  NOR2_X1 U18271 ( .A1(n15478), .A2(n19129), .ZN(n14970) );
  AOI211_X1 U18272 ( .C1(P2_EBX_REG_24__SCAN_IN), .C2(n19183), .A(n14971), .B(
        n14970), .ZN(n14972) );
  OAI211_X1 U18273 ( .C1(n19216), .C2(n14974), .A(n14973), .B(n14972), .ZN(
        P2_U2831) );
  INV_X1 U18274 ( .A(n14975), .ZN(n14991) );
  AOI21_X1 U18275 ( .B1(n10086), .B2(n15300), .A(n16312), .ZN(n14978) );
  OAI21_X1 U18276 ( .B1(n14978), .B2(n19167), .A(n14977), .ZN(n14990) );
  NOR2_X1 U18277 ( .A1(n15502), .A2(n14979), .ZN(n14980) );
  OR2_X1 U18278 ( .A1(n14981), .A2(n14980), .ZN(n15492) );
  INV_X1 U18279 ( .A(n15492), .ZN(n16335) );
  AOI22_X1 U18280 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n19221), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n19199), .ZN(n14986) );
  OR2_X1 U18281 ( .A1(n14982), .A2(n14983), .ZN(n14984) );
  AND2_X1 U18282 ( .A1(n14963), .A2(n14984), .ZN(n15489) );
  NAND2_X1 U18283 ( .A1(n19209), .A2(n15489), .ZN(n14985) );
  OAI211_X1 U18284 ( .C1(n19218), .C2(n14987), .A(n14986), .B(n14985), .ZN(
        n14988) );
  AOI21_X1 U18285 ( .B1(n16335), .B2(n19226), .A(n14988), .ZN(n14989) );
  OAI211_X1 U18286 ( .C1(n14991), .C2(n19216), .A(n14990), .B(n14989), .ZN(
        P2_U2832) );
  AOI21_X1 U18287 ( .B1(n19148), .B2(n9770), .A(n16312), .ZN(n14993) );
  INV_X1 U18288 ( .A(n19132), .ZN(n14992) );
  OAI21_X1 U18289 ( .B1(n19167), .B2(n14993), .A(n14992), .ZN(n15005) );
  NAND2_X1 U18290 ( .A1(n14351), .A2(n14995), .ZN(n14996) );
  AND2_X1 U18291 ( .A1(n14994), .A2(n14996), .ZN(n16360) );
  NAND2_X1 U18292 ( .A1(n19221), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14997) );
  OAI211_X1 U18293 ( .C1(n15355), .C2(n19215), .A(n14997), .B(n19214), .ZN(
        n15003) );
  NOR2_X1 U18294 ( .A1(n14998), .A2(n14999), .ZN(n15000) );
  OR2_X1 U18295 ( .A1(n15183), .A2(n15000), .ZN(n16346) );
  OAI22_X1 U18296 ( .A1(n16346), .A2(n19129), .B1(n19218), .B2(n15001), .ZN(
        n15002) );
  AOI211_X1 U18297 ( .C1(n16360), .C2(n19209), .A(n15003), .B(n15002), .ZN(
        n15004) );
  OAI211_X1 U18298 ( .C1(n19216), .C2(n15006), .A(n15005), .B(n15004), .ZN(
        P2_U2837) );
  AOI21_X1 U18299 ( .B1(n19227), .B2(n15016), .A(n19167), .ZN(n15024) );
  INV_X1 U18300 ( .A(n15007), .ZN(n15019) );
  OR2_X1 U18301 ( .A1(n15008), .A2(n13411), .ZN(n15010) );
  NAND2_X1 U18302 ( .A1(n15010), .A2(n15009), .ZN(n19235) );
  INV_X1 U18303 ( .A(n19235), .ZN(n15586) );
  INV_X1 U18304 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20033) );
  OAI21_X1 U18305 ( .B1(n19215), .B2(n20033), .A(n19214), .ZN(n15012) );
  INV_X1 U18306 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15372) );
  NOR2_X1 U18307 ( .A1(n19186), .A2(n15372), .ZN(n15011) );
  AOI211_X1 U18308 ( .C1(n19226), .C2(n15586), .A(n15012), .B(n15011), .ZN(
        n15013) );
  OAI21_X1 U18309 ( .B1(n19218), .B2(n15014), .A(n15013), .ZN(n15018) );
  INV_X1 U18310 ( .A(n15371), .ZN(n15015) );
  NOR3_X1 U18311 ( .A1(n15103), .A2(n15016), .A3(n15015), .ZN(n15017) );
  AOI211_X1 U18312 ( .C1(n19189), .C2(n15019), .A(n15018), .B(n15017), .ZN(
        n15023) );
  AOI21_X1 U18313 ( .B1(n15021), .B2(n15020), .A(n14352), .ZN(n19268) );
  NAND2_X1 U18314 ( .A1(n19268), .A2(n19209), .ZN(n15022) );
  OAI211_X1 U18315 ( .C1(n15371), .C2(n15024), .A(n15023), .B(n15022), .ZN(
        P2_U2839) );
  AOI21_X1 U18316 ( .B1(n19227), .B2(n15036), .A(n19167), .ZN(n15040) );
  OR2_X1 U18317 ( .A1(n15026), .A2(n15025), .ZN(n15028) );
  NAND2_X1 U18318 ( .A1(n15028), .A2(n15027), .ZN(n19239) );
  AOI21_X1 U18319 ( .B1(n15030), .B2(n15029), .A(n13408), .ZN(n19274) );
  AOI22_X1 U18320 ( .A1(n19209), .A2(n19274), .B1(n19221), .B2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15032) );
  AOI21_X1 U18321 ( .B1(n19199), .B2(P2_REIP_REG_14__SCAN_IN), .A(n19198), 
        .ZN(n15031) );
  OAI211_X1 U18322 ( .C1(n19129), .C2(n19239), .A(n15032), .B(n15031), .ZN(
        n15035) );
  NOR2_X1 U18323 ( .A1(n15033), .A2(n19216), .ZN(n15034) );
  AOI211_X1 U18324 ( .C1(P2_EBX_REG_14__SCAN_IN), .C2(n19183), .A(n15035), .B(
        n15034), .ZN(n15039) );
  OR2_X1 U18325 ( .A1(n15103), .A2(n15036), .ZN(n19160) );
  INV_X1 U18326 ( .A(n19160), .ZN(n15037) );
  NAND2_X1 U18327 ( .A1(n15037), .A2(n16400), .ZN(n15038) );
  OAI211_X1 U18328 ( .C1(n15040), .C2(n16400), .A(n15039), .B(n15038), .ZN(
        P2_U2841) );
  AOI21_X1 U18329 ( .B1(n19227), .B2(n15057), .A(n19167), .ZN(n15061) );
  INV_X1 U18330 ( .A(n15041), .ZN(n15042) );
  OR2_X1 U18331 ( .A1(n15043), .A2(n15042), .ZN(n15046) );
  INV_X1 U18332 ( .A(n15044), .ZN(n15045) );
  AND2_X1 U18333 ( .A1(n15046), .A2(n15045), .ZN(n19284) );
  AOI22_X1 U18334 ( .A1(n19209), .A2(n19284), .B1(n19221), .B2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15052) );
  OR2_X1 U18335 ( .A1(n15048), .A2(n15047), .ZN(n15050) );
  AND2_X1 U18336 ( .A1(n15050), .A2(n15049), .ZN(n19250) );
  AOI21_X1 U18337 ( .B1(n19250), .B2(n19226), .A(n19198), .ZN(n15051) );
  OAI211_X1 U18338 ( .C1(n19215), .C2(n15053), .A(n15052), .B(n15051), .ZN(
        n15056) );
  NOR2_X1 U18339 ( .A1(n15054), .A2(n19216), .ZN(n15055) );
  AOI211_X1 U18340 ( .C1(P2_EBX_REG_10__SCAN_IN), .C2(n19183), .A(n15056), .B(
        n15055), .ZN(n15060) );
  INV_X1 U18341 ( .A(n15057), .ZN(n15058) );
  NAND3_X1 U18342 ( .A1(n15133), .A2(n16435), .A3(n15058), .ZN(n15059) );
  OAI211_X1 U18343 ( .C1(n15061), .C2(n16435), .A(n15060), .B(n15059), .ZN(
        P2_U2845) );
  INV_X1 U18344 ( .A(n15073), .ZN(n15062) );
  AOI21_X1 U18345 ( .B1(n19227), .B2(n15062), .A(n19167), .ZN(n15076) );
  INV_X1 U18346 ( .A(n15063), .ZN(n16437) );
  OR2_X1 U18347 ( .A1(n15065), .A2(n15064), .ZN(n15066) );
  NAND2_X1 U18348 ( .A1(n15066), .A2(n15041), .ZN(n19288) );
  INV_X1 U18349 ( .A(n19288), .ZN(n15067) );
  AOI22_X1 U18350 ( .A1(n19209), .A2(n15067), .B1(n19221), .B2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15070) );
  OAI21_X1 U18351 ( .B1(n19215), .B2(n16436), .A(n19214), .ZN(n15068) );
  AOI21_X1 U18352 ( .B1(n19226), .B2(n16442), .A(n15068), .ZN(n15069) );
  OAI211_X1 U18353 ( .C1(n19218), .C2(n13838), .A(n15070), .B(n15069), .ZN(
        n15071) );
  AOI21_X1 U18354 ( .B1(n15072), .B2(n19189), .A(n15071), .ZN(n15075) );
  NAND3_X1 U18355 ( .A1(n15133), .A2(n15073), .A3(n16437), .ZN(n15074) );
  OAI211_X1 U18356 ( .C1(n15076), .C2(n16437), .A(n15075), .B(n15074), .ZN(
        P2_U2846) );
  AOI21_X1 U18357 ( .B1(n19227), .B2(n15085), .A(n19167), .ZN(n15089) );
  OR2_X1 U18358 ( .A1(n15077), .A2(n9783), .ZN(n15078) );
  NAND2_X1 U18359 ( .A1(n15078), .A2(n13832), .ZN(n19258) );
  AOI21_X1 U18360 ( .B1(n15079), .B2(n14275), .A(n15064), .ZN(n19289) );
  AOI22_X1 U18361 ( .A1(n19209), .A2(n19289), .B1(n19221), .B2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15081) );
  AOI21_X1 U18362 ( .B1(n19199), .B2(P2_REIP_REG_8__SCAN_IN), .A(n19198), .ZN(
        n15080) );
  OAI211_X1 U18363 ( .C1(n19129), .C2(n19258), .A(n15081), .B(n15080), .ZN(
        n15084) );
  NOR2_X1 U18364 ( .A1(n15082), .A2(n19216), .ZN(n15083) );
  AOI211_X1 U18365 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n19183), .A(n15084), .B(
        n15083), .ZN(n15088) );
  INV_X1 U18366 ( .A(n15085), .ZN(n15086) );
  NAND3_X1 U18367 ( .A1(n15133), .A2(n16459), .A3(n15086), .ZN(n15087) );
  OAI211_X1 U18368 ( .C1(n15089), .C2(n16459), .A(n15088), .B(n15087), .ZN(
        P2_U2847) );
  AOI21_X1 U18369 ( .B1(n19227), .B2(n15102), .A(n19167), .ZN(n15106) );
  INV_X1 U18370 ( .A(n19263), .ZN(n19398) );
  NOR2_X1 U18371 ( .A1(n19215), .A2(n19392), .ZN(n15090) );
  AOI211_X1 U18372 ( .C1(n15091), .C2(n19189), .A(n19198), .B(n15090), .ZN(
        n15093) );
  AOI22_X1 U18373 ( .A1(n19209), .A2(n19305), .B1(n19221), .B2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n15092) );
  OAI211_X1 U18374 ( .C1(n19218), .C2(n10627), .A(n15093), .B(n15092), .ZN(
        n15100) );
  NAND2_X1 U18375 ( .A1(n15095), .A2(n15094), .ZN(n15097) );
  NAND2_X1 U18376 ( .A1(n15097), .A2(n15096), .ZN(n19307) );
  NOR2_X1 U18377 ( .A1(n19307), .A2(n15098), .ZN(n15099) );
  AOI211_X1 U18378 ( .C1(n19398), .C2(n19226), .A(n15100), .B(n15099), .ZN(
        n15105) );
  INV_X1 U18379 ( .A(n19404), .ZN(n15101) );
  OR3_X1 U18380 ( .A1(n15103), .A2(n15102), .A3(n15101), .ZN(n15104) );
  OAI211_X1 U18381 ( .C1(n15106), .C2(n19404), .A(n15105), .B(n15104), .ZN(
        P2_U2851) );
  INV_X1 U18382 ( .A(n15117), .ZN(n15107) );
  AOI21_X1 U18383 ( .B1(n19227), .B2(n15107), .A(n19167), .ZN(n15121) );
  INV_X1 U18384 ( .A(n16472), .ZN(n15120) );
  XNOR2_X1 U18385 ( .A(n15108), .B(n15109), .ZN(n20078) );
  INV_X1 U18386 ( .A(n13743), .ZN(n15110) );
  INV_X1 U18387 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n15112) );
  OAI22_X1 U18388 ( .A1(n19218), .A2(n15112), .B1(n15111), .B2(n19216), .ZN(
        n15114) );
  OAI22_X1 U18389 ( .A1(n16484), .A2(n19186), .B1(n16471), .B2(n19215), .ZN(
        n15113) );
  AOI211_X1 U18390 ( .C1(n19226), .C2(n15110), .A(n15114), .B(n15113), .ZN(
        n15115) );
  OAI21_X1 U18391 ( .B1(n20078), .B2(n19231), .A(n15115), .ZN(n15116) );
  AOI21_X1 U18392 ( .B1(n20074), .B2(n15131), .A(n15116), .ZN(n15119) );
  NAND3_X1 U18393 ( .A1(n15133), .A2(n15117), .A3(n15120), .ZN(n15118) );
  OAI211_X1 U18394 ( .C1(n15121), .C2(n15120), .A(n15119), .B(n15118), .ZN(
        P2_U2852) );
  AOI21_X1 U18395 ( .B1(n19227), .B2(n15122), .A(n19167), .ZN(n15137) );
  OAI22_X1 U18396 ( .A1(n19218), .A2(n15123), .B1(n19298), .B2(n19231), .ZN(
        n15124) );
  AOI21_X1 U18397 ( .B1(n19189), .B2(n15125), .A(n15124), .ZN(n15126) );
  OAI21_X1 U18398 ( .B1(n20014), .B2(n19215), .A(n15126), .ZN(n15127) );
  AOI21_X1 U18399 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19221), .A(
        n15127), .ZN(n15128) );
  OAI21_X1 U18400 ( .B1(n15129), .B2(n19129), .A(n15128), .ZN(n15130) );
  AOI21_X1 U18401 ( .B1(n19540), .B2(n15131), .A(n15130), .ZN(n15135) );
  NAND3_X1 U18402 ( .A1(n15133), .A2(n15136), .A3(n15132), .ZN(n15134) );
  OAI211_X1 U18403 ( .C1(n15137), .C2(n15136), .A(n15135), .B(n15134), .ZN(
        P2_U2853) );
  NAND2_X1 U18404 ( .A1(n15138), .A2(n15139), .ZN(n15140) );
  XOR2_X1 U18405 ( .A(n15141), .B(n15140), .Z(n15199) );
  NAND2_X1 U18406 ( .A1(n15199), .A2(n19260), .ZN(n15143) );
  NAND2_X1 U18407 ( .A1(n19259), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15142) );
  OAI211_X1 U18408 ( .C1(n19259), .C2(n15144), .A(n15143), .B(n15142), .ZN(
        P2_U2859) );
  AOI21_X1 U18409 ( .B1(n15147), .B2(n15146), .A(n15145), .ZN(n15148) );
  INV_X1 U18410 ( .A(n15148), .ZN(n15206) );
  NAND2_X1 U18411 ( .A1(n19259), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15150) );
  NAND2_X1 U18412 ( .A1(n15438), .A2(n19252), .ZN(n15149) );
  OAI211_X1 U18413 ( .C1(n15206), .C2(n19254), .A(n15150), .B(n15149), .ZN(
        P2_U2860) );
  NAND2_X1 U18414 ( .A1(n14952), .A2(n15151), .ZN(n15152) );
  NAND2_X1 U18415 ( .A1(n15153), .A2(n15152), .ZN(n16322) );
  AOI21_X1 U18416 ( .B1(n15156), .B2(n15155), .A(n15154), .ZN(n15207) );
  NAND2_X1 U18417 ( .A1(n15207), .A2(n19260), .ZN(n15158) );
  NAND2_X1 U18418 ( .A1(n19259), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15157) );
  OAI211_X1 U18419 ( .C1(n16322), .C2(n19259), .A(n15158), .B(n15157), .ZN(
        P2_U2861) );
  OAI21_X1 U18420 ( .B1(n15160), .B2(n15162), .A(n15161), .ZN(n15219) );
  MUX2_X1 U18421 ( .A(n15458), .B(n15163), .S(n19259), .Z(n15164) );
  OAI21_X1 U18422 ( .B1(n15219), .B2(n19254), .A(n15164), .ZN(P2_U2862) );
  AOI21_X1 U18423 ( .B1(n9688), .B2(n15166), .A(n15165), .ZN(n15168) );
  XNOR2_X1 U18424 ( .A(n15168), .B(n15167), .ZN(n15225) );
  NAND2_X1 U18425 ( .A1(n15225), .A2(n19260), .ZN(n15170) );
  NAND2_X1 U18426 ( .A1(n19259), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n15169) );
  OAI211_X1 U18427 ( .C1(n15478), .C2(n19259), .A(n15170), .B(n15169), .ZN(
        P2_U2863) );
  OAI21_X1 U18428 ( .B1(n9737), .B2(n15173), .A(n15172), .ZN(n15243) );
  NAND2_X1 U18429 ( .A1(n15336), .A2(n15174), .ZN(n15175) );
  NAND2_X1 U18430 ( .A1(n15501), .A2(n15175), .ZN(n19106) );
  NOR2_X1 U18431 ( .A1(n19106), .A2(n19259), .ZN(n15176) );
  AOI21_X1 U18432 ( .B1(P2_EBX_REG_21__SCAN_IN), .B2(n19259), .A(n15176), .ZN(
        n15177) );
  OAI21_X1 U18433 ( .B1(n15243), .B2(n19254), .A(n15177), .ZN(P2_U2866) );
  OAI21_X1 U18434 ( .B1(n15178), .B2(n15180), .A(n15179), .ZN(n15255) );
  OR2_X1 U18435 ( .A1(n15183), .A2(n15182), .ZN(n15184) );
  NAND2_X1 U18436 ( .A1(n15181), .A2(n15184), .ZN(n19130) );
  NOR2_X1 U18437 ( .A1(n19259), .A2(n19130), .ZN(n15185) );
  AOI21_X1 U18438 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n19259), .A(n15185), .ZN(
        n15186) );
  OAI21_X1 U18439 ( .B1(n15255), .B2(n19254), .A(n15186), .ZN(P2_U2868) );
  OR2_X1 U18440 ( .A1(n15187), .A2(n19254), .ZN(n15191) );
  AND2_X1 U18441 ( .A1(n15009), .A2(n15188), .ZN(n15189) );
  OR2_X1 U18442 ( .A1(n15189), .A2(n14998), .ZN(n15569) );
  NAND2_X1 U18443 ( .A1(n19252), .A2(n19143), .ZN(n15190) );
  OAI211_X1 U18444 ( .C1(n19252), .C2(n19145), .A(n15191), .B(n15190), .ZN(
        P2_U2870) );
  INV_X1 U18445 ( .A(n16306), .ZN(n15192) );
  AOI22_X1 U18446 ( .A1(n15192), .A2(n19321), .B1(P2_EAX_REG_31__SCAN_IN), 
        .B2(n19320), .ZN(n15194) );
  NAND2_X1 U18447 ( .A1(n19266), .A2(BUF2_REG_31__SCAN_IN), .ZN(n15193) );
  OAI211_X1 U18448 ( .C1(n15248), .C2(n20371), .A(n15194), .B(n15193), .ZN(
        P2_U2888) );
  AOI22_X1 U18449 ( .A1(n19266), .A2(BUF2_REG_28__SCAN_IN), .B1(n19265), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n15196) );
  INV_X1 U18450 ( .A(n15247), .ZN(n19264) );
  MUX2_X1 U18451 ( .A(BUF1_REG_12__SCAN_IN), .B(BUF2_REG_12__SCAN_IN), .S(
        n15220), .Z(n19371) );
  AOI22_X1 U18452 ( .A1(n19264), .A2(n19371), .B1(P2_EAX_REG_28__SCAN_IN), 
        .B2(n19320), .ZN(n15195) );
  OAI211_X1 U18453 ( .C1(n15197), .C2(n15223), .A(n15196), .B(n15195), .ZN(
        n15198) );
  AOI21_X1 U18454 ( .B1(n15199), .B2(n19308), .A(n15198), .ZN(n15200) );
  INV_X1 U18455 ( .A(n15200), .ZN(P2_U2891) );
  INV_X1 U18456 ( .A(n15436), .ZN(n15203) );
  OAI22_X1 U18457 ( .A1(n15247), .A2(n19282), .B1(n19293), .B2(n15201), .ZN(
        n15202) );
  AOI21_X1 U18458 ( .B1(n19321), .B2(n15203), .A(n15202), .ZN(n15205) );
  AOI22_X1 U18459 ( .A1(n19266), .A2(BUF2_REG_27__SCAN_IN), .B1(n19265), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n15204) );
  OAI211_X1 U18460 ( .C1(n15206), .C2(n19325), .A(n15205), .B(n15204), .ZN(
        P2_U2892) );
  NAND2_X1 U18461 ( .A1(n15207), .A2(n19308), .ZN(n15214) );
  MUX2_X1 U18462 ( .A(BUF1_REG_10__SCAN_IN), .B(BUF2_REG_10__SCAN_IN), .S(
        n15220), .Z(n19367) );
  AOI22_X1 U18463 ( .A1(n19264), .A2(n19367), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n19320), .ZN(n15213) );
  AOI22_X1 U18464 ( .A1(n19266), .A2(BUF2_REG_26__SCAN_IN), .B1(n19265), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n15212) );
  OR2_X1 U18465 ( .A1(n15209), .A2(n15208), .ZN(n15210) );
  AND2_X1 U18466 ( .A1(n13449), .A2(n15210), .ZN(n16320) );
  NAND2_X1 U18467 ( .A1(n19321), .A2(n16320), .ZN(n15211) );
  NAND4_X1 U18468 ( .A1(n15214), .A2(n15213), .A3(n15212), .A4(n15211), .ZN(
        P2_U2893) );
  OAI22_X1 U18469 ( .A1(n15247), .A2(n19287), .B1(n19293), .B2(n15215), .ZN(
        n15216) );
  AOI21_X1 U18470 ( .B1(n19321), .B2(n15461), .A(n15216), .ZN(n15218) );
  AOI22_X1 U18471 ( .A1(n19266), .A2(BUF2_REG_25__SCAN_IN), .B1(n19265), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n15217) );
  OAI211_X1 U18472 ( .C1(n15219), .C2(n19325), .A(n15218), .B(n15217), .ZN(
        P2_U2894) );
  AOI22_X1 U18473 ( .A1(n19266), .A2(BUF2_REG_24__SCAN_IN), .B1(n19265), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n15222) );
  MUX2_X1 U18474 ( .A(BUF1_REG_8__SCAN_IN), .B(BUF2_REG_8__SCAN_IN), .S(n15220), .Z(n19363) );
  AOI22_X1 U18475 ( .A1(n19264), .A2(n19363), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n19320), .ZN(n15221) );
  OAI211_X1 U18476 ( .C1(n15223), .C2(n15479), .A(n15222), .B(n15221), .ZN(
        n15224) );
  AOI21_X1 U18477 ( .B1(n15225), .B2(n19308), .A(n15224), .ZN(n15226) );
  INV_X1 U18478 ( .A(n15226), .ZN(P2_U2895) );
  AOI21_X1 U18479 ( .B1(n15227), .B2(n15229), .A(n15228), .ZN(n16336) );
  INV_X1 U18480 ( .A(n16336), .ZN(n15234) );
  OAI22_X1 U18481 ( .A1(n15247), .A2(n19441), .B1(n15230), .B2(n19293), .ZN(
        n15231) );
  AOI21_X1 U18482 ( .B1(n19321), .B2(n15489), .A(n15231), .ZN(n15233) );
  AOI22_X1 U18483 ( .A1(n19266), .A2(BUF2_REG_23__SCAN_IN), .B1(n19265), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n15232) );
  OAI211_X1 U18484 ( .C1(n15234), .C2(n19325), .A(n15233), .B(n15232), .ZN(
        P2_U2896) );
  OR2_X1 U18485 ( .A1(n15530), .A2(n15235), .ZN(n15237) );
  INV_X1 U18486 ( .A(n15504), .ZN(n15236) );
  AND2_X1 U18487 ( .A1(n15237), .A2(n15236), .ZN(n19104) );
  OAI22_X1 U18488 ( .A1(n15247), .A2(n19424), .B1(n19293), .B2(n15238), .ZN(
        n15241) );
  INV_X1 U18489 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n15239) );
  OAI22_X1 U18490 ( .A1(n15250), .A2(n15239), .B1(n15248), .B2(n20355), .ZN(
        n15240) );
  AOI211_X1 U18491 ( .C1(n19321), .C2(n19104), .A(n15241), .B(n15240), .ZN(
        n15242) );
  OAI21_X1 U18492 ( .B1(n15243), .B2(n19325), .A(n15242), .ZN(P2_U2898) );
  NAND2_X1 U18493 ( .A1(n14994), .A2(n15244), .ZN(n15245) );
  NAND2_X1 U18494 ( .A1(n15529), .A2(n15245), .ZN(n19139) );
  INV_X1 U18495 ( .A(n19139), .ZN(n15253) );
  OAI22_X1 U18496 ( .A1(n15247), .A2(n19319), .B1(n19293), .B2(n15246), .ZN(
        n15252) );
  INV_X1 U18497 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n15249) );
  OAI22_X1 U18498 ( .A1(n15250), .A2(n15249), .B1(n15248), .B2(n20341), .ZN(
        n15251) );
  AOI211_X1 U18499 ( .C1(n19321), .C2(n15253), .A(n15252), .B(n15251), .ZN(
        n15254) );
  OAI21_X1 U18500 ( .B1(n15255), .B2(n19325), .A(n15254), .ZN(P2_U2900) );
  NAND2_X1 U18501 ( .A1(n15257), .A2(n15256), .ZN(n15259) );
  XOR2_X1 U18502 ( .A(n15259), .B(n15258), .Z(n15433) );
  AOI21_X1 U18503 ( .B1(n12339), .B2(n15422), .A(n15260), .ZN(n15431) );
  NOR2_X1 U18504 ( .A1(n16310), .A2(n19405), .ZN(n15263) );
  NAND2_X1 U18505 ( .A1(n19198), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15420) );
  NAND2_X1 U18506 ( .A1(n16447), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15261) );
  OAI211_X1 U18507 ( .C1(n16309), .C2(n16414), .A(n15420), .B(n15261), .ZN(
        n15262) );
  AOI211_X1 U18508 ( .C1(n15431), .C2(n19400), .A(n15263), .B(n15262), .ZN(
        n15264) );
  OAI21_X1 U18509 ( .B1(n15433), .B2(n16465), .A(n15264), .ZN(P2_U2985) );
  OR2_X1 U18510 ( .A1(n15265), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15266) );
  NAND2_X1 U18511 ( .A1(n12340), .A2(n15266), .ZN(n15445) );
  XNOR2_X1 U18512 ( .A(n15268), .B(n15267), .ZN(n15434) );
  NAND2_X1 U18513 ( .A1(n15434), .A2(n19397), .ZN(n15274) );
  NAND2_X1 U18514 ( .A1(n19198), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15435) );
  OAI21_X1 U18515 ( .B1(n19394), .B2(n15269), .A(n15435), .ZN(n15272) );
  NOR2_X1 U18516 ( .A1(n15270), .A2(n19405), .ZN(n15271) );
  AOI211_X1 U18517 ( .C1(n15438), .C2(n19399), .A(n15272), .B(n15271), .ZN(
        n15273) );
  OAI211_X1 U18518 ( .C1(n16463), .C2(n15445), .A(n15274), .B(n15273), .ZN(
        P2_U2987) );
  INV_X1 U18519 ( .A(n15284), .ZN(n15275) );
  OAI21_X1 U18520 ( .B1(n15286), .B2(n15285), .A(n15275), .ZN(n15276) );
  XOR2_X1 U18521 ( .A(n15277), .B(n15276), .Z(n15455) );
  AOI21_X1 U18522 ( .B1(n15446), .B2(n15278), .A(n15265), .ZN(n15453) );
  NOR2_X1 U18523 ( .A1(n19214), .A2(n20050), .ZN(n15448) );
  NOR2_X1 U18524 ( .A1(n16322), .A2(n16414), .ZN(n15279) );
  AOI211_X1 U18525 ( .C1(n16447), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15448), .B(n15279), .ZN(n15280) );
  OAI21_X1 U18526 ( .B1(n19405), .B2(n15281), .A(n15280), .ZN(n15282) );
  AOI21_X1 U18527 ( .B1(n15453), .B2(n19400), .A(n15282), .ZN(n15283) );
  OAI21_X1 U18528 ( .B1(n15455), .B2(n16465), .A(n15283), .ZN(P2_U2988) );
  NOR2_X1 U18529 ( .A1(n15285), .A2(n15284), .ZN(n15287) );
  XOR2_X1 U18530 ( .A(n15287), .B(n15286), .Z(n15468) );
  INV_X1 U18531 ( .A(n15278), .ZN(n15289) );
  AOI21_X1 U18532 ( .B1(n15456), .B2(n15288), .A(n15289), .ZN(n15466) );
  NAND2_X1 U18533 ( .A1(n15290), .A2(n16473), .ZN(n15292) );
  NOR2_X1 U18534 ( .A1(n19214), .A2(n20048), .ZN(n15460) );
  AOI21_X1 U18535 ( .B1(n16447), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15460), .ZN(n15291) );
  OAI211_X1 U18536 ( .C1(n15458), .C2(n16414), .A(n15292), .B(n15291), .ZN(
        n15293) );
  AOI21_X1 U18537 ( .B1(n15466), .B2(n19400), .A(n15293), .ZN(n15294) );
  OAI21_X1 U18538 ( .B1(n16465), .B2(n15468), .A(n15294), .ZN(P2_U2989) );
  AND2_X1 U18539 ( .A1(n15295), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15499) );
  OAI21_X1 U18540 ( .B1(n15499), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15296), .ZN(n15497) );
  OAI22_X1 U18541 ( .A1(n19394), .A2(n15297), .B1(n20044), .B2(n19214), .ZN(
        n15299) );
  NOR2_X1 U18542 ( .A1(n15492), .A2(n16414), .ZN(n15298) );
  AOI211_X1 U18543 ( .C1(n15300), .C2(n16473), .A(n15299), .B(n15298), .ZN(
        n15305) );
  OR2_X1 U18544 ( .A1(n15302), .A2(n15301), .ZN(n15494) );
  NAND3_X1 U18545 ( .A1(n15494), .A2(n15303), .A3(n19397), .ZN(n15304) );
  OAI211_X1 U18546 ( .C1(n15497), .C2(n16463), .A(n15305), .B(n15304), .ZN(
        P2_U2991) );
  INV_X1 U18547 ( .A(n16388), .ZN(n15306) );
  INV_X1 U18548 ( .A(n15379), .ZN(n15307) );
  INV_X1 U18549 ( .A(n15308), .ZN(n15369) );
  NAND2_X1 U18550 ( .A1(n15311), .A2(n15310), .ZN(n15363) );
  INV_X1 U18551 ( .A(n15311), .ZN(n15312) );
  INV_X1 U18552 ( .A(n15313), .ZN(n15351) );
  INV_X1 U18553 ( .A(n15327), .ZN(n15315) );
  INV_X1 U18554 ( .A(n15316), .ZN(n15318) );
  NAND2_X1 U18555 ( .A1(n15318), .A2(n15317), .ZN(n15319) );
  NAND2_X1 U18556 ( .A1(n15560), .A2(n15518), .ZN(n15331) );
  AOI21_X1 U18557 ( .B1(n15321), .B2(n15331), .A(n15295), .ZN(n15525) );
  NAND2_X1 U18558 ( .A1(n19198), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15522) );
  OAI21_X1 U18559 ( .B1(n19394), .B2(n15322), .A(n15522), .ZN(n15323) );
  AOI21_X1 U18560 ( .B1(n16473), .B2(n19099), .A(n15323), .ZN(n15324) );
  OAI21_X1 U18561 ( .B1(n16414), .B2(n19106), .A(n15324), .ZN(n15325) );
  AOI21_X1 U18562 ( .B1(n15525), .B2(n19400), .A(n15325), .ZN(n15326) );
  OAI21_X1 U18563 ( .B1(n15527), .B2(n16465), .A(n15326), .ZN(P2_U2993) );
  NAND2_X1 U18564 ( .A1(n15328), .A2(n15327), .ZN(n15330) );
  XOR2_X1 U18565 ( .A(n15330), .B(n15329), .Z(n15542) );
  INV_X1 U18566 ( .A(n15331), .ZN(n15333) );
  AOI21_X1 U18567 ( .B1(n15560), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15332) );
  NOR2_X1 U18568 ( .A1(n15333), .A2(n15332), .ZN(n15540) );
  NAND2_X1 U18569 ( .A1(n15181), .A2(n15334), .ZN(n15335) );
  NAND2_X1 U18570 ( .A1(n15336), .A2(n15335), .ZN(n19117) );
  NOR2_X1 U18571 ( .A1(n16414), .A2(n19117), .ZN(n15339) );
  NAND2_X1 U18572 ( .A1(n19198), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n15533) );
  NAND2_X1 U18573 ( .A1(n16447), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15337) );
  OAI211_X1 U18574 ( .C1(n19405), .C2(n19113), .A(n15533), .B(n15337), .ZN(
        n15338) );
  AOI211_X1 U18575 ( .C1(n15540), .C2(n19400), .A(n15339), .B(n15338), .ZN(
        n15340) );
  OAI21_X1 U18576 ( .B1(n15542), .B2(n16465), .A(n15340), .ZN(P2_U2994) );
  NAND2_X1 U18577 ( .A1(n15342), .A2(n15341), .ZN(n15346) );
  INV_X1 U18578 ( .A(n15343), .ZN(n15352) );
  NOR2_X1 U18579 ( .A1(n15344), .A2(n15352), .ZN(n15345) );
  XOR2_X1 U18580 ( .A(n15346), .B(n15345), .Z(n15553) );
  XNOR2_X1 U18581 ( .A(n15560), .B(n15549), .ZN(n15551) );
  NOR2_X1 U18582 ( .A1(n16414), .A2(n19130), .ZN(n15349) );
  NAND2_X1 U18583 ( .A1(n19198), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15544) );
  NAND2_X1 U18584 ( .A1(n16447), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15347) );
  OAI211_X1 U18585 ( .C1(n19131), .C2(n19405), .A(n15544), .B(n15347), .ZN(
        n15348) );
  AOI211_X1 U18586 ( .C1(n15551), .C2(n19400), .A(n15349), .B(n15348), .ZN(
        n15350) );
  OAI21_X1 U18587 ( .B1(n15553), .B2(n16465), .A(n15350), .ZN(P2_U2995) );
  NOR2_X1 U18588 ( .A1(n15352), .A2(n15351), .ZN(n15353) );
  XNOR2_X1 U18589 ( .A(n15354), .B(n15353), .ZN(n15567) );
  NOR2_X1 U18590 ( .A1(n19214), .A2(n15355), .ZN(n15558) );
  AOI21_X1 U18591 ( .B1(n16447), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15558), .ZN(n15356) );
  OAI21_X1 U18592 ( .B1(n16414), .B2(n16346), .A(n15356), .ZN(n15359) );
  INV_X1 U18593 ( .A(n15320), .ZN(n15357) );
  NOR2_X1 U18594 ( .A1(n15357), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15561) );
  NOR3_X1 U18595 ( .A1(n15561), .A2(n15560), .A3(n16463), .ZN(n15358) );
  AOI211_X1 U18596 ( .C1(n16473), .C2(n9770), .A(n15359), .B(n15358), .ZN(
        n15360) );
  OAI21_X1 U18597 ( .B1(n15567), .B2(n16465), .A(n15360), .ZN(P2_U2996) );
  AOI21_X1 U18598 ( .B1(n15363), .B2(n15362), .A(n15361), .ZN(n15585) );
  NAND2_X1 U18599 ( .A1(n19198), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15568) );
  NAND2_X1 U18600 ( .A1(n16447), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15364) );
  OAI211_X1 U18601 ( .C1(n19405), .C2(n19146), .A(n15568), .B(n15364), .ZN(
        n15365) );
  AOI21_X1 U18602 ( .B1(n19399), .B2(n19143), .A(n15365), .ZN(n15368) );
  NAND2_X1 U18603 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15571) );
  NOR2_X1 U18604 ( .A1(n16393), .A2(n15571), .ZN(n15577) );
  OAI211_X1 U18605 ( .C1(n15577), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n19400), .B(n15320), .ZN(n15367) );
  OAI211_X1 U18606 ( .C1(n15585), .C2(n16465), .A(n15368), .B(n15367), .ZN(
        P2_U2997) );
  XNOR2_X1 U18607 ( .A(n15370), .B(n15369), .ZN(n15595) );
  OAI22_X1 U18608 ( .A1(n19394), .A2(n15372), .B1(n19405), .B2(n15371), .ZN(
        n15374) );
  NOR2_X1 U18609 ( .A1(n19214), .A2(n20033), .ZN(n15373) );
  AOI211_X1 U18610 ( .C1(n19399), .C2(n15586), .A(n15374), .B(n15373), .ZN(
        n15378) );
  NOR2_X1 U18611 ( .A1(n16393), .A2(n15589), .ZN(n15376) );
  INV_X1 U18612 ( .A(n15577), .ZN(n15375) );
  OAI211_X1 U18613 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15376), .A(
        n15375), .B(n19400), .ZN(n15377) );
  OAI211_X1 U18614 ( .C1(n15595), .C2(n16465), .A(n15378), .B(n15377), .ZN(
        P2_U2998) );
  XNOR2_X1 U18615 ( .A(n16393), .B(n15589), .ZN(n15606) );
  NAND2_X1 U18616 ( .A1(n15380), .A2(n15379), .ZN(n15381) );
  XNOR2_X1 U18617 ( .A(n15382), .B(n15381), .ZN(n15596) );
  NAND2_X1 U18618 ( .A1(n15596), .A2(n19397), .ZN(n15388) );
  OAI22_X1 U18619 ( .A1(n19394), .A2(n15383), .B1(n19214), .B2(n20031), .ZN(
        n15386) );
  NOR2_X1 U18620 ( .A1(n19405), .A2(n15384), .ZN(n15385) );
  AOI211_X1 U18621 ( .C1(n15598), .C2(n19399), .A(n15386), .B(n15385), .ZN(
        n15387) );
  OAI211_X1 U18622 ( .C1(n15606), .C2(n16463), .A(n15388), .B(n15387), .ZN(
        P2_U2999) );
  XNOR2_X1 U18623 ( .A(n15390), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15391) );
  XNOR2_X1 U18624 ( .A(n15389), .B(n15391), .ZN(n16521) );
  NAND2_X1 U18625 ( .A1(n16473), .A2(n15392), .ZN(n15393) );
  NAND2_X1 U18626 ( .A1(n19198), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n16511) );
  OAI211_X1 U18627 ( .C1(n15394), .C2(n19394), .A(n15393), .B(n16511), .ZN(
        n15398) );
  NAND2_X1 U18628 ( .A1(n16450), .A2(n16452), .ZN(n15396) );
  XOR2_X1 U18629 ( .A(n15396), .B(n15395), .Z(n16516) );
  NOR2_X1 U18630 ( .A1(n16516), .A2(n16465), .ZN(n15397) );
  AOI211_X1 U18631 ( .C1(n19399), .C2(n16517), .A(n15398), .B(n15397), .ZN(
        n15399) );
  OAI21_X1 U18632 ( .B1(n16463), .B2(n16521), .A(n15399), .ZN(P2_U3007) );
  XNOR2_X1 U18633 ( .A(n15400), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15707) );
  XOR2_X1 U18634 ( .A(n15401), .B(n15402), .Z(n15694) );
  NOR2_X1 U18635 ( .A1(n15702), .A2(n16414), .ZN(n15405) );
  AOI22_X1 U18636 ( .A1(n16447), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n19198), .B2(P2_REIP_REG_6__SCAN_IN), .ZN(n15403) );
  OAI21_X1 U18637 ( .B1(n19205), .B2(n19405), .A(n15403), .ZN(n15404) );
  AOI211_X1 U18638 ( .C1(n15694), .C2(n19397), .A(n15405), .B(n15404), .ZN(
        n15406) );
  OAI21_X1 U18639 ( .B1(n15707), .B2(n16463), .A(n15406), .ZN(P2_U3008) );
  OAI211_X1 U18640 ( .C1(n15414), .C2(n11342), .A(n10246), .B(n10242), .ZN(
        n15415) );
  INV_X1 U18641 ( .A(n15415), .ZN(n15418) );
  OR2_X1 U18642 ( .A1(n15416), .A2(n16527), .ZN(n15417) );
  OAI211_X1 U18643 ( .C1(n15419), .C2(n16490), .A(n15418), .B(n15417), .ZN(
        P2_U3016) );
  OAI21_X1 U18644 ( .B1(n16522), .B2(n16317), .A(n15420), .ZN(n15429) );
  INV_X1 U18645 ( .A(n16309), .ZN(n15421) );
  OR2_X1 U18646 ( .A1(n15423), .A2(n15422), .ZN(n15425) );
  AOI21_X1 U18647 ( .B1(n15431), .B2(n10972), .A(n15430), .ZN(n15432) );
  OAI21_X1 U18648 ( .B1(n15433), .B2(n16490), .A(n15432), .ZN(P2_U3017) );
  NAND2_X1 U18649 ( .A1(n15434), .A2(n16530), .ZN(n15444) );
  OAI21_X1 U18650 ( .B1(n16522), .B2(n15436), .A(n15435), .ZN(n15437) );
  AOI21_X1 U18651 ( .B1(n15438), .B2(n16525), .A(n15437), .ZN(n15439) );
  OAI21_X1 U18652 ( .B1(n15440), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15439), .ZN(n15441) );
  AOI21_X1 U18653 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15442), .A(
        n15441), .ZN(n15443) );
  OAI211_X1 U18654 ( .C1(n15445), .C2(n16527), .A(n15444), .B(n15443), .ZN(
        P2_U3019) );
  NOR2_X1 U18655 ( .A1(n15457), .A2(n15446), .ZN(n15452) );
  XOR2_X1 U18656 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n15456), .Z(
        n15450) );
  NOR2_X1 U18657 ( .A1(n16322), .A2(n15710), .ZN(n15447) );
  AOI211_X1 U18658 ( .C1(n16502), .C2(n16320), .A(n15448), .B(n15447), .ZN(
        n15449) );
  OAI21_X1 U18659 ( .B1(n15463), .B2(n15450), .A(n15449), .ZN(n15451) );
  AOI211_X1 U18660 ( .C1(n15453), .C2(n10972), .A(n15452), .B(n15451), .ZN(
        n15454) );
  OAI21_X1 U18661 ( .B1(n15455), .B2(n16490), .A(n15454), .ZN(P2_U3020) );
  NOR2_X1 U18662 ( .A1(n15457), .A2(n15456), .ZN(n15465) );
  NOR2_X1 U18663 ( .A1(n15458), .A2(n15710), .ZN(n15459) );
  AOI211_X1 U18664 ( .C1(n16502), .C2(n15461), .A(n15460), .B(n15459), .ZN(
        n15462) );
  OAI21_X1 U18665 ( .B1(n15463), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15462), .ZN(n15464) );
  AOI211_X1 U18666 ( .C1(n15466), .C2(n10972), .A(n15465), .B(n15464), .ZN(
        n15467) );
  OAI21_X1 U18667 ( .B1(n16490), .B2(n15468), .A(n15467), .ZN(P2_U3021) );
  INV_X1 U18668 ( .A(n15469), .ZN(n15470) );
  OR2_X1 U18669 ( .A1(n15471), .A2(n15470), .ZN(n15472) );
  XNOR2_X1 U18670 ( .A(n15473), .B(n15472), .ZN(n16368) );
  NAND2_X1 U18671 ( .A1(n15296), .A2(n15474), .ZN(n15475) );
  NAND2_X1 U18672 ( .A1(n15288), .A2(n15475), .ZN(n16371) );
  OAI21_X1 U18673 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15477), .A(
        n15476), .ZN(n15482) );
  INV_X1 U18674 ( .A(n15478), .ZN(n16367) );
  NAND2_X1 U18675 ( .A1(n19198), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n16365) );
  OAI21_X1 U18676 ( .B1(n16522), .B2(n15479), .A(n16365), .ZN(n15480) );
  AOI21_X1 U18677 ( .B1(n16367), .B2(n16525), .A(n15480), .ZN(n15481) );
  OAI211_X1 U18678 ( .C1(n16371), .C2(n16527), .A(n15482), .B(n15481), .ZN(
        n15483) );
  AOI21_X1 U18679 ( .B1(n16530), .B2(n16368), .A(n15483), .ZN(n15484) );
  INV_X1 U18680 ( .A(n15484), .ZN(P2_U3022) );
  INV_X1 U18681 ( .A(n15520), .ZN(n15511) );
  AOI21_X1 U18682 ( .B1(n15486), .B2(n15485), .A(n15507), .ZN(n15488) );
  AOI22_X1 U18683 ( .A1(n15488), .A2(n15487), .B1(n19198), .B2(
        P2_REIP_REG_23__SCAN_IN), .ZN(n15491) );
  NAND2_X1 U18684 ( .A1(n16502), .A2(n15489), .ZN(n15490) );
  OAI211_X1 U18685 ( .C1(n15492), .C2(n15710), .A(n15491), .B(n15490), .ZN(
        n15493) );
  AOI21_X1 U18686 ( .B1(n15511), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15493), .ZN(n15496) );
  NAND3_X1 U18687 ( .A1(n15494), .A2(n15303), .A3(n16530), .ZN(n15495) );
  OAI211_X1 U18688 ( .C1(n15497), .C2(n16527), .A(n15496), .B(n15495), .ZN(
        P2_U3023) );
  NOR2_X1 U18689 ( .A1(n15295), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15498) );
  AND2_X1 U18690 ( .A1(n15501), .A2(n15500), .ZN(n15503) );
  OR2_X1 U18691 ( .A1(n15503), .A2(n15502), .ZN(n16340) );
  NOR2_X1 U18692 ( .A1(n15505), .A2(n15504), .ZN(n15506) );
  OR2_X1 U18693 ( .A1(n14982), .A2(n15506), .ZN(n15869) );
  INV_X1 U18694 ( .A(n15869), .ZN(n16348) );
  NAND2_X1 U18695 ( .A1(n19198), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n16376) );
  OAI21_X1 U18696 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15507), .A(
        n16376), .ZN(n15508) );
  AOI21_X1 U18697 ( .B1(n16502), .B2(n16348), .A(n15508), .ZN(n15509) );
  OAI21_X1 U18698 ( .B1(n16340), .B2(n15710), .A(n15509), .ZN(n15510) );
  AOI21_X1 U18699 ( .B1(n15511), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15510), .ZN(n15517) );
  NAND2_X1 U18700 ( .A1(n15513), .A2(n15512), .ZN(n15514) );
  XNOR2_X1 U18701 ( .A(n15515), .B(n15514), .ZN(n16378) );
  NAND2_X1 U18702 ( .A1(n16378), .A2(n16530), .ZN(n15516) );
  OAI211_X1 U18703 ( .C1(n16382), .C2(n16527), .A(n15517), .B(n15516), .ZN(
        P2_U3024) );
  AOI21_X1 U18704 ( .B1(n15547), .B2(n15518), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15519) );
  NOR2_X1 U18705 ( .A1(n15520), .A2(n15519), .ZN(n15524) );
  NAND2_X1 U18706 ( .A1(n16502), .A2(n19104), .ZN(n15521) );
  OAI211_X1 U18707 ( .C1(n15710), .C2(n19106), .A(n15522), .B(n15521), .ZN(
        n15523) );
  AOI211_X1 U18708 ( .C1(n15525), .C2(n10972), .A(n15524), .B(n15523), .ZN(
        n15526) );
  XNOR2_X1 U18709 ( .A(n15538), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15536) );
  AND2_X1 U18710 ( .A1(n15529), .A2(n15528), .ZN(n15531) );
  OR2_X1 U18711 ( .A1(n15531), .A2(n15530), .ZN(n16354) );
  INV_X1 U18712 ( .A(n19117), .ZN(n15532) );
  NAND2_X1 U18713 ( .A1(n15532), .A2(n16525), .ZN(n15534) );
  OAI211_X1 U18714 ( .C1(n16522), .C2(n16354), .A(n15534), .B(n15533), .ZN(
        n15535) );
  AOI21_X1 U18715 ( .B1(n15547), .B2(n15536), .A(n15535), .ZN(n15537) );
  OAI21_X1 U18716 ( .B1(n15554), .B2(n15538), .A(n15537), .ZN(n15539) );
  AOI21_X1 U18717 ( .B1(n15540), .B2(n10972), .A(n15539), .ZN(n15541) );
  OAI21_X1 U18718 ( .B1(n15542), .B2(n16490), .A(n15541), .ZN(P2_U3026) );
  INV_X1 U18719 ( .A(n19130), .ZN(n15543) );
  NAND2_X1 U18720 ( .A1(n16525), .A2(n15543), .ZN(n15545) );
  OAI211_X1 U18721 ( .C1(n16522), .C2(n19139), .A(n15545), .B(n15544), .ZN(
        n15546) );
  AOI21_X1 U18722 ( .B1(n15547), .B2(n15549), .A(n15546), .ZN(n15548) );
  OAI21_X1 U18723 ( .B1(n15554), .B2(n15549), .A(n15548), .ZN(n15550) );
  AOI21_X1 U18724 ( .B1(n15551), .B2(n10972), .A(n15550), .ZN(n15552) );
  OAI21_X1 U18725 ( .B1(n15553), .B2(n16490), .A(n15552), .ZN(P2_U3027) );
  INV_X1 U18726 ( .A(n15554), .ZN(n15565) );
  INV_X1 U18727 ( .A(n15692), .ZN(n15557) );
  OAI21_X1 U18728 ( .B1(n15557), .B2(n15556), .A(n15555), .ZN(n15564) );
  AOI21_X1 U18729 ( .B1(n16502), .B2(n16360), .A(n15558), .ZN(n15559) );
  OAI21_X1 U18730 ( .B1(n15710), .B2(n16346), .A(n15559), .ZN(n15563) );
  NOR3_X1 U18731 ( .A1(n15561), .A2(n15560), .A3(n16527), .ZN(n15562) );
  AOI211_X1 U18732 ( .C1(n15565), .C2(n15564), .A(n15563), .B(n15562), .ZN(
        n15566) );
  OAI21_X1 U18733 ( .B1(n15567), .B2(n16490), .A(n15566), .ZN(P2_U3028) );
  OAI21_X1 U18734 ( .B1(n15710), .B2(n15569), .A(n15568), .ZN(n15573) );
  INV_X1 U18735 ( .A(n15651), .ZN(n15570) );
  NAND2_X1 U18736 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15692), .ZN(
        n15668) );
  NOR2_X1 U18737 ( .A1(n15570), .A2(n15668), .ZN(n16494) );
  INV_X1 U18738 ( .A(n16494), .ZN(n15614) );
  NOR2_X1 U18739 ( .A1(n16493), .A2(n15614), .ZN(n15597) );
  AOI21_X1 U18740 ( .B1(n15366), .B2(n10972), .A(n15597), .ZN(n15590) );
  NOR3_X1 U18741 ( .A1(n15590), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15571), .ZN(n15572) );
  AOI211_X1 U18742 ( .C1(n16502), .C2(n15574), .A(n15573), .B(n15572), .ZN(
        n15584) );
  AND2_X1 U18743 ( .A1(n16527), .A2(n15575), .ZN(n15576) );
  OR2_X1 U18744 ( .A1(n15577), .A2(n15576), .ZN(n15580) );
  NAND2_X1 U18745 ( .A1(n15608), .A2(n15578), .ZN(n15579) );
  NAND2_X1 U18746 ( .A1(n15610), .A2(n15579), .ZN(n15601) );
  OAI211_X1 U18747 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15581), .A(
        n15580), .B(n15601), .ZN(n15593) );
  NOR2_X1 U18748 ( .A1(n16501), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15582) );
  OAI21_X1 U18749 ( .B1(n15593), .B2(n15582), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15583) );
  OAI211_X1 U18750 ( .C1(n15585), .C2(n16490), .A(n15584), .B(n15583), .ZN(
        P2_U3029) );
  INV_X1 U18751 ( .A(n19268), .ZN(n15588) );
  AOI22_X1 U18752 ( .A1(n16525), .A2(n15586), .B1(n19198), .B2(
        P2_REIP_REG_16__SCAN_IN), .ZN(n15587) );
  OAI21_X1 U18753 ( .B1(n15588), .B2(n16522), .A(n15587), .ZN(n15592) );
  NOR3_X1 U18754 ( .A1(n15590), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15589), .ZN(n15591) );
  AOI211_X1 U18755 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15593), .A(
        n15592), .B(n15591), .ZN(n15594) );
  OAI21_X1 U18756 ( .B1(n16490), .B2(n15595), .A(n15594), .ZN(P2_U3030) );
  NAND2_X1 U18757 ( .A1(n15596), .A2(n16530), .ZN(n15605) );
  INV_X1 U18758 ( .A(n19273), .ZN(n15603) );
  AOI22_X1 U18759 ( .A1(n15597), .A2(n15589), .B1(n19198), .B2(
        P2_REIP_REG_15__SCAN_IN), .ZN(n15600) );
  NAND2_X1 U18760 ( .A1(n16525), .A2(n15598), .ZN(n15599) );
  OAI211_X1 U18761 ( .C1(n15601), .C2(n15589), .A(n15600), .B(n15599), .ZN(
        n15602) );
  AOI21_X1 U18762 ( .B1(n15603), .B2(n16502), .A(n15602), .ZN(n15604) );
  OAI211_X1 U18763 ( .C1(n15606), .C2(n16527), .A(n15605), .B(n15604), .ZN(
        P2_U3031) );
  OR2_X1 U18764 ( .A1(n15607), .A2(n15635), .ZN(n16412) );
  XNOR2_X1 U18765 ( .A(n16412), .B(n16392), .ZN(n16405) );
  NAND2_X1 U18766 ( .A1(n15608), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15609) );
  NAND2_X1 U18767 ( .A1(n15610), .A2(n15609), .ZN(n15672) );
  OR2_X1 U18768 ( .A1(n16501), .A2(n15651), .ZN(n15611) );
  NAND2_X1 U18769 ( .A1(n15672), .A2(n15611), .ZN(n16485) );
  OR2_X1 U18770 ( .A1(n15612), .A2(n9762), .ZN(n15613) );
  NAND2_X1 U18771 ( .A1(n15613), .A2(n15029), .ZN(n19279) );
  NAND2_X1 U18772 ( .A1(n16525), .A2(n19165), .ZN(n15617) );
  AOI211_X1 U18773 ( .C1(n15635), .C2(n16392), .A(n16495), .B(n15614), .ZN(
        n15615) );
  AOI21_X1 U18774 ( .B1(n19198), .B2(P2_REIP_REG_13__SCAN_IN), .A(n15615), 
        .ZN(n15616) );
  OAI211_X1 U18775 ( .C1(n16522), .C2(n19279), .A(n15617), .B(n15616), .ZN(
        n15623) );
  NAND2_X1 U18776 ( .A1(n15620), .A2(n15619), .ZN(n15621) );
  XNOR2_X1 U18777 ( .A(n15618), .B(n15621), .ZN(n16404) );
  NOR2_X1 U18778 ( .A1(n16404), .A2(n16490), .ZN(n15622) );
  AOI211_X1 U18779 ( .C1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n16485), .A(
        n15623), .B(n15622), .ZN(n15624) );
  OAI21_X1 U18780 ( .B1(n16527), .B2(n16405), .A(n15624), .ZN(P2_U3033) );
  INV_X1 U18781 ( .A(n15626), .ZN(n15628) );
  NAND2_X1 U18782 ( .A1(n15628), .A2(n15627), .ZN(n15629) );
  XNOR2_X1 U18783 ( .A(n15625), .B(n15629), .ZN(n16416) );
  INV_X1 U18784 ( .A(n16416), .ZN(n15642) );
  NAND2_X1 U18785 ( .A1(n15607), .A2(n15635), .ZN(n16411) );
  NAND3_X1 U18786 ( .A1(n16412), .A2(n10972), .A3(n16411), .ZN(n15641) );
  XNOR2_X1 U18787 ( .A(n15630), .B(n15631), .ZN(n19281) );
  INV_X1 U18788 ( .A(n19281), .ZN(n15639) );
  OR2_X1 U18789 ( .A1(n15633), .A2(n15632), .ZN(n15634) );
  NAND2_X1 U18790 ( .A1(n15634), .A2(n13905), .ZN(n19245) );
  NAND2_X1 U18791 ( .A1(n16485), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15637) );
  AOI22_X1 U18792 ( .A1(n19198), .A2(P2_REIP_REG_12__SCAN_IN), .B1(n16494), 
        .B2(n15635), .ZN(n15636) );
  OAI211_X1 U18793 ( .C1(n19245), .C2(n15710), .A(n15637), .B(n15636), .ZN(
        n15638) );
  AOI21_X1 U18794 ( .B1(n15639), .B2(n16502), .A(n15638), .ZN(n15640) );
  OAI211_X1 U18795 ( .C1(n15642), .C2(n16490), .A(n15641), .B(n15640), .ZN(
        P2_U3034) );
  INV_X1 U18796 ( .A(n15643), .ZN(n15644) );
  NAND2_X1 U18797 ( .A1(n15645), .A2(n15644), .ZN(n15649) );
  NOR2_X1 U18798 ( .A1(n15647), .A2(n15646), .ZN(n15648) );
  XNOR2_X1 U18799 ( .A(n15649), .B(n15648), .ZN(n16421) );
  OAI21_X1 U18800 ( .B1(n15044), .B2(n15650), .A(n15630), .ZN(n19283) );
  INV_X1 U18801 ( .A(n19283), .ZN(n15660) );
  NAND2_X1 U18802 ( .A1(n19198), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n16419) );
  AOI211_X1 U18803 ( .C1(n15656), .C2(n15674), .A(n15651), .B(n15668), .ZN(
        n15652) );
  INV_X1 U18804 ( .A(n15652), .ZN(n15653) );
  NAND2_X1 U18805 ( .A1(n16419), .A2(n15653), .ZN(n15654) );
  AOI21_X1 U18806 ( .B1(n16525), .B2(n19194), .A(n15654), .ZN(n15655) );
  OAI21_X1 U18807 ( .B1(n15672), .B2(n15656), .A(n15655), .ZN(n15659) );
  OAI21_X1 U18808 ( .B1(n15657), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15607), .ZN(n16422) );
  NOR2_X1 U18809 ( .A1(n16422), .A2(n16527), .ZN(n15658) );
  AOI211_X1 U18810 ( .C1(n16502), .C2(n15660), .A(n15659), .B(n15658), .ZN(
        n15661) );
  OAI21_X1 U18811 ( .B1(n16421), .B2(n16490), .A(n15661), .ZN(P2_U3035) );
  INV_X1 U18812 ( .A(n15662), .ZN(n15679) );
  OR2_X1 U18813 ( .A1(n15663), .A2(n15679), .ZN(n15667) );
  NAND2_X1 U18814 ( .A1(n15665), .A2(n15664), .ZN(n15666) );
  XNOR2_X1 U18815 ( .A(n15667), .B(n15666), .ZN(n16428) );
  NAND2_X1 U18816 ( .A1(n19198), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n16426) );
  OAI21_X1 U18817 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n15668), .A(
        n16426), .ZN(n15669) );
  AOI21_X1 U18818 ( .B1(n16502), .B2(n19284), .A(n15669), .ZN(n15671) );
  NAND2_X1 U18819 ( .A1(n16525), .A2(n19250), .ZN(n15670) );
  OAI211_X1 U18820 ( .C1(n15672), .C2(n15674), .A(n15671), .B(n15670), .ZN(
        n15677) );
  AND2_X1 U18821 ( .A1(n15673), .A2(n15674), .ZN(n15675) );
  OR2_X1 U18822 ( .A1(n15657), .A2(n15675), .ZN(n16431) );
  NOR2_X1 U18823 ( .A1(n16431), .A2(n16527), .ZN(n15676) );
  AOI211_X1 U18824 ( .C1(n16530), .C2(n16428), .A(n15677), .B(n15676), .ZN(
        n15678) );
  INV_X1 U18825 ( .A(n15678), .ZN(P2_U3036) );
  OR2_X1 U18826 ( .A1(n15680), .A2(n15679), .ZN(n15681) );
  XNOR2_X1 U18827 ( .A(n15682), .B(n15681), .ZN(n16439) );
  INV_X1 U18828 ( .A(n16442), .ZN(n15687) );
  NAND2_X1 U18829 ( .A1(n15683), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15686) );
  OAI22_X1 U18830 ( .A1(n16522), .A2(n19288), .B1(n16436), .B2(n19214), .ZN(
        n15684) );
  INV_X1 U18831 ( .A(n15684), .ZN(n15685) );
  OAI211_X1 U18832 ( .C1(n15710), .C2(n15687), .A(n15686), .B(n15685), .ZN(
        n15690) );
  OAI21_X1 U18833 ( .B1(n15688), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15673), .ZN(n16440) );
  NOR2_X1 U18834 ( .A1(n16440), .A2(n16527), .ZN(n15689) );
  AOI211_X1 U18835 ( .C1(n15692), .C2(n15691), .A(n15690), .B(n15689), .ZN(
        n15693) );
  OAI21_X1 U18836 ( .B1(n16490), .B2(n16439), .A(n15693), .ZN(P2_U3037) );
  NAND2_X1 U18837 ( .A1(n15694), .A2(n16530), .ZN(n15706) );
  OAI21_X1 U18838 ( .B1(n16501), .B2(n15697), .A(n16533), .ZN(n15704) );
  NAND3_X1 U18839 ( .A1(n15697), .A2(n15696), .A3(n15695), .ZN(n15701) );
  XNOR2_X1 U18840 ( .A(n15698), .B(n15699), .ZN(n19294) );
  INV_X1 U18841 ( .A(n19294), .ZN(n19208) );
  AOI22_X1 U18842 ( .A1(n16502), .A2(n19208), .B1(n19198), .B2(
        P2_REIP_REG_6__SCAN_IN), .ZN(n15700) );
  OAI211_X1 U18843 ( .C1(n15710), .C2(n15702), .A(n15701), .B(n15700), .ZN(
        n15703) );
  AOI21_X1 U18844 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15704), .A(
        n15703), .ZN(n15705) );
  OAI211_X1 U18845 ( .C1(n15707), .C2(n16527), .A(n15706), .B(n15705), .ZN(
        P2_U3040) );
  OAI21_X1 U18846 ( .B1(n15710), .B2(n15709), .A(n15708), .ZN(n15711) );
  AOI21_X1 U18847 ( .B1(n16502), .B2(n15712), .A(n15711), .ZN(n15719) );
  INV_X1 U18848 ( .A(n15713), .ZN(n15715) );
  AOI22_X1 U18849 ( .A1(n10972), .A2(n15715), .B1(n16530), .B2(n15714), .ZN(
        n15718) );
  MUX2_X1 U18850 ( .A(n16501), .B(n15716), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n15717) );
  NAND3_X1 U18851 ( .A1(n15719), .A2(n15718), .A3(n15717), .ZN(P2_U3046) );
  MUX2_X1 U18852 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n15720), .S(
        n13426), .Z(n15725) );
  AOI22_X1 U18853 ( .A1(n15722), .A2(n16543), .B1(n15733), .B2(n15721), .ZN(
        n15723) );
  OAI21_X1 U18854 ( .B1(n15725), .B2(n11320), .A(n15723), .ZN(n15724) );
  MUX2_X1 U18855 ( .A(n15724), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n15737), .Z(P2_U3601) );
  NAND2_X1 U18856 ( .A1(n15725), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n15736) );
  OR2_X1 U18857 ( .A1(n13426), .A2(n13550), .ZN(n15726) );
  NAND2_X1 U18858 ( .A1(n15727), .A2(n15726), .ZN(n15731) );
  AOI22_X1 U18859 ( .A1(n20094), .A2(n16543), .B1(n15733), .B2(n15728), .ZN(
        n15729) );
  OAI21_X1 U18860 ( .B1(n15736), .B2(n15731), .A(n15729), .ZN(n15730) );
  MUX2_X1 U18861 ( .A(n15730), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n15737), .Z(P2_U3600) );
  INV_X1 U18862 ( .A(n15731), .ZN(n15735) );
  AOI22_X1 U18863 ( .A1(n19540), .A2(n16543), .B1(n15733), .B2(n15732), .ZN(
        n15734) );
  OAI21_X1 U18864 ( .B1(n15736), .B2(n15735), .A(n15734), .ZN(n15738) );
  MUX2_X1 U18865 ( .A(n15738), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15737), .Z(P2_U3599) );
  AOI22_X1 U18866 ( .A1(n17356), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17381), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15739) );
  OAI21_X1 U18867 ( .B1(n12918), .B2(n17418), .A(n15739), .ZN(n15749) );
  AOI22_X1 U18868 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17320), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15746) );
  OAI22_X1 U18869 ( .A1(n17367), .A2(n17205), .B1(n17358), .B2(n17302), .ZN(
        n15744) );
  AOI22_X1 U18870 ( .A1(n12945), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15742) );
  AOI22_X1 U18871 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15741) );
  AOI22_X1 U18872 ( .A1(n17321), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13039), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15740) );
  NAND3_X1 U18873 ( .A1(n15742), .A2(n15741), .A3(n15740), .ZN(n15743) );
  AOI211_X1 U18874 ( .C1(n17384), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n15744), .B(n15743), .ZN(n15745) );
  OAI211_X1 U18875 ( .C1(n17303), .C2(n15747), .A(n15746), .B(n15745), .ZN(
        n15748) );
  AOI211_X1 U18876 ( .C1(n17306), .C2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A(
        n15749), .B(n15748), .ZN(n17144) );
  AOI22_X1 U18877 ( .A1(n17381), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15750) );
  OAI21_X1 U18878 ( .B1(n12918), .B2(n17424), .A(n15750), .ZN(n15760) );
  AOI22_X1 U18879 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9665), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15758) );
  AOI22_X1 U18880 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15751) );
  OAI21_X1 U18881 ( .B1(n17358), .B2(n17232), .A(n15751), .ZN(n15756) );
  AOI22_X1 U18882 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12945), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15753) );
  AOI22_X1 U18883 ( .A1(n17356), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15752) );
  OAI211_X1 U18884 ( .C1(n17380), .C2(n15754), .A(n15753), .B(n15752), .ZN(
        n15755) );
  AOI211_X1 U18885 ( .C1(n17374), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n15756), .B(n15755), .ZN(n15757) );
  OAI211_X1 U18886 ( .C1(n17287), .C2(n17348), .A(n15758), .B(n15757), .ZN(
        n15759) );
  AOI211_X1 U18887 ( .C1(n17306), .C2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A(
        n15760), .B(n15759), .ZN(n17155) );
  AOI22_X1 U18888 ( .A1(n17356), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17352), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15761) );
  OAI21_X1 U18889 ( .B1(n14414), .B2(n17395), .A(n15761), .ZN(n15772) );
  AOI22_X1 U18890 ( .A1(n13117), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15769) );
  OAI22_X1 U18891 ( .A1(n17120), .A2(n15762), .B1(n17380), .B2(n17267), .ZN(
        n15767) );
  AOI22_X1 U18892 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15765) );
  AOI22_X1 U18893 ( .A1(n13080), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12945), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15764) );
  AOI22_X1 U18894 ( .A1(n13039), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17392), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15763) );
  NAND3_X1 U18895 ( .A1(n15765), .A2(n15764), .A3(n15763), .ZN(n15766) );
  AOI211_X1 U18896 ( .C1(n9653), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n15767), .B(n15766), .ZN(n15768) );
  OAI211_X1 U18897 ( .C1(n17287), .C2(n15770), .A(n15769), .B(n15768), .ZN(
        n15771) );
  AOI211_X1 U18898 ( .C1(n17306), .C2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A(
        n15772), .B(n15771), .ZN(n17165) );
  AOI22_X1 U18899 ( .A1(n13117), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15773) );
  OAI21_X1 U18900 ( .B1(n12928), .B2(n17119), .A(n15773), .ZN(n15783) );
  AOI22_X1 U18901 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15781) );
  AOI22_X1 U18902 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15774) );
  INV_X1 U18903 ( .A(n15774), .ZN(n15779) );
  AOI22_X1 U18904 ( .A1(n12945), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15777) );
  AOI22_X1 U18905 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15776) );
  AOI22_X1 U18906 ( .A1(n13039), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17392), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15775) );
  NAND3_X1 U18907 ( .A1(n15777), .A2(n15776), .A3(n15775), .ZN(n15778) );
  AOI211_X1 U18908 ( .C1(n17321), .C2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n15779), .B(n15778), .ZN(n15780) );
  OAI211_X1 U18909 ( .C1(n17367), .C2(n17406), .A(n15781), .B(n15780), .ZN(
        n15782) );
  AOI211_X1 U18910 ( .C1(n17306), .C2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A(
        n15783), .B(n15782), .ZN(n17166) );
  NOR2_X1 U18911 ( .A1(n17165), .A2(n17166), .ZN(n17164) );
  AOI22_X1 U18912 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17356), .B1(
        n17375), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15794) );
  AOI22_X1 U18913 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17384), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n14415), .ZN(n15793) );
  AOI22_X1 U18914 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n17392), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17321), .ZN(n15792) );
  OAI22_X1 U18915 ( .A1(n17396), .A2(n17247), .B1(n15784), .B2(n17354), .ZN(
        n15790) );
  AOI22_X1 U18916 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17382), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15788) );
  AOI22_X1 U18917 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n17376), .ZN(n15787) );
  AOI22_X1 U18918 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17352), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15786) );
  NAND2_X1 U18919 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n13039), .ZN(
        n15785) );
  NAND4_X1 U18920 ( .A1(n15788), .A2(n15787), .A3(n15786), .A4(n15785), .ZN(
        n15789) );
  AOI211_X1 U18921 ( .C1(n17320), .C2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A(
        n15790), .B(n15789), .ZN(n15791) );
  NAND4_X1 U18922 ( .A1(n15794), .A2(n15793), .A3(n15792), .A4(n15791), .ZN(
        n17160) );
  NAND2_X1 U18923 ( .A1(n17164), .A2(n17160), .ZN(n17159) );
  NOR2_X1 U18924 ( .A1(n17155), .A2(n17159), .ZN(n17154) );
  AOI22_X1 U18925 ( .A1(n17384), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17306), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15804) );
  AOI22_X1 U18926 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15796) );
  AOI22_X1 U18927 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17352), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15795) );
  OAI211_X1 U18928 ( .C1(n17380), .C2(n17218), .A(n15796), .B(n15795), .ZN(
        n15802) );
  AOI22_X1 U18929 ( .A1(n12945), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15800) );
  AOI22_X1 U18930 ( .A1(n13117), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15799) );
  AOI22_X1 U18931 ( .A1(n12938), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15798) );
  NAND2_X1 U18932 ( .A1(n17392), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n15797) );
  NAND4_X1 U18933 ( .A1(n15800), .A2(n15799), .A3(n15798), .A4(n15797), .ZN(
        n15801) );
  AOI211_X1 U18934 ( .C1(n17374), .C2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n15802), .B(n15801), .ZN(n15803) );
  OAI211_X1 U18935 ( .C1(n17287), .C2(n17330), .A(n15804), .B(n15803), .ZN(
        n17150) );
  NAND2_X1 U18936 ( .A1(n17154), .A2(n17150), .ZN(n17149) );
  NOR2_X1 U18937 ( .A1(n17144), .A2(n17149), .ZN(n17143) );
  AOI22_X1 U18938 ( .A1(n12945), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15815) );
  AOI22_X1 U18939 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17375), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15806) );
  AOI22_X1 U18940 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15805) );
  OAI211_X1 U18941 ( .C1(n17380), .C2(n15807), .A(n15806), .B(n15805), .ZN(
        n15813) );
  AOI22_X1 U18942 ( .A1(n17356), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17352), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15811) );
  AOI22_X1 U18943 ( .A1(n17384), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15810) );
  AOI22_X1 U18944 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15809) );
  NAND2_X1 U18945 ( .A1(n17374), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n15808) );
  NAND4_X1 U18946 ( .A1(n15811), .A2(n15810), .A3(n15809), .A4(n15808), .ZN(
        n15812) );
  AOI211_X1 U18947 ( .C1(n17392), .C2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n15813), .B(n15812), .ZN(n15814) );
  OAI211_X1 U18948 ( .C1(n17287), .C2(n15825), .A(n15815), .B(n15814), .ZN(
        n15816) );
  NAND2_X1 U18949 ( .A1(n17143), .A2(n15816), .ZN(n17136) );
  OAI21_X1 U18950 ( .B1(n17143), .B2(n15816), .A(n17136), .ZN(n17459) );
  AND2_X1 U18951 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17140) );
  NOR2_X1 U18952 ( .A1(n18449), .A2(n17263), .ZN(n17431) );
  INV_X1 U18953 ( .A(n17431), .ZN(n17429) );
  INV_X1 U18954 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17099) );
  INV_X1 U18955 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16806) );
  INV_X1 U18956 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16836) );
  INV_X1 U18957 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n16867) );
  INV_X1 U18958 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17260) );
  NAND4_X1 U18959 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .A4(P3_EBX_REG_4__SCAN_IN), .ZN(n15819) );
  NAND4_X1 U18960 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(P3_EBX_REG_11__SCAN_IN), .A4(P3_EBX_REG_10__SCAN_IN), .ZN(n15818)
         );
  INV_X1 U18961 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17404) );
  INV_X1 U18962 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17403) );
  NOR2_X1 U18963 ( .A1(n17404), .A2(n17403), .ZN(n17398) );
  NAND4_X1 U18964 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_15__SCAN_IN), 
        .A3(P3_EBX_REG_13__SCAN_IN), .A4(n17398), .ZN(n15817) );
  NOR4_X1 U18965 ( .A1(n15820), .A2(n15819), .A3(n15818), .A4(n15817), .ZN(
        n17261) );
  INV_X1 U18966 ( .A(n17261), .ZN(n17262) );
  NAND2_X1 U18967 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17246), .ZN(n17229) );
  INV_X1 U18968 ( .A(n17229), .ZN(n17202) );
  NAND2_X1 U18969 ( .A1(n17527), .A2(n17216), .ZN(n17201) );
  NAND2_X1 U18970 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17170), .ZN(n17163) );
  NAND2_X1 U18971 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17169), .ZN(n17153) );
  NAND2_X1 U18972 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17158), .ZN(n17148) );
  NAND2_X1 U18973 ( .A1(n17423), .A2(n17148), .ZN(n17146) );
  OAI21_X1 U18974 ( .B1(n17140), .B2(n17429), .A(n17146), .ZN(n17138) );
  INV_X1 U18975 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17147) );
  NOR3_X1 U18976 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17147), .A3(n17148), .ZN(
        n15821) );
  AOI21_X1 U18977 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17138), .A(n15821), .ZN(
        n15822) );
  OAI21_X1 U18978 ( .B1(n17459), .B2(n17423), .A(n15822), .ZN(P3_U2675) );
  INV_X1 U18979 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17190) );
  AOI22_X1 U18980 ( .A1(n17376), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15823) );
  OAI21_X1 U18981 ( .B1(n17396), .B2(n17190), .A(n15823), .ZN(n15835) );
  AOI22_X1 U18982 ( .A1(n9665), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17320), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15831) );
  AOI22_X1 U18983 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17374), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15824) );
  OAI21_X1 U18984 ( .B1(n12928), .B2(n15825), .A(n15824), .ZN(n15829) );
  INV_X1 U18985 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17414) );
  AOI22_X1 U18986 ( .A1(n12945), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15827) );
  AOI22_X1 U18987 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15826) );
  OAI211_X1 U18988 ( .C1(n17380), .C2(n17414), .A(n15827), .B(n15826), .ZN(
        n15828) );
  AOI211_X1 U18989 ( .C1(n17392), .C2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n15829), .B(n15828), .ZN(n15830) );
  OAI211_X1 U18990 ( .C1(n15833), .C2(n15832), .A(n15831), .B(n15830), .ZN(
        n15834) );
  AOI211_X1 U18991 ( .C1(n17336), .C2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n15835), .B(n15834), .ZN(n17536) );
  OAI21_X1 U18992 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17317), .A(n15836), .ZN(
        n15837) );
  AOI22_X1 U18993 ( .A1(n17432), .A2(n17536), .B1(n15837), .B2(n17423), .ZN(
        P3_U2690) );
  NOR2_X1 U18994 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19008), .ZN(
        n18458) );
  INV_X1 U18995 ( .A(n18458), .ZN(n15838) );
  NAND3_X1 U18996 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n19006)
         );
  AOI211_X1 U18997 ( .C1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(n18850), .A(
        n9653), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18402) );
  NOR2_X1 U18998 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19062) );
  AOI21_X1 U18999 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n19062), .ZN(n18914) );
  INV_X1 U19000 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n16697) );
  OR2_X1 U19001 ( .A1(n16697), .A2(n19006), .ZN(n15851) );
  OAI211_X1 U19002 ( .C1(n19006), .C2(n18402), .A(n18525), .B(n15851), .ZN(
        n18408) );
  NAND2_X1 U19003 ( .A1(n15838), .A2(n18408), .ZN(n15841) );
  INV_X1 U19004 ( .A(n15841), .ZN(n15840) );
  NAND3_X1 U19005 ( .A1(n19056), .A2(n19008), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18755) );
  NAND2_X1 U19006 ( .A1(n19056), .A2(n19008), .ZN(n16692) );
  AND2_X1 U19007 ( .A1(n19009), .A2(n16692), .ZN(n19053) );
  INV_X1 U19008 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16716) );
  NOR2_X1 U19009 ( .A1(n19018), .A2(n16716), .ZN(n18041) );
  OAI22_X1 U19010 ( .A1(n19053), .A2(n18041), .B1(n18414), .B2(n19008), .ZN(
        n15843) );
  NAND3_X1 U19011 ( .A1(n18864), .A2(n18408), .A3(n15843), .ZN(n15839) );
  OAI221_X1 U19012 ( .B1(n18864), .B2(n15840), .C1(n18864), .C2(n18755), .A(
        n15839), .ZN(P3_U2864) );
  NAND2_X1 U19013 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18589) );
  NOR2_X1 U19014 ( .A1(n19053), .A2(n18041), .ZN(n15842) );
  AOI221_X1 U19015 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18589), .C1(n15842), 
        .C2(n18589), .A(n15841), .ZN(n18407) );
  INV_X1 U19016 ( .A(n18755), .ZN(n18706) );
  OAI221_X1 U19017 ( .B1(n18706), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18706), .C2(n15843), .A(n18408), .ZN(n18405) );
  AOI22_X1 U19018 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18407), .B1(
        n18405), .B2(n18884), .ZN(P3_U2865) );
  NAND2_X1 U19019 ( .A1(n16690), .A2(n19050), .ZN(n15850) );
  NAND2_X1 U19020 ( .A1(n17658), .A2(n9661), .ZN(n18896) );
  NAND2_X1 U19021 ( .A1(n9970), .A2(n18896), .ZN(n15844) );
  INV_X1 U19022 ( .A(n16690), .ZN(n18841) );
  INV_X1 U19023 ( .A(n18872), .ZN(n15846) );
  NOR3_X1 U19024 ( .A1(n15941), .A2(n15848), .A3(n15847), .ZN(n15849) );
  NAND2_X1 U19025 ( .A1(n19059), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18409) );
  INV_X1 U19026 ( .A(n19009), .ZN(n19034) );
  AOI21_X1 U19027 ( .B1(n18850), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15853) );
  NOR2_X1 U19028 ( .A1(n15853), .A2(n15852), .ZN(n18894) );
  NAND3_X1 U19029 ( .A1(n19036), .A2(n19034), .A3(n18894), .ZN(n15854) );
  OAI21_X1 U19030 ( .B1(n19036), .B2(n18849), .A(n15854), .ZN(P3_U3284) );
  OAI22_X1 U19031 ( .A1(n16587), .A2(n18391), .B1(n16584), .B2(n18319), .ZN(
        n15855) );
  NOR2_X1 U19032 ( .A1(n15856), .A2(n15855), .ZN(n15919) );
  AOI211_X1 U19033 ( .C1(n18309), .C2(n15858), .A(n18386), .B(n15857), .ZN(
        n15860) );
  AOI22_X1 U19034 ( .A1(n15859), .A2(n16566), .B1(n18397), .B2(n16567), .ZN(
        n15923) );
  OAI21_X1 U19035 ( .B1(n18393), .B2(n15860), .A(n15923), .ZN(n15864) );
  NOR2_X1 U19036 ( .A1(n15862), .A2(n15861), .ZN(n15863) );
  XOR2_X1 U19037 ( .A(n15863), .B(n16586), .Z(n16590) );
  AOI22_X1 U19038 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15864), .B1(
        n18315), .B2(n16590), .ZN(n15865) );
  NAND2_X1 U19039 ( .A1(n18393), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16595) );
  OAI211_X1 U19040 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15919), .A(
        n15865), .B(n16595), .ZN(P3_U2833) );
  AOI22_X1 U19041 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19221), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19199), .ZN(n15876) );
  INV_X1 U19042 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15866) );
  OAI22_X1 U19043 ( .A1(n15867), .A2(n19216), .B1(n19218), .B2(n15866), .ZN(
        n15868) );
  INV_X1 U19044 ( .A(n15868), .ZN(n15875) );
  OAI22_X1 U19045 ( .A1(n16340), .A2(n19129), .B1(n15869), .B2(n19231), .ZN(
        n15870) );
  INV_X1 U19046 ( .A(n15870), .ZN(n15874) );
  NAND3_X1 U19047 ( .A1(n19100), .A2(n15871), .A3(n13426), .ZN(n15872) );
  NAND3_X1 U19048 ( .A1(n10086), .A2(n19227), .A3(n15872), .ZN(n15873) );
  NAND4_X1 U19049 ( .A1(n15876), .A2(n15875), .A3(n15874), .A4(n15873), .ZN(
        P2_U2833) );
  OAI22_X1 U19050 ( .A1(n15879), .A2(n15878), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15877), .ZN(n20949) );
  NAND2_X1 U19051 ( .A1(n15880), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n20957) );
  INV_X1 U19052 ( .A(n20957), .ZN(n15881) );
  NOR3_X1 U19053 ( .A1(n20949), .A2(n15881), .A3(n20751), .ZN(n15885) );
  NAND2_X1 U19054 ( .A1(n15885), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n15887) );
  INV_X1 U19055 ( .A(n15882), .ZN(n15883) );
  OAI22_X1 U19056 ( .A1(n15885), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n15884), .B2(n15883), .ZN(n15886) );
  NAND2_X1 U19057 ( .A1(n15887), .A2(n15886), .ZN(n15892) );
  INV_X1 U19058 ( .A(n15888), .ZN(n15890) );
  NAND2_X1 U19059 ( .A1(n15890), .A2(n15889), .ZN(n15891) );
  AOI222_X1 U19060 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n15892), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15891), .C1(n15892), 
        .C2(n15891), .ZN(n15893) );
  AOI222_X1 U19061 ( .A1(n20710), .A2(n15894), .B1(n20710), .B2(n15893), .C1(
        n15894), .C2(n15893), .ZN(n15902) );
  INV_X1 U19062 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n21056) );
  AOI21_X1 U19063 ( .B1(n21056), .B2(n21100), .A(n15895), .ZN(n15897) );
  NOR4_X1 U19064 ( .A1(n15899), .A2(n15898), .A3(n15897), .A4(n15896), .ZN(
        n15901) );
  OAI211_X1 U19065 ( .C1(n15902), .C2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n15901), .B(n15900), .ZN(n15903) );
  INV_X1 U19066 ( .A(n15903), .ZN(n15915) );
  AOI21_X1 U19067 ( .B1(n11516), .B2(n20892), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n16293) );
  NAND2_X1 U19068 ( .A1(n20892), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n16287) );
  INV_X1 U19069 ( .A(n15904), .ZN(n15907) );
  INV_X1 U19070 ( .A(n16287), .ZN(n20975) );
  INV_X1 U19071 ( .A(n15913), .ZN(n15905) );
  NOR2_X1 U19072 ( .A1(n15905), .A2(n20976), .ZN(n20883) );
  AOI211_X1 U19073 ( .C1(n15907), .C2(n15906), .A(n20975), .B(n20883), .ZN(
        n16290) );
  OAI221_X1 U19074 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n15915), 
        .A(n16290), .ZN(n15910) );
  NAND2_X1 U19075 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15910), .ZN(n16294) );
  AOI211_X1 U19076 ( .C1(n16293), .C2(n16287), .A(n15908), .B(n16294), .ZN(
        n15914) );
  AOI221_X1 U19077 ( .B1(n15911), .B2(n15910), .C1(n15909), .C2(n15910), .A(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n15912) );
  AOI221_X1 U19078 ( .B1(n15915), .B2(n15914), .C1(n15913), .C2(n15914), .A(
        n15912), .ZN(P1_U3161) );
  NAND2_X1 U19079 ( .A1(n15917), .A2(n15916), .ZN(n15918) );
  INV_X1 U19080 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18995) );
  NOR2_X1 U19081 ( .A1(n18380), .A2(n18995), .ZN(n16570) );
  NOR3_X1 U19082 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15919), .A3(
        n16586), .ZN(n15920) );
  AOI211_X1 U19083 ( .C1(n18315), .C2(n16577), .A(n16570), .B(n15920), .ZN(
        n15921) );
  OAI221_X1 U19084 ( .B1(n16579), .B2(n15923), .C1(n16579), .C2(n15922), .A(
        n15921), .ZN(P3_U2832) );
  INV_X1 U19085 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20885) );
  INV_X1 U19086 ( .A(HOLD), .ZN(n21115) );
  NOR2_X1 U19087 ( .A1(n20885), .A2(n21115), .ZN(n20888) );
  AOI22_X1 U19088 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n15926) );
  NAND2_X1 U19089 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n15924), .ZN(n20895) );
  OAI211_X1 U19090 ( .C1(n20888), .C2(n15926), .A(n15925), .B(n20895), .ZN(
        P1_U3195) );
  AND2_X1 U19091 ( .A1(n20218), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  INV_X1 U19092 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15934) );
  AOI211_X1 U19093 ( .C1(n15934), .C2(n11766), .A(n16273), .B(n16155), .ZN(
        n15932) );
  OR2_X1 U19094 ( .A1(n15927), .A2(n15934), .ZN(n15928) );
  OAI22_X1 U19095 ( .A1(n16068), .A2(n16225), .B1(n20288), .B2(n15995), .ZN(
        n15930) );
  AOI21_X1 U19096 ( .B1(n15932), .B2(n15931), .A(n15930), .ZN(n15933) );
  NAND2_X1 U19097 ( .A1(n20290), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n16072) );
  OAI211_X1 U19098 ( .C1(n16156), .C2(n15934), .A(n15933), .B(n16072), .ZN(
        P1_U3011) );
  AOI21_X1 U19099 ( .B1(n16540), .B2(n15936), .A(n15935), .ZN(n15937) );
  OR2_X1 U19100 ( .A1(n19936), .A2(n15937), .ZN(n20105) );
  NOR2_X1 U19101 ( .A1(n15938), .A2(n20105), .ZN(P2_U3047) );
  OAI21_X1 U19102 ( .B1(n15941), .B2(n15940), .A(n19054), .ZN(n15942) );
  NAND2_X1 U19104 ( .A1(n17527), .A2(n17593), .ZN(n17589) );
  INV_X1 U19105 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17655) );
  NOR2_X1 U19106 ( .A1(n17577), .A2(n18858), .ZN(n17587) );
  NOR2_X2 U19107 ( .A1(n15943), .A2(n15942), .ZN(n17586) );
  OAI221_X1 U19108 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17589), .C1(n17655), 
        .C2(n17593), .A(n15944), .ZN(P3_U2735) );
  INV_X1 U19109 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21055) );
  AOI21_X1 U19110 ( .B1(n20146), .B2(n21055), .A(n15957), .ZN(n15956) );
  NAND2_X1 U19111 ( .A1(n15945), .A2(n21116), .ZN(n15950) );
  NAND2_X1 U19112 ( .A1(n20173), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n15949) );
  INV_X1 U19113 ( .A(n15946), .ZN(n15947) );
  AOI22_X1 U19114 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n20186), .B1(
        n20171), .B2(n15947), .ZN(n15948) );
  OAI211_X1 U19115 ( .C1(n15950), .C2(n20175), .A(n15949), .B(n15948), .ZN(
        n15951) );
  INV_X1 U19116 ( .A(n15951), .ZN(n15955) );
  AOI22_X1 U19117 ( .A1(n15953), .A2(n20165), .B1(n15952), .B2(n20196), .ZN(
        n15954) );
  OAI211_X1 U19118 ( .C1(n15956), .C2(n21116), .A(n15955), .B(n15954), .ZN(
        P1_U2815) );
  AOI22_X1 U19119 ( .A1(n15957), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_EBX_REG_24__SCAN_IN), .B2(n20173), .ZN(n15965) );
  AND3_X1 U19120 ( .A1(n20146), .A2(n15958), .A3(n21055), .ZN(n15962) );
  OAI22_X1 U19121 ( .A1(n15960), .A2(n20148), .B1(n15959), .B2(n20162), .ZN(
        n15961) );
  AOI211_X1 U19122 ( .C1(n20171), .C2(n15963), .A(n15962), .B(n15961), .ZN(
        n15964) );
  OAI211_X1 U19123 ( .C1(n15966), .C2(n20141), .A(n15965), .B(n15964), .ZN(
        P1_U2816) );
  INV_X1 U19124 ( .A(n15967), .ZN(n15969) );
  OAI21_X1 U19125 ( .B1(n15969), .B2(n15968), .A(n16051), .ZN(n16020) );
  AOI21_X1 U19126 ( .B1(n15971), .B2(n15970), .A(n16020), .ZN(n16000) );
  OAI21_X1 U19127 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n20175), .A(n16000), 
        .ZN(n15972) );
  AOI22_X1 U19128 ( .A1(n15972), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_EBX_REG_22__SCAN_IN), .B2(n20173), .ZN(n15973) );
  OAI21_X1 U19129 ( .B1(n15974), .B2(n20141), .A(n15973), .ZN(n15978) );
  OAI22_X1 U19130 ( .A1(n15976), .A2(n20148), .B1(P1_REIP_REG_22__SCAN_IN), 
        .B2(n15975), .ZN(n15977) );
  AOI211_X1 U19131 ( .C1(n15979), .C2(n20171), .A(n15978), .B(n15977), .ZN(
        n15980) );
  OAI21_X1 U19132 ( .B1(n20162), .B2(n16146), .A(n15980), .ZN(P1_U2818) );
  INV_X1 U19133 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n15989) );
  NOR2_X1 U19134 ( .A1(n16000), .A2(n15989), .ZN(n15986) );
  INV_X1 U19135 ( .A(n15981), .ZN(n15982) );
  AOI22_X1 U19136 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n20186), .B1(
        n20171), .B2(n15982), .ZN(n15983) );
  OAI21_X1 U19137 ( .B1(n20190), .B2(n15984), .A(n15983), .ZN(n15985) );
  AOI211_X1 U19138 ( .C1(n15987), .C2(n20165), .A(n15986), .B(n15985), .ZN(
        n15993) );
  INV_X1 U19139 ( .A(n15988), .ZN(n15991) );
  AOI22_X1 U19140 ( .A1(n20196), .A2(n15991), .B1(n15990), .B2(n15989), .ZN(
        n15992) );
  NAND2_X1 U19141 ( .A1(n15993), .A2(n15992), .ZN(P1_U2819) );
  OAI22_X1 U19142 ( .A1(n20190), .A2(n15994), .B1(n16075), .B2(n20141), .ZN(
        n15997) );
  OAI22_X1 U19143 ( .A1(n16069), .A2(n20148), .B1(n20162), .B2(n15995), .ZN(
        n15996) );
  AOI211_X1 U19144 ( .C1(n16071), .C2(n20171), .A(n15997), .B(n15996), .ZN(
        n15998) );
  OAI221_X1 U19145 ( .B1(n16000), .B2(n21073), .C1(n16000), .C2(n15999), .A(
        n15998), .ZN(P1_U2820) );
  AOI21_X1 U19146 ( .B1(n20186), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n20177), .ZN(n16001) );
  INV_X1 U19147 ( .A(n16001), .ZN(n16004) );
  OAI22_X1 U19148 ( .A1(n20190), .A2(n16002), .B1(n20189), .B2(n16081), .ZN(
        n16003) );
  AOI211_X1 U19149 ( .C1(P1_REIP_REG_19__SCAN_IN), .C2(n16020), .A(n16004), 
        .B(n16003), .ZN(n16008) );
  AOI22_X1 U19150 ( .A1(n16078), .A2(n20165), .B1(n20196), .B2(n16159), .ZN(
        n16007) );
  NAND2_X1 U19151 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n16005) );
  OAI211_X1 U19152 ( .C1(P1_REIP_REG_19__SCAN_IN), .C2(P1_REIP_REG_18__SCAN_IN), .A(n16013), .B(n16005), .ZN(n16006) );
  NAND3_X1 U19153 ( .A1(n16008), .A2(n16007), .A3(n16006), .ZN(P1_U2821) );
  AOI22_X1 U19154 ( .A1(n20171), .A2(n16009), .B1(n20173), .B2(
        P1_EBX_REG_18__SCAN_IN), .ZN(n16010) );
  OAI211_X1 U19155 ( .C1(n20141), .C2(n16011), .A(n16010), .B(n20187), .ZN(
        n16012) );
  AOI221_X1 U19156 ( .B1(n16013), .B2(n14775), .C1(n16020), .C2(
        P1_REIP_REG_18__SCAN_IN), .A(n16012), .ZN(n16017) );
  INV_X1 U19157 ( .A(n16014), .ZN(n16015) );
  NAND2_X1 U19158 ( .A1(n16015), .A2(n20165), .ZN(n16016) );
  OAI211_X1 U19159 ( .C1(n16179), .C2(n20162), .A(n16017), .B(n16016), .ZN(
        P1_U2822) );
  AOI22_X1 U19160 ( .A1(n20173), .A2(P1_EBX_REG_17__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n20186), .ZN(n16025) );
  AOI21_X1 U19161 ( .B1(n20171), .B2(n16088), .A(n20177), .ZN(n16024) );
  INV_X1 U19162 ( .A(n16018), .ZN(n16089) );
  INV_X1 U19163 ( .A(n16019), .ZN(n16184) );
  AOI22_X1 U19164 ( .A1(n16089), .A2(n20165), .B1(n20196), .B2(n16184), .ZN(
        n16023) );
  NOR2_X1 U19165 ( .A1(n20923), .A2(n16195), .ZN(n16021) );
  OAI221_X1 U19166 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n16021), .C1(
        P1_REIP_REG_17__SCAN_IN), .C2(n16026), .A(n16020), .ZN(n16022) );
  NAND4_X1 U19167 ( .A1(n16025), .A2(n16024), .A3(n16023), .A4(n16022), .ZN(
        P1_U2823) );
  AOI22_X1 U19168 ( .A1(n16098), .A2(n20171), .B1(n20196), .B2(n16200), .ZN(
        n16030) );
  AOI22_X1 U19169 ( .A1(n20173), .A2(P1_EBX_REG_15__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n20186), .ZN(n16029) );
  AOI21_X1 U19170 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n16035), .A(n20177), 
        .ZN(n16028) );
  AOI22_X1 U19171 ( .A1(n16099), .A2(n20165), .B1(n16026), .B2(n16195), .ZN(
        n16027) );
  NAND4_X1 U19172 ( .A1(n16030), .A2(n16029), .A3(n16028), .A4(n16027), .ZN(
        P1_U2825) );
  INV_X1 U19173 ( .A(n16031), .ZN(n16032) );
  AOI22_X1 U19174 ( .A1(n20173), .A2(P1_EBX_REG_14__SCAN_IN), .B1(n16032), 
        .B2(n20171), .ZN(n16039) );
  AOI22_X1 U19175 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n20186), .B1(
        n20196), .B2(n16204), .ZN(n16038) );
  OAI21_X1 U19176 ( .B1(n16033), .B2(n16053), .A(n20919), .ZN(n16034) );
  AOI22_X1 U19177 ( .A1(n16036), .A2(n20165), .B1(n16035), .B2(n16034), .ZN(
        n16037) );
  NAND4_X1 U19178 ( .A1(n16039), .A2(n16038), .A3(n16037), .A4(n20187), .ZN(
        P1_U2826) );
  AOI22_X1 U19179 ( .A1(n20173), .A2(P1_EBX_REG_12__SCAN_IN), .B1(n16107), 
        .B2(n20171), .ZN(n16045) );
  AOI22_X1 U19180 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n20186), .B1(
        n20196), .B2(n16040), .ZN(n16044) );
  INV_X1 U19181 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n16052) );
  INV_X1 U19182 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20917) );
  OAI21_X1 U19183 ( .B1(n16052), .B2(n16053), .A(n20917), .ZN(n16041) );
  AOI22_X1 U19184 ( .A1(n20165), .A2(n16106), .B1(n16042), .B2(n16041), .ZN(
        n16043) );
  NAND4_X1 U19185 ( .A1(n16045), .A2(n16044), .A3(n16043), .A4(n20187), .ZN(
        P1_U2828) );
  AOI21_X1 U19186 ( .B1(n20186), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20177), .ZN(n16048) );
  INV_X1 U19187 ( .A(n16046), .ZN(n16234) );
  AOI22_X1 U19188 ( .A1(n16234), .A2(n20196), .B1(n20173), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n16047) );
  OAI211_X1 U19189 ( .C1(n16118), .C2(n20189), .A(n16048), .B(n16047), .ZN(
        n16049) );
  AOI21_X1 U19190 ( .B1(n20165), .B2(n16115), .A(n16049), .ZN(n16050) );
  OAI221_X1 U19191 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n16053), .C1(n16052), 
        .C2(n16051), .A(n16050), .ZN(P1_U2829) );
  AOI22_X1 U19192 ( .A1(n16059), .A2(n16054), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n16057), .ZN(n16055) );
  OAI21_X1 U19193 ( .B1(n14715), .B2(n16056), .A(n16055), .ZN(P1_U2892) );
  AOI22_X1 U19194 ( .A1(n16059), .A2(n16058), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n16057), .ZN(n16060) );
  OAI21_X1 U19195 ( .B1(n14715), .B2(n16061), .A(n16060), .ZN(P1_U2893) );
  AOI22_X1 U19196 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n20290), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n16066) );
  XNOR2_X1 U19197 ( .A(n16086), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16062) );
  XNOR2_X1 U19198 ( .A(n16063), .B(n16062), .ZN(n16140) );
  AOI22_X1 U19199 ( .A1(n16064), .A2(n20313), .B1(n20250), .B2(n16140), .ZN(
        n16065) );
  OAI211_X1 U19200 ( .C1(n20243), .C2(n16067), .A(n16066), .B(n16065), .ZN(
        P1_U2976) );
  OAI22_X1 U19201 ( .A1(n16069), .A2(n20254), .B1(n16068), .B2(n20115), .ZN(
        n16070) );
  AOI21_X1 U19202 ( .B1(n20249), .B2(n16071), .A(n16070), .ZN(n16073) );
  OAI211_X1 U19203 ( .C1(n16075), .C2(n16074), .A(n16073), .B(n16072), .ZN(
        P1_U2979) );
  AOI22_X1 U19204 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n20290), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16080) );
  MUX2_X1 U19205 ( .A(n16086), .B(n16076), .S(n16163), .Z(n16077) );
  XNOR2_X1 U19206 ( .A(n16077), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16158) );
  AOI22_X1 U19207 ( .A1(n16078), .A2(n20313), .B1(n16158), .B2(n20250), .ZN(
        n16079) );
  OAI211_X1 U19208 ( .C1(n20243), .C2(n16081), .A(n16080), .B(n16079), .ZN(
        P1_U2980) );
  INV_X1 U19209 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16182) );
  OAI21_X1 U19210 ( .B1(n16083), .B2(n16082), .A(n9720), .ZN(n16085) );
  INV_X1 U19211 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16194) );
  NAND3_X1 U19212 ( .A1(n16086), .A2(n16194), .A3(n16085), .ZN(n16084) );
  OAI21_X1 U19213 ( .B1(n16086), .B2(n16085), .A(n16084), .ZN(n16087) );
  XOR2_X1 U19214 ( .A(n16182), .B(n16087), .Z(n16187) );
  AOI22_X1 U19215 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n20290), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n16091) );
  AOI22_X1 U19216 ( .A1(n16089), .A2(n20313), .B1(n16088), .B2(n20249), .ZN(
        n16090) );
  OAI211_X1 U19217 ( .C1(n20115), .C2(n16187), .A(n16091), .B(n16090), .ZN(
        P1_U2982) );
  INV_X1 U19218 ( .A(n16092), .ZN(n16093) );
  NOR2_X1 U19219 ( .A1(n16094), .A2(n16093), .ZN(n16097) );
  OAI21_X1 U19220 ( .B1(n16202), .B2(n16110), .A(n16095), .ZN(n16096) );
  XNOR2_X1 U19221 ( .A(n16097), .B(n16096), .ZN(n16196) );
  AOI22_X1 U19222 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20290), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16101) );
  AOI22_X1 U19223 ( .A1(n16099), .A2(n20313), .B1(n16098), .B2(n20249), .ZN(
        n16100) );
  OAI211_X1 U19224 ( .C1(n16196), .C2(n20115), .A(n16101), .B(n16100), .ZN(
        P1_U2984) );
  INV_X1 U19225 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16223) );
  INV_X1 U19226 ( .A(n16102), .ZN(n16103) );
  OAI21_X1 U19227 ( .B1(n16223), .B2(n16110), .A(n16103), .ZN(n16104) );
  AOI21_X1 U19228 ( .B1(n16105), .B2(n16104), .A(n10237), .ZN(n16226) );
  AOI22_X1 U19229 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20290), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16109) );
  AOI22_X1 U19230 ( .A1(n20249), .A2(n16107), .B1(n20313), .B2(n16106), .ZN(
        n16108) );
  OAI211_X1 U19231 ( .C1(n16226), .C2(n20115), .A(n16109), .B(n16108), .ZN(
        P1_U2987) );
  AOI22_X1 U19232 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20290), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16117) );
  NAND2_X1 U19233 ( .A1(n16110), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16112) );
  OAI21_X1 U19234 ( .B1(n14781), .B2(n16112), .A(n16111), .ZN(n16114) );
  XNOR2_X1 U19235 ( .A(n16114), .B(n16113), .ZN(n16235) );
  AOI22_X1 U19236 ( .A1(n20250), .A2(n16235), .B1(n20313), .B2(n16115), .ZN(
        n16116) );
  OAI211_X1 U19237 ( .C1(n20243), .C2(n16118), .A(n16117), .B(n16116), .ZN(
        P1_U2988) );
  AOI22_X1 U19238 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20290), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16125) );
  NAND2_X1 U19239 ( .A1(n16120), .A2(n16119), .ZN(n16121) );
  XNOR2_X1 U19240 ( .A(n16122), .B(n16121), .ZN(n16268) );
  INV_X1 U19241 ( .A(n20149), .ZN(n16123) );
  AOI22_X1 U19242 ( .A1(n16268), .A2(n20250), .B1(n20313), .B2(n16123), .ZN(
        n16124) );
  OAI211_X1 U19243 ( .C1(n20243), .C2(n20156), .A(n16125), .B(n16124), .ZN(
        P1_U2992) );
  AOI22_X1 U19244 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20290), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16131) );
  XNOR2_X1 U19245 ( .A(n16127), .B(n16126), .ZN(n16128) );
  XNOR2_X1 U19246 ( .A(n16129), .B(n16128), .ZN(n16275) );
  AOI22_X1 U19247 ( .A1(n16275), .A2(n20250), .B1(n20313), .B2(n20166), .ZN(
        n16130) );
  OAI211_X1 U19248 ( .C1(n20243), .C2(n20158), .A(n16131), .B(n16130), .ZN(
        P1_U2993) );
  AOI22_X1 U19249 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20290), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16137) );
  OAI21_X1 U19250 ( .B1(n16134), .B2(n16133), .A(n16132), .ZN(n16135) );
  INV_X1 U19251 ( .A(n16135), .ZN(n16279) );
  AOI22_X1 U19252 ( .A1(n16279), .A2(n20250), .B1(n20313), .B2(n20179), .ZN(
        n16136) );
  OAI211_X1 U19253 ( .C1(n20243), .C2(n20170), .A(n16137), .B(n16136), .ZN(
        P1_U2994) );
  AOI22_X1 U19254 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n20290), .B1(n16138), 
        .B2(n16143), .ZN(n16142) );
  AOI22_X1 U19255 ( .A1(n16140), .A2(n20296), .B1(n20292), .B2(n16139), .ZN(
        n16141) );
  OAI211_X1 U19256 ( .C1(n16144), .C2(n16143), .A(n16142), .B(n16141), .ZN(
        P1_U3008) );
  INV_X1 U19257 ( .A(n16145), .ZN(n16147) );
  OAI22_X1 U19258 ( .A1(n9815), .A2(n16147), .B1(n20288), .B2(n16146), .ZN(
        n16148) );
  AOI21_X1 U19259 ( .B1(n20296), .B2(n16149), .A(n16148), .ZN(n16153) );
  OAI211_X1 U19260 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16151), .B(n16150), .ZN(
        n16152) );
  OAI211_X1 U19261 ( .C1(n16154), .C2(n10234), .A(n16153), .B(n16152), .ZN(
        P1_U3009) );
  OR2_X1 U19262 ( .A1(n16155), .A2(n16273), .ZN(n16162) );
  INV_X1 U19263 ( .A(n16156), .ZN(n16157) );
  AOI22_X1 U19264 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n16157), .B1(
        n20290), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16161) );
  AOI22_X1 U19265 ( .A1(n20292), .A2(n16159), .B1(n20296), .B2(n16158), .ZN(
        n16160) );
  OAI211_X1 U19266 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n16162), .A(
        n16161), .B(n16160), .ZN(P1_U3012) );
  AND3_X1 U19267 ( .A1(n16164), .A2(n16163), .A3(n20296), .ZN(n16177) );
  NAND4_X1 U19268 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A4(n16205), .ZN(n16181) );
  NOR3_X1 U19269 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16182), .A3(
        n16181), .ZN(n16176) );
  INV_X1 U19270 ( .A(n16169), .ZN(n16166) );
  AOI21_X1 U19271 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16211), .A(
        n16165), .ZN(n16210) );
  AOI211_X1 U19272 ( .C1(n20276), .C2(n16166), .A(n16210), .B(n20258), .ZN(
        n16171) );
  INV_X1 U19273 ( .A(n16211), .ZN(n16167) );
  NOR3_X1 U19274 ( .A1(n16168), .A2(n16172), .A3(n16167), .ZN(n16170) );
  OAI211_X1 U19275 ( .C1(n16170), .C2(n20276), .A(n16169), .B(n16213), .ZN(
        n16212) );
  OAI211_X1 U19276 ( .C1(n16211), .C2(n16172), .A(n16171), .B(n16212), .ZN(
        n16215) );
  AOI21_X1 U19277 ( .B1(n16188), .B2(n16173), .A(n16215), .ZN(n16180) );
  OAI22_X1 U19278 ( .A1(n16180), .A2(n16174), .B1(n14775), .B2(n10234), .ZN(
        n16175) );
  NOR3_X1 U19279 ( .A1(n16177), .A2(n16176), .A3(n16175), .ZN(n16178) );
  OAI21_X1 U19280 ( .B1(n20288), .B2(n16179), .A(n16178), .ZN(P1_U3013) );
  AOI21_X1 U19281 ( .B1(n16182), .B2(n16181), .A(n16180), .ZN(n16183) );
  AOI21_X1 U19282 ( .B1(n20292), .B2(n16184), .A(n16183), .ZN(n16186) );
  NAND2_X1 U19283 ( .A1(n20290), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16185) );
  OAI211_X1 U19284 ( .C1(n16187), .C2(n16225), .A(n16186), .B(n16185), .ZN(
        P1_U3014) );
  AOI21_X1 U19285 ( .B1(n10013), .B2(n16188), .A(n16215), .ZN(n16203) );
  NAND2_X1 U19286 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16205), .ZN(
        n16197) );
  AOI221_X1 U19287 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(n16202), .C2(n16194), .A(
        n16197), .ZN(n16191) );
  OAI22_X1 U19288 ( .A1(n10234), .A2(n20923), .B1(n20288), .B2(n16189), .ZN(
        n16190) );
  AOI211_X1 U19289 ( .C1(n20296), .C2(n16192), .A(n16191), .B(n16190), .ZN(
        n16193) );
  OAI21_X1 U19290 ( .B1(n16203), .B2(n16194), .A(n16193), .ZN(P1_U3015) );
  NOR2_X1 U19291 ( .A1(n10234), .A2(n16195), .ZN(n16199) );
  OAI22_X1 U19292 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n16197), .B1(
        n16196), .B2(n16225), .ZN(n16198) );
  AOI211_X1 U19293 ( .C1(n20292), .C2(n16200), .A(n16199), .B(n16198), .ZN(
        n16201) );
  OAI21_X1 U19294 ( .B1(n16203), .B2(n16202), .A(n16201), .ZN(P1_U3016) );
  INV_X1 U19295 ( .A(n16215), .ZN(n16209) );
  AOI22_X1 U19296 ( .A1(n20290), .A2(P1_REIP_REG_14__SCAN_IN), .B1(n20292), 
        .B2(n16204), .ZN(n16208) );
  AOI22_X1 U19297 ( .A1(n20296), .A2(n16206), .B1(n16205), .B2(n10013), .ZN(
        n16207) );
  OAI211_X1 U19298 ( .C1(n16209), .C2(n10013), .A(n16208), .B(n16207), .ZN(
        P1_U3017) );
  AOI22_X1 U19299 ( .A1(n20290), .A2(P1_REIP_REG_13__SCAN_IN), .B1(n16211), 
        .B2(n16210), .ZN(n16218) );
  NAND2_X1 U19300 ( .A1(n16213), .A2(n16212), .ZN(n16214) );
  AOI22_X1 U19301 ( .A1(n20296), .A2(n16216), .B1(n16215), .B2(n16214), .ZN(
        n16217) );
  OAI211_X1 U19302 ( .C1(n20288), .C2(n16219), .A(n16218), .B(n16217), .ZN(
        P1_U3018) );
  NOR2_X1 U19303 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16273), .ZN(
        n16229) );
  NOR2_X1 U19304 ( .A1(n16220), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16233) );
  AOI21_X1 U19305 ( .B1(n20276), .B2(n16280), .A(n20258), .ZN(n16256) );
  OAI21_X1 U19306 ( .B1(n16244), .B2(n16220), .A(n20260), .ZN(n16221) );
  OAI211_X1 U19307 ( .C1(n16228), .C2(n20261), .A(n16256), .B(n16221), .ZN(
        n16236) );
  AOI21_X1 U19308 ( .B1(n16222), .B2(n16233), .A(n16236), .ZN(n16224) );
  OAI22_X1 U19309 ( .A1(n16226), .A2(n16225), .B1(n16224), .B2(n16223), .ZN(
        n16227) );
  AOI21_X1 U19310 ( .B1(n16229), .B2(n16228), .A(n16227), .ZN(n16231) );
  NAND2_X1 U19311 ( .A1(n20290), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n16230) );
  OAI211_X1 U19312 ( .C1(n20288), .C2(n16232), .A(n16231), .B(n16230), .ZN(
        P1_U3019) );
  INV_X1 U19313 ( .A(n16233), .ZN(n16239) );
  AOI22_X1 U19314 ( .A1(n20290), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n20292), 
        .B2(n16234), .ZN(n16238) );
  AOI22_X1 U19315 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16236), .B1(
        n20296), .B2(n16235), .ZN(n16237) );
  OAI211_X1 U19316 ( .C1(n16273), .C2(n16239), .A(n16238), .B(n16237), .ZN(
        P1_U3020) );
  NAND3_X1 U19317 ( .A1(n16264), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n16265), .ZN(n16254) );
  AOI22_X1 U19318 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n16241), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16240), .ZN(n16249) );
  AOI22_X1 U19319 ( .A1(n20290), .A2(P1_REIP_REG_10__SCAN_IN), .B1(n20292), 
        .B2(n16242), .ZN(n16248) );
  AOI211_X1 U19320 ( .C1(n20260), .C2(n16244), .A(n16126), .B(n16243), .ZN(
        n16245) );
  AOI21_X1 U19321 ( .B1(n16256), .B2(n16245), .A(n16259), .ZN(n16250) );
  AOI22_X1 U19322 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n16250), .B1(
        n20296), .B2(n16246), .ZN(n16247) );
  OAI211_X1 U19323 ( .C1(n16254), .C2(n16249), .A(n16248), .B(n16247), .ZN(
        P1_U3021) );
  AOI22_X1 U19324 ( .A1(n20290), .A2(P1_REIP_REG_9__SCAN_IN), .B1(n20292), 
        .B2(n20130), .ZN(n16253) );
  AOI22_X1 U19325 ( .A1(n16251), .A2(n20296), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16250), .ZN(n16252) );
  OAI211_X1 U19326 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n16254), .A(
        n16253), .B(n16252), .ZN(P1_U3022) );
  OAI211_X1 U19327 ( .C1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n16265), .ZN(n16263) );
  AOI22_X1 U19328 ( .A1(n20290), .A2(P1_REIP_REG_8__SCAN_IN), .B1(n20292), 
        .B2(n16255), .ZN(n16262) );
  NOR4_X1 U19329 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20259), .A3(
        n20256), .A4(n20279), .ZN(n16284) );
  OAI21_X1 U19330 ( .B1(n16258), .B2(n16257), .A(n16256), .ZN(n16278) );
  NOR3_X1 U19331 ( .A1(n16284), .A2(n16278), .A3(n16126), .ZN(n16272) );
  NOR2_X1 U19332 ( .A1(n16259), .A2(n16272), .ZN(n16267) );
  AOI22_X1 U19333 ( .A1(n16260), .A2(n20296), .B1(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n16267), .ZN(n16261) );
  OAI211_X1 U19334 ( .C1(n16264), .C2(n16263), .A(n16262), .B(n16261), .ZN(
        P1_U3023) );
  NAND2_X1 U19335 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16265), .ZN(
        n16271) );
  INV_X1 U19336 ( .A(n16266), .ZN(n20153) );
  AOI22_X1 U19337 ( .A1(n20290), .A2(P1_REIP_REG_7__SCAN_IN), .B1(n20292), 
        .B2(n20153), .ZN(n16270) );
  AOI22_X1 U19338 ( .A1(n16268), .A2(n20296), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16267), .ZN(n16269) );
  OAI211_X1 U19339 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n16271), .A(
        n16270), .B(n16269), .ZN(P1_U3024) );
  AOI21_X1 U19340 ( .B1(n16273), .B2(n16126), .A(n16272), .ZN(n16274) );
  AOI21_X1 U19341 ( .B1(n16275), .B2(n20296), .A(n16274), .ZN(n16277) );
  NAND2_X1 U19342 ( .A1(n20290), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n16276) );
  OAI211_X1 U19343 ( .C1(n20288), .C2(n20161), .A(n16277), .B(n16276), .ZN(
        P1_U3025) );
  AOI22_X1 U19344 ( .A1(n16279), .A2(n20296), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n16278), .ZN(n16286) );
  INV_X1 U19345 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20908) );
  NAND2_X1 U19346 ( .A1(n20276), .A2(n16280), .ZN(n16281) );
  OAI22_X1 U19347 ( .A1(n10234), .A2(n20908), .B1(n16282), .B2(n16281), .ZN(
        n16283) );
  AOI211_X1 U19348 ( .C1(n20292), .C2(n20178), .A(n16284), .B(n16283), .ZN(
        n16285) );
  NAND2_X1 U19349 ( .A1(n16286), .A2(n16285), .ZN(P1_U3026) );
  NOR3_X1 U19350 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20971), .A3(n16287), 
        .ZN(n16288) );
  AOI21_X1 U19351 ( .B1(n16289), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n16288), 
        .ZN(n20882) );
  AOI21_X1 U19352 ( .B1(n20882), .B2(n16295), .A(n16290), .ZN(n16291) );
  AOI221_X1 U19353 ( .B1(n16293), .B2(n16292), .C1(n16294), .C2(n16292), .A(
        n16291), .ZN(P1_U3162) );
  INV_X1 U19354 ( .A(n16294), .ZN(n16296) );
  OAI22_X1 U19355 ( .A1(n16296), .A2(n11516), .B1(n20971), .B2(n16295), .ZN(
        P1_U3466) );
  INV_X1 U19356 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16333) );
  OAI22_X1 U19357 ( .A1(n16333), .A2(n16297), .B1(n10109), .B2(n19186), .ZN(
        n16298) );
  AOI21_X1 U19358 ( .B1(n19199), .B2(P2_REIP_REG_31__SCAN_IN), .A(n16298), 
        .ZN(n16299) );
  OAI21_X1 U19359 ( .B1(n16300), .B2(n19216), .A(n16299), .ZN(n16301) );
  AOI21_X1 U19360 ( .B1(n16302), .B2(n19226), .A(n16301), .ZN(n16305) );
  OR2_X1 U19361 ( .A1(n14922), .A2(n16303), .ZN(n16304) );
  OAI211_X1 U19362 ( .C1(n16306), .C2(n19231), .A(n16305), .B(n16304), .ZN(
        P2_U2824) );
  AOI22_X1 U19363 ( .A1(n19221), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B1(
        n19199), .B2(P2_REIP_REG_29__SCAN_IN), .ZN(n16308) );
  NAND2_X1 U19364 ( .A1(n19183), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n16307) );
  OAI211_X1 U19365 ( .C1(n16309), .C2(n19129), .A(n16308), .B(n16307), .ZN(
        n16314) );
  OAI21_X1 U19366 ( .B1(n16317), .B2(n19231), .A(n16316), .ZN(P2_U2826) );
  OAI22_X1 U19367 ( .A1(n16318), .A2(n19216), .B1(n20050), .B2(n19215), .ZN(
        n16319) );
  INV_X1 U19368 ( .A(n16319), .ZN(n16332) );
  AOI22_X1 U19369 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19221), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n19183), .ZN(n16331) );
  INV_X1 U19370 ( .A(n16320), .ZN(n16321) );
  OAI22_X1 U19371 ( .A1(n16322), .A2(n19129), .B1(n16321), .B2(n19231), .ZN(
        n16323) );
  INV_X1 U19372 ( .A(n16323), .ZN(n16330) );
  INV_X1 U19373 ( .A(n16324), .ZN(n16328) );
  NAND3_X1 U19374 ( .A1(n16326), .A2(n16325), .A3(n13426), .ZN(n16327) );
  NAND3_X1 U19375 ( .A1(n16328), .A2(n19227), .A3(n16327), .ZN(n16329) );
  NAND4_X1 U19376 ( .A1(n16332), .A2(n16331), .A3(n16330), .A4(n16329), .ZN(
        P2_U2829) );
  AOI22_X1 U19377 ( .A1(n19252), .A2(n16334), .B1(n16333), .B2(n19259), .ZN(
        P2_U2856) );
  AOI22_X1 U19378 ( .A1(n16336), .A2(n19260), .B1(n19252), .B2(n16335), .ZN(
        n16337) );
  OAI21_X1 U19379 ( .B1(n19252), .B2(n14987), .A(n16337), .ZN(P2_U2864) );
  AOI21_X1 U19380 ( .B1(n16339), .B2(n15172), .A(n16338), .ZN(n16349) );
  INV_X1 U19381 ( .A(n16340), .ZN(n16379) );
  AOI22_X1 U19382 ( .A1(n16349), .A2(n19260), .B1(n19252), .B2(n16379), .ZN(
        n16341) );
  OAI21_X1 U19383 ( .B1(n19252), .B2(n15866), .A(n16341), .ZN(P2_U2865) );
  AOI21_X1 U19384 ( .B1(n16342), .B2(n15179), .A(n9737), .ZN(n16355) );
  AOI22_X1 U19385 ( .A1(n16355), .A2(n19260), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n19259), .ZN(n16343) );
  OAI21_X1 U19386 ( .B1(n19259), .B2(n19117), .A(n16343), .ZN(P2_U2867) );
  AOI21_X1 U19387 ( .B1(n16344), .B2(n14349), .A(n15178), .ZN(n16361) );
  AOI22_X1 U19388 ( .A1(n16361), .A2(n19260), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n19259), .ZN(n16345) );
  OAI21_X1 U19389 ( .B1(n19259), .B2(n16346), .A(n16345), .ZN(P2_U2869) );
  AOI22_X1 U19390 ( .A1(n19264), .A2(n16347), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n19320), .ZN(n16352) );
  AOI22_X1 U19391 ( .A1(n19266), .A2(BUF2_REG_22__SCAN_IN), .B1(n19265), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n16351) );
  AOI22_X1 U19392 ( .A1(n16349), .A2(n19308), .B1(n19321), .B2(n16348), .ZN(
        n16350) );
  NAND3_X1 U19393 ( .A1(n16352), .A2(n16351), .A3(n16350), .ZN(P2_U2897) );
  AOI22_X1 U19394 ( .A1(n19264), .A2(n16353), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n19320), .ZN(n16358) );
  AOI22_X1 U19395 ( .A1(n19266), .A2(BUF2_REG_20__SCAN_IN), .B1(n19265), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n16357) );
  INV_X1 U19396 ( .A(n16354), .ZN(n19123) );
  AOI22_X1 U19397 ( .A1(n16355), .A2(n19308), .B1(n19321), .B2(n19123), .ZN(
        n16356) );
  NAND3_X1 U19398 ( .A1(n16358), .A2(n16357), .A3(n16356), .ZN(P2_U2899) );
  AOI22_X1 U19399 ( .A1(n19264), .A2(n16359), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n19320), .ZN(n16364) );
  AOI22_X1 U19400 ( .A1(n19266), .A2(BUF2_REG_18__SCAN_IN), .B1(n19265), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n16363) );
  AOI22_X1 U19401 ( .A1(n16361), .A2(n19308), .B1(n19321), .B2(n16360), .ZN(
        n16362) );
  NAND3_X1 U19402 ( .A1(n16364), .A2(n16363), .A3(n16362), .ZN(P2_U2901) );
  INV_X1 U19403 ( .A(n16365), .ZN(n16366) );
  AOI21_X1 U19404 ( .B1(n16447), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16366), .ZN(n16374) );
  NAND2_X1 U19405 ( .A1(n16367), .A2(n19399), .ZN(n16370) );
  NAND2_X1 U19406 ( .A1(n16368), .A2(n19397), .ZN(n16369) );
  OAI211_X1 U19407 ( .C1(n16371), .C2(n16463), .A(n16370), .B(n16369), .ZN(
        n16372) );
  INV_X1 U19408 ( .A(n16372), .ZN(n16373) );
  OAI211_X1 U19409 ( .C1(n19405), .C2(n16375), .A(n16374), .B(n16373), .ZN(
        P2_U2990) );
  INV_X1 U19410 ( .A(n16376), .ZN(n16377) );
  AOI21_X1 U19411 ( .B1(n16447), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16377), .ZN(n16385) );
  NAND2_X1 U19412 ( .A1(n16378), .A2(n19397), .ZN(n16381) );
  NAND2_X1 U19413 ( .A1(n16379), .A2(n19399), .ZN(n16380) );
  OAI211_X1 U19414 ( .C1(n16382), .C2(n16463), .A(n16381), .B(n16380), .ZN(
        n16383) );
  INV_X1 U19415 ( .A(n16383), .ZN(n16384) );
  OAI211_X1 U19416 ( .C1(n19405), .C2(n16386), .A(n16385), .B(n16384), .ZN(
        P2_U2992) );
  NAND2_X1 U19417 ( .A1(n19198), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n16497) );
  INV_X1 U19418 ( .A(n16497), .ZN(n16387) );
  AOI21_X1 U19419 ( .B1(n16447), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16387), .ZN(n16399) );
  NAND2_X1 U19420 ( .A1(n16389), .A2(n16388), .ZN(n16390) );
  XNOR2_X1 U19421 ( .A(n16391), .B(n16390), .ZN(n16491) );
  OAI21_X1 U19422 ( .B1(n16412), .B2(n16392), .A(n11230), .ZN(n16394) );
  NAND2_X1 U19423 ( .A1(n16394), .A2(n16393), .ZN(n16486) );
  OR2_X1 U19424 ( .A1(n16486), .A2(n16463), .ZN(n16396) );
  INV_X1 U19425 ( .A(n19239), .ZN(n16487) );
  NAND2_X1 U19426 ( .A1(n19399), .A2(n16487), .ZN(n16395) );
  OAI211_X1 U19427 ( .C1(n16491), .C2(n16465), .A(n16396), .B(n16395), .ZN(
        n16397) );
  INV_X1 U19428 ( .A(n16397), .ZN(n16398) );
  OAI211_X1 U19429 ( .C1(n19405), .C2(n16400), .A(n16399), .B(n16398), .ZN(
        P2_U3000) );
  INV_X1 U19430 ( .A(n19166), .ZN(n16402) );
  OAI22_X1 U19431 ( .A1(n19405), .A2(n16402), .B1(n19214), .B2(n16401), .ZN(
        n16403) );
  INV_X1 U19432 ( .A(n16403), .ZN(n16408) );
  OAI22_X1 U19433 ( .A1(n16405), .A2(n16463), .B1(n16465), .B2(n16404), .ZN(
        n16406) );
  AOI21_X1 U19434 ( .B1(n19399), .B2(n19165), .A(n16406), .ZN(n16407) );
  OAI211_X1 U19435 ( .C1(n19394), .C2(n16409), .A(n16408), .B(n16407), .ZN(
        P2_U3001) );
  OAI22_X1 U19436 ( .A1(n19394), .A2(n10120), .B1(n19214), .B2(n19170), .ZN(
        n16410) );
  INV_X1 U19437 ( .A(n16410), .ZN(n16418) );
  NAND3_X1 U19438 ( .A1(n16412), .A2(n19400), .A3(n16411), .ZN(n16413) );
  OAI21_X1 U19439 ( .B1(n16414), .B2(n19245), .A(n16413), .ZN(n16415) );
  AOI21_X1 U19440 ( .B1(n19397), .B2(n16416), .A(n16415), .ZN(n16417) );
  OAI211_X1 U19441 ( .C1(n19405), .C2(n19177), .A(n16418), .B(n16417), .ZN(
        P2_U3002) );
  INV_X1 U19442 ( .A(n16419), .ZN(n16420) );
  AOI21_X1 U19443 ( .B1(n16473), .B2(n19192), .A(n16420), .ZN(n16425) );
  OAI22_X1 U19444 ( .A1(n16422), .A2(n16463), .B1(n16421), .B2(n16465), .ZN(
        n16423) );
  AOI21_X1 U19445 ( .B1(n19399), .B2(n19194), .A(n16423), .ZN(n16424) );
  OAI211_X1 U19446 ( .C1(n19394), .C2(n19187), .A(n16425), .B(n16424), .ZN(
        P2_U3003) );
  INV_X1 U19447 ( .A(n16426), .ZN(n16427) );
  AOI21_X1 U19448 ( .B1(n16447), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16427), .ZN(n16434) );
  NAND2_X1 U19449 ( .A1(n16428), .A2(n19397), .ZN(n16430) );
  NAND2_X1 U19450 ( .A1(n19399), .A2(n19250), .ZN(n16429) );
  OAI211_X1 U19451 ( .C1(n16431), .C2(n16463), .A(n16430), .B(n16429), .ZN(
        n16432) );
  INV_X1 U19452 ( .A(n16432), .ZN(n16433) );
  OAI211_X1 U19453 ( .C1(n19405), .C2(n16435), .A(n16434), .B(n16433), .ZN(
        P2_U3004) );
  OAI22_X1 U19454 ( .A1(n19405), .A2(n16437), .B1(n19214), .B2(n16436), .ZN(
        n16438) );
  INV_X1 U19455 ( .A(n16438), .ZN(n16444) );
  OAI22_X1 U19456 ( .A1(n16440), .A2(n16463), .B1(n16465), .B2(n16439), .ZN(
        n16441) );
  AOI21_X1 U19457 ( .B1(n19399), .B2(n16442), .A(n16441), .ZN(n16443) );
  OAI211_X1 U19458 ( .C1(n19394), .C2(n16445), .A(n16444), .B(n16443), .ZN(
        P2_U3005) );
  NAND2_X1 U19459 ( .A1(n19198), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n16508) );
  INV_X1 U19460 ( .A(n16508), .ZN(n16446) );
  AOI21_X1 U19461 ( .B1(n16447), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16446), .ZN(n16458) );
  NAND2_X1 U19462 ( .A1(n16449), .A2(n16448), .ZN(n16454) );
  INV_X1 U19463 ( .A(n16450), .ZN(n16451) );
  AOI21_X1 U19464 ( .B1(n15395), .B2(n16452), .A(n16451), .ZN(n16453) );
  XOR2_X1 U19465 ( .A(n16454), .B(n16453), .Z(n16505) );
  INV_X1 U19466 ( .A(n19258), .ZN(n16504) );
  XOR2_X1 U19467 ( .A(n16455), .B(n16456), .Z(n16503) );
  AOI222_X1 U19468 ( .A1(n16505), .A2(n19397), .B1(n19399), .B2(n16504), .C1(
        n16503), .C2(n19400), .ZN(n16457) );
  OAI211_X1 U19469 ( .C1(n19405), .C2(n16459), .A(n16458), .B(n16457), .ZN(
        P2_U3006) );
  INV_X1 U19470 ( .A(n19223), .ZN(n16461) );
  OAI22_X1 U19471 ( .A1(n19405), .A2(n16461), .B1(n19214), .B2(n16460), .ZN(
        n16462) );
  INV_X1 U19472 ( .A(n16462), .ZN(n16469) );
  OAI22_X1 U19473 ( .A1(n16466), .A2(n16465), .B1(n16464), .B2(n16463), .ZN(
        n16467) );
  AOI21_X1 U19474 ( .B1(n19399), .B2(n19225), .A(n16467), .ZN(n16468) );
  OAI211_X1 U19475 ( .C1(n19394), .C2(n16470), .A(n16469), .B(n16468), .ZN(
        P2_U3009) );
  NOR2_X1 U19476 ( .A1(n19214), .A2(n16471), .ZN(n16524) );
  AOI21_X1 U19477 ( .B1(n16473), .B2(n16472), .A(n16524), .ZN(n16483) );
  NAND2_X1 U19478 ( .A1(n16475), .A2(n16474), .ZN(n16477) );
  XNOR2_X1 U19479 ( .A(n16477), .B(n16476), .ZN(n16531) );
  OAI21_X1 U19480 ( .B1(n16480), .B2(n16479), .A(n16478), .ZN(n16528) );
  INV_X1 U19481 ( .A(n16528), .ZN(n16481) );
  AOI222_X1 U19482 ( .A1(n16531), .A2(n19397), .B1(n19400), .B2(n16481), .C1(
        n15110), .C2(n19399), .ZN(n16482) );
  OAI211_X1 U19483 ( .C1(n16484), .C2(n19394), .A(n16483), .B(n16482), .ZN(
        P2_U3011) );
  AOI22_X1 U19484 ( .A1(n16485), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n16502), .B2(n19274), .ZN(n16499) );
  OR2_X1 U19485 ( .A1(n16486), .A2(n16527), .ZN(n16489) );
  NAND2_X1 U19486 ( .A1(n16525), .A2(n16487), .ZN(n16488) );
  OAI211_X1 U19487 ( .C1(n16491), .C2(n16490), .A(n16489), .B(n16488), .ZN(
        n16492) );
  INV_X1 U19488 ( .A(n16492), .ZN(n16498) );
  OAI211_X1 U19489 ( .C1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n16495), .A(
        n16494), .B(n16493), .ZN(n16496) );
  NAND4_X1 U19490 ( .A1(n16499), .A2(n16498), .A3(n16497), .A4(n16496), .ZN(
        P2_U3032) );
  INV_X1 U19491 ( .A(n16506), .ZN(n16500) );
  OAI21_X1 U19492 ( .B1(n16501), .B2(n16500), .A(n16533), .ZN(n16513) );
  AOI22_X1 U19493 ( .A1(n16513), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16502), .B2(n19289), .ZN(n16510) );
  AOI222_X1 U19494 ( .A1(n16505), .A2(n16530), .B1(n16525), .B2(n16504), .C1(
        n16503), .C2(n10972), .ZN(n16509) );
  NOR2_X1 U19495 ( .A1(n16506), .A2(n16535), .ZN(n16515) );
  OAI221_X1 U19496 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n11205), .C2(n16514), .A(
        n16515), .ZN(n16507) );
  NAND4_X1 U19497 ( .A1(n16510), .A2(n16509), .A3(n16508), .A4(n16507), .ZN(
        P2_U3038) );
  OAI21_X1 U19498 ( .B1(n16522), .B2(n19292), .A(n16511), .ZN(n16512) );
  AOI221_X1 U19499 ( .B1(n16515), .B2(n16514), .C1(n16513), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16512), .ZN(n16520) );
  INV_X1 U19500 ( .A(n16516), .ZN(n16518) );
  AOI22_X1 U19501 ( .A1(n16518), .A2(n16530), .B1(n16525), .B2(n16517), .ZN(
        n16519) );
  OAI211_X1 U19502 ( .C1(n16527), .C2(n16521), .A(n16520), .B(n16519), .ZN(
        P2_U3039) );
  NOR2_X1 U19503 ( .A1(n20078), .A2(n16522), .ZN(n16523) );
  AOI211_X1 U19504 ( .C1(n16525), .C2(n15110), .A(n16524), .B(n16523), .ZN(
        n16526) );
  OAI21_X1 U19505 ( .B1(n16528), .B2(n16527), .A(n16526), .ZN(n16529) );
  AOI21_X1 U19506 ( .B1(n16531), .B2(n16530), .A(n16529), .ZN(n16532) );
  OAI221_X1 U19507 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16535), .C1(
        n16534), .C2(n16533), .A(n16532), .ZN(P2_U3043) );
  INV_X1 U19508 ( .A(n16536), .ZN(n16537) );
  AOI211_X1 U19509 ( .C1(n16540), .C2(n16539), .A(n16538), .B(n16537), .ZN(
        n16547) );
  AOI21_X1 U19510 ( .B1(n16543), .B2(n16542), .A(n16541), .ZN(n16545) );
  OAI21_X1 U19511 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16545), .A(n16544), 
        .ZN(n16546) );
  OAI211_X1 U19512 ( .C1(n16549), .C2(n16548), .A(n16547), .B(n16546), .ZN(
        P2_U3176) );
  NOR2_X4 U19513 ( .A1(n9969), .A2(n16696), .ZN(n18070) );
  OAI21_X4 U19514 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19053), .A(n16696), 
        .ZN(n18080) );
  NOR2_X2 U19515 ( .A1(n18039), .A2(n18041), .ZN(n18078) );
  NAND2_X2 U19516 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18078), .ZN(n17926) );
  INV_X1 U19517 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16555) );
  INV_X1 U19518 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17939) );
  NAND2_X1 U19519 ( .A1(n17920), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17878) );
  NAND3_X1 U19520 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17834) );
  INV_X1 U19521 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17833) );
  INV_X1 U19522 ( .A(n17805), .ZN(n16552) );
  NAND3_X1 U19523 ( .A1(n17759), .A2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17749) );
  INV_X1 U19524 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17748) );
  INV_X1 U19525 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17711) );
  INV_X1 U19526 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18077) );
  NAND2_X1 U19527 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16591), .ZN(
        n16553) );
  XOR2_X2 U19528 ( .A(n16555), .B(n16553), .Z(n17018) );
  NAND2_X1 U19529 ( .A1(n19059), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18917) );
  INV_X1 U19530 ( .A(n18917), .ZN(n17757) );
  INV_X2 U19531 ( .A(n18786), .ZN(n18478) );
  OAI21_X2 U19532 ( .B1(n18077), .B2(n17830), .A(n18478), .ZN(n17918) );
  OR2_X1 U19533 ( .A1(n16554), .A2(n17879), .ZN(n16574) );
  XNOR2_X1 U19534 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16556) );
  NOR2_X1 U19535 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17830), .ZN(
        n16593) );
  NAND2_X1 U19536 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9790), .ZN(
        n16592) );
  INV_X1 U19537 ( .A(n16592), .ZN(n16717) );
  NAND2_X1 U19538 ( .A1(n18786), .A2(n16554), .ZN(n16580) );
  OAI211_X1 U19539 ( .C1(n16717), .C2(n18917), .A(n18080), .B(n16580), .ZN(
        n16582) );
  NOR2_X1 U19540 ( .A1(n16593), .A2(n16582), .ZN(n16572) );
  OAI22_X1 U19541 ( .A1(n16574), .A2(n16556), .B1(n16572), .B2(n16555), .ZN(
        n16557) );
  AOI211_X1 U19542 ( .C1(n17943), .C2(n17018), .A(n16558), .B(n16557), .ZN(
        n16564) );
  NOR2_X4 U19543 ( .A1(n16696), .A2(n17658), .ZN(n18074) );
  AOI21_X1 U19544 ( .B1(n16562), .B2(n17996), .A(n16561), .ZN(n16563) );
  OAI211_X1 U19545 ( .C1(n16565), .C2(n18084), .A(n16564), .B(n16563), .ZN(
        P3_U2799) );
  NAND2_X1 U19546 ( .A1(n17809), .A2(n16566), .ZN(n16583) );
  NAND2_X1 U19547 ( .A1(n18070), .A2(n16567), .ZN(n16585) );
  OAI22_X2 U19548 ( .A1(n18084), .A2(n18244), .B1(n17999), .B2(n18272), .ZN(
        n17980) );
  AND3_X1 U19549 ( .A1(n16579), .A2(n16569), .A3(n17742), .ZN(n16576) );
  INV_X1 U19550 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16573) );
  XNOR2_X1 U19551 ( .A(n16573), .B(n16591), .ZN(n16735) );
  AOI21_X1 U19552 ( .B1(n17943), .B2(n16735), .A(n16570), .ZN(n16571) );
  OAI221_X1 U19553 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16574), .C1(
        n16573), .C2(n16572), .A(n16571), .ZN(n16575) );
  AOI211_X1 U19554 ( .C1(n17996), .C2(n16577), .A(n16576), .B(n16575), .ZN(
        n16578) );
  OAI221_X1 U19555 ( .B1(n16579), .B2(n16583), .C1(n16579), .C2(n16585), .A(
        n16578), .ZN(P3_U2800) );
  INV_X1 U19556 ( .A(n16580), .ZN(n16581) );
  AOI22_X1 U19557 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n16582), .B1(
        n9790), .B2(n16581), .ZN(n16597) );
  AOI21_X1 U19558 ( .B1(n16586), .B2(n16584), .A(n16583), .ZN(n16589) );
  AOI21_X1 U19559 ( .B1(n16587), .B2(n16586), .A(n16585), .ZN(n16588) );
  AOI211_X1 U19560 ( .C1(n17996), .C2(n16590), .A(n16589), .B(n16588), .ZN(
        n16596) );
  AOI21_X1 U19561 ( .B1(n9951), .B2(n16592), .A(n16591), .ZN(n16746) );
  OAI21_X1 U19562 ( .B1(n16593), .B2(n17943), .A(n16746), .ZN(n16594) );
  NAND4_X1 U19563 ( .A1(n16597), .A2(n16596), .A3(n16595), .A4(n16594), .ZN(
        P3_U2801) );
  NOR3_X1 U19564 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16599) );
  NOR4_X1 U19565 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16598) );
  INV_X2 U19566 ( .A(n16682), .ZN(U215) );
  NAND4_X1 U19567 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16599), .A3(n16598), .A4(
        U215), .ZN(U213) );
  INV_X1 U19568 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16684) );
  INV_X2 U19569 ( .A(U214), .ZN(n16645) );
  INV_X1 U19570 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16685) );
  OAI222_X1 U19571 ( .A1(U212), .A2(n16684), .B1(n16647), .B2(n20371), .C1(
        U214), .C2(n16685), .ZN(U216) );
  INV_X1 U19572 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20360) );
  AOI22_X1 U19573 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16630), .ZN(n16601) );
  OAI21_X1 U19574 ( .B1(n20360), .B2(n16647), .A(n16601), .ZN(U217) );
  INV_X1 U19575 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20353) );
  AOI22_X1 U19576 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16630), .ZN(n16602) );
  OAI21_X1 U19577 ( .B1(n20353), .B2(n16647), .A(n16602), .ZN(U218) );
  INV_X1 U19578 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20346) );
  AOI22_X1 U19579 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16630), .ZN(n16603) );
  OAI21_X1 U19580 ( .B1(n20346), .B2(n16647), .A(n16603), .ZN(U219) );
  AOI22_X1 U19581 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16630), .ZN(n16604) );
  OAI21_X1 U19582 ( .B1(n20338), .B2(n16647), .A(n16604), .ZN(U220) );
  INV_X1 U19583 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20331) );
  AOI22_X1 U19584 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16630), .ZN(n16605) );
  OAI21_X1 U19585 ( .B1(n20331), .B2(n16647), .A(n16605), .ZN(U221) );
  AOI22_X1 U19586 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16630), .ZN(n16606) );
  OAI21_X1 U19587 ( .B1(n20325), .B2(n16647), .A(n16606), .ZN(U222) );
  INV_X1 U19588 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20314) );
  AOI22_X1 U19589 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16630), .ZN(n16607) );
  OAI21_X1 U19590 ( .B1(n20314), .B2(n16647), .A(n16607), .ZN(U223) );
  INV_X1 U19591 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20367) );
  AOI22_X1 U19592 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16630), .ZN(n16608) );
  OAI21_X1 U19593 ( .B1(n20367), .B2(n16647), .A(n16608), .ZN(U224) );
  INV_X1 U19594 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20362) );
  AOI22_X1 U19595 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16630), .ZN(n16609) );
  OAI21_X1 U19596 ( .B1(n20362), .B2(n16647), .A(n16609), .ZN(U225) );
  AOI22_X1 U19597 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16630), .ZN(n16610) );
  OAI21_X1 U19598 ( .B1(n20355), .B2(n16647), .A(n16610), .ZN(U226) );
  INV_X1 U19599 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20349) );
  AOI22_X1 U19600 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16630), .ZN(n16611) );
  OAI21_X1 U19601 ( .B1(n20349), .B2(n16647), .A(n16611), .ZN(U227) );
  AOI22_X1 U19602 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16630), .ZN(n16612) );
  OAI21_X1 U19603 ( .B1(n20341), .B2(n16647), .A(n16612), .ZN(U228) );
  INV_X1 U19604 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20333) );
  AOI22_X1 U19605 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16630), .ZN(n16613) );
  OAI21_X1 U19606 ( .B1(n20333), .B2(n16647), .A(n16613), .ZN(U229) );
  AOI22_X1 U19607 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16630), .ZN(n16614) );
  OAI21_X1 U19608 ( .B1(n14356), .B2(n16647), .A(n16614), .ZN(U230) );
  INV_X1 U19609 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20321) );
  AOI22_X1 U19610 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16630), .ZN(n16615) );
  OAI21_X1 U19611 ( .B1(n20321), .B2(n16647), .A(n16615), .ZN(U231) );
  AOI22_X1 U19612 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16630), .ZN(n16616) );
  OAI21_X1 U19613 ( .B1(n16617), .B2(n16647), .A(n16616), .ZN(U232) );
  INV_X1 U19614 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16619) );
  AOI22_X1 U19615 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16630), .ZN(n16618) );
  OAI21_X1 U19616 ( .B1(n16619), .B2(n16647), .A(n16618), .ZN(U233) );
  AOI22_X1 U19617 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16630), .ZN(n16620) );
  OAI21_X1 U19618 ( .B1(n16621), .B2(n16647), .A(n16620), .ZN(U234) );
  INV_X1 U19619 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16623) );
  AOI22_X1 U19620 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16630), .ZN(n16622) );
  OAI21_X1 U19621 ( .B1(n16623), .B2(n16647), .A(n16622), .ZN(U235) );
  AOI22_X1 U19622 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16630), .ZN(n16624) );
  OAI21_X1 U19623 ( .B1(n13510), .B2(n16647), .A(n16624), .ZN(U236) );
  INV_X1 U19624 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16626) );
  AOI22_X1 U19625 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16630), .ZN(n16625) );
  OAI21_X1 U19626 ( .B1(n16626), .B2(n16647), .A(n16625), .ZN(U237) );
  AOI22_X1 U19627 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16630), .ZN(n16627) );
  OAI21_X1 U19628 ( .B1(n13522), .B2(n16647), .A(n16627), .ZN(U238) );
  INV_X1 U19629 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16629) );
  AOI22_X1 U19630 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16630), .ZN(n16628) );
  OAI21_X1 U19631 ( .B1(n16629), .B2(n16647), .A(n16628), .ZN(U239) );
  AOI22_X1 U19632 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16630), .ZN(n16631) );
  OAI21_X1 U19633 ( .B1(n16632), .B2(n16647), .A(n16631), .ZN(U240) );
  AOI22_X1 U19634 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16630), .ZN(n16633) );
  OAI21_X1 U19635 ( .B1(n16634), .B2(n16647), .A(n16633), .ZN(U241) );
  AOI22_X1 U19636 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16630), .ZN(n16635) );
  OAI21_X1 U19637 ( .B1(n16636), .B2(n16647), .A(n16635), .ZN(U242) );
  AOI22_X1 U19638 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16630), .ZN(n16637) );
  OAI21_X1 U19639 ( .B1(n16638), .B2(n16647), .A(n16637), .ZN(U243) );
  INV_X1 U19640 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16640) );
  AOI22_X1 U19641 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16630), .ZN(n16639) );
  OAI21_X1 U19642 ( .B1(n16640), .B2(n16647), .A(n16639), .ZN(U244) );
  INV_X1 U19643 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16642) );
  AOI22_X1 U19644 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16630), .ZN(n16641) );
  OAI21_X1 U19645 ( .B1(n16642), .B2(n16647), .A(n16641), .ZN(U245) );
  INV_X1 U19646 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16644) );
  AOI22_X1 U19647 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16630), .ZN(n16643) );
  OAI21_X1 U19648 ( .B1(n16644), .B2(n16647), .A(n16643), .ZN(U246) );
  INV_X1 U19649 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16648) );
  AOI22_X1 U19650 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16645), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16630), .ZN(n16646) );
  OAI21_X1 U19651 ( .B1(n16648), .B2(n16647), .A(n16646), .ZN(U247) );
  OAI22_X1 U19652 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16682), .ZN(n16649) );
  INV_X1 U19653 ( .A(n16649), .ZN(U251) );
  OAI22_X1 U19654 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16682), .ZN(n16650) );
  INV_X1 U19655 ( .A(n16650), .ZN(U252) );
  OAI22_X1 U19656 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16682), .ZN(n16651) );
  INV_X1 U19657 ( .A(n16651), .ZN(U253) );
  OAI22_X1 U19658 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16682), .ZN(n16652) );
  INV_X1 U19659 ( .A(n16652), .ZN(U254) );
  OAI22_X1 U19660 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16682), .ZN(n16653) );
  INV_X1 U19661 ( .A(n16653), .ZN(U255) );
  OAI22_X1 U19662 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16682), .ZN(n16654) );
  INV_X1 U19663 ( .A(n16654), .ZN(U256) );
  OAI22_X1 U19664 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16682), .ZN(n16655) );
  INV_X1 U19665 ( .A(n16655), .ZN(U257) );
  OAI22_X1 U19666 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16682), .ZN(n16656) );
  INV_X1 U19667 ( .A(n16656), .ZN(U258) );
  OAI22_X1 U19668 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16682), .ZN(n16657) );
  INV_X1 U19669 ( .A(n16657), .ZN(U259) );
  OAI22_X1 U19670 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16676), .ZN(n16658) );
  INV_X1 U19671 ( .A(n16658), .ZN(U260) );
  OAI22_X1 U19672 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16676), .ZN(n16659) );
  INV_X1 U19673 ( .A(n16659), .ZN(U261) );
  OAI22_X1 U19674 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16682), .ZN(n16660) );
  INV_X1 U19675 ( .A(n16660), .ZN(U262) );
  OAI22_X1 U19676 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16682), .ZN(n16661) );
  INV_X1 U19677 ( .A(n16661), .ZN(U263) );
  OAI22_X1 U19678 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16682), .ZN(n16662) );
  INV_X1 U19679 ( .A(n16662), .ZN(U264) );
  OAI22_X1 U19680 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16682), .ZN(n16663) );
  INV_X1 U19681 ( .A(n16663), .ZN(U265) );
  OAI22_X1 U19682 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16676), .ZN(n16664) );
  INV_X1 U19683 ( .A(n16664), .ZN(U266) );
  OAI22_X1 U19684 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16676), .ZN(n16665) );
  INV_X1 U19685 ( .A(n16665), .ZN(U267) );
  OAI22_X1 U19686 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16676), .ZN(n16666) );
  INV_X1 U19687 ( .A(n16666), .ZN(U268) );
  OAI22_X1 U19688 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16676), .ZN(n16667) );
  INV_X1 U19689 ( .A(n16667), .ZN(U269) );
  OAI22_X1 U19690 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16676), .ZN(n16668) );
  INV_X1 U19691 ( .A(n16668), .ZN(U270) );
  OAI22_X1 U19692 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16676), .ZN(n16669) );
  INV_X1 U19693 ( .A(n16669), .ZN(U271) );
  OAI22_X1 U19694 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16682), .ZN(n16670) );
  INV_X1 U19695 ( .A(n16670), .ZN(U272) );
  OAI22_X1 U19696 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16682), .ZN(n16671) );
  INV_X1 U19697 ( .A(n16671), .ZN(U273) );
  OAI22_X1 U19698 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16676), .ZN(n16672) );
  INV_X1 U19699 ( .A(n16672), .ZN(U274) );
  OAI22_X1 U19700 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16682), .ZN(n16673) );
  INV_X1 U19701 ( .A(n16673), .ZN(U275) );
  OAI22_X1 U19702 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16682), .ZN(n16674) );
  INV_X1 U19703 ( .A(n16674), .ZN(U276) );
  OAI22_X1 U19704 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16682), .ZN(n16675) );
  INV_X1 U19705 ( .A(n16675), .ZN(U277) );
  OAI22_X1 U19706 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16676), .ZN(n16677) );
  INV_X1 U19707 ( .A(n16677), .ZN(U278) );
  OAI22_X1 U19708 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16682), .ZN(n16678) );
  INV_X1 U19709 ( .A(n16678), .ZN(U279) );
  OAI22_X1 U19710 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16682), .ZN(n16679) );
  INV_X1 U19711 ( .A(n16679), .ZN(U280) );
  OAI22_X1 U19712 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16682), .ZN(n16681) );
  INV_X1 U19713 ( .A(n16681), .ZN(U281) );
  INV_X1 U19714 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18452) );
  AOI22_X1 U19715 ( .A1(n16682), .A2(n16684), .B1(n18452), .B2(U215), .ZN(U282) );
  INV_X1 U19716 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16683) );
  AOI222_X1 U19717 ( .A1(n16685), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16684), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16683), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16686) );
  INV_X2 U19718 ( .A(n16688), .ZN(n16687) );
  INV_X1 U19719 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18952) );
  INV_X1 U19720 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20025) );
  AOI22_X1 U19721 ( .A1(n16687), .A2(n18952), .B1(n20025), .B2(n16688), .ZN(
        U347) );
  INV_X1 U19722 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18950) );
  INV_X1 U19723 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20024) );
  AOI22_X1 U19724 ( .A1(n16687), .A2(n18950), .B1(n20024), .B2(n16688), .ZN(
        U348) );
  INV_X1 U19725 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18947) );
  INV_X1 U19726 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20023) );
  AOI22_X1 U19727 ( .A1(n16687), .A2(n18947), .B1(n20023), .B2(n16688), .ZN(
        U349) );
  INV_X1 U19728 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18946) );
  INV_X1 U19729 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20022) );
  AOI22_X1 U19730 ( .A1(n16687), .A2(n18946), .B1(n20022), .B2(n16688), .ZN(
        U350) );
  INV_X1 U19731 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18944) );
  INV_X1 U19732 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20020) );
  AOI22_X1 U19733 ( .A1(n16687), .A2(n18944), .B1(n20020), .B2(n16688), .ZN(
        U351) );
  INV_X1 U19734 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18942) );
  INV_X1 U19735 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20018) );
  AOI22_X1 U19736 ( .A1(n16687), .A2(n18942), .B1(n20018), .B2(n16688), .ZN(
        U352) );
  INV_X1 U19737 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18940) );
  INV_X1 U19738 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20017) );
  AOI22_X1 U19739 ( .A1(n16687), .A2(n18940), .B1(n20017), .B2(n16688), .ZN(
        U353) );
  INV_X1 U19740 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18938) );
  AOI22_X1 U19741 ( .A1(n16687), .A2(n18938), .B1(n20016), .B2(n16688), .ZN(
        U354) );
  INV_X1 U19742 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18992) );
  INV_X1 U19743 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20057) );
  AOI22_X1 U19744 ( .A1(n16687), .A2(n18992), .B1(n20057), .B2(n16688), .ZN(
        U356) );
  INV_X1 U19745 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18988) );
  INV_X1 U19746 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20055) );
  AOI22_X1 U19747 ( .A1(n16687), .A2(n18988), .B1(n20055), .B2(n16688), .ZN(
        U357) );
  INV_X1 U19748 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18987) );
  INV_X1 U19749 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20052) );
  AOI22_X1 U19750 ( .A1(n16687), .A2(n18987), .B1(n20052), .B2(n16688), .ZN(
        U358) );
  INV_X1 U19751 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18984) );
  INV_X1 U19752 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20051) );
  AOI22_X1 U19753 ( .A1(n16687), .A2(n18984), .B1(n20051), .B2(n16688), .ZN(
        U359) );
  INV_X1 U19754 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18982) );
  INV_X1 U19755 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20049) );
  AOI22_X1 U19756 ( .A1(n16687), .A2(n18982), .B1(n20049), .B2(n16688), .ZN(
        U360) );
  INV_X1 U19757 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18980) );
  INV_X1 U19758 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20047) );
  AOI22_X1 U19759 ( .A1(n16687), .A2(n18980), .B1(n20047), .B2(n16688), .ZN(
        U361) );
  INV_X1 U19760 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18977) );
  INV_X1 U19761 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20045) );
  AOI22_X1 U19762 ( .A1(n16687), .A2(n18977), .B1(n20045), .B2(n16688), .ZN(
        U362) );
  INV_X1 U19763 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18976) );
  INV_X1 U19764 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20043) );
  AOI22_X1 U19765 ( .A1(n16687), .A2(n18976), .B1(n20043), .B2(n16688), .ZN(
        U363) );
  INV_X1 U19766 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18973) );
  INV_X1 U19767 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20042) );
  AOI22_X1 U19768 ( .A1(n16687), .A2(n18973), .B1(n20042), .B2(n16688), .ZN(
        U364) );
  INV_X1 U19769 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18936) );
  INV_X1 U19770 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20015) );
  AOI22_X1 U19771 ( .A1(n16687), .A2(n18936), .B1(n20015), .B2(n16688), .ZN(
        U365) );
  INV_X1 U19772 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18972) );
  INV_X1 U19773 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20040) );
  AOI22_X1 U19774 ( .A1(n16687), .A2(n18972), .B1(n20040), .B2(n16688), .ZN(
        U366) );
  INV_X1 U19775 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18969) );
  INV_X1 U19776 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20039) );
  AOI22_X1 U19777 ( .A1(n16687), .A2(n18969), .B1(n20039), .B2(n16688), .ZN(
        U367) );
  INV_X1 U19778 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18968) );
  INV_X1 U19779 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20037) );
  AOI22_X1 U19780 ( .A1(n16687), .A2(n18968), .B1(n20037), .B2(n16688), .ZN(
        U368) );
  INV_X1 U19781 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18966) );
  INV_X1 U19782 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20036) );
  AOI22_X1 U19783 ( .A1(n16687), .A2(n18966), .B1(n20036), .B2(n16688), .ZN(
        U369) );
  INV_X1 U19784 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18964) );
  INV_X1 U19785 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20034) );
  AOI22_X1 U19786 ( .A1(n16687), .A2(n18964), .B1(n20034), .B2(n16688), .ZN(
        U370) );
  INV_X1 U19787 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18962) );
  INV_X1 U19788 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20032) );
  AOI22_X1 U19789 ( .A1(n16687), .A2(n18962), .B1(n20032), .B2(n16688), .ZN(
        U371) );
  INV_X1 U19790 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18959) );
  INV_X1 U19791 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20030) );
  AOI22_X1 U19792 ( .A1(n16687), .A2(n18959), .B1(n20030), .B2(n16688), .ZN(
        U372) );
  INV_X1 U19793 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18958) );
  INV_X1 U19794 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20029) );
  AOI22_X1 U19795 ( .A1(n16687), .A2(n18958), .B1(n20029), .B2(n16688), .ZN(
        U373) );
  INV_X1 U19796 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18956) );
  INV_X1 U19797 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20028) );
  AOI22_X1 U19798 ( .A1(n16687), .A2(n18956), .B1(n20028), .B2(n16688), .ZN(
        U374) );
  INV_X1 U19799 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18954) );
  INV_X1 U19800 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20027) );
  AOI22_X1 U19801 ( .A1(n16687), .A2(n18954), .B1(n20027), .B2(n16688), .ZN(
        U375) );
  INV_X1 U19802 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18934) );
  INV_X1 U19803 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20012) );
  AOI22_X1 U19804 ( .A1(n16687), .A2(n18934), .B1(n20012), .B2(n16688), .ZN(
        U376) );
  INV_X1 U19805 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18933) );
  NAND2_X1 U19806 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18933), .ZN(n18922) );
  AOI22_X1 U19807 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18922), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18931), .ZN(n19005) );
  AOI21_X1 U19808 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n19005), .ZN(n16689) );
  INV_X1 U19809 ( .A(n16689), .ZN(P3_U2633) );
  OAI21_X1 U19810 ( .B1(n16695), .B2(n17659), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16691) );
  OAI21_X1 U19811 ( .B1(n16692), .B2(n18909), .A(n16691), .ZN(P3_U2634) );
  AOI21_X1 U19812 ( .B1(n18931), .B2(n18933), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16693) );
  AOI22_X1 U19813 ( .A1(n19000), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16693), 
        .B2(n19066), .ZN(P3_U2635) );
  OAI21_X1 U19814 ( .B1(n18919), .B2(BS16), .A(n19005), .ZN(n19003) );
  OAI21_X1 U19815 ( .B1(n19005), .B2(n16716), .A(n19003), .ZN(P3_U2636) );
  NOR3_X1 U19816 ( .A1(n16695), .A2(n18841), .A3(n16694), .ZN(n18846) );
  NOR2_X1 U19817 ( .A1(n18846), .A2(n18904), .ZN(n19048) );
  OAI21_X1 U19818 ( .B1(n19048), .B2(n16697), .A(n16696), .ZN(P3_U2637) );
  NOR4_X1 U19819 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16701) );
  NOR4_X1 U19820 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16700) );
  NOR4_X1 U19821 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16699) );
  NOR4_X1 U19822 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16698) );
  NAND4_X1 U19823 ( .A1(n16701), .A2(n16700), .A3(n16699), .A4(n16698), .ZN(
        n16707) );
  NOR4_X1 U19824 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16705) );
  AOI211_X1 U19825 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16704) );
  NOR4_X1 U19826 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16703) );
  NOR4_X1 U19827 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16702) );
  NAND4_X1 U19828 ( .A1(n16705), .A2(n16704), .A3(n16703), .A4(n16702), .ZN(
        n16706) );
  NOR2_X1 U19829 ( .A1(n16707), .A2(n16706), .ZN(n19046) );
  INV_X1 U19830 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16709) );
  NOR3_X1 U19831 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16710) );
  OAI21_X1 U19832 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16710), .A(n19046), .ZN(
        n16708) );
  OAI21_X1 U19833 ( .B1(n19046), .B2(n16709), .A(n16708), .ZN(P3_U2638) );
  INV_X1 U19834 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19039) );
  INV_X1 U19835 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19004) );
  AOI21_X1 U19836 ( .B1(n19039), .B2(n19004), .A(n16710), .ZN(n16712) );
  INV_X1 U19837 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16711) );
  INV_X1 U19838 ( .A(n19046), .ZN(n19041) );
  AOI22_X1 U19839 ( .A1(n19046), .A2(n16712), .B1(n16711), .B2(n19041), .ZN(
        P3_U2639) );
  INV_X1 U19840 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18989) );
  INV_X1 U19841 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18986) );
  INV_X1 U19842 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18981) );
  AOI211_X1 U19843 ( .C1(n18924), .C2(n17658), .A(n19057), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n16714) );
  INV_X1 U19844 ( .A(n16714), .ZN(n18897) );
  INV_X1 U19845 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18979) );
  INV_X1 U19846 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18974) );
  INV_X1 U19847 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18975) );
  INV_X1 U19848 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18955) );
  INV_X1 U19849 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18945) );
  INV_X1 U19850 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18941) );
  INV_X1 U19851 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18935) );
  NOR2_X1 U19852 ( .A1(n19039), .A2(n18935), .ZN(n17066) );
  NAND2_X1 U19853 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n17066), .ZN(n17030) );
  INV_X1 U19854 ( .A(n17030), .ZN(n17034) );
  NAND2_X1 U19855 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17034), .ZN(n17022) );
  NOR2_X1 U19856 ( .A1(n18941), .A2(n17022), .ZN(n16994) );
  NAND2_X1 U19857 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16994), .ZN(n16998) );
  NOR2_X1 U19858 ( .A1(n18945), .A2(n16998), .ZN(n16991) );
  NAND2_X1 U19859 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16991), .ZN(n16965) );
  NAND2_X1 U19860 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16966) );
  NOR2_X1 U19861 ( .A1(n16965), .A2(n16966), .ZN(n16944) );
  NAND2_X1 U19862 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16944), .ZN(n16935) );
  NOR2_X1 U19863 ( .A1(n18955), .A2(n16935), .ZN(n16919) );
  NAND3_X1 U19864 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n16919), .ZN(n16908) );
  INV_X1 U19865 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18970) );
  INV_X1 U19866 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18967) );
  NAND3_X1 U19867 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n16858) );
  NOR3_X1 U19868 ( .A1(n18970), .A2(n18967), .A3(n16858), .ZN(n16844) );
  NAND2_X1 U19869 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16844), .ZN(n16829) );
  NOR4_X1 U19870 ( .A1(n18974), .A2(n18975), .A3(n16908), .A4(n16829), .ZN(
        n16805) );
  NAND2_X1 U19871 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16805), .ZN(n16793) );
  NOR2_X1 U19872 ( .A1(n18979), .A2(n16793), .ZN(n16727) );
  NAND2_X1 U19873 ( .A1(n17086), .A2(n16727), .ZN(n16792) );
  NOR2_X1 U19874 ( .A1(n18981), .A2(n16792), .ZN(n16778) );
  NAND2_X1 U19875 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16778), .ZN(n16767) );
  NOR3_X1 U19876 ( .A1(n18989), .A2(n18986), .A3(n16767), .ZN(n16751) );
  NAND2_X1 U19877 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16751), .ZN(n16733) );
  NAND2_X1 U19878 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n18993), .ZN(n16732) );
  NAND2_X1 U19879 ( .A1(n19056), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18780) );
  NOR2_X1 U19880 ( .A1(n18393), .A2(n17070), .ZN(n16986) );
  AOI211_X4 U19881 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n9969), .A(n16714), .B(
        n19071), .ZN(n17093) );
  AOI22_X1 U19882 ( .A1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n17076), .B1(
        P3_EBX_REG_31__SCAN_IN), .B2(n17093), .ZN(n16731) );
  NAND2_X1 U19883 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n9969), .ZN(n16715) );
  AOI211_X4 U19884 ( .C1(n16716), .C2(n19050), .A(n19071), .B(n16715), .ZN(
        n17092) );
  NOR3_X1 U19885 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17064) );
  NAND2_X1 U19886 ( .A1(n17064), .A2(n17055), .ZN(n17054) );
  NOR2_X1 U19887 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17054), .ZN(n17031) );
  NAND2_X1 U19888 ( .A1(n17031), .A2(n17026), .ZN(n17025) );
  NOR2_X1 U19889 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17025), .ZN(n17006) );
  NAND2_X1 U19890 ( .A1(n17006), .A2(n17404), .ZN(n17001) );
  NOR2_X1 U19891 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17001), .ZN(n16982) );
  INV_X1 U19892 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16973) );
  NAND2_X1 U19893 ( .A1(n16982), .A2(n16973), .ZN(n16972) );
  NOR2_X1 U19894 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16972), .ZN(n16959) );
  INV_X1 U19895 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16951) );
  NAND2_X1 U19896 ( .A1(n16959), .A2(n16951), .ZN(n16950) );
  NOR2_X1 U19897 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16950), .ZN(n16933) );
  INV_X1 U19898 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16923) );
  NAND2_X1 U19899 ( .A1(n16933), .A2(n16923), .ZN(n16922) );
  NOR2_X1 U19900 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16922), .ZN(n16909) );
  INV_X1 U19901 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16905) );
  NAND2_X1 U19902 ( .A1(n16909), .A2(n16905), .ZN(n16904) );
  NOR2_X1 U19903 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16904), .ZN(n16886) );
  NAND2_X1 U19904 ( .A1(n16886), .A2(n17260), .ZN(n16877) );
  NOR2_X1 U19905 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16877), .ZN(n16866) );
  INV_X1 U19906 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16853) );
  NAND2_X1 U19907 ( .A1(n16866), .A2(n16853), .ZN(n16852) );
  NOR2_X1 U19908 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16852), .ZN(n16841) );
  NAND2_X1 U19909 ( .A1(n16841), .A2(n16836), .ZN(n16835) );
  NOR2_X1 U19910 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16835), .ZN(n16816) );
  NAND2_X1 U19911 ( .A1(n16816), .A2(n16806), .ZN(n16812) );
  NOR2_X1 U19912 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16812), .ZN(n16797) );
  NAND2_X1 U19913 ( .A1(n16797), .A2(n17099), .ZN(n16789) );
  NOR2_X1 U19914 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16789), .ZN(n16775) );
  NAND2_X1 U19915 ( .A1(n16775), .A2(n17147), .ZN(n16770) );
  NOR2_X1 U19916 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16770), .ZN(n16755) );
  INV_X1 U19917 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17139) );
  NAND2_X1 U19918 ( .A1(n16755), .A2(n17139), .ZN(n16736) );
  NOR2_X1 U19919 ( .A1(n17082), .A2(n16736), .ZN(n16739) );
  INV_X1 U19920 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17104) );
  OR2_X1 U19921 ( .A1(n18077), .A2(n17719), .ZN(n16718) );
  AOI21_X1 U19922 ( .B1(n17711), .B2(n16718), .A(n16717), .ZN(n17720) );
  NAND2_X1 U19923 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17759), .ZN(
        n16725) );
  INV_X1 U19924 ( .A(n16725), .ZN(n16726) );
  NAND3_X1 U19925 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A3(n16726), .ZN(n17715) );
  NOR2_X1 U19926 ( .A1(n17748), .A2(n17715), .ZN(n16719) );
  OAI21_X1 U19927 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16719), .A(
        n16718), .ZN(n17737) );
  INV_X1 U19928 ( .A(n17737), .ZN(n16765) );
  AOI21_X1 U19929 ( .B1(n17748), .B2(n17715), .A(n16719), .ZN(n17751) );
  INV_X1 U19930 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17772) );
  NOR2_X1 U19931 ( .A1(n17772), .A2(n16725), .ZN(n16720) );
  OAI21_X1 U19932 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16720), .A(
        n17715), .ZN(n17760) );
  INV_X1 U19933 ( .A(n17760), .ZN(n16785) );
  INV_X1 U19934 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17788) );
  INV_X1 U19935 ( .A(n17802), .ZN(n17804) );
  NOR2_X1 U19936 ( .A1(n18077), .A2(n17804), .ZN(n16724) );
  NAND3_X1 U19937 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A3(n16724), .ZN(n17756) );
  AOI21_X1 U19938 ( .B1(n17788), .B2(n17756), .A(n16726), .ZN(n17785) );
  NAND2_X1 U19939 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16724), .ZN(
        n16722) );
  INV_X1 U19940 ( .A(n16722), .ZN(n16721) );
  OAI21_X1 U19941 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n16721), .A(
        n17756), .ZN(n17807) );
  INV_X1 U19942 ( .A(n17807), .ZN(n16821) );
  OAI21_X1 U19943 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n16724), .A(
        n16722), .ZN(n17813) );
  INV_X1 U19944 ( .A(n17813), .ZN(n16832) );
  NOR3_X1 U19945 ( .A1(n18077), .A2(n16723), .A3(n17834), .ZN(n17801) );
  INV_X1 U19946 ( .A(n17801), .ZN(n16850) );
  AOI21_X1 U19947 ( .B1(n17833), .B2(n16850), .A(n16724), .ZN(n17836) );
  INV_X1 U19948 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16997) );
  INV_X1 U19949 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16911) );
  NAND2_X1 U19950 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17985), .ZN(
        n17009) );
  INV_X1 U19951 ( .A(n17009), .ZN(n16996) );
  NAND2_X1 U19952 ( .A1(n17923), .A2(n16996), .ZN(n16945) );
  INV_X1 U19953 ( .A(n16945), .ZN(n17921) );
  NAND2_X1 U19954 ( .A1(n17920), .A2(n17921), .ZN(n16920) );
  NOR2_X1 U19955 ( .A1(n16911), .A2(n16920), .ZN(n17876) );
  NAND2_X1 U19956 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17876), .ZN(
        n16898) );
  INV_X1 U19957 ( .A(n16898), .ZN(n16879) );
  NAND2_X1 U19958 ( .A1(n16997), .A2(n16879), .ZN(n16899) );
  INV_X1 U19959 ( .A(n16899), .ZN(n16887) );
  NOR2_X1 U19960 ( .A1(n17836), .A2(n16840), .ZN(n16839) );
  NOR2_X1 U19961 ( .A1(n16839), .A2(n17048), .ZN(n16831) );
  NOR2_X1 U19962 ( .A1(n17785), .A2(n16809), .ZN(n16808) );
  NOR2_X1 U19963 ( .A1(n16808), .A2(n17048), .ZN(n16796) );
  OAI22_X1 U19964 ( .A1(n17772), .A2(n16726), .B1(n16725), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17769) );
  NOR2_X1 U19965 ( .A1(n16765), .A2(n16764), .ZN(n16763) );
  NOR2_X1 U19966 ( .A1(n16763), .A2(n17048), .ZN(n16757) );
  NOR2_X1 U19967 ( .A1(n17720), .A2(n16757), .ZN(n16756) );
  NOR2_X1 U19968 ( .A1(n16756), .A2(n17048), .ZN(n16745) );
  INV_X1 U19969 ( .A(n17070), .ZN(n18913) );
  NOR2_X1 U19970 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16733), .ZN(n16738) );
  INV_X1 U19971 ( .A(n16738), .ZN(n16729) );
  NAND4_X1 U19972 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(P3_REIP_REG_26__SCAN_IN), 
        .A3(n16727), .A4(n17094), .ZN(n16779) );
  NAND3_X1 U19973 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16728) );
  NAND2_X1 U19974 ( .A1(n17065), .A2(n17094), .ZN(n17091) );
  OAI21_X1 U19975 ( .B1(n16779), .B2(n16728), .A(n17091), .ZN(n16754) );
  AOI21_X1 U19976 ( .B1(n16729), .B2(n16754), .A(n18993), .ZN(n16730) );
  XNOR2_X1 U19977 ( .A(n16735), .B(n16734), .ZN(n16742) );
  NAND2_X1 U19978 ( .A1(n17092), .A2(n16736), .ZN(n16747) );
  OAI22_X1 U19979 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16747), .B1(n18995), 
        .B2(n16754), .ZN(n16737) );
  AOI211_X1 U19980 ( .C1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .C2(n17076), .A(
        n16738), .B(n16737), .ZN(n16741) );
  OAI21_X1 U19981 ( .B1(n17093), .B2(n16739), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16740) );
  OAI211_X1 U19982 ( .C1(n18913), .C2(n16742), .A(n16741), .B(n16740), .ZN(
        P3_U2641) );
  INV_X1 U19983 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18991) );
  AOI22_X1 U19984 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17076), .B1(
        n17093), .B2(P3_EBX_REG_29__SCAN_IN), .ZN(n16753) );
  INV_X1 U19985 ( .A(n16743), .ZN(n16744) );
  AOI211_X1 U19986 ( .C1(n16746), .C2(n16745), .A(n16744), .B(n18913), .ZN(
        n16750) );
  INV_X1 U19987 ( .A(n16755), .ZN(n16748) );
  AOI21_X1 U19988 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16748), .A(n16747), .ZN(
        n16749) );
  AOI211_X1 U19989 ( .C1(n16751), .C2(n18991), .A(n16750), .B(n16749), .ZN(
        n16752) );
  OAI211_X1 U19990 ( .C1(n18991), .C2(n16754), .A(n16753), .B(n16752), .ZN(
        P3_U2642) );
  OAI21_X1 U19991 ( .B1(n18986), .B2(n16779), .A(n17091), .ZN(n16766) );
  AOI22_X1 U19992 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17076), .B1(
        n17093), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16762) );
  AOI211_X1 U19993 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16770), .A(n16755), .B(
        n17082), .ZN(n16760) );
  NOR3_X1 U19994 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n18986), .A3(n16767), 
        .ZN(n16759) );
  AOI211_X1 U19995 ( .C1(n17720), .C2(n16757), .A(n16756), .B(n18913), .ZN(
        n16758) );
  NOR3_X1 U19996 ( .A1(n16760), .A2(n16759), .A3(n16758), .ZN(n16761) );
  OAI211_X1 U19997 ( .C1(n18989), .C2(n16766), .A(n16762), .B(n16761), .ZN(
        P3_U2643) );
  AOI22_X1 U19998 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17076), .B1(
        n17093), .B2(P3_EBX_REG_27__SCAN_IN), .ZN(n16773) );
  AOI211_X1 U19999 ( .C1(n16765), .C2(n16764), .A(n16763), .B(n18913), .ZN(
        n16769) );
  AOI21_X1 U20000 ( .B1(n16767), .B2(n18986), .A(n16766), .ZN(n16768) );
  NOR2_X1 U20001 ( .A1(n16769), .A2(n16768), .ZN(n16772) );
  OAI211_X1 U20002 ( .C1(n16775), .C2(n17147), .A(n17092), .B(n16770), .ZN(
        n16771) );
  NAND3_X1 U20003 ( .A1(n16773), .A2(n16772), .A3(n16771), .ZN(P3_U2644) );
  AOI22_X1 U20004 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17076), .B1(
        n17093), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16782) );
  INV_X1 U20005 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18983) );
  AOI211_X1 U20006 ( .C1(n17751), .C2(n16774), .A(n9757), .B(n18913), .ZN(
        n16777) );
  AOI211_X1 U20007 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16789), .A(n16775), .B(
        n17082), .ZN(n16776) );
  AOI211_X1 U20008 ( .C1(n16778), .C2(n18983), .A(n16777), .B(n16776), .ZN(
        n16781) );
  NAND3_X1 U20009 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n17091), .A3(n16779), 
        .ZN(n16780) );
  NAND3_X1 U20010 ( .A1(n16782), .A2(n16781), .A3(n16780), .ZN(P3_U2645) );
  AOI21_X1 U20011 ( .B1(n17086), .B2(n16793), .A(n17029), .ZN(n16815) );
  OAI21_X1 U20012 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n17065), .A(n16815), 
        .ZN(n16788) );
  AOI211_X1 U20013 ( .C1(n16785), .C2(n16784), .A(n16783), .B(n18913), .ZN(
        n16787) );
  INV_X1 U20014 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17758) );
  OAI22_X1 U20015 ( .A1(n17758), .A2(n17050), .B1(n17083), .B2(n17099), .ZN(
        n16786) );
  AOI211_X1 U20016 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n16788), .A(n16787), 
        .B(n16786), .ZN(n16791) );
  OAI211_X1 U20017 ( .C1(n16797), .C2(n17099), .A(n17092), .B(n16789), .ZN(
        n16790) );
  OAI211_X1 U20018 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n16792), .A(n16791), 
        .B(n16790), .ZN(P3_U2646) );
  AOI22_X1 U20019 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17076), .B1(
        n17093), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n16802) );
  NOR2_X1 U20020 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17065), .ZN(n16800) );
  INV_X1 U20021 ( .A(n16793), .ZN(n16803) );
  INV_X1 U20022 ( .A(n16794), .ZN(n16795) );
  AOI211_X1 U20023 ( .C1(n17769), .C2(n16796), .A(n16795), .B(n18913), .ZN(
        n16799) );
  AOI211_X1 U20024 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16812), .A(n16797), .B(
        n17082), .ZN(n16798) );
  AOI211_X1 U20025 ( .C1(n16800), .C2(n16803), .A(n16799), .B(n16798), .ZN(
        n16801) );
  OAI211_X1 U20026 ( .C1(n16815), .C2(n18979), .A(n16802), .B(n16801), .ZN(
        P3_U2647) );
  INV_X1 U20027 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18978) );
  NOR2_X1 U20028 ( .A1(n16803), .A2(n17065), .ZN(n16804) );
  AOI22_X1 U20029 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17076), .B1(
        n16805), .B2(n16804), .ZN(n16814) );
  NOR2_X1 U20030 ( .A1(n16816), .A2(n16806), .ZN(n16807) );
  OAI22_X1 U20031 ( .A1(n17082), .A2(n16807), .B1(n17083), .B2(n16806), .ZN(
        n16811) );
  AOI211_X1 U20032 ( .C1(n17785), .C2(n16809), .A(n16808), .B(n18913), .ZN(
        n16810) );
  AOI21_X1 U20033 ( .B1(n16812), .B2(n16811), .A(n16810), .ZN(n16813) );
  OAI211_X1 U20034 ( .C1(n16815), .C2(n18978), .A(n16814), .B(n16813), .ZN(
        P3_U2648) );
  INV_X1 U20035 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16826) );
  AOI211_X1 U20036 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16835), .A(n16816), .B(
        n17082), .ZN(n16817) );
  AOI21_X1 U20037 ( .B1(n17076), .B2(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16817), .ZN(n16825) );
  NOR3_X1 U20038 ( .A1(n17029), .A2(n16829), .A3(n16908), .ZN(n16849) );
  INV_X1 U20039 ( .A(n17091), .ZN(n16818) );
  AOI21_X1 U20040 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n16849), .A(n16818), 
        .ZN(n16827) );
  NOR3_X1 U20041 ( .A1(n18974), .A2(n16829), .A3(n16897), .ZN(n16823) );
  AOI211_X1 U20042 ( .C1(n16821), .C2(n16820), .A(n16819), .B(n18913), .ZN(
        n16822) );
  AOI221_X1 U20043 ( .B1(n16827), .B2(P3_REIP_REG_22__SCAN_IN), .C1(n16823), 
        .C2(n18975), .A(n16822), .ZN(n16824) );
  OAI211_X1 U20044 ( .C1(n17083), .C2(n16826), .A(n16825), .B(n16824), .ZN(
        P3_U2649) );
  INV_X1 U20045 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17816) );
  INV_X1 U20046 ( .A(n16827), .ZN(n16828) );
  AOI221_X1 U20047 ( .B1(n16829), .B2(n18974), .C1(n16897), .C2(n18974), .A(
        n16828), .ZN(n16834) );
  AOI211_X1 U20048 ( .C1(n16832), .C2(n16831), .A(n16830), .B(n18913), .ZN(
        n16833) );
  AOI211_X1 U20049 ( .C1(P3_EBX_REG_21__SCAN_IN), .C2(n17093), .A(n16834), .B(
        n16833), .ZN(n16838) );
  OAI211_X1 U20050 ( .C1(n16841), .C2(n16836), .A(n17092), .B(n16835), .ZN(
        n16837) );
  OAI211_X1 U20051 ( .C1(n17050), .C2(n17816), .A(n16838), .B(n16837), .ZN(
        P3_U2650) );
  NAND2_X1 U20052 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n17091), .ZN(n16848) );
  AOI22_X1 U20053 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17076), .B1(
        n17093), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n16847) );
  NOR2_X1 U20054 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16897), .ZN(n16845) );
  AOI211_X1 U20055 ( .C1(n17836), .C2(n16840), .A(n16839), .B(n18913), .ZN(
        n16843) );
  AOI211_X1 U20056 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16852), .A(n16841), .B(
        n17082), .ZN(n16842) );
  AOI211_X1 U20057 ( .C1(n16845), .C2(n16844), .A(n16843), .B(n16842), .ZN(
        n16846) );
  OAI211_X1 U20058 ( .C1(n16849), .C2(n16848), .A(n16847), .B(n16846), .ZN(
        P3_U2651) );
  OAI21_X1 U20059 ( .B1(n16858), .B2(n16915), .A(n17091), .ZN(n16873) );
  NOR2_X1 U20060 ( .A1(n17083), .A2(n16853), .ZN(n16857) );
  NAND2_X1 U20061 ( .A1(n17831), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17843) );
  NOR2_X1 U20062 ( .A1(n18077), .A2(n17843), .ZN(n17842) );
  NAND2_X1 U20063 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17842), .ZN(
        n16862) );
  OAI21_X1 U20064 ( .B1(n16862), .B2(n16899), .A(n17018), .ZN(n16864) );
  INV_X1 U20065 ( .A(n16862), .ZN(n16851) );
  OAI21_X1 U20066 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16851), .A(
        n16850), .ZN(n17847) );
  XNOR2_X1 U20067 ( .A(n16864), .B(n17847), .ZN(n16855) );
  OAI211_X1 U20068 ( .C1(n16866), .C2(n16853), .A(n17092), .B(n16852), .ZN(
        n16854) );
  OAI211_X1 U20069 ( .C1(n18913), .C2(n16855), .A(n18380), .B(n16854), .ZN(
        n16856) );
  AOI211_X1 U20070 ( .C1(n17076), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16857), .B(n16856), .ZN(n16860) );
  NOR2_X1 U20071 ( .A1(n16858), .A2(n16897), .ZN(n16861) );
  OAI221_X1 U20072 ( .B1(P3_REIP_REG_19__SCAN_IN), .B2(P3_REIP_REG_18__SCAN_IN), .C1(n18970), .C2(n18967), .A(n16861), .ZN(n16859) );
  OAI211_X1 U20073 ( .C1(n16873), .C2(n18970), .A(n16860), .B(n16859), .ZN(
        P3_U2652) );
  INV_X1 U20074 ( .A(n16861), .ZN(n16872) );
  INV_X1 U20075 ( .A(n16986), .ZN(n16964) );
  OAI21_X1 U20076 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17842), .A(
        n16862), .ZN(n17853) );
  INV_X1 U20077 ( .A(n17853), .ZN(n16865) );
  INV_X1 U20078 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17856) );
  AOI21_X1 U20079 ( .B1(n16887), .B2(n17856), .A(n17048), .ZN(n16863) );
  OAI221_X1 U20080 ( .B1(n16865), .B2(n16864), .C1(n17853), .C2(n16863), .A(
        n18380), .ZN(n16870) );
  AOI211_X1 U20081 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16877), .A(n16866), .B(
        n17082), .ZN(n16869) );
  OAI22_X1 U20082 ( .A1(n17856), .A2(n17050), .B1(n17083), .B2(n16867), .ZN(
        n16868) );
  AOI211_X1 U20083 ( .C1(n16964), .C2(n16870), .A(n16869), .B(n16868), .ZN(
        n16871) );
  OAI221_X1 U20084 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16872), .C1(n18967), 
        .C2(n16873), .A(n16871), .ZN(P3_U2653) );
  INV_X1 U20085 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18963) );
  INV_X1 U20086 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18961) );
  NOR3_X1 U20087 ( .A1(n18963), .A2(n18961), .A3(n16897), .ZN(n16876) );
  INV_X1 U20088 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18965) );
  INV_X1 U20089 ( .A(n16873), .ZN(n16875) );
  INV_X1 U20090 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17865) );
  OAI22_X1 U20091 ( .A1(n17865), .A2(n17050), .B1(n17083), .B2(n17260), .ZN(
        n16874) );
  AOI221_X1 U20092 ( .B1(n16876), .B2(n18965), .C1(n16875), .C2(
        P3_REIP_REG_17__SCAN_IN), .A(n16874), .ZN(n16884) );
  OAI211_X1 U20093 ( .C1(n16886), .C2(n17260), .A(n17092), .B(n16877), .ZN(
        n16883) );
  NAND2_X1 U20094 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17831), .ZN(
        n16878) );
  AOI21_X1 U20095 ( .B1(n17865), .B2(n16878), .A(n17842), .ZN(n17867) );
  OAI21_X1 U20096 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16879), .A(
        n16878), .ZN(n17883) );
  AOI21_X1 U20097 ( .B1(n16887), .B2(n17883), .A(n17048), .ZN(n16881) );
  AOI21_X1 U20098 ( .B1(n17867), .B2(n16881), .A(n18913), .ZN(n16880) );
  OAI21_X1 U20099 ( .B1(n17867), .B2(n16881), .A(n16880), .ZN(n16882) );
  NAND4_X1 U20100 ( .A1(n16884), .A2(n18380), .A3(n16883), .A4(n16882), .ZN(
        P3_U2654) );
  NAND2_X1 U20101 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16885), .ZN(n16895) );
  AOI22_X1 U20102 ( .A1(n16885), .A2(n18961), .B1(n17091), .B2(n16915), .ZN(
        n16896) );
  AOI211_X1 U20103 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16904), .A(n16886), .B(
        n17082), .ZN(n16893) );
  NAND2_X1 U20104 ( .A1(n17018), .A2(n16899), .ZN(n16889) );
  OAI21_X1 U20105 ( .B1(n16887), .B2(n17048), .A(n17883), .ZN(n16888) );
  OAI211_X1 U20106 ( .C1(n16889), .C2(n17883), .A(n17070), .B(n16888), .ZN(
        n16890) );
  OAI211_X1 U20107 ( .C1(n16891), .C2(n17050), .A(n18380), .B(n16890), .ZN(
        n16892) );
  AOI211_X1 U20108 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17093), .A(n16893), .B(
        n16892), .ZN(n16894) );
  OAI221_X1 U20109 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(n16895), .C1(n18963), 
        .C2(n16896), .A(n16894), .ZN(P3_U2655) );
  AOI21_X1 U20110 ( .B1(n18961), .B2(n16897), .A(n16896), .ZN(n16903) );
  NOR2_X1 U20111 ( .A1(n18913), .A2(n17018), .ZN(n16978) );
  INV_X1 U20112 ( .A(n16978), .ZN(n17062) );
  OAI21_X1 U20113 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17876), .A(
        n16898), .ZN(n17894) );
  NAND2_X1 U20114 ( .A1(n17018), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16957) );
  NAND2_X1 U20115 ( .A1(n17070), .A2(n16957), .ZN(n17088) );
  AOI211_X1 U20116 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n17062), .A(
        n17894), .B(n17088), .ZN(n16902) );
  NOR2_X1 U20117 ( .A1(n17048), .A2(n18913), .ZN(n17077) );
  NAND3_X1 U20118 ( .A1(n17077), .A2(n16899), .A3(n17894), .ZN(n16900) );
  OAI211_X1 U20119 ( .C1(n17083), .C2(n16905), .A(n18380), .B(n16900), .ZN(
        n16901) );
  NOR3_X1 U20120 ( .A1(n16903), .A2(n16902), .A3(n16901), .ZN(n16907) );
  OAI211_X1 U20121 ( .C1(n16909), .C2(n16905), .A(n17092), .B(n16904), .ZN(
        n16906) );
  OAI211_X1 U20122 ( .C1(n17050), .C2(n17897), .A(n16907), .B(n16906), .ZN(
        P3_U2656) );
  AOI21_X1 U20123 ( .B1(n17086), .B2(n16908), .A(n17029), .ZN(n16918) );
  INV_X1 U20124 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18960) );
  AOI211_X1 U20125 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16922), .A(n16909), .B(
        n17082), .ZN(n16914) );
  AOI21_X1 U20126 ( .B1(n16911), .B2(n16920), .A(n17876), .ZN(n17906) );
  OAI21_X1 U20127 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16920), .A(
        n17018), .ZN(n16926) );
  OAI21_X1 U20128 ( .B1(n17906), .B2(n16926), .A(n18380), .ZN(n16910) );
  AOI21_X1 U20129 ( .B1(n17906), .B2(n16926), .A(n16910), .ZN(n16912) );
  OAI22_X1 U20130 ( .A1(n16986), .A2(n16912), .B1(n16911), .B2(n17050), .ZN(
        n16913) );
  AOI211_X1 U20131 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17093), .A(n16914), .B(
        n16913), .ZN(n16917) );
  NAND4_X1 U20132 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17086), .A3(n16919), 
        .A4(n16915), .ZN(n16916) );
  OAI211_X1 U20133 ( .C1(n16918), .C2(n18960), .A(n16917), .B(n16916), .ZN(
        P3_U2657) );
  NAND2_X1 U20134 ( .A1(n17086), .A2(n16919), .ZN(n16932) );
  AOI22_X1 U20135 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17076), .B1(
        n17093), .B2(P3_EBX_REG_13__SCAN_IN), .ZN(n16931) );
  AOI21_X1 U20136 ( .B1(n17086), .B2(n16935), .A(n17029), .ZN(n16954) );
  OAI21_X1 U20137 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n17065), .A(n16954), 
        .ZN(n16929) );
  NAND2_X1 U20138 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17921), .ZN(
        n16921) );
  INV_X1 U20139 ( .A(n16921), .ZN(n16938) );
  OAI21_X1 U20140 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16938), .A(
        n16920), .ZN(n17925) );
  AOI211_X1 U20141 ( .C1(n17018), .C2(n16921), .A(n17925), .B(n17088), .ZN(
        n16928) );
  NAND2_X1 U20142 ( .A1(n17070), .A2(n17925), .ZN(n16925) );
  OAI211_X1 U20143 ( .C1(n16933), .C2(n16923), .A(n17092), .B(n16922), .ZN(
        n16924) );
  OAI211_X1 U20144 ( .C1(n16926), .C2(n16925), .A(n18380), .B(n16924), .ZN(
        n16927) );
  AOI211_X1 U20145 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16929), .A(n16928), 
        .B(n16927), .ZN(n16930) );
  OAI211_X1 U20146 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16932), .A(n16931), 
        .B(n16930), .ZN(P3_U2658) );
  AOI211_X1 U20147 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16950), .A(n16933), .B(
        n17082), .ZN(n16937) );
  NAND2_X1 U20148 ( .A1(n17086), .A2(n18955), .ZN(n16934) );
  OAI22_X1 U20149 ( .A1(n18955), .A2(n16954), .B1(n16935), .B2(n16934), .ZN(
        n16936) );
  AOI211_X1 U20150 ( .C1(n17076), .C2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16937), .B(n16936), .ZN(n16942) );
  AOI21_X1 U20151 ( .B1(n17939), .B2(n16945), .A(n16938), .ZN(n17942) );
  INV_X1 U20152 ( .A(n17877), .ZN(n17919) );
  NAND2_X1 U20153 ( .A1(n16997), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17035) );
  INV_X1 U20154 ( .A(n17035), .ZN(n17071) );
  AOI21_X1 U20155 ( .B1(n17919), .B2(n17071), .A(n17048), .ZN(n16939) );
  XOR2_X1 U20156 ( .A(n17942), .B(n16939), .Z(n16940) );
  AOI21_X1 U20157 ( .B1(n16940), .B2(n17070), .A(n18393), .ZN(n16941) );
  OAI211_X1 U20158 ( .C1(n16943), .C2(n17083), .A(n16942), .B(n16941), .ZN(
        P3_U2659) );
  AOI21_X1 U20159 ( .B1(n17086), .B2(n16944), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16955) );
  INV_X1 U20160 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16975) );
  NAND2_X1 U20161 ( .A1(n17986), .A2(n16996), .ZN(n16983) );
  NOR2_X1 U20162 ( .A1(n16975), .A2(n16983), .ZN(n16974) );
  NAND2_X1 U20163 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16974), .ZN(
        n16956) );
  OAI21_X1 U20164 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16956), .A(
        n17018), .ZN(n16947) );
  INV_X1 U20165 ( .A(n16956), .ZN(n16946) );
  OAI21_X1 U20166 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16946), .A(
        n16945), .ZN(n17952) );
  XNOR2_X1 U20167 ( .A(n16947), .B(n17952), .ZN(n16948) );
  OAI22_X1 U20168 ( .A1(n17083), .A2(n16951), .B1(n18913), .B2(n16948), .ZN(
        n16949) );
  AOI211_X1 U20169 ( .C1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n17076), .A(
        n18393), .B(n16949), .ZN(n16953) );
  OAI211_X1 U20170 ( .C1(n16959), .C2(n16951), .A(n17092), .B(n16950), .ZN(
        n16952) );
  OAI211_X1 U20171 ( .C1(n16955), .C2(n16954), .A(n16953), .B(n16952), .ZN(
        P3_U2660) );
  AOI21_X1 U20172 ( .B1(n17086), .B2(n16965), .A(n17029), .ZN(n16969) );
  INV_X1 U20173 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18951) );
  OAI21_X1 U20174 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16974), .A(
        n16956), .ZN(n17971) );
  OAI21_X1 U20175 ( .B1(n16974), .B2(n17048), .A(n16957), .ZN(n16976) );
  AOI21_X1 U20176 ( .B1(n17971), .B2(n16976), .A(n18393), .ZN(n16958) );
  OAI21_X1 U20177 ( .B1(n17971), .B2(n16976), .A(n16958), .ZN(n16963) );
  AOI211_X1 U20178 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16972), .A(n16959), .B(
        n17082), .ZN(n16962) );
  INV_X1 U20179 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17965) );
  OAI22_X1 U20180 ( .A1(n17965), .A2(n17050), .B1(n17083), .B2(n16960), .ZN(
        n16961) );
  AOI211_X1 U20181 ( .C1(n16964), .C2(n16963), .A(n16962), .B(n16961), .ZN(
        n16968) );
  NOR2_X1 U20182 ( .A1(n17065), .A2(n16965), .ZN(n16971) );
  OAI211_X1 U20183 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(P3_REIP_REG_9__SCAN_IN), 
        .A(n16971), .B(n16966), .ZN(n16967) );
  OAI211_X1 U20184 ( .C1(n16969), .C2(n18951), .A(n16968), .B(n16967), .ZN(
        P3_U2661) );
  INV_X1 U20185 ( .A(n16969), .ZN(n16990) );
  INV_X1 U20186 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18949) );
  OAI22_X1 U20187 ( .A1(n16975), .A2(n17050), .B1(n17083), .B2(n16973), .ZN(
        n16970) );
  AOI221_X1 U20188 ( .B1(n16990), .B2(P3_REIP_REG_9__SCAN_IN), .C1(n16971), 
        .C2(n18949), .A(n16970), .ZN(n16981) );
  OAI211_X1 U20189 ( .C1(n16982), .C2(n16973), .A(n17092), .B(n16972), .ZN(
        n16980) );
  AOI21_X1 U20190 ( .B1(n16975), .B2(n16983), .A(n16974), .ZN(n17974) );
  AND3_X1 U20191 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17985), .A3(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16995) );
  NAND2_X1 U20192 ( .A1(n16995), .A2(n16997), .ZN(n16984) );
  AOI221_X1 U20193 ( .B1(n17988), .B2(n17974), .C1(n16984), .C2(n17974), .A(
        n18913), .ZN(n16977) );
  OAI22_X1 U20194 ( .A1(n16978), .A2(n16977), .B1(n17974), .B2(n16976), .ZN(
        n16979) );
  NAND4_X1 U20195 ( .A1(n16981), .A2(n18380), .A3(n16980), .A4(n16979), .ZN(
        P3_U2662) );
  AOI211_X1 U20196 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17001), .A(n16982), .B(
        n17082), .ZN(n16989) );
  OAI21_X1 U20197 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16995), .A(
        n16983), .ZN(n17989) );
  NAND2_X1 U20198 ( .A1(n17018), .A2(n16984), .ZN(n16985) );
  XNOR2_X1 U20199 ( .A(n17989), .B(n16985), .ZN(n16987) );
  AOI21_X1 U20200 ( .B1(n16987), .B2(n18380), .A(n16986), .ZN(n16988) );
  AOI211_X1 U20201 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17093), .A(n16989), .B(
        n16988), .ZN(n16993) );
  OAI221_X1 U20202 ( .B1(P3_REIP_REG_8__SCAN_IN), .B2(n17086), .C1(
        P3_REIP_REG_8__SCAN_IN), .C2(n16991), .A(n16990), .ZN(n16992) );
  OAI211_X1 U20203 ( .C1(n17050), .C2(n17988), .A(n16993), .B(n16992), .ZN(
        P3_U2663) );
  INV_X1 U20204 ( .A(n16994), .ZN(n17016) );
  NOR3_X1 U20205 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17065), .A3(n17016), .ZN(
        n17008) );
  OAI21_X1 U20206 ( .B1(n16994), .B2(n17065), .A(n17094), .ZN(n17024) );
  AOI21_X1 U20207 ( .B1(n18004), .B2(n17009), .A(n16995), .ZN(n18008) );
  AOI21_X1 U20208 ( .B1(n16997), .B2(n16996), .A(n17048), .ZN(n17010) );
  XOR2_X1 U20209 ( .A(n18008), .B(n17010), .Z(n17000) );
  NOR3_X1 U20210 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n17065), .A3(n16998), .ZN(
        n16999) );
  AOI211_X1 U20211 ( .C1(n17070), .C2(n17000), .A(n18393), .B(n16999), .ZN(
        n17003) );
  OAI211_X1 U20212 ( .C1(n17006), .C2(n17404), .A(n17092), .B(n17001), .ZN(
        n17002) );
  OAI211_X1 U20213 ( .C1(n17404), .C2(n17083), .A(n17003), .B(n17002), .ZN(
        n17004) );
  AOI221_X1 U20214 ( .B1(n17008), .B2(P3_REIP_REG_7__SCAN_IN), .C1(n17024), 
        .C2(P3_REIP_REG_7__SCAN_IN), .A(n17004), .ZN(n17005) );
  OAI21_X1 U20215 ( .B1(n18004), .B2(n17050), .A(n17005), .ZN(P3_U2664) );
  AOI211_X1 U20216 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17025), .A(n17006), .B(
        n17082), .ZN(n17007) );
  AOI211_X1 U20217 ( .C1(n17076), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n17008), .B(n17007), .ZN(n17015) );
  NOR2_X1 U20218 ( .A1(n18077), .A2(n18014), .ZN(n17017) );
  OAI21_X1 U20219 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17017), .A(
        n17009), .ZN(n18023) );
  AOI211_X1 U20220 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n17018), .A(
        n18023), .B(n17088), .ZN(n17013) );
  NAND3_X1 U20221 ( .A1(n17070), .A2(n17010), .A3(n18023), .ZN(n17011) );
  OAI211_X1 U20222 ( .C1(n17083), .C2(n17403), .A(n18380), .B(n17011), .ZN(
        n17012) );
  AOI211_X1 U20223 ( .C1(P3_REIP_REG_6__SCAN_IN), .C2(n17024), .A(n17013), .B(
        n17012), .ZN(n17014) );
  NAND2_X1 U20224 ( .A1(n17015), .A2(n17014), .ZN(P3_U2665) );
  NAND2_X1 U20225 ( .A1(n17086), .A2(n17016), .ZN(n17021) );
  NAND2_X1 U20226 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18024), .ZN(
        n17032) );
  AOI21_X1 U20227 ( .B1(n9946), .B2(n17032), .A(n17017), .ZN(n18029) );
  OAI21_X1 U20228 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17032), .A(
        n17018), .ZN(n17036) );
  XNOR2_X1 U20229 ( .A(n18029), .B(n17036), .ZN(n17019) );
  AOI22_X1 U20230 ( .A1(n17093), .A2(P3_EBX_REG_5__SCAN_IN), .B1(n17070), .B2(
        n17019), .ZN(n17020) );
  OAI211_X1 U20231 ( .C1(n17022), .C2(n17021), .A(n17020), .B(n18380), .ZN(
        n17023) );
  AOI21_X1 U20232 ( .B1(P3_REIP_REG_5__SCAN_IN), .B2(n17024), .A(n17023), .ZN(
        n17028) );
  OAI211_X1 U20233 ( .C1(n17031), .C2(n17026), .A(n17092), .B(n17025), .ZN(
        n17027) );
  OAI211_X1 U20234 ( .C1(n17050), .C2(n9946), .A(n17028), .B(n17027), .ZN(
        P3_U2666) );
  INV_X1 U20235 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18939) );
  AOI21_X1 U20236 ( .B1(n17086), .B2(n17030), .A(n17029), .ZN(n17058) );
  AOI211_X1 U20237 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17054), .A(n17031), .B(
        n17082), .ZN(n17043) );
  NOR2_X1 U20238 ( .A1(n18077), .A2(n18040), .ZN(n17047) );
  OAI21_X1 U20239 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17047), .A(
        n17032), .ZN(n18043) );
  NOR2_X1 U20240 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17065), .ZN(n17033) );
  AOI22_X1 U20241 ( .A1(n17093), .A2(P3_EBX_REG_4__SCAN_IN), .B1(n17034), .B2(
        n17033), .ZN(n17041) );
  INV_X1 U20242 ( .A(n18043), .ZN(n17037) );
  OR2_X1 U20243 ( .A1(n18040), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18047) );
  OAI22_X1 U20244 ( .A1(n17037), .A2(n17036), .B1(n17035), .B2(n18047), .ZN(
        n17039) );
  NOR2_X1 U20245 ( .A1(n18411), .A2(n19069), .ZN(n17090) );
  INV_X1 U20246 ( .A(n17090), .ZN(n17079) );
  AOI21_X1 U20247 ( .B1(n17268), .B2(n18849), .A(n17079), .ZN(n17038) );
  AOI211_X1 U20248 ( .C1(n17070), .C2(n17039), .A(n18393), .B(n17038), .ZN(
        n17040) );
  OAI211_X1 U20249 ( .C1(n18043), .C2(n17062), .A(n17041), .B(n17040), .ZN(
        n17042) );
  AOI211_X1 U20250 ( .C1(n17076), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n17043), .B(n17042), .ZN(n17044) );
  OAI21_X1 U20251 ( .B1(n18939), .B2(n17058), .A(n17044), .ZN(P3_U2667) );
  AOI21_X1 U20252 ( .B1(n17086), .B2(n17066), .A(P3_REIP_REG_3__SCAN_IN), .ZN(
        n17059) );
  INV_X1 U20253 ( .A(n18850), .ZN(n18869) );
  NOR2_X1 U20254 ( .A1(n17045), .A2(n18869), .ZN(n18854) );
  INV_X1 U20255 ( .A(n18854), .ZN(n17046) );
  AOI21_X1 U20256 ( .B1(n19014), .B2(n17046), .A(n13117), .ZN(n19012) );
  INV_X1 U20257 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17051) );
  NAND2_X1 U20258 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17061) );
  AOI21_X1 U20259 ( .B1(n17051), .B2(n17061), .A(n17047), .ZN(n18054) );
  AOI21_X1 U20260 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17071), .A(
        n17048), .ZN(n17069) );
  OAI21_X1 U20261 ( .B1(n18054), .B2(n17069), .A(n17070), .ZN(n17049) );
  AOI21_X1 U20262 ( .B1(n18054), .B2(n17069), .A(n17049), .ZN(n17053) );
  OAI22_X1 U20263 ( .A1(n17051), .A2(n17050), .B1(n17083), .B2(n17055), .ZN(
        n17052) );
  AOI211_X1 U20264 ( .C1(n19012), .C2(n17090), .A(n17053), .B(n17052), .ZN(
        n17057) );
  OAI211_X1 U20265 ( .C1(n17064), .C2(n17055), .A(n17092), .B(n17054), .ZN(
        n17056) );
  OAI211_X1 U20266 ( .C1(n17059), .C2(n17058), .A(n17057), .B(n17056), .ZN(
        P3_U2668) );
  NAND2_X1 U20267 ( .A1(n19025), .A2(n17060), .ZN(n18852) );
  OAI21_X1 U20268 ( .B1(n18869), .B2(n17045), .A(n18852), .ZN(n18879) );
  INV_X1 U20269 ( .A(n18879), .ZN(n19021) );
  AOI22_X1 U20270 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n17076), .B1(
        n19021), .B2(n17090), .ZN(n17075) );
  OAI21_X1 U20271 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17061), .ZN(n18064) );
  OAI22_X1 U20272 ( .A1(n18935), .A2(n17094), .B1(n18064), .B2(n17062), .ZN(
        n17063) );
  INV_X1 U20273 ( .A(n17063), .ZN(n17074) );
  INV_X1 U20274 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17434) );
  INV_X1 U20275 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17428) );
  NAND2_X1 U20276 ( .A1(n17434), .A2(n17428), .ZN(n17081) );
  AOI211_X1 U20277 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17081), .A(n17064), .B(
        n17082), .ZN(n17068) );
  AOI211_X1 U20278 ( .C1(n19039), .C2(n18935), .A(n17066), .B(n17065), .ZN(
        n17067) );
  AOI211_X1 U20279 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17093), .A(n17068), .B(
        n17067), .ZN(n17073) );
  OAI211_X1 U20280 ( .C1(n17071), .C2(n18064), .A(n17070), .B(n17069), .ZN(
        n17072) );
  NAND4_X1 U20281 ( .A1(n17075), .A2(n17074), .A3(n17073), .A4(n17072), .ZN(
        P3_U2669) );
  AOI211_X1 U20282 ( .C1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n17077), .A(
        n17076), .B(n18077), .ZN(n17089) );
  NOR2_X1 U20283 ( .A1(n10055), .A2(n17078), .ZN(n19028) );
  INV_X1 U20284 ( .A(n19028), .ZN(n18862) );
  OAI22_X1 U20285 ( .A1(n19039), .A2(n17094), .B1(n18862), .B2(n17079), .ZN(
        n17085) );
  NOR2_X1 U20286 ( .A1(n17434), .A2(n17428), .ZN(n17421) );
  INV_X1 U20287 ( .A(n17421), .ZN(n17080) );
  NAND2_X1 U20288 ( .A1(n17081), .A2(n17080), .ZN(n17430) );
  OAI22_X1 U20289 ( .A1(n17083), .A2(n17428), .B1(n17082), .B2(n17430), .ZN(
        n17084) );
  AOI211_X1 U20290 ( .C1(n17086), .C2(n19039), .A(n17085), .B(n17084), .ZN(
        n17087) );
  OAI221_X1 U20291 ( .B1(n17089), .B2(n18077), .C1(n17089), .C2(n17088), .A(
        n17087), .ZN(P3_U2670) );
  AOI22_X1 U20292 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n17091), .B1(n17090), 
        .B2(n17045), .ZN(n17097) );
  OAI21_X1 U20293 ( .B1(n17093), .B2(n17092), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n17096) );
  NAND3_X1 U20294 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19009), .A3(
        n17094), .ZN(n17095) );
  NAND3_X1 U20295 ( .A1(n17097), .A2(n17096), .A3(n17095), .ZN(P3_U2671) );
  NAND4_X1 U20296 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n17098)
         );
  NOR3_X1 U20297 ( .A1(n17139), .A2(n17099), .A3(n17098), .ZN(n17100) );
  NAND4_X1 U20298 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17216), .A3(n17140), 
        .A4(n17100), .ZN(n17103) );
  NOR2_X1 U20299 ( .A1(n17104), .A2(n17103), .ZN(n17134) );
  NAND2_X1 U20300 ( .A1(n17423), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17102) );
  NAND2_X1 U20301 ( .A1(n17134), .A2(n17527), .ZN(n17101) );
  OAI22_X1 U20302 ( .A1(n17134), .A2(n17102), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17101), .ZN(P3_U2672) );
  NAND2_X1 U20303 ( .A1(n17104), .A2(n17103), .ZN(n17105) );
  NAND2_X1 U20304 ( .A1(n17105), .A2(n17423), .ZN(n17133) );
  OAI22_X1 U20305 ( .A1(n17396), .A2(n17106), .B1(n17367), .B2(n17175), .ZN(
        n17117) );
  AOI22_X1 U20306 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17375), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17115) );
  AOI22_X1 U20307 ( .A1(n17384), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17114) );
  OAI22_X1 U20308 ( .A1(n17380), .A2(n17107), .B1(n12918), .B2(n17179), .ZN(
        n17112) );
  AOI22_X1 U20309 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17110) );
  AOI22_X1 U20310 ( .A1(n12945), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17381), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17109) );
  AOI22_X1 U20311 ( .A1(n13039), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17392), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17108) );
  NAND3_X1 U20312 ( .A1(n17110), .A2(n17109), .A3(n17108), .ZN(n17111) );
  AOI211_X1 U20313 ( .C1(n17320), .C2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n17112), .B(n17111), .ZN(n17113) );
  NAND3_X1 U20314 ( .A1(n17115), .A2(n17114), .A3(n17113), .ZN(n17116) );
  AOI211_X1 U20315 ( .C1(n17306), .C2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        n17117), .B(n17116), .ZN(n17137) );
  NOR2_X1 U20316 ( .A1(n17137), .A2(n17136), .ZN(n17135) );
  AOI22_X1 U20317 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17131) );
  AOI22_X1 U20318 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12945), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17118) );
  OAI21_X1 U20319 ( .B1(n17120), .B2(n17119), .A(n17118), .ZN(n17129) );
  AOI22_X1 U20320 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17126) );
  INV_X1 U20321 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17123) );
  AOI22_X1 U20322 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17122) );
  AOI22_X1 U20323 ( .A1(n17352), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17121) );
  OAI211_X1 U20324 ( .C1(n17380), .C2(n17123), .A(n17122), .B(n17121), .ZN(
        n17124) );
  AOI21_X1 U20325 ( .B1(n17374), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A(
        n17124), .ZN(n17125) );
  OAI211_X1 U20326 ( .C1(n17358), .C2(n17127), .A(n17126), .B(n17125), .ZN(
        n17128) );
  AOI211_X1 U20327 ( .C1(n17217), .C2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n17129), .B(n17128), .ZN(n17130) );
  OAI211_X1 U20328 ( .C1(n17287), .C2(n17284), .A(n17131), .B(n17130), .ZN(
        n17132) );
  XNOR2_X1 U20329 ( .A(n17135), .B(n17132), .ZN(n17447) );
  OAI22_X1 U20330 ( .A1(n17134), .A2(n17133), .B1(n17447), .B2(n17423), .ZN(
        P3_U2673) );
  AOI21_X1 U20331 ( .B1(n17137), .B2(n17136), .A(n17135), .ZN(n17451) );
  AOI22_X1 U20332 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17138), .B1(n17451), 
        .B2(n17432), .ZN(n17142) );
  NAND4_X1 U20333 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17158), .A3(n17140), 
        .A4(n17139), .ZN(n17141) );
  NAND2_X1 U20334 ( .A1(n17142), .A2(n17141), .ZN(P3_U2674) );
  AOI21_X1 U20335 ( .B1(n17144), .B2(n17149), .A(n17143), .ZN(n17460) );
  NAND2_X1 U20336 ( .A1(n17460), .A2(n17432), .ZN(n17145) );
  OAI221_X1 U20337 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17148), .C1(n17147), 
        .C2(n17146), .A(n17145), .ZN(P3_U2676) );
  INV_X1 U20338 ( .A(n17148), .ZN(n17152) );
  AOI21_X1 U20339 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17423), .A(n17158), .ZN(
        n17151) );
  OAI21_X1 U20340 ( .B1(n17154), .B2(n17150), .A(n17149), .ZN(n17467) );
  OAI22_X1 U20341 ( .A1(n17152), .A2(n17151), .B1(n17467), .B2(n17423), .ZN(
        P3_U2677) );
  INV_X1 U20342 ( .A(n17153), .ZN(n17162) );
  AOI21_X1 U20343 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17423), .A(n17162), .ZN(
        n17157) );
  AOI21_X1 U20344 ( .B1(n17155), .B2(n17159), .A(n17154), .ZN(n17468) );
  INV_X1 U20345 ( .A(n17468), .ZN(n17156) );
  OAI22_X1 U20346 ( .A1(n17158), .A2(n17157), .B1(n17156), .B2(n17423), .ZN(
        P3_U2678) );
  AOI21_X1 U20347 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17423), .A(n17169), .ZN(
        n17161) );
  OAI21_X1 U20348 ( .B1(n17164), .B2(n17160), .A(n17159), .ZN(n17478) );
  OAI22_X1 U20349 ( .A1(n17162), .A2(n17161), .B1(n17478), .B2(n17423), .ZN(
        P3_U2679) );
  INV_X1 U20350 ( .A(n17163), .ZN(n17187) );
  AOI21_X1 U20351 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17423), .A(n17187), .ZN(
        n17168) );
  AOI21_X1 U20352 ( .B1(n17166), .B2(n17165), .A(n17164), .ZN(n17482) );
  INV_X1 U20353 ( .A(n17482), .ZN(n17167) );
  OAI22_X1 U20354 ( .A1(n17169), .A2(n17168), .B1(n17167), .B2(n17423), .ZN(
        P3_U2680) );
  AOI21_X1 U20355 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17423), .A(n17170), .ZN(
        n17186) );
  AOI22_X1 U20356 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17183) );
  AOI22_X1 U20357 ( .A1(n12945), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17171) );
  OAI21_X1 U20358 ( .B1(n17355), .B2(n17172), .A(n17171), .ZN(n17181) );
  AOI22_X1 U20359 ( .A1(n13039), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17381), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17178) );
  AOI22_X1 U20360 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17375), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17174) );
  AOI22_X1 U20361 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17173) );
  OAI211_X1 U20362 ( .C1(n17380), .C2(n17175), .A(n17174), .B(n17173), .ZN(
        n17176) );
  AOI21_X1 U20363 ( .B1(n17392), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n17176), .ZN(n17177) );
  OAI211_X1 U20364 ( .C1(n17367), .C2(n17179), .A(n17178), .B(n17177), .ZN(
        n17180) );
  AOI211_X1 U20365 ( .C1(n9665), .C2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n17181), .B(n17180), .ZN(n17182) );
  OAI211_X1 U20366 ( .C1(n17396), .C2(n17184), .A(n17183), .B(n17182), .ZN(
        n17485) );
  INV_X1 U20367 ( .A(n17485), .ZN(n17185) );
  OAI22_X1 U20368 ( .A1(n17187), .A2(n17186), .B1(n17185), .B2(n17423), .ZN(
        P3_U2681) );
  AOI22_X1 U20369 ( .A1(n12945), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17374), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17198) );
  AOI22_X1 U20370 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17381), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17189) );
  AOI22_X1 U20371 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17188) );
  OAI211_X1 U20372 ( .C1(n17358), .C2(n17190), .A(n17189), .B(n17188), .ZN(
        n17196) );
  AOI22_X1 U20373 ( .A1(n17384), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17194) );
  AOI22_X1 U20374 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17193) );
  AOI22_X1 U20375 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17192) );
  NAND2_X1 U20376 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n17191) );
  NAND4_X1 U20377 ( .A1(n17194), .A2(n17193), .A3(n17192), .A4(n17191), .ZN(
        n17195) );
  AOI211_X1 U20378 ( .C1(n17321), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n17196), .B(n17195), .ZN(n17197) );
  OAI211_X1 U20379 ( .C1(n17367), .C2(n17414), .A(n17198), .B(n17197), .ZN(
        n17492) );
  INV_X1 U20380 ( .A(n17492), .ZN(n17200) );
  NAND3_X1 U20381 ( .A1(n17201), .A2(P3_EBX_REG_21__SCAN_IN), .A3(n17423), 
        .ZN(n17199) );
  OAI221_X1 U20382 ( .B1(n17201), .B2(P3_EBX_REG_21__SCAN_IN), .C1(n17423), 
        .C2(n17200), .A(n17199), .ZN(P3_U2682) );
  OAI21_X1 U20383 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17202), .A(n17423), .ZN(
        n17215) );
  AOI22_X1 U20384 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17213) );
  AOI22_X1 U20385 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17204) );
  AOI22_X1 U20386 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17203) );
  OAI211_X1 U20387 ( .C1(n17380), .C2(n17205), .A(n17204), .B(n17203), .ZN(
        n17211) );
  AOI22_X1 U20388 ( .A1(n17384), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17381), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17209) );
  AOI22_X1 U20389 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12945), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17208) );
  AOI22_X1 U20390 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17320), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17207) );
  NAND2_X1 U20391 ( .A1(n17374), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n17206) );
  NAND4_X1 U20392 ( .A1(n17209), .A2(n17208), .A3(n17207), .A4(n17206), .ZN(
        n17210) );
  AOI211_X1 U20393 ( .C1(n17392), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n17211), .B(n17210), .ZN(n17212) );
  OAI211_X1 U20394 ( .C1(n17303), .C2(n17305), .A(n17213), .B(n17212), .ZN(
        n17495) );
  INV_X1 U20395 ( .A(n17495), .ZN(n17214) );
  OAI22_X1 U20396 ( .A1(n17216), .A2(n17215), .B1(n17214), .B2(n17423), .ZN(
        P3_U2683) );
  AOI22_X1 U20397 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17228) );
  AOI22_X1 U20398 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17227) );
  AOI22_X1 U20399 ( .A1(n17321), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17374), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17226) );
  OAI22_X1 U20400 ( .A1(n17367), .A2(n17420), .B1(n17268), .B2(n17218), .ZN(
        n17224) );
  AOI22_X1 U20401 ( .A1(n17384), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12945), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17222) );
  AOI22_X1 U20402 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17381), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17221) );
  AOI22_X1 U20403 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17320), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17220) );
  NAND2_X1 U20404 ( .A1(n17392), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n17219) );
  NAND4_X1 U20405 ( .A1(n17222), .A2(n17221), .A3(n17220), .A4(n17219), .ZN(
        n17223) );
  AOI211_X1 U20406 ( .C1(n17375), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n17224), .B(n17223), .ZN(n17225) );
  NAND4_X1 U20407 ( .A1(n17228), .A2(n17227), .A3(n17226), .A4(n17225), .ZN(
        n17499) );
  INV_X1 U20408 ( .A(n17499), .ZN(n17231) );
  OAI21_X1 U20409 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17246), .A(n17229), .ZN(
        n17230) );
  AOI22_X1 U20410 ( .A1(n17432), .A2(n17231), .B1(n17230), .B2(n17423), .ZN(
        P3_U2684) );
  NAND2_X1 U20411 ( .A1(n17423), .A2(P3_EBX_REG_18__SCAN_IN), .ZN(n17245) );
  AOI22_X1 U20412 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17356), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17242) );
  AOI22_X1 U20413 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17241) );
  AOI22_X1 U20414 ( .A1(n17321), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17392), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17240) );
  OAI22_X1 U20415 ( .A1(n17396), .A2(n17232), .B1(n17367), .B2(n17424), .ZN(
        n17238) );
  AOI22_X1 U20416 ( .A1(n17381), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17236) );
  AOI22_X1 U20417 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17235) );
  AOI22_X1 U20418 ( .A1(n17384), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17320), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17234) );
  NAND2_X1 U20419 ( .A1(n17374), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n17233) );
  NAND4_X1 U20420 ( .A1(n17236), .A2(n17235), .A3(n17234), .A4(n17233), .ZN(
        n17237) );
  AOI211_X1 U20421 ( .C1(n12945), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n17238), .B(n17237), .ZN(n17239) );
  NAND4_X1 U20422 ( .A1(n17242), .A2(n17241), .A3(n17240), .A4(n17239), .ZN(
        n17505) );
  NOR4_X1 U20423 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17260), .A3(n17262), .A4(
        n17429), .ZN(n17243) );
  AOI21_X1 U20424 ( .B1(n17432), .B2(n17505), .A(n17243), .ZN(n17244) );
  OAI21_X1 U20425 ( .B1(n17246), .B2(n17245), .A(n17244), .ZN(P3_U2685) );
  OAI22_X1 U20426 ( .A1(n17248), .A2(n17287), .B1(n17303), .B2(n17247), .ZN(
        n17259) );
  AOI22_X1 U20427 ( .A1(n12945), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n13117), .ZN(n17257) );
  AOI22_X1 U20428 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n17381), .ZN(n17256) );
  OAI22_X1 U20429 ( .A1(n17354), .A2(n17249), .B1(n12918), .B2(n17366), .ZN(
        n17254) );
  AOI22_X1 U20430 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17384), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17252) );
  AOI22_X1 U20431 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17251) );
  AOI22_X1 U20432 ( .A1(n17321), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17392), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17250) );
  NAND3_X1 U20433 ( .A1(n17252), .A2(n17251), .A3(n17250), .ZN(n17253) );
  AOI211_X1 U20434 ( .C1(n9653), .C2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A(
        n17254), .B(n17253), .ZN(n17255) );
  NAND3_X1 U20435 ( .A1(n17257), .A2(n17256), .A3(n17255), .ZN(n17258) );
  AOI211_X1 U20436 ( .C1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .C2(n14415), .A(
        n17259), .B(n17258), .ZN(n17515) );
  NAND3_X1 U20437 ( .A1(n17261), .A2(n17431), .A3(n17260), .ZN(n17266) );
  NAND2_X1 U20438 ( .A1(n17527), .A2(n17262), .ZN(n17282) );
  INV_X1 U20439 ( .A(n17282), .ZN(n17264) );
  OAI21_X1 U20440 ( .B1(n17264), .B2(n17263), .A(P3_EBX_REG_17__SCAN_IN), .ZN(
        n17265) );
  OAI211_X1 U20441 ( .C1(n17515), .C2(n17423), .A(n17266), .B(n17265), .ZN(
        P3_U2686) );
  NAND2_X1 U20442 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17297), .ZN(n17281) );
  OAI22_X1 U20443 ( .A1(n17367), .A2(n17379), .B1(n17268), .B2(n17267), .ZN(
        n17279) );
  AOI22_X1 U20444 ( .A1(n12945), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17382), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17277) );
  AOI22_X1 U20445 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17276) );
  INV_X1 U20446 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17270) );
  AOI22_X1 U20447 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17320), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17269) );
  OAI21_X1 U20448 ( .B1(n17380), .B2(n17270), .A(n17269), .ZN(n17274) );
  AOI22_X1 U20449 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17272) );
  AOI22_X1 U20450 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17381), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17271) );
  OAI211_X1 U20451 ( .C1(n17358), .C2(n17395), .A(n17272), .B(n17271), .ZN(
        n17273) );
  AOI211_X1 U20452 ( .C1(n17374), .C2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n17274), .B(n17273), .ZN(n17275) );
  NAND3_X1 U20453 ( .A1(n17277), .A2(n17276), .A3(n17275), .ZN(n17278) );
  AOI211_X1 U20454 ( .C1(n17384), .C2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A(
        n17279), .B(n17278), .ZN(n17522) );
  INV_X1 U20455 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17280) );
  NAND2_X1 U20456 ( .A1(n17423), .A2(n17281), .ZN(n17298) );
  OAI222_X1 U20457 ( .A1(n17282), .A2(n17281), .B1(n17423), .B2(n17522), .C1(
        n17280), .C2(n17298), .ZN(P3_U2687) );
  AOI22_X1 U20458 ( .A1(n12945), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17283) );
  OAI21_X1 U20459 ( .B1(n12928), .B2(n17284), .A(n17283), .ZN(n17296) );
  INV_X1 U20460 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17294) );
  AOI22_X1 U20461 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17293) );
  INV_X1 U20462 ( .A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17286) );
  AOI22_X1 U20463 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17374), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17285) );
  OAI21_X1 U20464 ( .B1(n17287), .B2(n17286), .A(n17285), .ZN(n17291) );
  AOI22_X1 U20465 ( .A1(n17384), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17289) );
  AOI22_X1 U20466 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17288) );
  OAI211_X1 U20467 ( .C1(n17380), .C2(n17406), .A(n17289), .B(n17288), .ZN(
        n17290) );
  AOI211_X1 U20468 ( .C1(n17392), .C2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n17291), .B(n17290), .ZN(n17292) );
  OAI211_X1 U20469 ( .C1(n17367), .C2(n17294), .A(n17293), .B(n17292), .ZN(
        n17295) );
  AOI211_X1 U20470 ( .C1(n12938), .C2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n17296), .B(n17295), .ZN(n17525) );
  NOR2_X1 U20471 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17297), .ZN(n17299) );
  OAI22_X1 U20472 ( .A1(n17525), .A2(n17423), .B1(n17299), .B2(n17298), .ZN(
        P3_U2688) );
  NOR2_X1 U20473 ( .A1(n18449), .A2(n17333), .ZN(n17300) );
  AOI21_X1 U20474 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17423), .A(n17300), .ZN(
        n17316) );
  AOI22_X1 U20475 ( .A1(n17381), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17301) );
  OAI21_X1 U20476 ( .B1(n17303), .B2(n17302), .A(n17301), .ZN(n17315) );
  AOI22_X1 U20477 ( .A1(n17384), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17320), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17312) );
  AOI22_X1 U20478 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17392), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17304) );
  OAI21_X1 U20479 ( .B1(n12918), .B2(n17305), .A(n17304), .ZN(n17310) );
  AOI22_X1 U20480 ( .A1(n17306), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17308) );
  AOI22_X1 U20481 ( .A1(n9662), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17307) );
  OAI211_X1 U20482 ( .C1(n17380), .C2(n17418), .A(n17308), .B(n17307), .ZN(
        n17309) );
  AOI211_X1 U20483 ( .C1(n17374), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n17310), .B(n17309), .ZN(n17311) );
  OAI211_X1 U20484 ( .C1(n14414), .C2(n17313), .A(n17312), .B(n17311), .ZN(
        n17314) );
  AOI211_X1 U20485 ( .C1(n12945), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n17315), .B(n17314), .ZN(n17539) );
  OAI22_X1 U20486 ( .A1(n17317), .A2(n17316), .B1(n17539), .B2(n17423), .ZN(
        P3_U2691) );
  AOI22_X1 U20487 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17318) );
  OAI21_X1 U20488 ( .B1(n12918), .B2(n17319), .A(n17318), .ZN(n17332) );
  AOI22_X1 U20489 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17329) );
  AOI22_X1 U20490 ( .A1(n17321), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17320), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17322) );
  INV_X1 U20491 ( .A(n17322), .ZN(n17327) );
  AOI22_X1 U20492 ( .A1(n17384), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12945), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17325) );
  AOI22_X1 U20493 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17324) );
  AOI22_X1 U20494 ( .A1(n13039), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17392), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17323) );
  NAND3_X1 U20495 ( .A1(n17325), .A2(n17324), .A3(n17323), .ZN(n17326) );
  AOI211_X1 U20496 ( .C1(n17375), .C2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n17327), .B(n17326), .ZN(n17328) );
  OAI211_X1 U20497 ( .C1(n12928), .C2(n17330), .A(n17329), .B(n17328), .ZN(
        n17331) );
  AOI211_X1 U20498 ( .C1(n17217), .C2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n17332), .B(n17331), .ZN(n17543) );
  OAI21_X1 U20499 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17351), .A(n17333), .ZN(
        n17334) );
  AOI22_X1 U20500 ( .A1(n17432), .A2(n17543), .B1(n17334), .B2(n17423), .ZN(
        P3_U2692) );
  INV_X1 U20501 ( .A(n17370), .ZN(n17335) );
  AOI22_X1 U20502 ( .A1(n17527), .A2(n17335), .B1(P3_EBX_REG_10__SCAN_IN), 
        .B2(n17423), .ZN(n17350) );
  AOI22_X1 U20503 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17347) );
  AOI22_X1 U20504 ( .A1(n17217), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12945), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17338) );
  AOI22_X1 U20505 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17337) );
  OAI211_X1 U20506 ( .C1(n17380), .C2(n17424), .A(n17338), .B(n17337), .ZN(
        n17345) );
  AOI22_X1 U20507 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17385), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17343) );
  AOI22_X1 U20508 ( .A1(n17384), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17342) );
  AOI22_X1 U20509 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17341) );
  NAND2_X1 U20510 ( .A1(n17374), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n17340) );
  NAND4_X1 U20511 ( .A1(n17343), .A2(n17342), .A3(n17341), .A4(n17340), .ZN(
        n17344) );
  AOI211_X1 U20512 ( .C1(n17392), .C2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n17345), .B(n17344), .ZN(n17346) );
  OAI211_X1 U20513 ( .C1(n12928), .C2(n17348), .A(n17347), .B(n17346), .ZN(
        n17546) );
  INV_X1 U20514 ( .A(n17546), .ZN(n17349) );
  OAI22_X1 U20515 ( .A1(n17351), .A2(n17350), .B1(n17349), .B2(n17423), .ZN(
        P3_U2693) );
  AOI22_X1 U20516 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17336), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17352), .ZN(n17353) );
  OAI21_X1 U20517 ( .B1(n17355), .B2(n17354), .A(n17353), .ZN(n17369) );
  AOI22_X1 U20518 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17356), .B1(
        n12945), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17365) );
  AOI22_X1 U20519 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n13117), .ZN(n17357) );
  OAI21_X1 U20520 ( .B1(n17359), .B2(n17358), .A(n17357), .ZN(n17363) );
  AOI22_X1 U20521 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n17382), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n14415), .ZN(n17361) );
  AOI22_X1 U20522 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n9665), .B1(
        n17375), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17360) );
  OAI211_X1 U20523 ( .C1(n17427), .C2(n17380), .A(n17361), .B(n17360), .ZN(
        n17362) );
  AOI211_X1 U20524 ( .C1(n17374), .C2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n17363), .B(n17362), .ZN(n17364) );
  OAI211_X1 U20525 ( .C1(n17367), .C2(n17366), .A(n17365), .B(n17364), .ZN(
        n17368) );
  AOI211_X1 U20526 ( .C1(n17217), .C2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n17369), .B(n17368), .ZN(n17551) );
  OAI21_X1 U20527 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17371), .A(n17370), .ZN(
        n17372) );
  AOI22_X1 U20528 ( .A1(n17432), .A2(n17551), .B1(n17372), .B2(n17423), .ZN(
        P3_U2694) );
  NAND2_X1 U20529 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17373), .ZN(n17401) );
  AOI22_X1 U20530 ( .A1(n17320), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17374), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17394) );
  AOI22_X1 U20531 ( .A1(n17375), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13117), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17378) );
  AOI22_X1 U20532 ( .A1(n17336), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17376), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17377) );
  OAI211_X1 U20533 ( .C1(n17380), .C2(n17379), .A(n17378), .B(n17377), .ZN(
        n17391) );
  AOI22_X1 U20534 ( .A1(n17382), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17381), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17389) );
  AOI22_X1 U20535 ( .A1(n17384), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12945), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17388) );
  AOI22_X1 U20536 ( .A1(n17385), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14415), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17387) );
  NAND2_X1 U20537 ( .A1(n9653), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n17386) );
  NAND4_X1 U20538 ( .A1(n17389), .A2(n17388), .A3(n17387), .A4(n17386), .ZN(
        n17390) );
  AOI211_X1 U20539 ( .C1(n17392), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n17391), .B(n17390), .ZN(n17393) );
  OAI211_X1 U20540 ( .C1(n17396), .C2(n17395), .A(n17394), .B(n17393), .ZN(
        n17554) );
  INV_X1 U20541 ( .A(n17554), .ZN(n17400) );
  NAND4_X1 U20542 ( .A1(n17527), .A2(n17408), .A3(n17398), .A4(n17397), .ZN(
        n17399) );
  OAI221_X1 U20543 ( .B1(n17432), .B2(n17401), .C1(n17423), .C2(n17400), .A(
        n17399), .ZN(P3_U2695) );
  INV_X1 U20544 ( .A(n17408), .ZN(n17402) );
  OAI21_X1 U20545 ( .B1(n17403), .B2(n17402), .A(P3_EBX_REG_7__SCAN_IN), .ZN(
        n17407) );
  NAND4_X1 U20546 ( .A1(n17527), .A2(P3_EBX_REG_6__SCAN_IN), .A3(n17408), .A4(
        n17404), .ZN(n17405) );
  OAI221_X1 U20547 ( .B1(n17432), .B2(n17407), .C1(n17423), .C2(n17406), .A(
        n17405), .ZN(P3_U2696) );
  NAND2_X1 U20548 ( .A1(n17527), .A2(n17408), .ZN(n17410) );
  NOR2_X1 U20549 ( .A1(n17432), .A2(n17408), .ZN(n17411) );
  AOI22_X1 U20550 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n17432), .B1(
        P3_EBX_REG_6__SCAN_IN), .B2(n17411), .ZN(n17409) );
  OAI21_X1 U20551 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17410), .A(n17409), .ZN(
        P3_U2697) );
  INV_X1 U20552 ( .A(n17415), .ZN(n17412) );
  OAI21_X1 U20553 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17412), .A(n17411), .ZN(
        n17413) );
  OAI21_X1 U20554 ( .B1(n17423), .B2(n17414), .A(n17413), .ZN(P3_U2698) );
  OAI21_X1 U20555 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17416), .A(n17415), .ZN(
        n17417) );
  AOI22_X1 U20556 ( .A1(n17432), .A2(n17418), .B1(n17417), .B2(n17423), .ZN(
        P3_U2699) );
  NAND3_X1 U20557 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17421), .A3(n17431), .ZN(
        n17422) );
  NAND3_X1 U20558 ( .A1(n17422), .A2(P3_EBX_REG_3__SCAN_IN), .A3(n17423), .ZN(
        n17419) );
  OAI221_X1 U20559 ( .B1(n17422), .B2(P3_EBX_REG_3__SCAN_IN), .C1(n17423), 
        .C2(n17420), .A(n17419), .ZN(P3_U2700) );
  AOI21_X1 U20560 ( .B1(n17435), .B2(n17421), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n17426) );
  NAND2_X1 U20561 ( .A1(n17423), .A2(n17422), .ZN(n17425) );
  OAI22_X1 U20562 ( .A1(n17426), .A2(n17425), .B1(n17424), .B2(n17423), .ZN(
        P3_U2701) );
  OAI222_X1 U20563 ( .A1(n17430), .A2(n17429), .B1(n17428), .B2(n17435), .C1(
        n17427), .C2(n17423), .ZN(P3_U2702) );
  AOI22_X1 U20564 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17432), .B1(
        n17431), .B2(n17434), .ZN(n17433) );
  OAI21_X1 U20565 ( .B1(n17435), .B2(n17434), .A(n17433), .ZN(P3_U2703) );
  NOR2_X1 U20566 ( .A1(n17577), .A2(n17436), .ZN(n17516) );
  INV_X1 U20567 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17604) );
  INV_X1 U20568 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17608) );
  NAND4_X1 U20569 ( .A1(n17593), .A2(P3_EAX_REG_7__SCAN_IN), .A3(
        P3_EAX_REG_6__SCAN_IN), .A4(P3_EAX_REG_3__SCAN_IN), .ZN(n17439) );
  NAND3_X1 U20570 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .A3(P3_EAX_REG_0__SCAN_IN), .ZN(n17558) );
  INV_X1 U20571 ( .A(n17558), .ZN(n17437) );
  NAND3_X1 U20572 ( .A1(n17437), .A2(P3_EAX_REG_4__SCAN_IN), .A3(
        P3_EAX_REG_5__SCAN_IN), .ZN(n17438) );
  NAND2_X1 U20573 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .ZN(n17528) );
  NAND3_X1 U20574 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .ZN(n17530) );
  NOR2_X1 U20575 ( .A1(n17528), .A2(n17530), .ZN(n17440) );
  AND2_X1 U20576 ( .A1(n17440), .A2(n10226), .ZN(n17441) );
  NAND2_X1 U20577 ( .A1(n17526), .A2(n17441), .ZN(n17532) );
  INV_X1 U20578 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17707) );
  NAND3_X1 U20579 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .ZN(n17489) );
  INV_X1 U20580 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17612) );
  INV_X1 U20581 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17662) );
  INV_X1 U20582 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17606) );
  INV_X1 U20583 ( .A(n17442), .ZN(n17474) );
  INV_X1 U20584 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17601) );
  NOR2_X1 U20585 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n17452), .ZN(n17444) );
  OAI21_X1 U20586 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17589), .A(n17450), .ZN(
        n17443) );
  AOI22_X1 U20587 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17444), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17443), .ZN(n17445) );
  OAI21_X1 U20588 ( .B1(n18452), .B2(n17504), .A(n17445), .ZN(P3_U2704) );
  INV_X1 U20589 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17676) );
  NAND2_X1 U20590 ( .A1(n17446), .A2(n17555), .ZN(n17510) );
  INV_X1 U20591 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n19429) );
  OAI22_X1 U20592 ( .A1(n17447), .A2(n17579), .B1(n19429), .B2(n17504), .ZN(
        n17448) );
  AOI21_X1 U20593 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17517), .A(n17448), .ZN(
        n17449) );
  OAI221_X1 U20594 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17452), .C1(n17676), 
        .C2(n17450), .A(n17449), .ZN(P3_U2705) );
  INV_X1 U20595 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18440) );
  AOI22_X1 U20596 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17517), .B1(n17586), .B2(
        n17451), .ZN(n17455) );
  OAI211_X1 U20597 ( .C1(n17453), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17577), .B(
        n17452), .ZN(n17454) );
  OAI211_X1 U20598 ( .C1(n17504), .C2(n18440), .A(n17455), .B(n17454), .ZN(
        P3_U2706) );
  AOI22_X1 U20599 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17517), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17516), .ZN(n17458) );
  OAI211_X1 U20600 ( .C1(n9709), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17577), .B(
        n17456), .ZN(n17457) );
  OAI211_X1 U20601 ( .C1(n17459), .C2(n17579), .A(n17458), .B(n17457), .ZN(
        P3_U2707) );
  AOI22_X1 U20602 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17517), .B1(n17586), .B2(
        n17460), .ZN(n17463) );
  AOI211_X1 U20603 ( .C1(n17601), .C2(n17464), .A(n9709), .B(n17555), .ZN(
        n17461) );
  INV_X1 U20604 ( .A(n17461), .ZN(n17462) );
  OAI211_X1 U20605 ( .C1(n17504), .C2(n18430), .A(n17463), .B(n17462), .ZN(
        P3_U2708) );
  AOI22_X1 U20606 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17517), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17516), .ZN(n17466) );
  OAI211_X1 U20607 ( .C1(n17469), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17577), .B(
        n17464), .ZN(n17465) );
  OAI211_X1 U20608 ( .C1(n17467), .C2(n17579), .A(n17466), .B(n17465), .ZN(
        P3_U2709) );
  AOI22_X1 U20609 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17517), .B1(n17586), .B2(
        n17468), .ZN(n17472) );
  AOI211_X1 U20610 ( .C1(n17604), .C2(n17474), .A(n17469), .B(n17555), .ZN(
        n17470) );
  INV_X1 U20611 ( .A(n17470), .ZN(n17471) );
  OAI211_X1 U20612 ( .C1(n17504), .C2(n18421), .A(n17472), .B(n17471), .ZN(
        P3_U2710) );
  AOI22_X1 U20613 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17517), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17516), .ZN(n17477) );
  OAI21_X1 U20614 ( .B1(n17606), .B2(n17555), .A(n17473), .ZN(n17475) );
  NAND2_X1 U20615 ( .A1(n17475), .A2(n17474), .ZN(n17476) );
  OAI211_X1 U20616 ( .C1(n17478), .C2(n17579), .A(n17477), .B(n17476), .ZN(
        P3_U2711) );
  AOI22_X1 U20617 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17517), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17516), .ZN(n17484) );
  AOI211_X1 U20618 ( .C1(n17608), .C2(n17480), .A(n17555), .B(n17479), .ZN(
        n17481) );
  AOI21_X1 U20619 ( .B1(n17482), .B2(n17586), .A(n17481), .ZN(n17483) );
  NAND2_X1 U20620 ( .A1(n17484), .A2(n17483), .ZN(P3_U2712) );
  NAND2_X1 U20621 ( .A1(n17527), .A2(n10240), .ZN(n17491) );
  AOI22_X1 U20622 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17516), .B1(n17586), .B2(
        n17485), .ZN(n17488) );
  NOR2_X1 U20623 ( .A1(n17555), .A2(n10240), .ZN(n17486) );
  AOI22_X1 U20624 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17517), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17486), .ZN(n17487) );
  OAI211_X1 U20625 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n17491), .A(n17488), .B(
        n17487), .ZN(P3_U2713) );
  INV_X1 U20626 ( .A(n17507), .ZN(n17511) );
  OR2_X1 U20627 ( .A1(n17489), .A2(n17511), .ZN(n17496) );
  OAI21_X1 U20628 ( .B1(n17555), .B2(n17612), .A(n17496), .ZN(n17490) );
  AOI22_X1 U20629 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n17516), .B1(n17491), .B2(
        n17490), .ZN(n17494) );
  AOI22_X1 U20630 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17517), .B1(n17586), .B2(
        n17492), .ZN(n17493) );
  NAND2_X1 U20631 ( .A1(n17494), .A2(n17493), .ZN(P3_U2714) );
  INV_X1 U20632 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n18435) );
  AOI22_X1 U20633 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17517), .B1(n17586), .B2(
        n17495), .ZN(n17498) );
  INV_X1 U20634 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17616) );
  NAND2_X1 U20635 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17507), .ZN(n17506) );
  NOR2_X1 U20636 ( .A1(n17616), .A2(n17506), .ZN(n17500) );
  OAI211_X1 U20637 ( .C1(n17500), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17577), .B(
        n17496), .ZN(n17497) );
  OAI211_X1 U20638 ( .C1(n17504), .C2(n18435), .A(n17498), .B(n17497), .ZN(
        P3_U2715) );
  AOI22_X1 U20639 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17517), .B1(n17586), .B2(
        n17499), .ZN(n17503) );
  AOI211_X1 U20640 ( .C1(n17616), .C2(n17506), .A(n17500), .B(n17555), .ZN(
        n17501) );
  INV_X1 U20641 ( .A(n17501), .ZN(n17502) );
  OAI211_X1 U20642 ( .C1(n17504), .C2(n15249), .A(n17503), .B(n17502), .ZN(
        P3_U2716) );
  INV_X1 U20643 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18426) );
  AOI22_X1 U20644 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n17516), .B1(n17586), .B2(
        n17505), .ZN(n17509) );
  OAI211_X1 U20645 ( .C1(n17507), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17577), .B(
        n17506), .ZN(n17508) );
  OAI211_X1 U20646 ( .C1(n17510), .C2(n18426), .A(n17509), .B(n17508), .ZN(
        P3_U2717) );
  AOI22_X1 U20647 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17517), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17516), .ZN(n17514) );
  INV_X1 U20648 ( .A(n17519), .ZN(n17512) );
  OAI211_X1 U20649 ( .C1(n17512), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17577), .B(
        n17511), .ZN(n17513) );
  OAI211_X1 U20650 ( .C1(n17515), .C2(n17579), .A(n17514), .B(n17513), .ZN(
        P3_U2718) );
  AOI22_X1 U20651 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17517), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17516), .ZN(n17521) );
  OAI211_X1 U20652 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17518), .A(n17577), .B(
        n17519), .ZN(n17520) );
  OAI211_X1 U20653 ( .C1(n17522), .C2(n17579), .A(n17521), .B(n17520), .ZN(
        P3_U2719) );
  AOI211_X1 U20654 ( .C1(n17707), .C2(n17532), .A(n17555), .B(n17518), .ZN(
        n17523) );
  AOI21_X1 U20655 ( .B1(n17587), .B2(BUF2_REG_15__SCAN_IN), .A(n17523), .ZN(
        n17524) );
  OAI21_X1 U20656 ( .B1(n17525), .B2(n17579), .A(n17524), .ZN(P3_U2720) );
  NAND2_X1 U20657 ( .A1(n17527), .A2(n17526), .ZN(n17550) );
  INV_X1 U20658 ( .A(n17553), .ZN(n17529) );
  NOR2_X1 U20659 ( .A1(n17530), .A2(n17529), .ZN(n17541) );
  NAND2_X1 U20660 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17541), .ZN(n17535) );
  AOI22_X1 U20661 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17587), .B1(n17586), .B2(
        n17531), .ZN(n17534) );
  NAND3_X1 U20662 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17577), .A3(n17532), 
        .ZN(n17533) );
  OAI211_X1 U20663 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n17535), .A(n17534), .B(
        n17533), .ZN(P3_U2721) );
  INV_X1 U20664 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17700) );
  INV_X1 U20665 ( .A(n17535), .ZN(n17538) );
  AOI21_X1 U20666 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17577), .A(n17541), .ZN(
        n17537) );
  OAI222_X1 U20667 ( .A1(n17580), .A2(n17700), .B1(n17538), .B2(n17537), .C1(
        n17579), .C2(n17536), .ZN(P3_U2722) );
  INV_X1 U20668 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17697) );
  INV_X1 U20669 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17632) );
  NAND2_X1 U20670 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17553), .ZN(n17547) );
  NOR2_X1 U20671 ( .A1(n17632), .A2(n17547), .ZN(n17545) );
  AOI21_X1 U20672 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17577), .A(n17545), .ZN(
        n17540) );
  OAI222_X1 U20673 ( .A1(n17580), .A2(n17697), .B1(n17541), .B2(n17540), .C1(
        n17579), .C2(n17539), .ZN(P3_U2723) );
  INV_X1 U20674 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17694) );
  INV_X1 U20675 ( .A(n17547), .ZN(n17542) );
  AOI21_X1 U20676 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17577), .A(n17542), .ZN(
        n17544) );
  OAI222_X1 U20677 ( .A1(n17580), .A2(n17694), .B1(n17545), .B2(n17544), .C1(
        n17579), .C2(n17543), .ZN(P3_U2724) );
  AOI22_X1 U20678 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17587), .B1(n17586), .B2(
        n17546), .ZN(n17549) );
  OAI211_X1 U20679 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n17553), .A(n17577), .B(
        n17547), .ZN(n17548) );
  NAND2_X1 U20680 ( .A1(n17549), .A2(n17548), .ZN(P3_U2725) );
  INV_X1 U20681 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17689) );
  INV_X1 U20682 ( .A(n17550), .ZN(n17561) );
  AOI22_X1 U20683 ( .A1(n17561), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n17577), .ZN(n17552) );
  OAI222_X1 U20684 ( .A1(n17580), .A2(n17689), .B1(n17553), .B2(n17552), .C1(
        n17579), .C2(n17551), .ZN(P3_U2726) );
  INV_X1 U20685 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17687) );
  INV_X1 U20686 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17638) );
  AOI22_X1 U20687 ( .A1(n17586), .A2(n17554), .B1(n17561), .B2(n17638), .ZN(
        n17557) );
  OR3_X1 U20688 ( .A1(n17638), .A2(n17555), .A3(n17526), .ZN(n17556) );
  OAI211_X1 U20689 ( .C1(n17580), .C2(n17687), .A(n17557), .B(n17556), .ZN(
        P3_U2727) );
  INV_X1 U20690 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18451) );
  INV_X1 U20691 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17642) );
  INV_X1 U20692 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17646) );
  NAND2_X1 U20693 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17584), .ZN(n17570) );
  NOR2_X1 U20694 ( .A1(n17646), .A2(n17570), .ZN(n17573) );
  NAND2_X1 U20695 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17573), .ZN(n17562) );
  NOR2_X1 U20696 ( .A1(n17642), .A2(n17562), .ZN(n17565) );
  AOI21_X1 U20697 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17577), .A(n17565), .ZN(
        n17560) );
  OAI222_X1 U20698 ( .A1(n17580), .A2(n18451), .B1(n17561), .B2(n17560), .C1(
        n17579), .C2(n17559), .ZN(P3_U2728) );
  INV_X1 U20699 ( .A(n17562), .ZN(n17569) );
  AOI21_X1 U20700 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17577), .A(n17569), .ZN(
        n17564) );
  OAI222_X1 U20701 ( .A1(n18446), .A2(n17580), .B1(n17565), .B2(n17564), .C1(
        n17579), .C2(n17563), .ZN(P3_U2729) );
  INV_X1 U20702 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18441) );
  AOI21_X1 U20703 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17577), .A(n17573), .ZN(
        n17568) );
  INV_X1 U20704 ( .A(n17566), .ZN(n17567) );
  OAI222_X1 U20705 ( .A1(n18441), .A2(n17580), .B1(n17569), .B2(n17568), .C1(
        n17579), .C2(n17567), .ZN(P3_U2730) );
  INV_X1 U20706 ( .A(n17570), .ZN(n17576) );
  AOI21_X1 U20707 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17577), .A(n17576), .ZN(
        n17572) );
  OAI222_X1 U20708 ( .A1(n18436), .A2(n17580), .B1(n17573), .B2(n17572), .C1(
        n17579), .C2(n17571), .ZN(P3_U2731) );
  INV_X1 U20709 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18431) );
  AOI21_X1 U20710 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17577), .A(n17584), .ZN(
        n17575) );
  OAI222_X1 U20711 ( .A1(n18431), .A2(n17580), .B1(n17576), .B2(n17575), .C1(
        n17579), .C2(n17574), .ZN(P3_U2732) );
  INV_X1 U20712 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17679) );
  NOR2_X1 U20713 ( .A1(n17679), .A2(n17655), .ZN(n17588) );
  OAI221_X1 U20714 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17593), .C1(
        P3_EAX_REG_2__SCAN_IN), .C2(n17588), .A(n17577), .ZN(n17583) );
  OAI22_X1 U20715 ( .A1(n17580), .A2(n18426), .B1(n17579), .B2(n17578), .ZN(
        n17581) );
  INV_X1 U20716 ( .A(n17581), .ZN(n17582) );
  OAI21_X1 U20717 ( .B1(n17584), .B2(n17583), .A(n17582), .ZN(P3_U2733) );
  AOI22_X1 U20718 ( .A1(n17587), .A2(BUF2_REG_1__SCAN_IN), .B1(n17586), .B2(
        n17585), .ZN(n17592) );
  AOI211_X1 U20719 ( .C1(n17679), .C2(n17655), .A(n17589), .B(n17588), .ZN(
        n17590) );
  INV_X1 U20720 ( .A(n17590), .ZN(n17591) );
  OAI211_X1 U20721 ( .C1(n17593), .C2(n17679), .A(n17592), .B(n17591), .ZN(
        P3_U2734) );
  NOR2_X2 U20722 ( .A1(n19018), .A2(n18917), .ZN(n19051) );
  NOR2_X4 U20723 ( .A1(n19051), .A2(n17624), .ZN(n17620) );
  AND2_X1 U20724 ( .A1(n17620), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  AOI22_X1 U20725 ( .A1(n19051), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17620), .ZN(n17595) );
  OAI21_X1 U20726 ( .B1(n17676), .B2(n17622), .A(n17595), .ZN(P3_U2737) );
  INV_X1 U20727 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17597) );
  AOI22_X1 U20728 ( .A1(n19051), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17596) );
  OAI21_X1 U20729 ( .B1(n17597), .B2(n17622), .A(n17596), .ZN(P3_U2738) );
  INV_X1 U20730 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17599) );
  AOI22_X1 U20731 ( .A1(n19051), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17598) );
  OAI21_X1 U20732 ( .B1(n17599), .B2(n17622), .A(n17598), .ZN(P3_U2739) );
  AOI22_X1 U20733 ( .A1(n19051), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17600) );
  OAI21_X1 U20734 ( .B1(n17601), .B2(n17622), .A(n17600), .ZN(P3_U2740) );
  AOI22_X1 U20735 ( .A1(n19051), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17602) );
  OAI21_X1 U20736 ( .B1(n9972), .B2(n17622), .A(n17602), .ZN(P3_U2741) );
  AOI22_X1 U20737 ( .A1(n19051), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17603) );
  OAI21_X1 U20738 ( .B1(n17604), .B2(n17622), .A(n17603), .ZN(P3_U2742) );
  AOI22_X1 U20739 ( .A1(n19051), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17605) );
  OAI21_X1 U20740 ( .B1(n17606), .B2(n17622), .A(n17605), .ZN(P3_U2743) );
  CLKBUF_X1 U20741 ( .A(n19051), .Z(n17652) );
  AOI22_X1 U20742 ( .A1(n17652), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17607) );
  OAI21_X1 U20743 ( .B1(n17608), .B2(n17622), .A(n17607), .ZN(P3_U2744) );
  INV_X1 U20744 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17610) );
  AOI22_X1 U20745 ( .A1(n17652), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17609) );
  OAI21_X1 U20746 ( .B1(n17610), .B2(n17622), .A(n17609), .ZN(P3_U2745) );
  AOI22_X1 U20747 ( .A1(n17652), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17611) );
  OAI21_X1 U20748 ( .B1(n17612), .B2(n17622), .A(n17611), .ZN(P3_U2746) );
  INV_X1 U20749 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17614) );
  AOI22_X1 U20750 ( .A1(n17652), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17613) );
  OAI21_X1 U20751 ( .B1(n17614), .B2(n17622), .A(n17613), .ZN(P3_U2747) );
  AOI22_X1 U20752 ( .A1(n17652), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17615) );
  OAI21_X1 U20753 ( .B1(n17616), .B2(n17622), .A(n17615), .ZN(P3_U2748) );
  INV_X1 U20754 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17618) );
  AOI22_X1 U20755 ( .A1(n17652), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17617) );
  OAI21_X1 U20756 ( .B1(n17618), .B2(n17622), .A(n17617), .ZN(P3_U2749) );
  AOI22_X1 U20757 ( .A1(n17652), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17619) );
  OAI21_X1 U20758 ( .B1(n17662), .B2(n17622), .A(n17619), .ZN(P3_U2750) );
  INV_X1 U20759 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17623) );
  AOI22_X1 U20760 ( .A1(n17652), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17621) );
  OAI21_X1 U20761 ( .B1(n17623), .B2(n17622), .A(n17621), .ZN(P3_U2751) );
  AOI22_X1 U20762 ( .A1(n17652), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17625) );
  OAI21_X1 U20763 ( .B1(n17707), .B2(n17654), .A(n17625), .ZN(P3_U2752) );
  INV_X1 U20764 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17702) );
  AOI22_X1 U20765 ( .A1(n17652), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17626) );
  OAI21_X1 U20766 ( .B1(n17702), .B2(n17654), .A(n17626), .ZN(P3_U2753) );
  INV_X1 U20767 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17628) );
  AOI22_X1 U20768 ( .A1(n17652), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17627) );
  OAI21_X1 U20769 ( .B1(n17628), .B2(n17654), .A(n17627), .ZN(P3_U2754) );
  INV_X1 U20770 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17630) );
  AOI22_X1 U20771 ( .A1(n17652), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17629) );
  OAI21_X1 U20772 ( .B1(n17630), .B2(n17654), .A(n17629), .ZN(P3_U2755) );
  AOI22_X1 U20773 ( .A1(n17652), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17631) );
  OAI21_X1 U20774 ( .B1(n17632), .B2(n17654), .A(n17631), .ZN(P3_U2756) );
  INV_X1 U20775 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17634) );
  AOI22_X1 U20776 ( .A1(n17652), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17633) );
  OAI21_X1 U20777 ( .B1(n17634), .B2(n17654), .A(n17633), .ZN(P3_U2757) );
  INV_X1 U20778 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17636) );
  AOI22_X1 U20779 ( .A1(n17652), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17635) );
  OAI21_X1 U20780 ( .B1(n17636), .B2(n17654), .A(n17635), .ZN(P3_U2758) );
  AOI22_X1 U20781 ( .A1(n17652), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17637) );
  OAI21_X1 U20782 ( .B1(n17638), .B2(n17654), .A(n17637), .ZN(P3_U2759) );
  INV_X1 U20783 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17640) );
  AOI22_X1 U20784 ( .A1(n17652), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17639) );
  OAI21_X1 U20785 ( .B1(n17640), .B2(n17654), .A(n17639), .ZN(P3_U2760) );
  AOI22_X1 U20786 ( .A1(n17652), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17641) );
  OAI21_X1 U20787 ( .B1(n17642), .B2(n17654), .A(n17641), .ZN(P3_U2761) );
  INV_X1 U20788 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17644) );
  AOI22_X1 U20789 ( .A1(n17652), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17643) );
  OAI21_X1 U20790 ( .B1(n17644), .B2(n17654), .A(n17643), .ZN(P3_U2762) );
  AOI22_X1 U20791 ( .A1(n17652), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17645) );
  OAI21_X1 U20792 ( .B1(n17646), .B2(n17654), .A(n17645), .ZN(P3_U2763) );
  INV_X1 U20793 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17648) );
  AOI22_X1 U20794 ( .A1(n17652), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17647) );
  OAI21_X1 U20795 ( .B1(n17648), .B2(n17654), .A(n17647), .ZN(P3_U2764) );
  INV_X1 U20796 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17650) );
  AOI22_X1 U20797 ( .A1(n17652), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17649) );
  OAI21_X1 U20798 ( .B1(n17650), .B2(n17654), .A(n17649), .ZN(P3_U2765) );
  AOI22_X1 U20799 ( .A1(n17652), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17651) );
  OAI21_X1 U20800 ( .B1(n17679), .B2(n17654), .A(n17651), .ZN(P3_U2766) );
  AOI22_X1 U20801 ( .A1(n17652), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17620), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17653) );
  OAI21_X1 U20802 ( .B1(n17655), .B2(n17654), .A(n17653), .ZN(P3_U2767) );
  INV_X1 U20803 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18413) );
  INV_X2 U20804 ( .A(n17704), .ZN(n17699) );
  OR2_X1 U20805 ( .A1(n18896), .A2(n17659), .ZN(n17706) );
  AOI22_X1 U20806 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17695), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17703), .ZN(n17660) );
  OAI21_X1 U20807 ( .B1(n18413), .B2(n17699), .A(n17660), .ZN(P3_U2768) );
  AOI22_X1 U20808 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17704), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17703), .ZN(n17661) );
  OAI21_X1 U20809 ( .B1(n17662), .B2(n17706), .A(n17661), .ZN(P3_U2769) );
  AOI22_X1 U20810 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17695), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17703), .ZN(n17663) );
  OAI21_X1 U20811 ( .B1(n18426), .B2(n17699), .A(n17663), .ZN(P3_U2770) );
  AOI22_X1 U20812 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17695), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17703), .ZN(n17664) );
  OAI21_X1 U20813 ( .B1(n18431), .B2(n17699), .A(n17664), .ZN(P3_U2771) );
  AOI22_X1 U20814 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17695), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17703), .ZN(n17665) );
  OAI21_X1 U20815 ( .B1(n18436), .B2(n17699), .A(n17665), .ZN(P3_U2772) );
  AOI22_X1 U20816 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17695), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17703), .ZN(n17666) );
  OAI21_X1 U20817 ( .B1(n18441), .B2(n17699), .A(n17666), .ZN(P3_U2773) );
  AOI22_X1 U20818 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17695), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17703), .ZN(n17667) );
  OAI21_X1 U20819 ( .B1(n18446), .B2(n17699), .A(n17667), .ZN(P3_U2774) );
  AOI22_X1 U20820 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17695), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17703), .ZN(n17668) );
  OAI21_X1 U20821 ( .B1(n18451), .B2(n17699), .A(n17668), .ZN(P3_U2775) );
  AOI22_X1 U20822 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17695), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17703), .ZN(n17669) );
  OAI21_X1 U20823 ( .B1(n17687), .B2(n17699), .A(n17669), .ZN(P3_U2776) );
  AOI22_X1 U20824 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17695), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17703), .ZN(n17670) );
  OAI21_X1 U20825 ( .B1(n17689), .B2(n17699), .A(n17670), .ZN(P3_U2777) );
  INV_X1 U20826 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17691) );
  AOI22_X1 U20827 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17695), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17703), .ZN(n17671) );
  OAI21_X1 U20828 ( .B1(n17691), .B2(n17699), .A(n17671), .ZN(P3_U2778) );
  AOI22_X1 U20829 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17695), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17703), .ZN(n17672) );
  OAI21_X1 U20830 ( .B1(n17694), .B2(n17699), .A(n17672), .ZN(P3_U2779) );
  AOI22_X1 U20831 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17695), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17703), .ZN(n17673) );
  OAI21_X1 U20832 ( .B1(n17697), .B2(n17699), .A(n17673), .ZN(P3_U2780) );
  INV_X2 U20833 ( .A(n17706), .ZN(n17695) );
  AOI22_X1 U20834 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17695), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17703), .ZN(n17674) );
  OAI21_X1 U20835 ( .B1(n17700), .B2(n17699), .A(n17674), .ZN(P3_U2781) );
  AOI22_X1 U20836 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17704), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17703), .ZN(n17675) );
  OAI21_X1 U20837 ( .B1(n17676), .B2(n17706), .A(n17675), .ZN(P3_U2782) );
  AOI22_X1 U20838 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17695), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17703), .ZN(n17677) );
  OAI21_X1 U20839 ( .B1(n18413), .B2(n17699), .A(n17677), .ZN(P3_U2783) );
  AOI22_X1 U20840 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17704), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17703), .ZN(n17678) );
  OAI21_X1 U20841 ( .B1(n17679), .B2(n17706), .A(n17678), .ZN(P3_U2784) );
  AOI22_X1 U20842 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17695), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17692), .ZN(n17680) );
  OAI21_X1 U20843 ( .B1(n18426), .B2(n17699), .A(n17680), .ZN(P3_U2785) );
  AOI22_X1 U20844 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17695), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17692), .ZN(n17681) );
  OAI21_X1 U20845 ( .B1(n18431), .B2(n17699), .A(n17681), .ZN(P3_U2786) );
  AOI22_X1 U20846 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17695), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17692), .ZN(n17682) );
  OAI21_X1 U20847 ( .B1(n18436), .B2(n17699), .A(n17682), .ZN(P3_U2787) );
  AOI22_X1 U20848 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17695), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17692), .ZN(n17683) );
  OAI21_X1 U20849 ( .B1(n18441), .B2(n17699), .A(n17683), .ZN(P3_U2788) );
  AOI22_X1 U20850 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17695), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17692), .ZN(n17684) );
  OAI21_X1 U20851 ( .B1(n18446), .B2(n17699), .A(n17684), .ZN(P3_U2789) );
  AOI22_X1 U20852 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17695), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17692), .ZN(n17685) );
  OAI21_X1 U20853 ( .B1(n18451), .B2(n17699), .A(n17685), .ZN(P3_U2790) );
  AOI22_X1 U20854 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17695), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17692), .ZN(n17686) );
  OAI21_X1 U20855 ( .B1(n17687), .B2(n17699), .A(n17686), .ZN(P3_U2791) );
  AOI22_X1 U20856 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17695), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17692), .ZN(n17688) );
  OAI21_X1 U20857 ( .B1(n17689), .B2(n17699), .A(n17688), .ZN(P3_U2792) );
  AOI22_X1 U20858 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17695), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17692), .ZN(n17690) );
  OAI21_X1 U20859 ( .B1(n17691), .B2(n17699), .A(n17690), .ZN(P3_U2793) );
  AOI22_X1 U20860 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17695), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17692), .ZN(n17693) );
  OAI21_X1 U20861 ( .B1(n17694), .B2(n17699), .A(n17693), .ZN(P3_U2794) );
  AOI22_X1 U20862 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17695), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17703), .ZN(n17696) );
  OAI21_X1 U20863 ( .B1(n17697), .B2(n17699), .A(n17696), .ZN(P3_U2795) );
  AOI22_X1 U20864 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17695), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17703), .ZN(n17698) );
  OAI21_X1 U20865 ( .B1(n17700), .B2(n17699), .A(n17698), .ZN(P3_U2796) );
  AOI22_X1 U20866 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17704), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17703), .ZN(n17701) );
  OAI21_X1 U20867 ( .B1(n17702), .B2(n17706), .A(n17701), .ZN(P3_U2797) );
  AOI22_X1 U20868 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17704), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17703), .ZN(n17705) );
  OAI21_X1 U20869 ( .B1(n17707), .B2(n17706), .A(n17705), .ZN(P3_U2798) );
  INV_X1 U20870 ( .A(n17742), .ZN(n17731) );
  AOI21_X1 U20871 ( .B1(n17709), .B2(n17708), .A(n17984), .ZN(n17725) );
  INV_X1 U20872 ( .A(n17710), .ZN(n17724) );
  NAND2_X1 U20873 ( .A1(n17711), .A2(n17918), .ZN(n17718) );
  INV_X1 U20874 ( .A(n17713), .ZN(n17712) );
  NOR3_X1 U20875 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17879), .A3(
        n17712), .ZN(n17739) );
  INV_X1 U20876 ( .A(n18041), .ZN(n17922) );
  OAI21_X1 U20877 ( .B1(n17713), .B2(n17922), .A(n18080), .ZN(n17714) );
  AOI21_X1 U20878 ( .B1(n17757), .B2(n17715), .A(n17714), .ZN(n17747) );
  OAI21_X1 U20879 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17830), .A(
        n17747), .ZN(n17740) );
  OAI21_X1 U20880 ( .B1(n17739), .B2(n17740), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17717) );
  OAI211_X1 U20881 ( .C1(n17719), .C2(n17718), .A(n17717), .B(n17716), .ZN(
        n17722) );
  AND2_X1 U20882 ( .A1(n17943), .A2(n17720), .ZN(n17721) );
  NOR2_X1 U20883 ( .A1(n18070), .A2(n17809), .ZN(n17827) );
  INV_X1 U20884 ( .A(n17827), .ZN(n17728) );
  OAI22_X1 U20885 ( .A1(n18084), .A2(n17726), .B1(n17999), .B2(n18090), .ZN(
        n17752) );
  OR2_X1 U20886 ( .A1(n17727), .A2(n17752), .ZN(n17741) );
  NAND3_X1 U20887 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17728), .A3(
        n17741), .ZN(n17729) );
  OAI211_X1 U20888 ( .C1(n17732), .C2(n17731), .A(n17730), .B(n17729), .ZN(
        P3_U2802) );
  INV_X1 U20889 ( .A(n17733), .ZN(n17734) );
  NAND2_X1 U20890 ( .A1(n17735), .A2(n17734), .ZN(n17736) );
  XOR2_X1 U20891 ( .A(n17819), .B(n17736), .Z(n18098) );
  OAI22_X1 U20892 ( .A1(n18380), .A2(n18986), .B1(n17926), .B2(n17737), .ZN(
        n17738) );
  AOI211_X1 U20893 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17740), .A(
        n17739), .B(n17738), .ZN(n17744) );
  OAI21_X1 U20894 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17742), .A(
        n17741), .ZN(n17743) );
  OAI211_X1 U20895 ( .C1(n18098), .C2(n17984), .A(n17744), .B(n17743), .ZN(
        P3_U2803) );
  AOI21_X1 U20896 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17746), .A(
        n17745), .ZN(n18105) );
  NAND2_X1 U20897 ( .A1(n17926), .A2(n17830), .ZN(n18073) );
  NOR2_X1 U20898 ( .A1(n18380), .A2(n18983), .ZN(n18102) );
  AOI221_X1 U20899 ( .B1(n17749), .B2(n17748), .C1(n18478), .C2(n17748), .A(
        n17747), .ZN(n17750) );
  AOI211_X1 U20900 ( .C1(n17751), .C2(n18073), .A(n18102), .B(n17750), .ZN(
        n17754) );
  NOR4_X1 U20901 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18112), .A3(
        n18152), .A4(n18115), .ZN(n18103) );
  AOI22_X1 U20902 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17752), .B1(
        n17812), .B2(n18103), .ZN(n17753) );
  OAI211_X1 U20903 ( .C1(n18105), .C2(n17984), .A(n17754), .B(n17753), .ZN(
        P3_U2804) );
  NAND2_X1 U20904 ( .A1(n17899), .A2(n17774), .ZN(n18125) );
  NOR2_X1 U20905 ( .A1(n10067), .A2(n18125), .ZN(n17755) );
  XOR2_X1 U20906 ( .A(n18115), .B(n17755), .Z(n18122) );
  NOR2_X1 U20907 ( .A1(n17759), .A2(n18478), .ZN(n17795) );
  AOI211_X1 U20908 ( .C1(n17757), .C2(n17756), .A(n18039), .B(n17795), .ZN(
        n17789) );
  OAI21_X1 U20909 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17830), .A(
        n17789), .ZN(n17771) );
  NOR2_X1 U20910 ( .A1(n18380), .A2(n18981), .ZN(n18117) );
  NOR2_X1 U20911 ( .A1(n17772), .A2(n17758), .ZN(n17762) );
  OAI211_X1 U20912 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17759), .B(n17918), .ZN(n17761) );
  OAI22_X1 U20913 ( .A1(n17762), .A2(n17761), .B1(n17760), .B2(n17926), .ZN(
        n17763) );
  AOI211_X1 U20914 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17771), .A(
        n18117), .B(n17763), .ZN(n17768) );
  INV_X1 U20915 ( .A(n18227), .ZN(n17900) );
  NAND3_X1 U20916 ( .A1(n17900), .A2(n17774), .A3(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17764) );
  XOR2_X1 U20917 ( .A(n17764), .B(n18115), .Z(n18119) );
  AOI21_X1 U20918 ( .B1(n10068), .B2(n17819), .A(n17765), .ZN(n17766) );
  XOR2_X1 U20919 ( .A(n17766), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18118) );
  AOI22_X1 U20920 ( .A1(n18070), .A2(n18119), .B1(n17996), .B2(n18118), .ZN(
        n17767) );
  OAI211_X1 U20921 ( .C1(n17999), .C2(n18122), .A(n17768), .B(n17767), .ZN(
        P3_U2805) );
  INV_X1 U20922 ( .A(n17769), .ZN(n17780) );
  NOR2_X1 U20923 ( .A1(n17879), .A2(n17770), .ZN(n17773) );
  NOR2_X1 U20924 ( .A1(n18380), .A2(n18979), .ZN(n18123) );
  AOI221_X1 U20925 ( .B1(n17773), .B2(n17772), .C1(n17771), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18123), .ZN(n17779) );
  AND2_X1 U20926 ( .A1(n10067), .A2(n17774), .ZN(n18124) );
  NAND2_X1 U20927 ( .A1(n17900), .A2(n17774), .ZN(n18126) );
  AOI22_X1 U20928 ( .A1(n18070), .A2(n18126), .B1(n17809), .B2(n18125), .ZN(
        n17790) );
  AOI21_X1 U20929 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17776), .A(
        n17775), .ZN(n18135) );
  OAI22_X1 U20930 ( .A1(n17790), .A2(n10067), .B1(n18135), .B2(n17984), .ZN(
        n17777) );
  AOI21_X1 U20931 ( .B1(n17812), .B2(n18124), .A(n17777), .ZN(n17778) );
  OAI211_X1 U20932 ( .C1(n17926), .C2(n17780), .A(n17779), .B(n17778), .ZN(
        P3_U2806) );
  AOI22_X1 U20933 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17819), .B1(
        n17782), .B2(n17797), .ZN(n17783) );
  NAND2_X1 U20934 ( .A1(n17781), .A2(n17783), .ZN(n17784) );
  XOR2_X1 U20935 ( .A(n17784), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(
        n18141) );
  NAND2_X1 U20936 ( .A1(n18393), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n18140) );
  INV_X1 U20937 ( .A(n17830), .ZN(n17786) );
  OAI21_X1 U20938 ( .B1(n17943), .B2(n17786), .A(n17785), .ZN(n17787) );
  OAI211_X1 U20939 ( .C1(n17789), .C2(n17788), .A(n18140), .B(n17787), .ZN(
        n17794) );
  NOR2_X1 U20940 ( .A1(n18152), .A2(n17887), .ZN(n17792) );
  INV_X1 U20941 ( .A(n17790), .ZN(n17791) );
  MUX2_X1 U20942 ( .A(n17792), .B(n17791), .S(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(n17793) );
  AOI211_X1 U20943 ( .C1(n9714), .C2(n17795), .A(n17794), .B(n17793), .ZN(
        n17796) );
  OAI21_X1 U20944 ( .B1(n17984), .B2(n18141), .A(n17796), .ZN(P3_U2807) );
  INV_X1 U20945 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18153) );
  INV_X1 U20946 ( .A(n17797), .ZN(n17799) );
  OAI221_X1 U20947 ( .B1(n17799), .B2(n17798), .C1(n17799), .C2(n18148), .A(
        n17781), .ZN(n17800) );
  XNOR2_X1 U20948 ( .A(n18153), .B(n17800), .ZN(n18160) );
  OAI22_X1 U20949 ( .A1(n17802), .A2(n17922), .B1(n17801), .B2(n18917), .ZN(
        n17803) );
  NOR2_X1 U20950 ( .A1(n18039), .A2(n17803), .ZN(n17832) );
  OAI21_X1 U20951 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17830), .A(
        n17832), .ZN(n17815) );
  NOR2_X1 U20952 ( .A1(n17879), .A2(n17804), .ZN(n17817) );
  OAI211_X1 U20953 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17817), .B(n17805), .ZN(n17806) );
  NAND2_X1 U20954 ( .A1(n18393), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18158) );
  OAI211_X1 U20955 ( .C1(n17926), .C2(n17807), .A(n17806), .B(n18158), .ZN(
        n17808) );
  AOI21_X1 U20956 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n17815), .A(
        n17808), .ZN(n17811) );
  AOI22_X1 U20957 ( .A1(n18070), .A2(n18227), .B1(n17809), .B2(n18218), .ZN(
        n17886) );
  OAI21_X1 U20958 ( .B1(n18148), .B2(n17827), .A(n17886), .ZN(n17824) );
  OAI222_X1 U20959 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18148), 
        .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17812), .C1(n18153), 
        .C2(n17824), .ZN(n17810) );
  OAI211_X1 U20960 ( .C1(n17984), .C2(n18160), .A(n17811), .B(n17810), .ZN(
        P3_U2808) );
  NAND2_X1 U20961 ( .A1(n18164), .A2(n17823), .ZN(n18168) );
  INV_X1 U20962 ( .A(n18162), .ZN(n18143) );
  NAND2_X1 U20963 ( .A1(n18143), .A2(n17812), .ZN(n17851) );
  OAI22_X1 U20964 ( .A1(n18380), .A2(n18974), .B1(n17926), .B2(n17813), .ZN(
        n17814) );
  AOI221_X1 U20965 ( .B1(n17817), .B2(n17816), .C1(n17815), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17814), .ZN(n17826) );
  INV_X1 U20966 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17852) );
  NOR3_X1 U20967 ( .A1(n17852), .A2(n17819), .A3(n17818), .ZN(n17840) );
  INV_X1 U20968 ( .A(n17820), .ZN(n17859) );
  AOI22_X1 U20969 ( .A1(n18164), .A2(n17840), .B1(n17859), .B2(n17821), .ZN(
        n17822) );
  XOR2_X1 U20970 ( .A(n17823), .B(n17822), .Z(n18161) );
  AOI22_X1 U20971 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17824), .B1(
        n17996), .B2(n18161), .ZN(n17825) );
  OAI211_X1 U20972 ( .C1(n18168), .C2(n17851), .A(n17826), .B(n17825), .ZN(
        P3_U2809) );
  NAND2_X1 U20973 ( .A1(n18143), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n18146) );
  INV_X1 U20974 ( .A(n18146), .ZN(n18172) );
  OAI21_X1 U20975 ( .B1(n17827), .B2(n18172), .A(n17886), .ZN(n17828) );
  INV_X1 U20976 ( .A(n17828), .ZN(n17850) );
  OAI221_X1 U20977 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17858), 
        .C1(n18183), .C2(n17840), .A(n17781), .ZN(n17829) );
  XOR2_X1 U20978 ( .A(n18150), .B(n17829), .Z(n18175) );
  NAND2_X1 U20979 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18150), .ZN(
        n18179) );
  NAND2_X1 U20980 ( .A1(n17831), .A2(n18786), .ZN(n17864) );
  AOI221_X1 U20981 ( .B1(n17834), .B2(n17833), .C1(n17864), .C2(n17833), .A(
        n17832), .ZN(n17835) );
  AOI221_X1 U20982 ( .B1(n17943), .B2(n17836), .C1(n17786), .C2(n17836), .A(
        n17835), .ZN(n17837) );
  NAND2_X1 U20983 ( .A1(n18393), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n18177) );
  OAI211_X1 U20984 ( .C1(n17851), .C2(n18179), .A(n17837), .B(n18177), .ZN(
        n17838) );
  AOI21_X1 U20985 ( .B1(n17996), .B2(n18175), .A(n17838), .ZN(n17839) );
  OAI21_X1 U20986 ( .B1(n17850), .B2(n18150), .A(n17839), .ZN(P3_U2810) );
  AOI21_X1 U20987 ( .B1(n17858), .B2(n17859), .A(n17840), .ZN(n17841) );
  XOR2_X1 U20988 ( .A(n18183), .B(n17841), .Z(n18180) );
  INV_X1 U20989 ( .A(n18078), .ZN(n18013) );
  OAI21_X1 U20990 ( .B1(n18039), .B2(n17843), .A(n18013), .ZN(n17863) );
  OAI21_X1 U20991 ( .B1(n17842), .B2(n18917), .A(n17863), .ZN(n17855) );
  AOI22_X1 U20992 ( .A1(n18393), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17855), .ZN(n17846) );
  NOR2_X1 U20993 ( .A1(n17879), .A2(n17843), .ZN(n17857) );
  NAND2_X1 U20994 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17844) );
  OAI211_X1 U20995 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17857), .B(n17844), .ZN(n17845) );
  OAI211_X1 U20996 ( .C1(n17926), .C2(n17847), .A(n17846), .B(n17845), .ZN(
        n17848) );
  AOI21_X1 U20997 ( .B1(n17996), .B2(n18180), .A(n17848), .ZN(n17849) );
  OAI221_X1 U20998 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17851), 
        .C1(n18183), .C2(n17850), .A(n17849), .ZN(P3_U2811) );
  NAND2_X1 U20999 ( .A1(n18193), .A2(n17852), .ZN(n18199) );
  OAI22_X1 U21000 ( .A1(n18380), .A2(n18967), .B1(n17926), .B2(n17853), .ZN(
        n17854) );
  AOI221_X1 U21001 ( .B1(n17857), .B2(n17856), .C1(n17855), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17854), .ZN(n17862) );
  OAI21_X1 U21002 ( .B1(n18193), .B2(n17887), .A(n17886), .ZN(n17870) );
  AOI21_X1 U21003 ( .B1(n10059), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17858), .ZN(n17860) );
  XOR2_X1 U21004 ( .A(n17860), .B(n17859), .Z(n18195) );
  AOI22_X1 U21005 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17870), .B1(
        n17996), .B2(n18195), .ZN(n17861) );
  OAI211_X1 U21006 ( .C1(n17887), .C2(n18199), .A(n17862), .B(n17861), .ZN(
        P3_U2812) );
  NAND2_X1 U21007 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18200), .ZN(
        n18204) );
  NOR2_X1 U21008 ( .A1(n18380), .A2(n18965), .ZN(n18202) );
  AOI21_X1 U21009 ( .B1(n17865), .B2(n17864), .A(n17863), .ZN(n17866) );
  AOI211_X1 U21010 ( .C1(n17867), .C2(n18073), .A(n18202), .B(n17866), .ZN(
        n17872) );
  OAI21_X1 U21011 ( .B1(n17869), .B2(n18200), .A(n17868), .ZN(n18203) );
  AOI22_X1 U21012 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17870), .B1(
        n17996), .B2(n18203), .ZN(n17871) );
  OAI211_X1 U21013 ( .C1(n17887), .C2(n18204), .A(n17872), .B(n17871), .ZN(
        P3_U2813) );
  AOI21_X1 U21014 ( .B1(n10059), .B2(n13026), .A(n17873), .ZN(n17874) );
  XOR2_X1 U21015 ( .A(n17874), .B(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .Z(
        n18210) );
  AOI21_X1 U21016 ( .B1(n18041), .B2(n17875), .A(n18039), .ZN(n17917) );
  OAI21_X1 U21017 ( .B1(n17876), .B2(n18917), .A(n17917), .ZN(n17896) );
  AOI22_X1 U21018 ( .A1(n18393), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17896), .ZN(n17882) );
  NOR3_X1 U21019 ( .A1(n17879), .A2(n17878), .A3(n17877), .ZN(n17898) );
  NAND2_X1 U21020 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17880) );
  OAI211_X1 U21021 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17898), .B(n17880), .ZN(n17881) );
  OAI211_X1 U21022 ( .C1(n17926), .C2(n17883), .A(n17882), .B(n17881), .ZN(
        n17884) );
  AOI21_X1 U21023 ( .B1(n17996), .B2(n18210), .A(n17884), .ZN(n17885) );
  OAI221_X1 U21024 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17887), 
        .C1(n18213), .C2(n17886), .A(n17885), .ZN(P3_U2814) );
  INV_X1 U21025 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17909) );
  INV_X1 U21026 ( .A(n18262), .ZN(n18246) );
  INV_X1 U21027 ( .A(n17910), .ZN(n17889) );
  INV_X1 U21028 ( .A(n17931), .ZN(n17888) );
  NAND3_X1 U21029 ( .A1(n18246), .A2(n17889), .A3(n17888), .ZN(n17890) );
  NAND2_X1 U21030 ( .A1(n17891), .A2(n17890), .ZN(n17892) );
  OAI221_X1 U21031 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17909), 
        .C1(n18261), .C2(n10059), .A(n17892), .ZN(n17893) );
  XOR2_X1 U21032 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17893), .Z(
        n18230) );
  OAI22_X1 U21033 ( .A1(n18380), .A2(n18961), .B1(n17926), .B2(n17894), .ZN(
        n17895) );
  AOI221_X1 U21034 ( .B1(n17898), .B2(n17897), .C1(n17896), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17895), .ZN(n17904) );
  NOR2_X1 U21035 ( .A1(n17899), .A2(n17999), .ZN(n17902) );
  INV_X1 U21036 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18223) );
  NAND2_X1 U21037 ( .A1(n18208), .A2(n17955), .ZN(n17912) );
  NAND2_X1 U21038 ( .A1(n18223), .A2(n17912), .ZN(n18217) );
  NOR2_X1 U21039 ( .A1(n17900), .A2(n18084), .ZN(n17901) );
  NOR2_X1 U21040 ( .A1(n18258), .A2(n18244), .ZN(n17930) );
  INV_X1 U21041 ( .A(n17930), .ZN(n18251) );
  OAI21_X1 U21042 ( .B1(n17910), .B2(n18251), .A(n18223), .ZN(n18226) );
  AOI22_X1 U21043 ( .A1(n17902), .A2(n18217), .B1(n17901), .B2(n18226), .ZN(
        n17903) );
  OAI211_X1 U21044 ( .C1(n17984), .C2(n18230), .A(n17904), .B(n17903), .ZN(
        P3_U2815) );
  NAND2_X1 U21045 ( .A1(n17985), .A2(n18786), .ZN(n17951) );
  NOR2_X1 U21046 ( .A1(n17905), .A2(n17951), .ZN(n17954) );
  AOI21_X1 U21047 ( .B1(n17920), .B2(n17954), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17916) );
  AOI22_X1 U21048 ( .A1(n18393), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n17906), 
        .B2(n18073), .ZN(n17915) );
  NOR2_X1 U21049 ( .A1(n18258), .A2(n17933), .ZN(n18232) );
  NAND2_X1 U21050 ( .A1(n10059), .A2(n17955), .ZN(n17949) );
  INV_X1 U21051 ( .A(n17949), .ZN(n17972) );
  AOI21_X1 U21052 ( .B1(n18232), .B2(n17972), .A(n17907), .ZN(n17908) );
  XOR2_X1 U21053 ( .A(n17909), .B(n17908), .Z(n18239) );
  NOR2_X1 U21054 ( .A1(n17933), .A2(n18251), .ZN(n17911) );
  OAI22_X1 U21055 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17911), .B1(
        n17910), .B2(n18251), .ZN(n18237) );
  OAI221_X1 U21056 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17955), 
        .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18232), .A(n17912), .ZN(
        n18236) );
  OAI22_X1 U21057 ( .A1(n18084), .A2(n18237), .B1(n17999), .B2(n18236), .ZN(
        n17913) );
  AOI21_X1 U21058 ( .B1(n17996), .B2(n18239), .A(n17913), .ZN(n17914) );
  OAI211_X1 U21059 ( .C1(n17917), .C2(n17916), .A(n17915), .B(n17914), .ZN(
        P3_U2816) );
  INV_X1 U21060 ( .A(n17980), .ZN(n17967) );
  NAND2_X1 U21061 ( .A1(n18231), .A2(n17933), .ZN(n18257) );
  NAND2_X1 U21062 ( .A1(n17919), .A2(n17918), .ZN(n17940) );
  AOI211_X1 U21063 ( .C1(n17939), .C2(n17927), .A(n17920), .B(n17940), .ZN(
        n17929) );
  OAI21_X1 U21064 ( .B1(n17985), .B2(n17922), .A(n18080), .ZN(n18003) );
  OAI22_X1 U21065 ( .A1(n17923), .A2(n17922), .B1(n17921), .B2(n18917), .ZN(
        n17924) );
  NOR2_X1 U21066 ( .A1(n18003), .A2(n17924), .ZN(n17938) );
  OAI22_X1 U21067 ( .A1(n17938), .A2(n17927), .B1(n17926), .B2(n17925), .ZN(
        n17928) );
  AOI211_X1 U21068 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n18393), .A(n17929), 
        .B(n17928), .ZN(n17936) );
  NOR2_X1 U21069 ( .A1(n18258), .A2(n18272), .ZN(n18249) );
  OAI22_X1 U21070 ( .A1(n17930), .A2(n18084), .B1(n18249), .B2(n17999), .ZN(
        n17944) );
  OAI22_X1 U21071 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n10059), .B1(
        n17931), .B2(n18258), .ZN(n17932) );
  OAI21_X1 U21072 ( .B1(n10059), .B2(n9739), .A(n17932), .ZN(n17934) );
  XOR2_X1 U21073 ( .A(n17934), .B(n17933), .Z(n18245) );
  AOI22_X1 U21074 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17944), .B1(
        n17996), .B2(n18245), .ZN(n17935) );
  OAI211_X1 U21075 ( .C1(n17967), .C2(n18257), .A(n17936), .B(n17935), .ZN(
        P3_U2817) );
  AOI21_X1 U21076 ( .B1(n17972), .B2(n18246), .A(n9739), .ZN(n17937) );
  XNOR2_X1 U21077 ( .A(n18261), .B(n17937), .ZN(n18267) );
  NAND2_X1 U21078 ( .A1(n18393), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18265) );
  OAI221_X1 U21079 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17940), .C1(
        n17939), .C2(n17938), .A(n18265), .ZN(n17941) );
  AOI21_X1 U21080 ( .B1(n17943), .B2(n17942), .A(n17941), .ZN(n17947) );
  OAI21_X1 U21081 ( .B1(n18262), .B2(n17967), .A(n18261), .ZN(n17945) );
  NAND2_X1 U21082 ( .A1(n17945), .A2(n17944), .ZN(n17946) );
  OAI211_X1 U21083 ( .C1(n18267), .C2(n17984), .A(n17947), .B(n17946), .ZN(
        P3_U2818) );
  INV_X1 U21084 ( .A(n17963), .ZN(n18280) );
  OAI21_X1 U21085 ( .B1(n18280), .B2(n17949), .A(n17948), .ZN(n17950) );
  XOR2_X1 U21086 ( .A(n17950), .B(n10080), .Z(n18268) );
  INV_X1 U21087 ( .A(n17951), .ZN(n18005) );
  NAND3_X1 U21088 ( .A1(n17986), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        n18005), .ZN(n17975) );
  NOR2_X1 U21089 ( .A1(n17965), .A2(n17975), .ZN(n17964) );
  AOI21_X1 U21090 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18013), .A(
        n17964), .ZN(n17953) );
  OAI22_X1 U21091 ( .A1(n17954), .A2(n17953), .B1(n18065), .B2(n17952), .ZN(
        n17957) );
  NAND2_X1 U21092 ( .A1(n17963), .A2(n10080), .ZN(n18285) );
  OAI22_X1 U21093 ( .A1(n17955), .A2(n17999), .B1(n18084), .B2(n18277), .ZN(
        n17982) );
  AOI21_X1 U21094 ( .B1(n18280), .B2(n17980), .A(n17982), .ZN(n17966) );
  OAI22_X1 U21095 ( .A1(n17967), .A2(n18285), .B1(n17966), .B2(n10080), .ZN(
        n17956) );
  AOI211_X1 U21096 ( .C1(n18393), .C2(P3_REIP_REG_11__SCAN_IN), .A(n17957), 
        .B(n17956), .ZN(n17958) );
  OAI21_X1 U21097 ( .B1(n18268), .B2(n17984), .A(n17958), .ZN(P3_U2819) );
  NOR4_X1 U21098 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n10059), .A3(
        n18286), .A4(n17959), .ZN(n17962) );
  AOI221_X1 U21099 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17972), .C1(
        n17981), .C2(n17960), .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17961) );
  AOI211_X1 U21100 ( .C1(n17972), .C2(n17963), .A(n17962), .B(n17961), .ZN(
        n18289) );
  AOI211_X1 U21101 ( .C1(n17975), .C2(n17965), .A(n18078), .B(n17964), .ZN(
        n17969) );
  AOI221_X1 U21102 ( .B1(n17967), .B2(n18286), .C1(n17981), .C2(n18286), .A(
        n17966), .ZN(n17968) );
  AOI211_X1 U21103 ( .C1(n17996), .C2(n18289), .A(n17969), .B(n17968), .ZN(
        n17970) );
  NAND2_X1 U21104 ( .A1(n18393), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n18291) );
  OAI211_X1 U21105 ( .C1(n18065), .C2(n17971), .A(n17970), .B(n18291), .ZN(
        P3_U2820) );
  NOR2_X1 U21106 ( .A1(n17972), .A2(n17960), .ZN(n17973) );
  XOR2_X1 U21107 ( .A(n17973), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n18303) );
  INV_X1 U21108 ( .A(n17974), .ZN(n17978) );
  AND2_X1 U21109 ( .A1(n17986), .A2(n18005), .ZN(n17976) );
  OAI211_X1 U21110 ( .C1(n17976), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n18013), .B(n17975), .ZN(n17977) );
  NAND2_X1 U21111 ( .A1(n18393), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n18300) );
  OAI211_X1 U21112 ( .C1(n18065), .C2(n17978), .A(n17977), .B(n18300), .ZN(
        n17979) );
  AOI221_X1 U21113 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17982), .C1(
        n17981), .C2(n17980), .A(n17979), .ZN(n17983) );
  OAI21_X1 U21114 ( .B1(n18303), .B2(n17984), .A(n17983), .ZN(P3_U2821) );
  NAND2_X1 U21115 ( .A1(n17985), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17987) );
  AOI211_X1 U21116 ( .C1(n17988), .C2(n17987), .A(n17986), .B(n18478), .ZN(
        n17991) );
  INV_X1 U21117 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18948) );
  OAI22_X1 U21118 ( .A1(n18065), .A2(n17989), .B1(n18380), .B2(n18948), .ZN(
        n17990) );
  AOI211_X1 U21119 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n18003), .A(
        n17991), .B(n17990), .ZN(n17998) );
  AOI21_X1 U21120 ( .B1(n17993), .B2(n18312), .A(n17992), .ZN(n18316) );
  OAI21_X1 U21121 ( .B1(n10059), .B2(n17995), .A(n17994), .ZN(n18314) );
  AOI22_X1 U21122 ( .A1(n18070), .A2(n18316), .B1(n17996), .B2(n18314), .ZN(
        n17997) );
  OAI211_X1 U21123 ( .C1(n17999), .C2(n18320), .A(n17998), .B(n17997), .ZN(
        P3_U2822) );
  NAND2_X1 U21124 ( .A1(n18001), .A2(n18000), .ZN(n18002) );
  XOR2_X1 U21125 ( .A(n18002), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18329) );
  NOR2_X1 U21126 ( .A1(n18380), .A2(n18945), .ZN(n18321) );
  AOI221_X1 U21127 ( .B1(n18005), .B2(n18004), .C1(n18003), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18321), .ZN(n18010) );
  AOI21_X1 U21128 ( .B1(n18324), .B2(n18007), .A(n18006), .ZN(n18325) );
  AOI22_X1 U21129 ( .A1(n18074), .A2(n18325), .B1(n18008), .B2(n18073), .ZN(
        n18009) );
  OAI211_X1 U21130 ( .C1(n18084), .C2(n18329), .A(n18010), .B(n18009), .ZN(
        P3_U2823) );
  AOI21_X1 U21131 ( .B1(n18012), .B2(n18336), .A(n18011), .ZN(n18333) );
  OR2_X1 U21132 ( .A1(n18014), .A2(n18478), .ZN(n18020) );
  OAI21_X1 U21133 ( .B1(n18478), .B2(n18014), .A(n18013), .ZN(n18032) );
  AOI21_X1 U21134 ( .B1(n18017), .B2(n18016), .A(n18015), .ZN(n18331) );
  AOI22_X1 U21135 ( .A1(n18074), .A2(n18331), .B1(n18393), .B2(
        P3_REIP_REG_6__SCAN_IN), .ZN(n18018) );
  OAI221_X1 U21136 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18020), .C1(
        n18019), .C2(n18032), .A(n18018), .ZN(n18021) );
  AOI21_X1 U21137 ( .B1(n18070), .B2(n18333), .A(n18021), .ZN(n18022) );
  OAI21_X1 U21138 ( .B1(n18065), .B2(n18023), .A(n18022), .ZN(P3_U2824) );
  AOI21_X1 U21139 ( .B1(n18024), .B2(n18080), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18033) );
  AOI21_X1 U21140 ( .B1(n18344), .B2(n18026), .A(n18025), .ZN(n18337) );
  AOI22_X1 U21141 ( .A1(n18074), .A2(n18337), .B1(n18393), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n18031) );
  AOI21_X1 U21142 ( .B1(n18344), .B2(n18028), .A(n18027), .ZN(n18340) );
  AOI22_X1 U21143 ( .A1(n18070), .A2(n18340), .B1(n18029), .B2(n18073), .ZN(
        n18030) );
  OAI211_X1 U21144 ( .C1(n18033), .C2(n18032), .A(n18031), .B(n18030), .ZN(
        P3_U2825) );
  AOI21_X1 U21145 ( .B1(n18035), .B2(n18034), .A(n9792), .ZN(n18345) );
  AOI22_X1 U21146 ( .A1(n18074), .A2(n18345), .B1(n18393), .B2(
        P3_REIP_REG_4__SCAN_IN), .ZN(n18046) );
  AOI21_X1 U21147 ( .B1(n18038), .B2(n18037), .A(n18036), .ZN(n18349) );
  AOI21_X1 U21148 ( .B1(n18041), .B2(n18040), .A(n18039), .ZN(n18058) );
  OAI22_X1 U21149 ( .A1(n18065), .A2(n18043), .B1(n18058), .B2(n18042), .ZN(
        n18044) );
  AOI21_X1 U21150 ( .B1(n18070), .B2(n18349), .A(n18044), .ZN(n18045) );
  OAI211_X1 U21151 ( .C1(n18478), .C2(n18047), .A(n18046), .B(n18045), .ZN(
        P3_U2826) );
  AOI21_X1 U21152 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18080), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18057) );
  AOI21_X1 U21153 ( .B1(n18050), .B2(n18049), .A(n18048), .ZN(n18355) );
  AOI22_X1 U21154 ( .A1(n18074), .A2(n18355), .B1(n18393), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n18056) );
  AOI21_X1 U21155 ( .B1(n18053), .B2(n18052), .A(n18051), .ZN(n18356) );
  AOI22_X1 U21156 ( .A1(n18070), .A2(n18356), .B1(n18054), .B2(n18073), .ZN(
        n18055) );
  OAI211_X1 U21157 ( .C1(n18058), .C2(n18057), .A(n18056), .B(n18055), .ZN(
        P3_U2827) );
  INV_X1 U21158 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18068) );
  AOI21_X1 U21159 ( .B1(n18061), .B2(n18060), .A(n18059), .ZN(n18364) );
  NOR2_X1 U21160 ( .A1(n18380), .A2(n18935), .ZN(n18363) );
  INV_X1 U21161 ( .A(n18074), .ZN(n18083) );
  XNOR2_X1 U21162 ( .A(n18063), .B(n18062), .ZN(n18361) );
  OAI22_X1 U21163 ( .A1(n18065), .A2(n18064), .B1(n18083), .B2(n18361), .ZN(
        n18066) );
  AOI211_X1 U21164 ( .C1(n18070), .C2(n18364), .A(n18363), .B(n18066), .ZN(
        n18067) );
  OAI221_X1 U21165 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18478), .C1(
        n18068), .C2(n18080), .A(n18067), .ZN(P3_U2828) );
  XNOR2_X1 U21166 ( .A(n18069), .B(n18072), .ZN(n18379) );
  AOI22_X1 U21167 ( .A1(n18070), .A2(n18379), .B1(n18393), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18076) );
  AOI21_X1 U21168 ( .B1(n18072), .B2(n18079), .A(n18071), .ZN(n18385) );
  AOI22_X1 U21169 ( .A1(n18074), .A2(n18385), .B1(n18077), .B2(n18073), .ZN(
        n18075) );
  OAI211_X1 U21170 ( .C1(n18078), .C2(n18077), .A(n18076), .B(n18075), .ZN(
        P3_U2829) );
  INV_X1 U21171 ( .A(n18400), .ZN(n18085) );
  NAND3_X1 U21172 ( .A1(n19018), .A2(n18917), .A3(n18080), .ZN(n18081) );
  AOI22_X1 U21173 ( .A1(n18393), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18081), .ZN(n18082) );
  OAI221_X1 U21174 ( .B1(n18085), .B2(n18084), .C1(n18400), .C2(n18083), .A(
        n18082), .ZN(P3_U2830) );
  NAND2_X1 U21175 ( .A1(n18857), .A2(n19035), .ZN(n18368) );
  NAND2_X1 U21176 ( .A1(n18086), .A2(n18368), .ZN(n18189) );
  OAI21_X1 U21177 ( .B1(n18152), .B2(n18189), .A(n18306), .ZN(n18127) );
  OAI21_X1 U21178 ( .B1(n18108), .B2(n18367), .A(n18127), .ZN(n18110) );
  NAND2_X1 U21179 ( .A1(n18087), .A2(n18306), .ZN(n18088) );
  OAI211_X1 U21180 ( .C1(n18090), .C2(n18248), .A(n18089), .B(n18088), .ZN(
        n18091) );
  AOI211_X1 U21181 ( .C1(n18252), .C2(n18092), .A(n18110), .B(n18091), .ZN(
        n18100) );
  AOI22_X1 U21182 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18100), .B1(
        n18094), .B2(n18093), .ZN(n18095) );
  AOI21_X1 U21183 ( .B1(n18388), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n18095), .ZN(n18097) );
  NAND2_X1 U21184 ( .A1(n18393), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n18096) );
  OAI211_X1 U21185 ( .C1(n18098), .C2(n18302), .A(n18097), .B(n18096), .ZN(
        P3_U2835) );
  INV_X1 U21186 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18099) );
  AOI211_X1 U21187 ( .C1(n18394), .C2(n18100), .A(n18393), .B(n18099), .ZN(
        n18101) );
  AOI211_X1 U21188 ( .C1(n18103), .C2(n18142), .A(n18102), .B(n18101), .ZN(
        n18104) );
  OAI21_X1 U21189 ( .B1(n18105), .B2(n18302), .A(n18104), .ZN(P3_U2836) );
  NAND2_X1 U21190 ( .A1(n18155), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18107) );
  INV_X1 U21191 ( .A(n18190), .ZN(n18106) );
  AOI21_X1 U21192 ( .B1(n18143), .B2(n18106), .A(n18844), .ZN(n18145) );
  AOI21_X1 U21193 ( .B1(n18880), .B2(n18107), .A(n18145), .ZN(n18131) );
  OAI211_X1 U21194 ( .C1(n18108), .C2(n18844), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n18131), .ZN(n18109) );
  OAI21_X1 U21195 ( .B1(n18110), .B2(n18109), .A(n18394), .ZN(n18114) );
  OR2_X1 U21196 ( .A1(n18112), .A2(n18111), .ZN(n18113) );
  AOI222_X1 U21197 ( .A1(n18115), .A2(n18114), .B1(n18115), .B2(n18113), .C1(
        n18114), .C2(n18378), .ZN(n18116) );
  AOI211_X1 U21198 ( .C1(n18118), .C2(n18315), .A(n18117), .B(n18116), .ZN(
        n18121) );
  NAND2_X1 U21199 ( .A1(n18397), .A2(n18119), .ZN(n18120) );
  OAI211_X1 U21200 ( .C1(n18122), .C2(n18319), .A(n18121), .B(n18120), .ZN(
        P3_U2837) );
  AOI21_X1 U21201 ( .B1(n18124), .B2(n18142), .A(n18123), .ZN(n18134) );
  INV_X1 U21202 ( .A(n18248), .ZN(n18273) );
  AOI22_X1 U21203 ( .A1(n18252), .A2(n18126), .B1(n18273), .B2(n18125), .ZN(
        n18128) );
  NAND3_X1 U21204 ( .A1(n18128), .A2(n18378), .A3(n18127), .ZN(n18132) );
  NOR2_X1 U21205 ( .A1(n18129), .A2(n18132), .ZN(n18130) );
  AOI21_X1 U21206 ( .B1(n18131), .B2(n18130), .A(n18393), .ZN(n18137) );
  OAI211_X1 U21207 ( .C1(n18309), .C2(n18132), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n18137), .ZN(n18133) );
  OAI211_X1 U21208 ( .C1(n18135), .C2(n18302), .A(n18134), .B(n18133), .ZN(
        P3_U2838) );
  NOR3_X1 U21209 ( .A1(n18388), .A2(n18136), .A3(n18152), .ZN(n18138) );
  OAI21_X1 U21210 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18138), .A(
        n18137), .ZN(n18139) );
  OAI211_X1 U21211 ( .C1(n18141), .C2(n18302), .A(n18140), .B(n18139), .ZN(
        P3_U2839) );
  NAND2_X1 U21212 ( .A1(n18143), .A2(n18142), .ZN(n18184) );
  OAI22_X1 U21213 ( .A1(n18144), .A2(n18184), .B1(n18153), .B2(n18386), .ZN(
        n18157) );
  NAND2_X1 U21214 ( .A1(n18843), .A2(n18248), .ZN(n18279) );
  INV_X1 U21215 ( .A(n18279), .ZN(n18191) );
  AOI22_X1 U21216 ( .A1(n18252), .A2(n18227), .B1(n18273), .B2(n18218), .ZN(
        n18169) );
  AOI221_X1 U21217 ( .B1(n18147), .B2(n18851), .C1(n18146), .C2(n18851), .A(
        n18145), .ZN(n18171) );
  OAI211_X1 U21218 ( .C1(n18148), .C2(n18191), .A(n18169), .B(n18171), .ZN(
        n18149) );
  AOI21_X1 U21219 ( .B1(n18851), .B2(n18150), .A(n18149), .ZN(n18163) );
  NAND2_X1 U21220 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18151), .ZN(
        n18296) );
  INV_X1 U21221 ( .A(n18296), .ZN(n18270) );
  NAND2_X1 U21222 ( .A1(n18187), .A2(n18270), .ZN(n18206) );
  OAI22_X1 U21223 ( .A1(n18857), .A2(n18153), .B1(n18152), .B2(n18206), .ZN(
        n18154) );
  OAI211_X1 U21224 ( .C1(n18155), .C2(n18287), .A(n18163), .B(n18154), .ZN(
        n18156) );
  AOI22_X1 U21225 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18388), .B1(
        n18157), .B2(n18156), .ZN(n18159) );
  OAI211_X1 U21226 ( .C1(n18302), .C2(n18160), .A(n18159), .B(n18158), .ZN(
        P3_U2840) );
  AOI22_X1 U21227 ( .A1(n18393), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18315), 
        .B2(n18161), .ZN(n18167) );
  OAI21_X1 U21228 ( .B1(n18162), .B2(n18206), .A(n18857), .ZN(n18170) );
  OAI211_X1 U21229 ( .C1(n18387), .C2(n18164), .A(n18170), .B(n18163), .ZN(
        n18165) );
  OAI211_X1 U21230 ( .C1(n18386), .C2(n18165), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18380), .ZN(n18166) );
  OAI211_X1 U21231 ( .C1(n18168), .C2(n18184), .A(n18167), .B(n18166), .ZN(
        P3_U2841) );
  NAND2_X1 U21232 ( .A1(n18183), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18174) );
  NAND2_X1 U21233 ( .A1(n18394), .A2(n18169), .ZN(n18209) );
  OAI211_X1 U21234 ( .C1(n18172), .C2(n18191), .A(n18171), .B(n18170), .ZN(
        n18173) );
  OAI21_X1 U21235 ( .B1(n18209), .B2(n18173), .A(n18380), .ZN(n18182) );
  OAI21_X1 U21236 ( .B1(n18387), .B2(n18174), .A(n18182), .ZN(n18176) );
  AOI22_X1 U21237 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18176), .B1(
        n18315), .B2(n18175), .ZN(n18178) );
  OAI211_X1 U21238 ( .C1(n18184), .C2(n18179), .A(n18178), .B(n18177), .ZN(
        P3_U2842) );
  AOI22_X1 U21239 ( .A1(n18393), .A2(P3_REIP_REG_19__SCAN_IN), .B1(n18315), 
        .B2(n18180), .ZN(n18181) );
  OAI221_X1 U21240 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18184), 
        .C1(n18183), .C2(n18182), .A(n18181), .ZN(P3_U2843) );
  OAI22_X1 U21241 ( .A1(n18348), .A2(n18844), .B1(n18366), .B2(n18185), .ZN(
        n18354) );
  NAND2_X1 U21242 ( .A1(n18186), .A2(n18354), .ZN(n18323) );
  NOR2_X1 U21243 ( .A1(n18243), .A2(n18323), .ZN(n18215) );
  OAI211_X1 U21244 ( .C1(n18188), .C2(n18215), .A(n18187), .B(n18394), .ZN(
        n18214) );
  NAND2_X1 U21245 ( .A1(n18880), .A2(n18190), .ZN(n18192) );
  AOI22_X1 U21246 ( .A1(n18193), .A2(n18192), .B1(n18191), .B2(n18844), .ZN(
        n18194) );
  AOI221_X1 U21247 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18201), 
        .C1(n18367), .C2(n18201), .A(n18393), .ZN(n18196) );
  AOI22_X1 U21248 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18196), .B1(
        n18315), .B2(n18195), .ZN(n18198) );
  NAND2_X1 U21249 ( .A1(n18393), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18197) );
  OAI211_X1 U21250 ( .C1(n18199), .C2(n18214), .A(n18198), .B(n18197), .ZN(
        P3_U2844) );
  NOR2_X1 U21251 ( .A1(n18205), .A2(n18844), .ZN(n18271) );
  AOI21_X1 U21252 ( .B1(n18851), .B2(n18274), .A(n18271), .ZN(n18247) );
  OAI21_X1 U21253 ( .B1(n18223), .B2(n18857), .A(n18206), .ZN(n18207) );
  OAI211_X1 U21254 ( .C1(n18208), .C2(n18287), .A(n18247), .B(n18207), .ZN(
        n18216) );
  OAI221_X1 U21255 ( .B1(n18209), .B2(n18309), .C1(n18209), .C2(n18216), .A(
        n18380), .ZN(n18212) );
  AOI22_X1 U21256 ( .A1(n18393), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18315), 
        .B2(n18210), .ZN(n18211) );
  OAI221_X1 U21257 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18214), 
        .C1(n18213), .C2(n18212), .A(n18211), .ZN(P3_U2846) );
  AND2_X1 U21258 ( .A1(n18215), .A2(n18232), .ZN(n18234) );
  OAI21_X1 U21259 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18234), .A(
        n18216), .ZN(n18221) );
  INV_X1 U21260 ( .A(n18217), .ZN(n18220) );
  NAND2_X1 U21261 ( .A1(n18273), .A2(n18218), .ZN(n18219) );
  OAI22_X1 U21262 ( .A1(n18222), .A2(n18221), .B1(n18220), .B2(n18219), .ZN(
        n18225) );
  OAI22_X1 U21263 ( .A1(n18223), .A2(n18378), .B1(n18380), .B2(n18961), .ZN(
        n18224) );
  AOI21_X1 U21264 ( .B1(n18394), .B2(n18225), .A(n18224), .ZN(n18229) );
  NAND3_X1 U21265 ( .A1(n18397), .A2(n18227), .A3(n18226), .ZN(n18228) );
  OAI211_X1 U21266 ( .C1(n18230), .C2(n18302), .A(n18229), .B(n18228), .ZN(
        P3_U2847) );
  AOI21_X1 U21267 ( .B1(n18231), .B2(n18270), .A(n18871), .ZN(n18254) );
  OAI211_X1 U21268 ( .C1(n18233), .C2(n18232), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18247), .ZN(n18235) );
  OAI22_X1 U21269 ( .A1(n18254), .A2(n18235), .B1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18234), .ZN(n18242) );
  AOI22_X1 U21270 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18388), .B1(
        n18393), .B2(P3_REIP_REG_14__SCAN_IN), .ZN(n18241) );
  OAI22_X1 U21271 ( .A1(n18391), .A2(n18237), .B1(n18319), .B2(n18236), .ZN(
        n18238) );
  AOI21_X1 U21272 ( .B1(n18315), .B2(n18239), .A(n18238), .ZN(n18240) );
  OAI211_X1 U21273 ( .C1(n18386), .C2(n18242), .A(n18241), .B(n18240), .ZN(
        P3_U2848) );
  NOR2_X1 U21274 ( .A1(n18386), .A2(n18323), .ZN(n18332) );
  INV_X1 U21275 ( .A(n18332), .ZN(n18304) );
  OAI222_X1 U21276 ( .A1(n18244), .A2(n18391), .B1(n18272), .B2(n18319), .C1(
        n18243), .C2(n18304), .ZN(n18299) );
  INV_X1 U21277 ( .A(n18299), .ZN(n18294) );
  AOI22_X1 U21278 ( .A1(n18393), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18315), 
        .B2(n18245), .ZN(n18256) );
  NOR2_X1 U21279 ( .A1(n18246), .A2(n18287), .ZN(n18282) );
  OAI21_X1 U21280 ( .B1(n18249), .B2(n18248), .A(n18247), .ZN(n18250) );
  AOI211_X1 U21281 ( .C1(n18252), .C2(n18251), .A(n18282), .B(n18250), .ZN(
        n18259) );
  OAI211_X1 U21282 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18287), .A(
        n18394), .B(n18259), .ZN(n18253) );
  OAI211_X1 U21283 ( .C1(n18254), .C2(n18253), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18380), .ZN(n18255) );
  OAI211_X1 U21284 ( .C1(n18294), .C2(n18257), .A(n18256), .B(n18255), .ZN(
        P3_U2849) );
  NOR2_X1 U21285 ( .A1(n18258), .A2(n18296), .ZN(n18260) );
  OAI211_X1 U21286 ( .C1(n18260), .C2(n18871), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n18259), .ZN(n18264) );
  OAI22_X1 U21287 ( .A1(n18294), .A2(n18262), .B1(n18261), .B2(n18386), .ZN(
        n18263) );
  AOI22_X1 U21288 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18388), .B1(
        n18264), .B2(n18263), .ZN(n18266) );
  OAI211_X1 U21289 ( .C1(n18267), .C2(n18302), .A(n18266), .B(n18265), .ZN(
        P3_U2850) );
  INV_X1 U21290 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18953) );
  OAI22_X1 U21291 ( .A1(n18380), .A2(n18953), .B1(n18302), .B2(n18268), .ZN(
        n18269) );
  INV_X1 U21292 ( .A(n18269), .ZN(n18284) );
  AOI21_X1 U21293 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18270), .A(
        n18871), .ZN(n18278) );
  AOI211_X1 U21294 ( .C1(n18273), .C2(n18272), .A(n18271), .B(n18386), .ZN(
        n18276) );
  NAND2_X1 U21295 ( .A1(n18851), .A2(n18274), .ZN(n18275) );
  OAI211_X1 U21296 ( .C1(n18277), .C2(n18843), .A(n18276), .B(n18275), .ZN(
        n18295) );
  AOI211_X1 U21297 ( .C1(n18280), .C2(n18279), .A(n18278), .B(n18295), .ZN(
        n18288) );
  OAI21_X1 U21298 ( .B1(n18871), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18288), .ZN(n18281) );
  OAI211_X1 U21299 ( .C1(n18282), .C2(n18281), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18380), .ZN(n18283) );
  OAI211_X1 U21300 ( .C1(n18294), .C2(n18285), .A(n18284), .B(n18283), .ZN(
        P3_U2851) );
  NAND2_X1 U21301 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18286), .ZN(
        n18293) );
  AOI221_X1 U21302 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18288), .C1(
        n18287), .C2(n18288), .A(n18393), .ZN(n18290) );
  AOI22_X1 U21303 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18290), .B1(
        n18315), .B2(n18289), .ZN(n18292) );
  OAI211_X1 U21304 ( .C1(n18294), .C2(n18293), .A(n18292), .B(n18291), .ZN(
        P3_U2852) );
  AOI21_X1 U21305 ( .B1(n18857), .B2(n18296), .A(n18295), .ZN(n18297) );
  OAI21_X1 U21306 ( .B1(n18393), .B2(n18297), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18298) );
  OAI21_X1 U21307 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18299), .A(
        n18298), .ZN(n18301) );
  OAI211_X1 U21308 ( .C1(n18303), .C2(n18302), .A(n18301), .B(n18300), .ZN(
        P3_U2853) );
  NOR3_X1 U21309 ( .A1(n18324), .A2(n18336), .A3(n18304), .ZN(n18313) );
  AOI22_X1 U21310 ( .A1(n18880), .A2(n18307), .B1(n18306), .B2(n18305), .ZN(
        n18308) );
  NAND2_X1 U21311 ( .A1(n18308), .A2(n18368), .ZN(n18330) );
  AOI211_X1 U21312 ( .C1(n18309), .C2(n18336), .A(n18324), .B(n18330), .ZN(
        n18322) );
  OAI21_X1 U21313 ( .B1(n18322), .B2(n18381), .A(n18378), .ZN(n18311) );
  NOR2_X1 U21314 ( .A1(n18380), .A2(n18948), .ZN(n18310) );
  AOI221_X1 U21315 ( .B1(n18313), .B2(n18312), .C1(n18311), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18310), .ZN(n18318) );
  AOI22_X1 U21316 ( .A1(n18397), .A2(n18316), .B1(n18315), .B2(n18314), .ZN(
        n18317) );
  OAI211_X1 U21317 ( .C1(n18320), .C2(n18319), .A(n18318), .B(n18317), .ZN(
        P3_U2854) );
  AOI21_X1 U21318 ( .B1(n18388), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18321), .ZN(n18328) );
  AOI221_X1 U21319 ( .B1(n18336), .B2(n18324), .C1(n18323), .C2(n18324), .A(
        n18322), .ZN(n18326) );
  AOI22_X1 U21320 ( .A1(n18394), .A2(n18326), .B1(n18384), .B2(n18325), .ZN(
        n18327) );
  OAI211_X1 U21321 ( .C1(n18391), .C2(n18329), .A(n18328), .B(n18327), .ZN(
        P3_U2855) );
  OAI21_X1 U21322 ( .B1(n18386), .B2(n18330), .A(n18380), .ZN(n18343) );
  AOI22_X1 U21323 ( .A1(n18393), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n18384), 
        .B2(n18331), .ZN(n18335) );
  AOI22_X1 U21324 ( .A1(n18333), .A2(n18397), .B1(n18332), .B2(n18336), .ZN(
        n18334) );
  OAI211_X1 U21325 ( .C1(n18336), .C2(n18343), .A(n18335), .B(n18334), .ZN(
        P3_U2856) );
  AOI22_X1 U21326 ( .A1(n18393), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18384), 
        .B2(n18337), .ZN(n18342) );
  NAND3_X1 U21327 ( .A1(n18394), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18354), .ZN(n18353) );
  NOR3_X1 U21328 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18338), .A3(
        n18353), .ZN(n18339) );
  AOI21_X1 U21329 ( .B1(n18340), .B2(n18397), .A(n18339), .ZN(n18341) );
  OAI211_X1 U21330 ( .C1(n18344), .C2(n18343), .A(n18342), .B(n18341), .ZN(
        P3_U2857) );
  AOI22_X1 U21331 ( .A1(n18393), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18384), 
        .B2(n18345), .ZN(n18352) );
  OAI211_X1 U21332 ( .C1(n18367), .C2(n18346), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n18368), .ZN(n18347) );
  AOI21_X1 U21333 ( .B1(n18880), .B2(n18348), .A(n18347), .ZN(n18360) );
  OAI21_X1 U21334 ( .B1(n18360), .B2(n18381), .A(n18378), .ZN(n18350) );
  AOI22_X1 U21335 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18350), .B1(
        n18397), .B2(n18349), .ZN(n18351) );
  OAI211_X1 U21336 ( .C1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n18353), .A(
        n18352), .B(n18351), .ZN(P3_U2858) );
  OAI21_X1 U21337 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18354), .A(
        n18394), .ZN(n18359) );
  AOI22_X1 U21338 ( .A1(n18393), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n18384), 
        .B2(n18355), .ZN(n18358) );
  AOI22_X1 U21339 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18388), .B1(
        n18397), .B2(n18356), .ZN(n18357) );
  OAI211_X1 U21340 ( .C1(n18360), .C2(n18359), .A(n18358), .B(n18357), .ZN(
        P3_U2859) );
  NOR2_X1 U21341 ( .A1(n18401), .A2(n18361), .ZN(n18362) );
  AOI211_X1 U21342 ( .C1(n18397), .C2(n18364), .A(n18363), .B(n18362), .ZN(
        n18377) );
  NOR2_X1 U21343 ( .A1(n18844), .A2(n18365), .ZN(n18375) );
  NOR2_X1 U21344 ( .A1(n19020), .A2(n18366), .ZN(n18373) );
  NOR2_X1 U21345 ( .A1(n19035), .A2(n19020), .ZN(n18370) );
  AOI21_X1 U21346 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18368), .A(
        n18367), .ZN(n18369) );
  AOI21_X1 U21347 ( .B1(n18370), .B2(n18880), .A(n18369), .ZN(n18371) );
  INV_X1 U21348 ( .A(n18371), .ZN(n18372) );
  MUX2_X1 U21349 ( .A(n18373), .B(n18372), .S(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n18374) );
  OAI21_X1 U21350 ( .B1(n18375), .B2(n18374), .A(n18394), .ZN(n18376) );
  OAI211_X1 U21351 ( .C1(n18378), .C2(n13001), .A(n18377), .B(n18376), .ZN(
        P3_U2860) );
  INV_X1 U21352 ( .A(n18379), .ZN(n18392) );
  NOR2_X1 U21353 ( .A1(n18380), .A2(n19039), .ZN(n18383) );
  AOI211_X1 U21354 ( .C1(n18859), .C2(n19035), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18381), .ZN(n18382) );
  AOI211_X1 U21355 ( .C1(n18385), .C2(n18384), .A(n18383), .B(n18382), .ZN(
        n18390) );
  NOR3_X1 U21356 ( .A1(n18387), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n18386), .ZN(n18396) );
  OAI21_X1 U21357 ( .B1(n18388), .B2(n18396), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18389) );
  OAI211_X1 U21358 ( .C1(n18392), .C2(n18391), .A(n18390), .B(n18389), .ZN(
        P3_U2861) );
  AOI211_X1 U21359 ( .C1(n18859), .C2(n18394), .A(n18393), .B(n19035), .ZN(
        n18395) );
  AOI211_X1 U21360 ( .C1(n18397), .C2(n18400), .A(n18396), .B(n18395), .ZN(
        n18399) );
  NAND2_X1 U21361 ( .A1(n18393), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18398) );
  OAI211_X1 U21362 ( .C1(n18401), .C2(n18400), .A(n18399), .B(n18398), .ZN(
        P3_U2862) );
  OAI211_X1 U21363 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n18402), .A(
        P3_STATE2_REG_2__SCAN_IN), .B(P3_STATE2_REG_1__SCAN_IN), .ZN(n18403)
         );
  INV_X1 U21364 ( .A(n18403), .ZN(n18898) );
  OAI21_X1 U21365 ( .B1(n18898), .B2(n18458), .A(n18408), .ZN(n18404) );
  OAI221_X1 U21366 ( .B1(n18414), .B2(n19053), .C1(n18414), .C2(n18408), .A(
        n18404), .ZN(P3_U2863) );
  NAND2_X1 U21367 ( .A1(n18884), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18682) );
  INV_X1 U21368 ( .A(n18682), .ZN(n18705) );
  NAND2_X1 U21369 ( .A1(n18887), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18567) );
  INV_X1 U21370 ( .A(n18567), .ZN(n18592) );
  NOR2_X1 U21371 ( .A1(n18705), .A2(n18592), .ZN(n18406) );
  OAI22_X1 U21372 ( .A1(n18407), .A2(n18887), .B1(n18406), .B2(n18405), .ZN(
        P3_U2866) );
  INV_X1 U21373 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18888) );
  NOR2_X1 U21374 ( .A1(n18888), .A2(n18408), .ZN(P3_U2867) );
  NOR2_X1 U21375 ( .A1(n18410), .A2(n18409), .ZN(n18450) );
  NAND2_X1 U21376 ( .A1(n18450), .A2(n18411), .ZN(n18790) );
  NAND2_X1 U21377 ( .A1(n18864), .A2(n18414), .ZN(n18866) );
  NAND2_X1 U21378 ( .A1(n18884), .A2(n18887), .ZN(n18501) );
  NOR2_X2 U21379 ( .A1(n18866), .A2(n18501), .ZN(n18520) );
  INV_X1 U21380 ( .A(n18520), .ZN(n18457) );
  INV_X1 U21381 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18412) );
  NOR2_X2 U21382 ( .A1(n18478), .A2(n18412), .ZN(n18782) );
  NAND2_X1 U21383 ( .A1(n18414), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18658) );
  INV_X1 U21384 ( .A(n18658), .ZN(n18415) );
  NOR2_X1 U21385 ( .A1(n18884), .A2(n18887), .ZN(n18732) );
  NAND2_X1 U21386 ( .A1(n18415), .A2(n18732), .ZN(n18779) );
  INV_X1 U21387 ( .A(n18779), .ZN(n18759) );
  NOR2_X2 U21388 ( .A1(n18525), .A2(n18413), .ZN(n18781) );
  INV_X1 U21389 ( .A(n18780), .ZN(n18907) );
  NOR2_X1 U21390 ( .A1(n18887), .A2(n18589), .ZN(n18784) );
  NAND2_X1 U21391 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18784), .ZN(
        n18836) );
  INV_X1 U21392 ( .A(n18836), .ZN(n18495) );
  NOR2_X1 U21393 ( .A1(n18495), .A2(n18520), .ZN(n18479) );
  NOR2_X1 U21394 ( .A1(n18907), .A2(n18479), .ZN(n18453) );
  AOI22_X1 U21395 ( .A1(n18782), .A2(n18759), .B1(n18781), .B2(n18453), .ZN(
        n18420) );
  NOR2_X1 U21396 ( .A1(n18414), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18636) );
  NOR2_X1 U21397 ( .A1(n18415), .A2(n18636), .ZN(n18708) );
  INV_X1 U21398 ( .A(n18708), .ZN(n18477) );
  NAND2_X1 U21399 ( .A1(n18477), .A2(n18732), .ZN(n18754) );
  INV_X1 U21400 ( .A(n18754), .ZN(n18417) );
  AOI211_X1 U21401 ( .C1(P3_STATE2_REG_3__SCAN_IN), .C2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18479), .B(n18525), .ZN(
        n18416) );
  AOI21_X1 U21402 ( .B1(n18417), .B2(n18786), .A(n18416), .ZN(n18454) );
  AND2_X1 U21403 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18786), .ZN(n18787) );
  INV_X1 U21404 ( .A(n18732), .ZN(n18418) );
  NOR2_X1 U21405 ( .A1(n18418), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18785) );
  NAND2_X1 U21406 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18785), .ZN(
        n18753) );
  INV_X1 U21407 ( .A(n18753), .ZN(n18829) );
  AOI22_X1 U21408 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18454), .B1(
        n18787), .B2(n18829), .ZN(n18419) );
  OAI211_X1 U21409 ( .C1(n18790), .C2(n18457), .A(n18420), .B(n18419), .ZN(
        P3_U2868) );
  NAND2_X1 U21410 ( .A1(n18450), .A2(n9969), .ZN(n18796) );
  AND2_X1 U21411 ( .A1(n18786), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18792) );
  AND2_X1 U21412 ( .A1(n18758), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18791) );
  AOI22_X1 U21413 ( .A1(n18792), .A2(n18759), .B1(n18791), .B2(n18453), .ZN(
        n18423) );
  NOR2_X2 U21414 ( .A1(n18421), .A2(n18478), .ZN(n18793) );
  AOI22_X1 U21415 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18454), .B1(
        n18793), .B2(n18829), .ZN(n18422) );
  OAI211_X1 U21416 ( .C1(n18796), .C2(n18457), .A(n18423), .B(n18422), .ZN(
        P3_U2869) );
  NAND2_X1 U21417 ( .A1(n18450), .A2(n18424), .ZN(n18802) );
  INV_X1 U21418 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n18425) );
  NOR2_X2 U21419 ( .A1(n18425), .A2(n18478), .ZN(n18799) );
  NOR2_X2 U21420 ( .A1(n18525), .A2(n18426), .ZN(n18797) );
  AOI22_X1 U21421 ( .A1(n18799), .A2(n18829), .B1(n18797), .B2(n18453), .ZN(
        n18428) );
  AND2_X1 U21422 ( .A1(n18786), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18798) );
  AOI22_X1 U21423 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18454), .B1(
        n18798), .B2(n18759), .ZN(n18427) );
  OAI211_X1 U21424 ( .C1(n18802), .C2(n18457), .A(n18428), .B(n18427), .ZN(
        P3_U2870) );
  NAND2_X1 U21425 ( .A1(n18450), .A2(n18429), .ZN(n18808) );
  NOR2_X2 U21426 ( .A1(n18430), .A2(n18478), .ZN(n18804) );
  NOR2_X2 U21427 ( .A1(n18525), .A2(n18431), .ZN(n18803) );
  AOI22_X1 U21428 ( .A1(n18804), .A2(n18829), .B1(n18803), .B2(n18453), .ZN(
        n18433) );
  NOR2_X2 U21429 ( .A1(n18478), .A2(n15249), .ZN(n18805) );
  AOI22_X1 U21430 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18454), .B1(
        n18805), .B2(n18759), .ZN(n18432) );
  OAI211_X1 U21431 ( .C1(n18808), .C2(n18457), .A(n18433), .B(n18432), .ZN(
        P3_U2871) );
  NAND2_X1 U21432 ( .A1(n18450), .A2(n18434), .ZN(n18814) );
  NOR2_X2 U21433 ( .A1(n18478), .A2(n18435), .ZN(n18811) );
  NOR2_X2 U21434 ( .A1(n18525), .A2(n18436), .ZN(n18809) );
  AOI22_X1 U21435 ( .A1(n18811), .A2(n18759), .B1(n18809), .B2(n18453), .ZN(
        n18438) );
  AND2_X1 U21436 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18786), .ZN(n18810) );
  AOI22_X1 U21437 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18454), .B1(
        n18810), .B2(n18829), .ZN(n18437) );
  OAI211_X1 U21438 ( .C1(n18814), .C2(n18457), .A(n18438), .B(n18437), .ZN(
        P3_U2872) );
  NAND2_X1 U21439 ( .A1(n18450), .A2(n18439), .ZN(n18820) );
  NOR2_X2 U21440 ( .A1(n18440), .A2(n18478), .ZN(n18816) );
  NOR2_X2 U21441 ( .A1(n18525), .A2(n18441), .ZN(n18815) );
  AOI22_X1 U21442 ( .A1(n18816), .A2(n18829), .B1(n18815), .B2(n18453), .ZN(
        n18443) );
  AND2_X1 U21443 ( .A1(n18786), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18817) );
  AOI22_X1 U21444 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18454), .B1(
        n18817), .B2(n18759), .ZN(n18442) );
  OAI211_X1 U21445 ( .C1(n18820), .C2(n18457), .A(n18443), .B(n18442), .ZN(
        P3_U2873) );
  NAND2_X1 U21446 ( .A1(n18450), .A2(n18444), .ZN(n18826) );
  INV_X1 U21447 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n18445) );
  NOR2_X2 U21448 ( .A1(n18478), .A2(n18445), .ZN(n18822) );
  NOR2_X2 U21449 ( .A1(n18525), .A2(n18446), .ZN(n18821) );
  AOI22_X1 U21450 ( .A1(n18822), .A2(n18759), .B1(n18821), .B2(n18453), .ZN(
        n18448) );
  NOR2_X2 U21451 ( .A1(n19429), .A2(n18478), .ZN(n18823) );
  AOI22_X1 U21452 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18454), .B1(
        n18823), .B2(n18829), .ZN(n18447) );
  OAI211_X1 U21453 ( .C1(n18826), .C2(n18457), .A(n18448), .B(n18447), .ZN(
        P3_U2874) );
  NAND2_X1 U21454 ( .A1(n18450), .A2(n18449), .ZN(n18837) );
  NOR2_X2 U21455 ( .A1(n18451), .A2(n18525), .ZN(n18828) );
  NOR2_X2 U21456 ( .A1(n18478), .A2(n18452), .ZN(n18832) );
  AOI22_X1 U21457 ( .A1(n18828), .A2(n18453), .B1(n18832), .B2(n18829), .ZN(
        n18456) );
  AND2_X1 U21458 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18786), .ZN(n18830) );
  AOI22_X1 U21459 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18454), .B1(
        n18830), .B2(n18759), .ZN(n18455) );
  OAI211_X1 U21460 ( .C1(n18837), .C2(n18457), .A(n18456), .B(n18455), .ZN(
        P3_U2875) );
  INV_X1 U21461 ( .A(n18501), .ZN(n18502) );
  NAND2_X1 U21462 ( .A1(n18636), .A2(n18502), .ZN(n18503) );
  NAND2_X1 U21463 ( .A1(n18864), .A2(n18780), .ZN(n18637) );
  NOR2_X1 U21464 ( .A1(n18501), .A2(n18637), .ZN(n18473) );
  AOI22_X1 U21465 ( .A1(n18787), .A2(n18759), .B1(n18781), .B2(n18473), .ZN(
        n18460) );
  NOR2_X1 U21466 ( .A1(n18525), .A2(n18458), .ZN(n18783) );
  AND2_X1 U21467 ( .A1(n18864), .A2(n18783), .ZN(n18731) );
  AOI22_X1 U21468 ( .A1(n18786), .A2(n18784), .B1(n18502), .B2(n18731), .ZN(
        n18474) );
  AOI22_X1 U21469 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18474), .B1(
        n18782), .B2(n18495), .ZN(n18459) );
  OAI211_X1 U21470 ( .C1(n18790), .C2(n18503), .A(n18460), .B(n18459), .ZN(
        P3_U2876) );
  AOI22_X1 U21471 ( .A1(n18792), .A2(n18495), .B1(n18791), .B2(n18473), .ZN(
        n18462) );
  AOI22_X1 U21472 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18474), .B1(
        n18793), .B2(n18759), .ZN(n18461) );
  OAI211_X1 U21473 ( .C1(n18796), .C2(n18503), .A(n18462), .B(n18461), .ZN(
        P3_U2877) );
  AOI22_X1 U21474 ( .A1(n18799), .A2(n18759), .B1(n18797), .B2(n18473), .ZN(
        n18464) );
  AOI22_X1 U21475 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18474), .B1(
        n18798), .B2(n18495), .ZN(n18463) );
  OAI211_X1 U21476 ( .C1(n18802), .C2(n18503), .A(n18464), .B(n18463), .ZN(
        P3_U2878) );
  AOI22_X1 U21477 ( .A1(n18804), .A2(n18759), .B1(n18803), .B2(n18473), .ZN(
        n18466) );
  AOI22_X1 U21478 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18474), .B1(
        n18805), .B2(n18495), .ZN(n18465) );
  OAI211_X1 U21479 ( .C1(n18808), .C2(n18503), .A(n18466), .B(n18465), .ZN(
        P3_U2879) );
  AOI22_X1 U21480 ( .A1(n18811), .A2(n18495), .B1(n18809), .B2(n18473), .ZN(
        n18468) );
  AOI22_X1 U21481 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18474), .B1(
        n18810), .B2(n18759), .ZN(n18467) );
  OAI211_X1 U21482 ( .C1(n18814), .C2(n18503), .A(n18468), .B(n18467), .ZN(
        P3_U2880) );
  AOI22_X1 U21483 ( .A1(n18817), .A2(n18495), .B1(n18815), .B2(n18473), .ZN(
        n18470) );
  AOI22_X1 U21484 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18474), .B1(
        n18816), .B2(n18759), .ZN(n18469) );
  OAI211_X1 U21485 ( .C1(n18820), .C2(n18503), .A(n18470), .B(n18469), .ZN(
        P3_U2881) );
  AOI22_X1 U21486 ( .A1(n18822), .A2(n18495), .B1(n18821), .B2(n18473), .ZN(
        n18472) );
  AOI22_X1 U21487 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18474), .B1(
        n18823), .B2(n18759), .ZN(n18471) );
  OAI211_X1 U21488 ( .C1(n18826), .C2(n18503), .A(n18472), .B(n18471), .ZN(
        P3_U2882) );
  AOI22_X1 U21489 ( .A1(n18830), .A2(n18495), .B1(n18828), .B2(n18473), .ZN(
        n18476) );
  AOI22_X1 U21490 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18474), .B1(
        n18832), .B2(n18759), .ZN(n18475) );
  OAI211_X1 U21491 ( .C1(n18837), .C2(n18503), .A(n18476), .B(n18475), .ZN(
        P3_U2883) );
  NOR2_X2 U21492 ( .A1(n18658), .A2(n18501), .ZN(n18563) );
  INV_X1 U21493 ( .A(n18563), .ZN(n18500) );
  NAND2_X1 U21494 ( .A1(n18780), .A2(n18477), .ZN(n18659) );
  NOR2_X1 U21495 ( .A1(n18501), .A2(n18659), .ZN(n18496) );
  AOI22_X1 U21496 ( .A1(n18787), .A2(n18495), .B1(n18781), .B2(n18496), .ZN(
        n18482) );
  NAND3_X1 U21497 ( .A1(n18502), .A2(n18758), .A3(n18477), .ZN(n18524) );
  OAI21_X1 U21498 ( .B1(n18479), .B2(n18478), .A(n18524), .ZN(n18480) );
  OAI21_X1 U21499 ( .B1(n18563), .B2(n19008), .A(n18480), .ZN(n18497) );
  AOI22_X1 U21500 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18497), .B1(
        n18782), .B2(n18520), .ZN(n18481) );
  OAI211_X1 U21501 ( .C1(n18790), .C2(n18500), .A(n18482), .B(n18481), .ZN(
        P3_U2884) );
  AOI22_X1 U21502 ( .A1(n18791), .A2(n18496), .B1(n18793), .B2(n18495), .ZN(
        n18484) );
  AOI22_X1 U21503 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18497), .B1(
        n18792), .B2(n18520), .ZN(n18483) );
  OAI211_X1 U21504 ( .C1(n18796), .C2(n18500), .A(n18484), .B(n18483), .ZN(
        P3_U2885) );
  AOI22_X1 U21505 ( .A1(n18798), .A2(n18520), .B1(n18797), .B2(n18496), .ZN(
        n18486) );
  AOI22_X1 U21506 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18497), .B1(
        n18799), .B2(n18495), .ZN(n18485) );
  OAI211_X1 U21507 ( .C1(n18802), .C2(n18500), .A(n18486), .B(n18485), .ZN(
        P3_U2886) );
  AOI22_X1 U21508 ( .A1(n18804), .A2(n18495), .B1(n18803), .B2(n18496), .ZN(
        n18488) );
  AOI22_X1 U21509 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18497), .B1(
        n18805), .B2(n18520), .ZN(n18487) );
  OAI211_X1 U21510 ( .C1(n18808), .C2(n18500), .A(n18488), .B(n18487), .ZN(
        P3_U2887) );
  AOI22_X1 U21511 ( .A1(n18811), .A2(n18520), .B1(n18809), .B2(n18496), .ZN(
        n18490) );
  AOI22_X1 U21512 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18497), .B1(
        n18810), .B2(n18495), .ZN(n18489) );
  OAI211_X1 U21513 ( .C1(n18814), .C2(n18500), .A(n18490), .B(n18489), .ZN(
        P3_U2888) );
  AOI22_X1 U21514 ( .A1(n18816), .A2(n18495), .B1(n18815), .B2(n18496), .ZN(
        n18492) );
  AOI22_X1 U21515 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18497), .B1(
        n18817), .B2(n18520), .ZN(n18491) );
  OAI211_X1 U21516 ( .C1(n18820), .C2(n18500), .A(n18492), .B(n18491), .ZN(
        P3_U2889) );
  AOI22_X1 U21517 ( .A1(n18823), .A2(n18495), .B1(n18821), .B2(n18496), .ZN(
        n18494) );
  AOI22_X1 U21518 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18497), .B1(
        n18822), .B2(n18520), .ZN(n18493) );
  OAI211_X1 U21519 ( .C1(n18826), .C2(n18500), .A(n18494), .B(n18493), .ZN(
        P3_U2890) );
  AOI22_X1 U21520 ( .A1(n18828), .A2(n18496), .B1(n18832), .B2(n18495), .ZN(
        n18499) );
  AOI22_X1 U21521 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18497), .B1(
        n18830), .B2(n18520), .ZN(n18498) );
  OAI211_X1 U21522 ( .C1(n18837), .C2(n18500), .A(n18499), .B(n18498), .ZN(
        P3_U2891) );
  NOR2_X1 U21523 ( .A1(n18864), .A2(n18501), .ZN(n18547) );
  NAND2_X1 U21524 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18547), .ZN(
        n18523) );
  AND2_X1 U21525 ( .A1(n18780), .A2(n18547), .ZN(n18518) );
  AOI22_X1 U21526 ( .A1(n18787), .A2(n18520), .B1(n18781), .B2(n18518), .ZN(
        n18505) );
  AOI21_X1 U21527 ( .B1(n18864), .B2(n18755), .A(n18525), .ZN(n18591) );
  OAI211_X1 U21528 ( .C1(n18584), .C2(n19008), .A(n18502), .B(n18591), .ZN(
        n18519) );
  INV_X1 U21529 ( .A(n18503), .ZN(n18541) );
  AOI22_X1 U21530 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18519), .B1(
        n18782), .B2(n18541), .ZN(n18504) );
  OAI211_X1 U21531 ( .C1(n18523), .C2(n18790), .A(n18505), .B(n18504), .ZN(
        P3_U2892) );
  AOI22_X1 U21532 ( .A1(n18791), .A2(n18518), .B1(n18793), .B2(n18520), .ZN(
        n18507) );
  AOI22_X1 U21533 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18519), .B1(
        n18792), .B2(n18541), .ZN(n18506) );
  OAI211_X1 U21534 ( .C1(n18523), .C2(n18796), .A(n18507), .B(n18506), .ZN(
        P3_U2893) );
  AOI22_X1 U21535 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18519), .B1(
        n18797), .B2(n18518), .ZN(n18509) );
  AOI22_X1 U21536 ( .A1(n18799), .A2(n18520), .B1(n18798), .B2(n18541), .ZN(
        n18508) );
  OAI211_X1 U21537 ( .C1(n18523), .C2(n18802), .A(n18509), .B(n18508), .ZN(
        P3_U2894) );
  AOI22_X1 U21538 ( .A1(n18803), .A2(n18518), .B1(n18805), .B2(n18541), .ZN(
        n18511) );
  AOI22_X1 U21539 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18519), .B1(
        n18804), .B2(n18520), .ZN(n18510) );
  OAI211_X1 U21540 ( .C1(n18523), .C2(n18808), .A(n18511), .B(n18510), .ZN(
        P3_U2895) );
  AOI22_X1 U21541 ( .A1(n18811), .A2(n18541), .B1(n18809), .B2(n18518), .ZN(
        n18513) );
  AOI22_X1 U21542 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18519), .B1(
        n18810), .B2(n18520), .ZN(n18512) );
  OAI211_X1 U21543 ( .C1(n18523), .C2(n18814), .A(n18513), .B(n18512), .ZN(
        P3_U2896) );
  AOI22_X1 U21544 ( .A1(n18817), .A2(n18541), .B1(n18815), .B2(n18518), .ZN(
        n18515) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18519), .B1(
        n18816), .B2(n18520), .ZN(n18514) );
  OAI211_X1 U21546 ( .C1(n18523), .C2(n18820), .A(n18515), .B(n18514), .ZN(
        P3_U2897) );
  AOI22_X1 U21547 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18519), .B1(
        n18821), .B2(n18518), .ZN(n18517) );
  AOI22_X1 U21548 ( .A1(n18822), .A2(n18541), .B1(n18823), .B2(n18520), .ZN(
        n18516) );
  OAI211_X1 U21549 ( .C1(n18523), .C2(n18826), .A(n18517), .B(n18516), .ZN(
        P3_U2898) );
  AOI22_X1 U21550 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18519), .B1(
        n18828), .B2(n18518), .ZN(n18522) );
  AOI22_X1 U21551 ( .A1(n18830), .A2(n18541), .B1(n18832), .B2(n18520), .ZN(
        n18521) );
  OAI211_X1 U21552 ( .C1(n18523), .C2(n18837), .A(n18522), .B(n18521), .ZN(
        P3_U2899) );
  NOR2_X2 U21553 ( .A1(n18866), .A2(n18567), .ZN(n18609) );
  INV_X1 U21554 ( .A(n18609), .ZN(n18546) );
  NOR2_X1 U21555 ( .A1(n18609), .A2(n18584), .ZN(n18568) );
  NOR2_X1 U21556 ( .A1(n18907), .A2(n18568), .ZN(n18542) );
  AOI22_X1 U21557 ( .A1(n18782), .A2(n18563), .B1(n18781), .B2(n18542), .ZN(
        n18528) );
  OAI22_X1 U21558 ( .A1(n18568), .A2(n18525), .B1(n18755), .B2(n18524), .ZN(
        n18526) );
  OAI21_X1 U21559 ( .B1(n18609), .B2(n19008), .A(n18526), .ZN(n18543) );
  AOI22_X1 U21560 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18543), .B1(
        n18787), .B2(n18541), .ZN(n18527) );
  OAI211_X1 U21561 ( .C1(n18546), .C2(n18790), .A(n18528), .B(n18527), .ZN(
        P3_U2900) );
  AOI22_X1 U21562 ( .A1(n18791), .A2(n18542), .B1(n18793), .B2(n18541), .ZN(
        n18530) );
  AOI22_X1 U21563 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18543), .B1(
        n18792), .B2(n18563), .ZN(n18529) );
  OAI211_X1 U21564 ( .C1(n18546), .C2(n18796), .A(n18530), .B(n18529), .ZN(
        P3_U2901) );
  AOI22_X1 U21565 ( .A1(n18798), .A2(n18563), .B1(n18797), .B2(n18542), .ZN(
        n18532) );
  AOI22_X1 U21566 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18543), .B1(
        n18799), .B2(n18541), .ZN(n18531) );
  OAI211_X1 U21567 ( .C1(n18546), .C2(n18802), .A(n18532), .B(n18531), .ZN(
        P3_U2902) );
  AOI22_X1 U21568 ( .A1(n18803), .A2(n18542), .B1(n18805), .B2(n18563), .ZN(
        n18534) );
  AOI22_X1 U21569 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18543), .B1(
        n18804), .B2(n18541), .ZN(n18533) );
  OAI211_X1 U21570 ( .C1(n18546), .C2(n18808), .A(n18534), .B(n18533), .ZN(
        P3_U2903) );
  AOI22_X1 U21571 ( .A1(n18811), .A2(n18563), .B1(n18809), .B2(n18542), .ZN(
        n18536) );
  AOI22_X1 U21572 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18543), .B1(
        n18810), .B2(n18541), .ZN(n18535) );
  OAI211_X1 U21573 ( .C1(n18546), .C2(n18814), .A(n18536), .B(n18535), .ZN(
        P3_U2904) );
  AOI22_X1 U21574 ( .A1(n18816), .A2(n18541), .B1(n18815), .B2(n18542), .ZN(
        n18538) );
  AOI22_X1 U21575 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18543), .B1(
        n18817), .B2(n18563), .ZN(n18537) );
  OAI211_X1 U21576 ( .C1(n18546), .C2(n18820), .A(n18538), .B(n18537), .ZN(
        P3_U2905) );
  AOI22_X1 U21577 ( .A1(n18822), .A2(n18563), .B1(n18821), .B2(n18542), .ZN(
        n18540) );
  AOI22_X1 U21578 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18543), .B1(
        n18823), .B2(n18541), .ZN(n18539) );
  OAI211_X1 U21579 ( .C1(n18546), .C2(n18826), .A(n18540), .B(n18539), .ZN(
        P3_U2906) );
  AOI22_X1 U21580 ( .A1(n18828), .A2(n18542), .B1(n18832), .B2(n18541), .ZN(
        n18545) );
  AOI22_X1 U21581 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18543), .B1(
        n18830), .B2(n18563), .ZN(n18544) );
  OAI211_X1 U21582 ( .C1(n18546), .C2(n18837), .A(n18545), .B(n18544), .ZN(
        P3_U2907) );
  NAND2_X1 U21583 ( .A1(n18592), .A2(n18636), .ZN(n18590) );
  NOR2_X1 U21584 ( .A1(n18567), .A2(n18637), .ZN(n18562) );
  AOI22_X1 U21585 ( .A1(n18584), .A2(n18782), .B1(n18781), .B2(n18562), .ZN(
        n18549) );
  AOI22_X1 U21586 ( .A1(n18786), .A2(n18547), .B1(n18592), .B2(n18731), .ZN(
        n18564) );
  AOI22_X1 U21587 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18564), .B1(
        n18787), .B2(n18563), .ZN(n18548) );
  OAI211_X1 U21588 ( .C1(n18590), .C2(n18790), .A(n18549), .B(n18548), .ZN(
        P3_U2908) );
  AOI22_X1 U21589 ( .A1(n18791), .A2(n18562), .B1(n18793), .B2(n18563), .ZN(
        n18551) );
  AOI22_X1 U21590 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18564), .B1(
        n18584), .B2(n18792), .ZN(n18550) );
  OAI211_X1 U21591 ( .C1(n18590), .C2(n18796), .A(n18551), .B(n18550), .ZN(
        P3_U2909) );
  AOI22_X1 U21592 ( .A1(n18584), .A2(n18798), .B1(n18797), .B2(n18562), .ZN(
        n18553) );
  AOI22_X1 U21593 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18564), .B1(
        n18799), .B2(n18563), .ZN(n18552) );
  OAI211_X1 U21594 ( .C1(n18590), .C2(n18802), .A(n18553), .B(n18552), .ZN(
        P3_U2910) );
  AOI22_X1 U21595 ( .A1(n18584), .A2(n18805), .B1(n18803), .B2(n18562), .ZN(
        n18555) );
  AOI22_X1 U21596 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18564), .B1(
        n18804), .B2(n18563), .ZN(n18554) );
  OAI211_X1 U21597 ( .C1(n18590), .C2(n18808), .A(n18555), .B(n18554), .ZN(
        P3_U2911) );
  AOI22_X1 U21598 ( .A1(n18810), .A2(n18563), .B1(n18809), .B2(n18562), .ZN(
        n18557) );
  AOI22_X1 U21599 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18564), .B1(
        n18584), .B2(n18811), .ZN(n18556) );
  OAI211_X1 U21600 ( .C1(n18590), .C2(n18814), .A(n18557), .B(n18556), .ZN(
        P3_U2912) );
  AOI22_X1 U21601 ( .A1(n18816), .A2(n18563), .B1(n18815), .B2(n18562), .ZN(
        n18559) );
  AOI22_X1 U21602 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18564), .B1(
        n18584), .B2(n18817), .ZN(n18558) );
  OAI211_X1 U21603 ( .C1(n18590), .C2(n18820), .A(n18559), .B(n18558), .ZN(
        P3_U2913) );
  AOI22_X1 U21604 ( .A1(n18584), .A2(n18822), .B1(n18821), .B2(n18562), .ZN(
        n18561) );
  AOI22_X1 U21605 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18564), .B1(
        n18823), .B2(n18563), .ZN(n18560) );
  OAI211_X1 U21606 ( .C1(n18590), .C2(n18826), .A(n18561), .B(n18560), .ZN(
        P3_U2914) );
  AOI22_X1 U21607 ( .A1(n18584), .A2(n18830), .B1(n18828), .B2(n18562), .ZN(
        n18566) );
  AOI22_X1 U21608 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18564), .B1(
        n18832), .B2(n18563), .ZN(n18565) );
  OAI211_X1 U21609 ( .C1(n18590), .C2(n18837), .A(n18566), .B(n18565), .ZN(
        P3_U2915) );
  NOR2_X2 U21610 ( .A1(n18658), .A2(n18567), .ZN(n18654) );
  INV_X1 U21611 ( .A(n18654), .ZN(n18588) );
  NOR2_X1 U21612 ( .A1(n18567), .A2(n18659), .ZN(n18613) );
  AOI22_X1 U21613 ( .A1(n18584), .A2(n18787), .B1(n18781), .B2(n18613), .ZN(
        n18571) );
  AOI221_X1 U21614 ( .B1(n18568), .B2(n18590), .C1(n18755), .C2(n18590), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18569) );
  OAI21_X1 U21615 ( .B1(n18654), .B2(n18569), .A(n18758), .ZN(n18585) );
  AOI22_X1 U21616 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18585), .B1(
        n18609), .B2(n18782), .ZN(n18570) );
  OAI211_X1 U21617 ( .C1(n18588), .C2(n18790), .A(n18571), .B(n18570), .ZN(
        P3_U2916) );
  AOI22_X1 U21618 ( .A1(n18584), .A2(n18793), .B1(n18613), .B2(n18791), .ZN(
        n18573) );
  AOI22_X1 U21619 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18585), .B1(
        n18609), .B2(n18792), .ZN(n18572) );
  OAI211_X1 U21620 ( .C1(n18588), .C2(n18796), .A(n18573), .B(n18572), .ZN(
        P3_U2917) );
  AOI22_X1 U21621 ( .A1(n18609), .A2(n18798), .B1(n18613), .B2(n18797), .ZN(
        n18575) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18585), .B1(
        n18584), .B2(n18799), .ZN(n18574) );
  OAI211_X1 U21623 ( .C1(n18588), .C2(n18802), .A(n18575), .B(n18574), .ZN(
        P3_U2918) );
  AOI22_X1 U21624 ( .A1(n18609), .A2(n18805), .B1(n18613), .B2(n18803), .ZN(
        n18577) );
  AOI22_X1 U21625 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18585), .B1(
        n18584), .B2(n18804), .ZN(n18576) );
  OAI211_X1 U21626 ( .C1(n18588), .C2(n18808), .A(n18577), .B(n18576), .ZN(
        P3_U2919) );
  AOI22_X1 U21627 ( .A1(n18609), .A2(n18811), .B1(n18613), .B2(n18809), .ZN(
        n18579) );
  AOI22_X1 U21628 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18585), .B1(
        n18584), .B2(n18810), .ZN(n18578) );
  OAI211_X1 U21629 ( .C1(n18588), .C2(n18814), .A(n18579), .B(n18578), .ZN(
        P3_U2920) );
  AOI22_X1 U21630 ( .A1(n18584), .A2(n18816), .B1(n18613), .B2(n18815), .ZN(
        n18581) );
  AOI22_X1 U21631 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18585), .B1(
        n18609), .B2(n18817), .ZN(n18580) );
  OAI211_X1 U21632 ( .C1(n18588), .C2(n18820), .A(n18581), .B(n18580), .ZN(
        P3_U2921) );
  AOI22_X1 U21633 ( .A1(n18584), .A2(n18823), .B1(n18613), .B2(n18821), .ZN(
        n18583) );
  AOI22_X1 U21634 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18585), .B1(
        n18609), .B2(n18822), .ZN(n18582) );
  OAI211_X1 U21635 ( .C1(n18588), .C2(n18826), .A(n18583), .B(n18582), .ZN(
        P3_U2922) );
  AOI22_X1 U21636 ( .A1(n18584), .A2(n18832), .B1(n18613), .B2(n18828), .ZN(
        n18587) );
  AOI22_X1 U21637 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18585), .B1(
        n18609), .B2(n18830), .ZN(n18586) );
  OAI211_X1 U21638 ( .C1(n18588), .C2(n18837), .A(n18587), .B(n18586), .ZN(
        P3_U2923) );
  NOR2_X1 U21639 ( .A1(n18589), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18638) );
  NAND2_X1 U21640 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18638), .ZN(
        n18612) );
  INV_X1 U21641 ( .A(n18590), .ZN(n18631) );
  AND2_X1 U21642 ( .A1(n18780), .A2(n18638), .ZN(n18607) );
  AOI22_X1 U21643 ( .A1(n18631), .A2(n18782), .B1(n18781), .B2(n18607), .ZN(
        n18594) );
  INV_X1 U21644 ( .A(n18612), .ZN(n18677) );
  OAI211_X1 U21645 ( .C1(n18677), .C2(n19008), .A(n18592), .B(n18591), .ZN(
        n18608) );
  AOI22_X1 U21646 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18608), .B1(
        n18609), .B2(n18787), .ZN(n18593) );
  OAI211_X1 U21647 ( .C1(n18790), .C2(n18612), .A(n18594), .B(n18593), .ZN(
        P3_U2924) );
  AOI22_X1 U21648 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18608), .B1(
        n18791), .B2(n18607), .ZN(n18596) );
  AOI22_X1 U21649 ( .A1(n18631), .A2(n18792), .B1(n18609), .B2(n18793), .ZN(
        n18595) );
  OAI211_X1 U21650 ( .C1(n18796), .C2(n18612), .A(n18596), .B(n18595), .ZN(
        P3_U2925) );
  AOI22_X1 U21651 ( .A1(n18631), .A2(n18798), .B1(n18797), .B2(n18607), .ZN(
        n18598) );
  AOI22_X1 U21652 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18608), .B1(
        n18609), .B2(n18799), .ZN(n18597) );
  OAI211_X1 U21653 ( .C1(n18802), .C2(n18612), .A(n18598), .B(n18597), .ZN(
        P3_U2926) );
  AOI22_X1 U21654 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18608), .B1(
        n18803), .B2(n18607), .ZN(n18600) );
  AOI22_X1 U21655 ( .A1(n18631), .A2(n18805), .B1(n18609), .B2(n18804), .ZN(
        n18599) );
  OAI211_X1 U21656 ( .C1(n18808), .C2(n18612), .A(n18600), .B(n18599), .ZN(
        P3_U2927) );
  AOI22_X1 U21657 ( .A1(n18609), .A2(n18810), .B1(n18809), .B2(n18607), .ZN(
        n18602) );
  AOI22_X1 U21658 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18608), .B1(
        n18631), .B2(n18811), .ZN(n18601) );
  OAI211_X1 U21659 ( .C1(n18814), .C2(n18612), .A(n18602), .B(n18601), .ZN(
        P3_U2928) );
  AOI22_X1 U21660 ( .A1(n18609), .A2(n18816), .B1(n18815), .B2(n18607), .ZN(
        n18604) );
  AOI22_X1 U21661 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18608), .B1(
        n18631), .B2(n18817), .ZN(n18603) );
  OAI211_X1 U21662 ( .C1(n18820), .C2(n18612), .A(n18604), .B(n18603), .ZN(
        P3_U2929) );
  AOI22_X1 U21663 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18608), .B1(
        n18821), .B2(n18607), .ZN(n18606) );
  AOI22_X1 U21664 ( .A1(n18631), .A2(n18822), .B1(n18609), .B2(n18823), .ZN(
        n18605) );
  OAI211_X1 U21665 ( .C1(n18826), .C2(n18612), .A(n18606), .B(n18605), .ZN(
        P3_U2930) );
  AOI22_X1 U21666 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18608), .B1(
        n18828), .B2(n18607), .ZN(n18611) );
  AOI22_X1 U21667 ( .A1(n18631), .A2(n18830), .B1(n18609), .B2(n18832), .ZN(
        n18610) );
  OAI211_X1 U21668 ( .C1(n18837), .C2(n18612), .A(n18611), .B(n18610), .ZN(
        P3_U2931) );
  NOR2_X2 U21669 ( .A1(n18866), .A2(n18682), .ZN(n18699) );
  INV_X1 U21670 ( .A(n18699), .ZN(n18635) );
  NOR2_X1 U21671 ( .A1(n18677), .A2(n18699), .ZN(n18660) );
  NOR2_X1 U21672 ( .A1(n18907), .A2(n18660), .ZN(n18630) );
  AOI22_X1 U21673 ( .A1(n18654), .A2(n18782), .B1(n18781), .B2(n18630), .ZN(
        n18617) );
  INV_X1 U21674 ( .A(n18613), .ZN(n18614) );
  OAI21_X1 U21675 ( .B1(n18755), .B2(n18614), .A(n18660), .ZN(n18615) );
  OAI211_X1 U21676 ( .C1(n18699), .C2(n19008), .A(n18758), .B(n18615), .ZN(
        n18632) );
  AOI22_X1 U21677 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18632), .B1(
        n18631), .B2(n18787), .ZN(n18616) );
  OAI211_X1 U21678 ( .C1(n18790), .C2(n18635), .A(n18617), .B(n18616), .ZN(
        P3_U2932) );
  AOI22_X1 U21679 ( .A1(n18631), .A2(n18793), .B1(n18791), .B2(n18630), .ZN(
        n18619) );
  AOI22_X1 U21680 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18632), .B1(
        n18654), .B2(n18792), .ZN(n18618) );
  OAI211_X1 U21681 ( .C1(n18796), .C2(n18635), .A(n18619), .B(n18618), .ZN(
        P3_U2933) );
  AOI22_X1 U21682 ( .A1(n18654), .A2(n18798), .B1(n18797), .B2(n18630), .ZN(
        n18621) );
  AOI22_X1 U21683 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18632), .B1(
        n18631), .B2(n18799), .ZN(n18620) );
  OAI211_X1 U21684 ( .C1(n18802), .C2(n18635), .A(n18621), .B(n18620), .ZN(
        P3_U2934) );
  AOI22_X1 U21685 ( .A1(n18631), .A2(n18804), .B1(n18803), .B2(n18630), .ZN(
        n18623) );
  AOI22_X1 U21686 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18632), .B1(
        n18654), .B2(n18805), .ZN(n18622) );
  OAI211_X1 U21687 ( .C1(n18808), .C2(n18635), .A(n18623), .B(n18622), .ZN(
        P3_U2935) );
  AOI22_X1 U21688 ( .A1(n18654), .A2(n18811), .B1(n18809), .B2(n18630), .ZN(
        n18625) );
  AOI22_X1 U21689 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18632), .B1(
        n18631), .B2(n18810), .ZN(n18624) );
  OAI211_X1 U21690 ( .C1(n18814), .C2(n18635), .A(n18625), .B(n18624), .ZN(
        P3_U2936) );
  AOI22_X1 U21691 ( .A1(n18631), .A2(n18816), .B1(n18815), .B2(n18630), .ZN(
        n18627) );
  AOI22_X1 U21692 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18632), .B1(
        n18654), .B2(n18817), .ZN(n18626) );
  OAI211_X1 U21693 ( .C1(n18820), .C2(n18635), .A(n18627), .B(n18626), .ZN(
        P3_U2937) );
  AOI22_X1 U21694 ( .A1(n18654), .A2(n18822), .B1(n18821), .B2(n18630), .ZN(
        n18629) );
  AOI22_X1 U21695 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18632), .B1(
        n18631), .B2(n18823), .ZN(n18628) );
  OAI211_X1 U21696 ( .C1(n18826), .C2(n18635), .A(n18629), .B(n18628), .ZN(
        P3_U2938) );
  AOI22_X1 U21697 ( .A1(n18654), .A2(n18830), .B1(n18828), .B2(n18630), .ZN(
        n18634) );
  AOI22_X1 U21698 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18632), .B1(
        n18631), .B2(n18832), .ZN(n18633) );
  OAI211_X1 U21699 ( .C1(n18837), .C2(n18635), .A(n18634), .B(n18633), .ZN(
        P3_U2939) );
  NAND2_X1 U21700 ( .A1(n18636), .A2(n18705), .ZN(n18684) );
  NOR2_X1 U21701 ( .A1(n18682), .A2(n18637), .ZN(n18653) );
  AOI22_X1 U21702 ( .A1(n18782), .A2(n18677), .B1(n18781), .B2(n18653), .ZN(
        n18640) );
  NOR2_X1 U21703 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18682), .ZN(
        n18683) );
  AOI22_X1 U21704 ( .A1(n18786), .A2(n18638), .B1(n18783), .B2(n18683), .ZN(
        n18655) );
  AOI22_X1 U21705 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18655), .B1(
        n18654), .B2(n18787), .ZN(n18639) );
  OAI211_X1 U21706 ( .C1(n18790), .C2(n18684), .A(n18640), .B(n18639), .ZN(
        P3_U2940) );
  AOI22_X1 U21707 ( .A1(n18654), .A2(n18793), .B1(n18791), .B2(n18653), .ZN(
        n18642) );
  AOI22_X1 U21708 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18655), .B1(
        n18792), .B2(n18677), .ZN(n18641) );
  OAI211_X1 U21709 ( .C1(n18796), .C2(n18684), .A(n18642), .B(n18641), .ZN(
        P3_U2941) );
  AOI22_X1 U21710 ( .A1(n18798), .A2(n18677), .B1(n18797), .B2(n18653), .ZN(
        n18644) );
  AOI22_X1 U21711 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18655), .B1(
        n18654), .B2(n18799), .ZN(n18643) );
  OAI211_X1 U21712 ( .C1(n18802), .C2(n18684), .A(n18644), .B(n18643), .ZN(
        P3_U2942) );
  AOI22_X1 U21713 ( .A1(n18654), .A2(n18804), .B1(n18803), .B2(n18653), .ZN(
        n18646) );
  AOI22_X1 U21714 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18655), .B1(
        n18805), .B2(n18677), .ZN(n18645) );
  OAI211_X1 U21715 ( .C1(n18808), .C2(n18684), .A(n18646), .B(n18645), .ZN(
        P3_U2943) );
  AOI22_X1 U21716 ( .A1(n18811), .A2(n18677), .B1(n18809), .B2(n18653), .ZN(
        n18648) );
  AOI22_X1 U21717 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18655), .B1(
        n18654), .B2(n18810), .ZN(n18647) );
  OAI211_X1 U21718 ( .C1(n18814), .C2(n18684), .A(n18648), .B(n18647), .ZN(
        P3_U2944) );
  AOI22_X1 U21719 ( .A1(n18817), .A2(n18677), .B1(n18815), .B2(n18653), .ZN(
        n18650) );
  AOI22_X1 U21720 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18655), .B1(
        n18654), .B2(n18816), .ZN(n18649) );
  OAI211_X1 U21721 ( .C1(n18820), .C2(n18684), .A(n18650), .B(n18649), .ZN(
        P3_U2945) );
  AOI22_X1 U21722 ( .A1(n18822), .A2(n18677), .B1(n18821), .B2(n18653), .ZN(
        n18652) );
  AOI22_X1 U21723 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18655), .B1(
        n18654), .B2(n18823), .ZN(n18651) );
  OAI211_X1 U21724 ( .C1(n18826), .C2(n18684), .A(n18652), .B(n18651), .ZN(
        P3_U2946) );
  AOI22_X1 U21725 ( .A1(n18830), .A2(n18677), .B1(n18828), .B2(n18653), .ZN(
        n18657) );
  AOI22_X1 U21726 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18655), .B1(
        n18654), .B2(n18832), .ZN(n18656) );
  OAI211_X1 U21727 ( .C1(n18837), .C2(n18684), .A(n18657), .B(n18656), .ZN(
        P3_U2947) );
  NOR2_X2 U21728 ( .A1(n18658), .A2(n18682), .ZN(n18748) );
  INV_X1 U21729 ( .A(n18748), .ZN(n18681) );
  NOR2_X1 U21730 ( .A1(n18659), .A2(n18682), .ZN(n18676) );
  AOI22_X1 U21731 ( .A1(n18782), .A2(n18699), .B1(n18781), .B2(n18676), .ZN(
        n18663) );
  AOI221_X1 U21732 ( .B1(n18660), .B2(n18684), .C1(n18755), .C2(n18684), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18661) );
  OAI21_X1 U21733 ( .B1(n18748), .B2(n18661), .A(n18758), .ZN(n18678) );
  AOI22_X1 U21734 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18678), .B1(
        n18787), .B2(n18677), .ZN(n18662) );
  OAI211_X1 U21735 ( .C1(n18790), .C2(n18681), .A(n18663), .B(n18662), .ZN(
        P3_U2948) );
  AOI22_X1 U21736 ( .A1(n18791), .A2(n18676), .B1(n18793), .B2(n18677), .ZN(
        n18665) );
  AOI22_X1 U21737 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18678), .B1(
        n18792), .B2(n18699), .ZN(n18664) );
  OAI211_X1 U21738 ( .C1(n18796), .C2(n18681), .A(n18665), .B(n18664), .ZN(
        P3_U2949) );
  AOI22_X1 U21739 ( .A1(n18798), .A2(n18699), .B1(n18797), .B2(n18676), .ZN(
        n18667) );
  AOI22_X1 U21740 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18678), .B1(
        n18799), .B2(n18677), .ZN(n18666) );
  OAI211_X1 U21741 ( .C1(n18802), .C2(n18681), .A(n18667), .B(n18666), .ZN(
        P3_U2950) );
  AOI22_X1 U21742 ( .A1(n18803), .A2(n18676), .B1(n18805), .B2(n18699), .ZN(
        n18669) );
  AOI22_X1 U21743 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18678), .B1(
        n18804), .B2(n18677), .ZN(n18668) );
  OAI211_X1 U21744 ( .C1(n18808), .C2(n18681), .A(n18669), .B(n18668), .ZN(
        P3_U2951) );
  AOI22_X1 U21745 ( .A1(n18811), .A2(n18699), .B1(n18809), .B2(n18676), .ZN(
        n18671) );
  AOI22_X1 U21746 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18678), .B1(
        n18810), .B2(n18677), .ZN(n18670) );
  OAI211_X1 U21747 ( .C1(n18814), .C2(n18681), .A(n18671), .B(n18670), .ZN(
        P3_U2952) );
  AOI22_X1 U21748 ( .A1(n18817), .A2(n18699), .B1(n18815), .B2(n18676), .ZN(
        n18673) );
  AOI22_X1 U21749 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18678), .B1(
        n18816), .B2(n18677), .ZN(n18672) );
  OAI211_X1 U21750 ( .C1(n18820), .C2(n18681), .A(n18673), .B(n18672), .ZN(
        P3_U2953) );
  AOI22_X1 U21751 ( .A1(n18823), .A2(n18677), .B1(n18821), .B2(n18676), .ZN(
        n18675) );
  AOI22_X1 U21752 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18678), .B1(
        n18822), .B2(n18699), .ZN(n18674) );
  OAI211_X1 U21753 ( .C1(n18826), .C2(n18681), .A(n18675), .B(n18674), .ZN(
        P3_U2954) );
  AOI22_X1 U21754 ( .A1(n18830), .A2(n18699), .B1(n18828), .B2(n18676), .ZN(
        n18680) );
  AOI22_X1 U21755 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18678), .B1(
        n18832), .B2(n18677), .ZN(n18679) );
  OAI211_X1 U21756 ( .C1(n18837), .C2(n18681), .A(n18680), .B(n18679), .ZN(
        P3_U2955) );
  NOR2_X1 U21757 ( .A1(n18864), .A2(n18682), .ZN(n18733) );
  NAND2_X1 U21758 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18733), .ZN(
        n18704) );
  AND2_X1 U21759 ( .A1(n18780), .A2(n18733), .ZN(n18700) );
  AOI22_X1 U21760 ( .A1(n18787), .A2(n18699), .B1(n18781), .B2(n18700), .ZN(
        n18686) );
  AOI22_X1 U21761 ( .A1(n18786), .A2(n18683), .B1(n18783), .B2(n18733), .ZN(
        n18701) );
  INV_X1 U21762 ( .A(n18684), .ZN(n18725) );
  AOI22_X1 U21763 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18701), .B1(
        n18782), .B2(n18725), .ZN(n18685) );
  OAI211_X1 U21764 ( .C1(n18790), .C2(n18704), .A(n18686), .B(n18685), .ZN(
        P3_U2956) );
  AOI22_X1 U21765 ( .A1(n18792), .A2(n18725), .B1(n18791), .B2(n18700), .ZN(
        n18688) );
  AOI22_X1 U21766 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18701), .B1(
        n18793), .B2(n18699), .ZN(n18687) );
  OAI211_X1 U21767 ( .C1(n18796), .C2(n18704), .A(n18688), .B(n18687), .ZN(
        P3_U2957) );
  AOI22_X1 U21768 ( .A1(n18798), .A2(n18725), .B1(n18797), .B2(n18700), .ZN(
        n18690) );
  AOI22_X1 U21769 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18701), .B1(
        n18799), .B2(n18699), .ZN(n18689) );
  OAI211_X1 U21770 ( .C1(n18802), .C2(n18704), .A(n18690), .B(n18689), .ZN(
        P3_U2958) );
  AOI22_X1 U21771 ( .A1(n18803), .A2(n18700), .B1(n18805), .B2(n18725), .ZN(
        n18692) );
  AOI22_X1 U21772 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18701), .B1(
        n18804), .B2(n18699), .ZN(n18691) );
  OAI211_X1 U21773 ( .C1(n18808), .C2(n18704), .A(n18692), .B(n18691), .ZN(
        P3_U2959) );
  AOI22_X1 U21774 ( .A1(n18810), .A2(n18699), .B1(n18809), .B2(n18700), .ZN(
        n18694) );
  AOI22_X1 U21775 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18701), .B1(
        n18811), .B2(n18725), .ZN(n18693) );
  OAI211_X1 U21776 ( .C1(n18814), .C2(n18704), .A(n18694), .B(n18693), .ZN(
        P3_U2960) );
  AOI22_X1 U21777 ( .A1(n18817), .A2(n18725), .B1(n18815), .B2(n18700), .ZN(
        n18696) );
  AOI22_X1 U21778 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18701), .B1(
        n18816), .B2(n18699), .ZN(n18695) );
  OAI211_X1 U21779 ( .C1(n18820), .C2(n18704), .A(n18696), .B(n18695), .ZN(
        P3_U2961) );
  AOI22_X1 U21780 ( .A1(n18822), .A2(n18725), .B1(n18821), .B2(n18700), .ZN(
        n18698) );
  AOI22_X1 U21781 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18701), .B1(
        n18823), .B2(n18699), .ZN(n18697) );
  OAI211_X1 U21782 ( .C1(n18826), .C2(n18704), .A(n18698), .B(n18697), .ZN(
        P3_U2962) );
  AOI22_X1 U21783 ( .A1(n18828), .A2(n18700), .B1(n18832), .B2(n18699), .ZN(
        n18703) );
  AOI22_X1 U21784 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18701), .B1(
        n18830), .B2(n18725), .ZN(n18702) );
  OAI211_X1 U21785 ( .C1(n18837), .C2(n18704), .A(n18703), .B(n18702), .ZN(
        P3_U2963) );
  INV_X1 U21786 ( .A(n18785), .ZN(n18730) );
  NOR2_X2 U21787 ( .A1(n18730), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18831) );
  INV_X1 U21788 ( .A(n18831), .ZN(n18729) );
  INV_X1 U21789 ( .A(n18704), .ZN(n18774) );
  NOR2_X1 U21790 ( .A1(n18774), .A2(n18831), .ZN(n18756) );
  NOR2_X1 U21791 ( .A1(n18907), .A2(n18756), .ZN(n18724) );
  AOI22_X1 U21792 ( .A1(n18787), .A2(n18725), .B1(n18781), .B2(n18724), .ZN(
        n18711) );
  NAND2_X1 U21793 ( .A1(n18706), .A2(n18705), .ZN(n18707) );
  OAI21_X1 U21794 ( .B1(n18708), .B2(n18707), .A(n18756), .ZN(n18709) );
  OAI211_X1 U21795 ( .C1(n18831), .C2(n19008), .A(n18758), .B(n18709), .ZN(
        n18726) );
  AOI22_X1 U21796 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18726), .B1(
        n18782), .B2(n18748), .ZN(n18710) );
  OAI211_X1 U21797 ( .C1(n18790), .C2(n18729), .A(n18711), .B(n18710), .ZN(
        P3_U2964) );
  AOI22_X1 U21798 ( .A1(n18792), .A2(n18748), .B1(n18791), .B2(n18724), .ZN(
        n18713) );
  AOI22_X1 U21799 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18726), .B1(
        n18793), .B2(n18725), .ZN(n18712) );
  OAI211_X1 U21800 ( .C1(n18796), .C2(n18729), .A(n18713), .B(n18712), .ZN(
        P3_U2965) );
  AOI22_X1 U21801 ( .A1(n18799), .A2(n18725), .B1(n18797), .B2(n18724), .ZN(
        n18715) );
  AOI22_X1 U21802 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18726), .B1(
        n18798), .B2(n18748), .ZN(n18714) );
  OAI211_X1 U21803 ( .C1(n18802), .C2(n18729), .A(n18715), .B(n18714), .ZN(
        P3_U2966) );
  AOI22_X1 U21804 ( .A1(n18804), .A2(n18725), .B1(n18803), .B2(n18724), .ZN(
        n18717) );
  AOI22_X1 U21805 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18726), .B1(
        n18805), .B2(n18748), .ZN(n18716) );
  OAI211_X1 U21806 ( .C1(n18808), .C2(n18729), .A(n18717), .B(n18716), .ZN(
        P3_U2967) );
  AOI22_X1 U21807 ( .A1(n18810), .A2(n18725), .B1(n18809), .B2(n18724), .ZN(
        n18719) );
  AOI22_X1 U21808 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18726), .B1(
        n18811), .B2(n18748), .ZN(n18718) );
  OAI211_X1 U21809 ( .C1(n18814), .C2(n18729), .A(n18719), .B(n18718), .ZN(
        P3_U2968) );
  AOI22_X1 U21810 ( .A1(n18817), .A2(n18748), .B1(n18815), .B2(n18724), .ZN(
        n18721) );
  AOI22_X1 U21811 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18726), .B1(
        n18816), .B2(n18725), .ZN(n18720) );
  OAI211_X1 U21812 ( .C1(n18820), .C2(n18729), .A(n18721), .B(n18720), .ZN(
        P3_U2969) );
  AOI22_X1 U21813 ( .A1(n18822), .A2(n18748), .B1(n18821), .B2(n18724), .ZN(
        n18723) );
  AOI22_X1 U21814 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18726), .B1(
        n18823), .B2(n18725), .ZN(n18722) );
  OAI211_X1 U21815 ( .C1(n18826), .C2(n18729), .A(n18723), .B(n18722), .ZN(
        P3_U2970) );
  AOI22_X1 U21816 ( .A1(n18830), .A2(n18748), .B1(n18828), .B2(n18724), .ZN(
        n18728) );
  AOI22_X1 U21817 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18726), .B1(
        n18832), .B2(n18725), .ZN(n18727) );
  OAI211_X1 U21818 ( .C1(n18837), .C2(n18729), .A(n18728), .B(n18727), .ZN(
        P3_U2971) );
  NOR2_X1 U21819 ( .A1(n18907), .A2(n18730), .ZN(n18749) );
  AOI22_X1 U21820 ( .A1(n18782), .A2(n18774), .B1(n18781), .B2(n18749), .ZN(
        n18735) );
  AOI22_X1 U21821 ( .A1(n18786), .A2(n18733), .B1(n18732), .B2(n18731), .ZN(
        n18750) );
  AOI22_X1 U21822 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18750), .B1(
        n18787), .B2(n18748), .ZN(n18734) );
  OAI211_X1 U21823 ( .C1(n18790), .C2(n18753), .A(n18735), .B(n18734), .ZN(
        P3_U2972) );
  AOI22_X1 U21824 ( .A1(n18791), .A2(n18749), .B1(n18793), .B2(n18748), .ZN(
        n18737) );
  AOI22_X1 U21825 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18750), .B1(
        n18792), .B2(n18774), .ZN(n18736) );
  OAI211_X1 U21826 ( .C1(n18796), .C2(n18753), .A(n18737), .B(n18736), .ZN(
        P3_U2973) );
  AOI22_X1 U21827 ( .A1(n18798), .A2(n18774), .B1(n18797), .B2(n18749), .ZN(
        n18739) );
  AOI22_X1 U21828 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18750), .B1(
        n18799), .B2(n18748), .ZN(n18738) );
  OAI211_X1 U21829 ( .C1(n18802), .C2(n18753), .A(n18739), .B(n18738), .ZN(
        P3_U2974) );
  AOI22_X1 U21830 ( .A1(n18803), .A2(n18749), .B1(n18805), .B2(n18774), .ZN(
        n18741) );
  AOI22_X1 U21831 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18750), .B1(
        n18804), .B2(n18748), .ZN(n18740) );
  OAI211_X1 U21832 ( .C1(n18808), .C2(n18753), .A(n18741), .B(n18740), .ZN(
        P3_U2975) );
  AOI22_X1 U21833 ( .A1(n18810), .A2(n18748), .B1(n18809), .B2(n18749), .ZN(
        n18743) );
  AOI22_X1 U21834 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18750), .B1(
        n18811), .B2(n18774), .ZN(n18742) );
  OAI211_X1 U21835 ( .C1(n18814), .C2(n18753), .A(n18743), .B(n18742), .ZN(
        P3_U2976) );
  AOI22_X1 U21836 ( .A1(n18816), .A2(n18748), .B1(n18815), .B2(n18749), .ZN(
        n18745) );
  AOI22_X1 U21837 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18750), .B1(
        n18817), .B2(n18774), .ZN(n18744) );
  OAI211_X1 U21838 ( .C1(n18820), .C2(n18753), .A(n18745), .B(n18744), .ZN(
        P3_U2977) );
  AOI22_X1 U21839 ( .A1(n18823), .A2(n18748), .B1(n18821), .B2(n18749), .ZN(
        n18747) );
  AOI22_X1 U21840 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18750), .B1(
        n18822), .B2(n18774), .ZN(n18746) );
  OAI211_X1 U21841 ( .C1(n18826), .C2(n18753), .A(n18747), .B(n18746), .ZN(
        P3_U2978) );
  AOI22_X1 U21842 ( .A1(n18828), .A2(n18749), .B1(n18832), .B2(n18748), .ZN(
        n18752) );
  AOI22_X1 U21843 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18750), .B1(
        n18830), .B2(n18774), .ZN(n18751) );
  OAI211_X1 U21844 ( .C1(n18837), .C2(n18753), .A(n18752), .B(n18751), .ZN(
        P3_U2979) );
  NOR2_X1 U21845 ( .A1(n18907), .A2(n18754), .ZN(n18775) );
  AOI22_X1 U21846 ( .A1(n18787), .A2(n18774), .B1(n18781), .B2(n18775), .ZN(
        n18761) );
  OAI21_X1 U21847 ( .B1(n18756), .B2(n18755), .A(n18754), .ZN(n18757) );
  OAI211_X1 U21848 ( .C1(n18759), .C2(n19008), .A(n18758), .B(n18757), .ZN(
        n18776) );
  AOI22_X1 U21849 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18776), .B1(
        n18782), .B2(n18831), .ZN(n18760) );
  OAI211_X1 U21850 ( .C1(n18790), .C2(n18779), .A(n18761), .B(n18760), .ZN(
        P3_U2980) );
  AOI22_X1 U21851 ( .A1(n18791), .A2(n18775), .B1(n18793), .B2(n18774), .ZN(
        n18763) );
  AOI22_X1 U21852 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18776), .B1(
        n18792), .B2(n18831), .ZN(n18762) );
  OAI211_X1 U21853 ( .C1(n18796), .C2(n18779), .A(n18763), .B(n18762), .ZN(
        P3_U2981) );
  AOI22_X1 U21854 ( .A1(n18799), .A2(n18774), .B1(n18797), .B2(n18775), .ZN(
        n18765) );
  AOI22_X1 U21855 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18776), .B1(
        n18798), .B2(n18831), .ZN(n18764) );
  OAI211_X1 U21856 ( .C1(n18802), .C2(n18779), .A(n18765), .B(n18764), .ZN(
        P3_U2982) );
  AOI22_X1 U21857 ( .A1(n18804), .A2(n18774), .B1(n18803), .B2(n18775), .ZN(
        n18767) );
  AOI22_X1 U21858 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18776), .B1(
        n18805), .B2(n18831), .ZN(n18766) );
  OAI211_X1 U21859 ( .C1(n18808), .C2(n18779), .A(n18767), .B(n18766), .ZN(
        P3_U2983) );
  AOI22_X1 U21860 ( .A1(n18811), .A2(n18831), .B1(n18809), .B2(n18775), .ZN(
        n18769) );
  AOI22_X1 U21861 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18776), .B1(
        n18810), .B2(n18774), .ZN(n18768) );
  OAI211_X1 U21862 ( .C1(n18814), .C2(n18779), .A(n18769), .B(n18768), .ZN(
        P3_U2984) );
  AOI22_X1 U21863 ( .A1(n18816), .A2(n18774), .B1(n18815), .B2(n18775), .ZN(
        n18771) );
  AOI22_X1 U21864 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18776), .B1(
        n18817), .B2(n18831), .ZN(n18770) );
  OAI211_X1 U21865 ( .C1(n18820), .C2(n18779), .A(n18771), .B(n18770), .ZN(
        P3_U2985) );
  AOI22_X1 U21866 ( .A1(n18822), .A2(n18831), .B1(n18821), .B2(n18775), .ZN(
        n18773) );
  AOI22_X1 U21867 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18776), .B1(
        n18823), .B2(n18774), .ZN(n18772) );
  OAI211_X1 U21868 ( .C1(n18826), .C2(n18779), .A(n18773), .B(n18772), .ZN(
        P3_U2986) );
  AOI22_X1 U21869 ( .A1(n18828), .A2(n18775), .B1(n18832), .B2(n18774), .ZN(
        n18778) );
  AOI22_X1 U21870 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18776), .B1(
        n18830), .B2(n18831), .ZN(n18777) );
  OAI211_X1 U21871 ( .C1(n18837), .C2(n18779), .A(n18778), .B(n18777), .ZN(
        P3_U2987) );
  AND2_X1 U21872 ( .A1(n18780), .A2(n18784), .ZN(n18827) );
  AOI22_X1 U21873 ( .A1(n18782), .A2(n18829), .B1(n18781), .B2(n18827), .ZN(
        n18789) );
  AOI22_X1 U21874 ( .A1(n18786), .A2(n18785), .B1(n18784), .B2(n18783), .ZN(
        n18833) );
  AOI22_X1 U21875 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18833), .B1(
        n18787), .B2(n18831), .ZN(n18788) );
  OAI211_X1 U21876 ( .C1(n18790), .C2(n18836), .A(n18789), .B(n18788), .ZN(
        P3_U2988) );
  AOI22_X1 U21877 ( .A1(n18792), .A2(n18829), .B1(n18791), .B2(n18827), .ZN(
        n18795) );
  AOI22_X1 U21878 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18833), .B1(
        n18793), .B2(n18831), .ZN(n18794) );
  OAI211_X1 U21879 ( .C1(n18796), .C2(n18836), .A(n18795), .B(n18794), .ZN(
        P3_U2989) );
  AOI22_X1 U21880 ( .A1(n18798), .A2(n18829), .B1(n18797), .B2(n18827), .ZN(
        n18801) );
  AOI22_X1 U21881 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18833), .B1(
        n18799), .B2(n18831), .ZN(n18800) );
  OAI211_X1 U21882 ( .C1(n18802), .C2(n18836), .A(n18801), .B(n18800), .ZN(
        P3_U2990) );
  AOI22_X1 U21883 ( .A1(n18804), .A2(n18831), .B1(n18803), .B2(n18827), .ZN(
        n18807) );
  AOI22_X1 U21884 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18833), .B1(
        n18805), .B2(n18829), .ZN(n18806) );
  OAI211_X1 U21885 ( .C1(n18808), .C2(n18836), .A(n18807), .B(n18806), .ZN(
        P3_U2991) );
  AOI22_X1 U21886 ( .A1(n18810), .A2(n18831), .B1(n18809), .B2(n18827), .ZN(
        n18813) );
  AOI22_X1 U21887 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18833), .B1(
        n18811), .B2(n18829), .ZN(n18812) );
  OAI211_X1 U21888 ( .C1(n18814), .C2(n18836), .A(n18813), .B(n18812), .ZN(
        P3_U2992) );
  AOI22_X1 U21889 ( .A1(n18816), .A2(n18831), .B1(n18815), .B2(n18827), .ZN(
        n18819) );
  AOI22_X1 U21890 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18833), .B1(
        n18817), .B2(n18829), .ZN(n18818) );
  OAI211_X1 U21891 ( .C1(n18820), .C2(n18836), .A(n18819), .B(n18818), .ZN(
        P3_U2993) );
  AOI22_X1 U21892 ( .A1(n18822), .A2(n18829), .B1(n18821), .B2(n18827), .ZN(
        n18825) );
  AOI22_X1 U21893 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18833), .B1(
        n18823), .B2(n18831), .ZN(n18824) );
  OAI211_X1 U21894 ( .C1(n18826), .C2(n18836), .A(n18825), .B(n18824), .ZN(
        P3_U2994) );
  AOI22_X1 U21895 ( .A1(n18830), .A2(n18829), .B1(n18828), .B2(n18827), .ZN(
        n18835) );
  AOI22_X1 U21896 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18833), .B1(
        n18832), .B2(n18831), .ZN(n18834) );
  OAI211_X1 U21897 ( .C1(n18837), .C2(n18836), .A(n18835), .B(n18834), .ZN(
        P3_U2995) );
  AOI22_X1 U21898 ( .A1(n18841), .A2(n18840), .B1(n18839), .B2(n18838), .ZN(
        n18842) );
  OAI221_X1 U21899 ( .B1(n18845), .B2(n18844), .C1(n18845), .C2(n18843), .A(
        n18842), .ZN(n19049) );
  OAI21_X1 U21900 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18846), .ZN(n18847) );
  OAI211_X1 U21901 ( .C1(n18849), .C2(n18881), .A(n18848), .B(n18847), .ZN(
        n18893) );
  NAND2_X1 U21902 ( .A1(n18859), .A2(n17045), .ZN(n18860) );
  AOI22_X1 U21903 ( .A1(n18850), .A2(n18860), .B1(n18880), .B2(n18852), .ZN(
        n19010) );
  NOR2_X1 U21904 ( .A1(n18882), .A2(n19010), .ZN(n18856) );
  AOI21_X1 U21905 ( .B1(n18869), .B2(n18851), .A(n18868), .ZN(n18853) );
  OAI21_X1 U21906 ( .B1(n18854), .B2(n18853), .A(n18852), .ZN(n19013) );
  OR2_X1 U21907 ( .A1(n19014), .A2(n19013), .ZN(n18855) );
  OAI22_X1 U21908 ( .A1(n18856), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n18882), .B2(n18855), .ZN(n18891) );
  NOR2_X1 U21909 ( .A1(n18858), .A2(n18857), .ZN(n18863) );
  AOI22_X1 U21910 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18859), .B1(
        n18863), .B2(n17045), .ZN(n19033) );
  NOR2_X1 U21911 ( .A1(n19033), .A2(n18864), .ZN(n18867) );
  INV_X1 U21912 ( .A(n18860), .ZN(n18861) );
  OAI22_X1 U21913 ( .A1(n18863), .A2(n18862), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18861), .ZN(n19029) );
  OAI221_X1 U21914 ( .B1(n19029), .B2(n19033), .C1(n19029), .C2(n18864), .A(
        n18881), .ZN(n18865) );
  AOI22_X1 U21915 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18867), .B1(
        n18866), .B2(n18865), .ZN(n18885) );
  AOI21_X1 U21916 ( .B1(n19031), .B2(n18872), .A(n18868), .ZN(n18877) );
  NAND2_X1 U21917 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n17060), .ZN(
        n18876) );
  OAI211_X1 U21918 ( .C1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n18870), .B(n18869), .ZN(
        n18875) );
  NOR2_X1 U21919 ( .A1(n18871), .A2(n17045), .ZN(n18873) );
  OAI211_X1 U21920 ( .C1(n18873), .C2(n18872), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n19025), .ZN(n18874) );
  OAI211_X1 U21921 ( .C1(n18877), .C2(n18876), .A(n18875), .B(n18874), .ZN(
        n18878) );
  AOI21_X1 U21922 ( .B1(n18880), .B2(n18879), .A(n18878), .ZN(n19017) );
  AOI22_X1 U21923 ( .A1(n18882), .A2(n19025), .B1(n19017), .B2(n18881), .ZN(
        n18886) );
  AND2_X1 U21924 ( .A1(n18885), .A2(n18886), .ZN(n18883) );
  OAI221_X1 U21925 ( .B1(n18885), .B2(n18886), .C1(n18884), .C2(n18883), .A(
        n18888), .ZN(n18890) );
  AOI21_X1 U21926 ( .B1(n18888), .B2(n18887), .A(n18886), .ZN(n18889) );
  AOI222_X1 U21927 ( .A1(n18891), .A2(n18890), .B1(n18891), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18890), .C2(n18889), .ZN(
        n18892) );
  NOR4_X1 U21928 ( .A1(n18894), .A2(n19049), .A3(n18893), .A4(n18892), .ZN(
        n18905) );
  AOI22_X1 U21929 ( .A1(n19032), .A2(n19062), .B1(n19057), .B2(n19051), .ZN(
        n18895) );
  INV_X1 U21930 ( .A(n18895), .ZN(n18900) );
  OAI211_X1 U21931 ( .C1(n18897), .C2(n18896), .A(n19054), .B(n18905), .ZN(
        n19007) );
  NAND2_X1 U21932 ( .A1(n19057), .A2(n19056), .ZN(n18906) );
  NAND2_X1 U21933 ( .A1(n19007), .A2(n18906), .ZN(n18908) );
  NOR2_X1 U21934 ( .A1(n18898), .A2(n18908), .ZN(n18899) );
  MUX2_X1 U21935 ( .A(n18900), .B(n18899), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18903) );
  INV_X1 U21936 ( .A(n18909), .ZN(n18901) );
  NAND2_X1 U21937 ( .A1(n18901), .A2(n18907), .ZN(n18902) );
  OAI211_X1 U21938 ( .C1(n18905), .C2(n18904), .A(n18903), .B(n18902), .ZN(
        P3_U2996) );
  NAND2_X1 U21939 ( .A1(n19057), .A2(n19051), .ZN(n18912) );
  NOR3_X1 U21940 ( .A1(n19018), .A2(n19059), .A3(n18906), .ZN(n18915) );
  INV_X1 U21941 ( .A(n18915), .ZN(n18911) );
  NAND4_X1 U21942 ( .A1(n18913), .A2(n18912), .A3(n18911), .A4(n18910), .ZN(
        P3_U2997) );
  OAI21_X1 U21943 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18914), .ZN(n18916) );
  AOI21_X1 U21944 ( .B1(n18917), .B2(n18916), .A(n18915), .ZN(P3_U2998) );
  AND2_X1 U21945 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18918), .ZN(
        P3_U2999) );
  AND2_X1 U21946 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18918), .ZN(
        P3_U3000) );
  AND2_X1 U21947 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18918), .ZN(
        P3_U3001) );
  AND2_X1 U21948 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18918), .ZN(
        P3_U3002) );
  AND2_X1 U21949 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18918), .ZN(
        P3_U3003) );
  AND2_X1 U21950 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18918), .ZN(
        P3_U3004) );
  AND2_X1 U21951 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18918), .ZN(
        P3_U3005) );
  AND2_X1 U21952 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18918), .ZN(
        P3_U3006) );
  AND2_X1 U21953 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18918), .ZN(
        P3_U3007) );
  AND2_X1 U21954 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18918), .ZN(
        P3_U3008) );
  AND2_X1 U21955 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18918), .ZN(
        P3_U3009) );
  AND2_X1 U21956 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18918), .ZN(
        P3_U3010) );
  AND2_X1 U21957 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18918), .ZN(
        P3_U3011) );
  AND2_X1 U21958 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18918), .ZN(
        P3_U3012) );
  AND2_X1 U21959 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18918), .ZN(
        P3_U3013) );
  AND2_X1 U21960 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18918), .ZN(
        P3_U3014) );
  AND2_X1 U21961 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18918), .ZN(
        P3_U3015) );
  AND2_X1 U21962 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18918), .ZN(
        P3_U3016) );
  AND2_X1 U21963 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18918), .ZN(
        P3_U3017) );
  AND2_X1 U21964 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18918), .ZN(
        P3_U3018) );
  AND2_X1 U21965 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18918), .ZN(
        P3_U3019) );
  AND2_X1 U21966 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18918), .ZN(
        P3_U3020) );
  AND2_X1 U21967 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18918), .ZN(P3_U3021) );
  AND2_X1 U21968 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18918), .ZN(P3_U3022) );
  AND2_X1 U21969 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18918), .ZN(P3_U3023) );
  AND2_X1 U21970 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18918), .ZN(P3_U3024) );
  AND2_X1 U21971 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18918), .ZN(P3_U3025) );
  AND2_X1 U21972 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18918), .ZN(P3_U3026) );
  AND2_X1 U21973 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18918), .ZN(P3_U3027) );
  AND2_X1 U21974 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18918), .ZN(P3_U3028) );
  OAI21_X1 U21975 ( .B1(n18919), .B2(n21115), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18920) );
  AOI22_X1 U21976 ( .A1(n18931), .A2(n18933), .B1(n19066), .B2(n18920), .ZN(
        n18921) );
  INV_X1 U21977 ( .A(NA), .ZN(n20898) );
  OR3_X1 U21978 ( .A1(n20898), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n18926) );
  OAI211_X1 U21979 ( .C1(n18922), .C2(n19050), .A(n18921), .B(n18926), .ZN(
        P3_U3029) );
  NOR2_X1 U21980 ( .A1(n18933), .A2(n21115), .ZN(n18929) );
  INV_X1 U21981 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19064) );
  OAI22_X1 U21982 ( .A1(n18929), .A2(n19064), .B1(n21115), .B2(n18922), .ZN(
        n18923) );
  AOI22_X1 U21983 ( .A1(n19057), .A2(P3_STATE_REG_1__SCAN_IN), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n18923), .ZN(n18925) );
  NAND2_X1 U21984 ( .A1(n18925), .A2(n18924), .ZN(P3_U3030) );
  AOI22_X1 U21985 ( .A1(n19057), .A2(P3_STATE_REG_1__SCAN_IN), .B1(n18931), 
        .B2(n18926), .ZN(n18932) );
  NAND2_X1 U21986 ( .A1(n19057), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18927) );
  OAI22_X1 U21987 ( .A1(NA), .A2(n18927), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18928) );
  OAI22_X1 U21988 ( .A1(n18929), .A2(n18928), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18930) );
  OAI22_X1 U21989 ( .A1(n18932), .A2(n18933), .B1(n18931), .B2(n18930), .ZN(
        P3_U3031) );
  OAI222_X1 U21990 ( .A1(n19039), .A2(n18990), .B1(n18934), .B2(n19000), .C1(
        n18935), .C2(n18985), .ZN(P3_U3032) );
  INV_X1 U21991 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18937) );
  OAI222_X1 U21992 ( .A1(n18985), .A2(n18937), .B1(n18936), .B2(n19000), .C1(
        n18935), .C2(n18990), .ZN(P3_U3033) );
  OAI222_X1 U21993 ( .A1(n18985), .A2(n18939), .B1(n18938), .B2(n19000), .C1(
        n18937), .C2(n18990), .ZN(P3_U3034) );
  OAI222_X1 U21994 ( .A1(n18985), .A2(n18941), .B1(n18940), .B2(n19000), .C1(
        n18939), .C2(n18990), .ZN(P3_U3035) );
  INV_X1 U21995 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18943) );
  OAI222_X1 U21996 ( .A1(n18985), .A2(n18943), .B1(n18942), .B2(n19000), .C1(
        n18941), .C2(n18990), .ZN(P3_U3036) );
  OAI222_X1 U21997 ( .A1(n18985), .A2(n18945), .B1(n18944), .B2(n19000), .C1(
        n18943), .C2(n18990), .ZN(P3_U3037) );
  OAI222_X1 U21998 ( .A1(n18985), .A2(n18948), .B1(n18946), .B2(n19000), .C1(
        n18945), .C2(n18990), .ZN(P3_U3038) );
  OAI222_X1 U21999 ( .A1(n18948), .A2(n18990), .B1(n18947), .B2(n19000), .C1(
        n18949), .C2(n18985), .ZN(P3_U3039) );
  OAI222_X1 U22000 ( .A1(n18985), .A2(n18951), .B1(n18950), .B2(n19000), .C1(
        n18949), .C2(n18990), .ZN(P3_U3040) );
  OAI222_X1 U22001 ( .A1(n18985), .A2(n18953), .B1(n18952), .B2(n19000), .C1(
        n18951), .C2(n18990), .ZN(P3_U3041) );
  OAI222_X1 U22002 ( .A1(n18985), .A2(n18955), .B1(n18954), .B2(n19000), .C1(
        n18953), .C2(n18990), .ZN(P3_U3042) );
  INV_X1 U22003 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18957) );
  OAI222_X1 U22004 ( .A1(n18985), .A2(n18957), .B1(n18956), .B2(n19000), .C1(
        n18955), .C2(n18990), .ZN(P3_U3043) );
  OAI222_X1 U22005 ( .A1(n18985), .A2(n18960), .B1(n18958), .B2(n19000), .C1(
        n18957), .C2(n18996), .ZN(P3_U3044) );
  OAI222_X1 U22006 ( .A1(n18960), .A2(n18990), .B1(n18959), .B2(n19000), .C1(
        n18961), .C2(n18985), .ZN(P3_U3045) );
  OAI222_X1 U22007 ( .A1(n18985), .A2(n18963), .B1(n18962), .B2(n19000), .C1(
        n18961), .C2(n18996), .ZN(P3_U3046) );
  OAI222_X1 U22008 ( .A1(n18985), .A2(n18965), .B1(n18964), .B2(n19000), .C1(
        n18963), .C2(n18996), .ZN(P3_U3047) );
  OAI222_X1 U22009 ( .A1(n18985), .A2(n18967), .B1(n18966), .B2(n19000), .C1(
        n18965), .C2(n18996), .ZN(P3_U3048) );
  OAI222_X1 U22010 ( .A1(n18985), .A2(n18970), .B1(n18968), .B2(n19000), .C1(
        n18967), .C2(n18996), .ZN(P3_U3049) );
  INV_X1 U22011 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18971) );
  OAI222_X1 U22012 ( .A1(n18970), .A2(n18990), .B1(n18969), .B2(n19000), .C1(
        n18971), .C2(n18985), .ZN(P3_U3050) );
  OAI222_X1 U22013 ( .A1(n18985), .A2(n18974), .B1(n18972), .B2(n19000), .C1(
        n18971), .C2(n18996), .ZN(P3_U3051) );
  OAI222_X1 U22014 ( .A1(n18974), .A2(n18990), .B1(n18973), .B2(n19000), .C1(
        n18975), .C2(n18985), .ZN(P3_U3052) );
  OAI222_X1 U22015 ( .A1(n18985), .A2(n18978), .B1(n18976), .B2(n19000), .C1(
        n18975), .C2(n18996), .ZN(P3_U3053) );
  OAI222_X1 U22016 ( .A1(n18978), .A2(n18990), .B1(n18977), .B2(n19000), .C1(
        n18979), .C2(n18985), .ZN(P3_U3054) );
  OAI222_X1 U22017 ( .A1(n18985), .A2(n18981), .B1(n18980), .B2(n19000), .C1(
        n18979), .C2(n18996), .ZN(P3_U3055) );
  OAI222_X1 U22018 ( .A1(n18985), .A2(n18983), .B1(n18982), .B2(n19000), .C1(
        n18981), .C2(n18996), .ZN(P3_U3056) );
  OAI222_X1 U22019 ( .A1(n18985), .A2(n18986), .B1(n18984), .B2(n19000), .C1(
        n18983), .C2(n18990), .ZN(P3_U3057) );
  OAI222_X1 U22020 ( .A1(n18985), .A2(n18989), .B1(n18987), .B2(n19000), .C1(
        n18986), .C2(n18990), .ZN(P3_U3058) );
  OAI222_X1 U22021 ( .A1(n18989), .A2(n18990), .B1(n18988), .B2(n19000), .C1(
        n18991), .C2(n18985), .ZN(P3_U3059) );
  OAI222_X1 U22022 ( .A1(n18985), .A2(n18995), .B1(n18992), .B2(n19000), .C1(
        n18991), .C2(n18990), .ZN(P3_U3060) );
  INV_X1 U22023 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18994) );
  OAI222_X1 U22024 ( .A1(n18996), .A2(n18995), .B1(n18994), .B2(n19000), .C1(
        n18993), .C2(n18985), .ZN(P3_U3061) );
  OAI22_X1 U22025 ( .A1(n19066), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n19000), .ZN(n18997) );
  INV_X1 U22026 ( .A(n18997), .ZN(P3_U3274) );
  OAI22_X1 U22027 ( .A1(n19066), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n19000), .ZN(n18998) );
  INV_X1 U22028 ( .A(n18998), .ZN(P3_U3275) );
  OAI22_X1 U22029 ( .A1(n19066), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n19000), .ZN(n18999) );
  INV_X1 U22030 ( .A(n18999), .ZN(P3_U3276) );
  OAI22_X1 U22031 ( .A1(n19066), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n19000), .ZN(n19001) );
  INV_X1 U22032 ( .A(n19001), .ZN(P3_U3277) );
  OAI21_X1 U22033 ( .B1(n19005), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n19003), 
        .ZN(n19002) );
  INV_X1 U22034 ( .A(n19002), .ZN(P3_U3280) );
  OAI21_X1 U22035 ( .B1(n19005), .B2(n19004), .A(n19003), .ZN(P3_U3281) );
  OAI221_X1 U22036 ( .B1(n19008), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19008), 
        .C2(n19007), .A(n19006), .ZN(P3_U3282) );
  NOR3_X1 U22037 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19010), .A3(
        n19009), .ZN(n19011) );
  AOI21_X1 U22038 ( .B1(n19012), .B2(n19032), .A(n19011), .ZN(n19016) );
  AOI21_X1 U22039 ( .B1(n19034), .B2(n19013), .A(n19038), .ZN(n19015) );
  OAI22_X1 U22040 ( .A1(n19038), .A2(n19016), .B1(n19015), .B2(n19014), .ZN(
        P3_U3285) );
  INV_X1 U22041 ( .A(n19017), .ZN(n19023) );
  NOR2_X1 U22042 ( .A1(n19018), .A2(n19035), .ZN(n19026) );
  OAI22_X1 U22043 ( .A1(n19020), .A2(n19019), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19027) );
  INV_X1 U22044 ( .A(n19027), .ZN(n19022) );
  AOI222_X1 U22045 ( .A1(n19023), .A2(n19034), .B1(n19026), .B2(n19022), .C1(
        n19032), .C2(n19021), .ZN(n19024) );
  AOI22_X1 U22046 ( .A1(n19038), .A2(n19025), .B1(n19024), .B2(n19036), .ZN(
        P3_U3288) );
  AOI222_X1 U22047 ( .A1(n19029), .A2(n19034), .B1(n19032), .B2(n19028), .C1(
        n19027), .C2(n19026), .ZN(n19030) );
  AOI22_X1 U22048 ( .A1(n19038), .A2(n19031), .B1(n19030), .B2(n19036), .ZN(
        P3_U3289) );
  AOI222_X1 U22049 ( .A1(n19035), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n19034), 
        .B2(n19033), .C1(n17045), .C2(n19032), .ZN(n19037) );
  AOI22_X1 U22050 ( .A1(n19038), .A2(n17045), .B1(n19037), .B2(n19036), .ZN(
        P3_U3290) );
  AOI21_X1 U22051 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19040) );
  AOI22_X1 U22052 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n19040), .B2(n19039), .ZN(n19043) );
  INV_X1 U22053 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19042) );
  AOI22_X1 U22054 ( .A1(n19046), .A2(n19043), .B1(n19042), .B2(n19041), .ZN(
        P3_U3292) );
  INV_X1 U22055 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19045) );
  OAI21_X1 U22056 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n19046), .ZN(n19044) );
  OAI21_X1 U22057 ( .B1(n19046), .B2(n19045), .A(n19044), .ZN(P3_U3293) );
  INV_X1 U22058 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19047) );
  AOI22_X1 U22059 ( .A1(n19000), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19047), 
        .B2(n19066), .ZN(P3_U3294) );
  MUX2_X1 U22060 ( .A(P3_MORE_REG_SCAN_IN), .B(n19049), .S(n19048), .Z(
        P3_U3295) );
  AOI21_X1 U22061 ( .B1(n19051), .B2(n19050), .A(n19073), .ZN(n19052) );
  OAI21_X1 U22062 ( .B1(n19054), .B2(n19053), .A(n19052), .ZN(n19065) );
  OAI21_X1 U22063 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n9969), .A(n19055), 
        .ZN(n19058) );
  AOI211_X1 U22064 ( .C1(n19068), .C2(n19058), .A(n19057), .B(n19056), .ZN(
        n19060) );
  NOR2_X1 U22065 ( .A1(n19060), .A2(n19059), .ZN(n19061) );
  OAI21_X1 U22066 ( .B1(n19062), .B2(n19061), .A(n19065), .ZN(n19063) );
  OAI21_X1 U22067 ( .B1(n19065), .B2(n19064), .A(n19063), .ZN(P3_U3296) );
  MUX2_X1 U22068 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .B(P3_M_IO_N_REG_SCAN_IN), 
        .S(n19066), .Z(P3_U3297) );
  OAI21_X1 U22069 ( .B1(n19070), .B2(P3_READREQUEST_REG_SCAN_IN), .A(n19069), 
        .ZN(n19067) );
  OAI21_X1 U22070 ( .B1(n19069), .B2(n19068), .A(n19067), .ZN(P3_U3298) );
  NOR2_X1 U22071 ( .A1(n19070), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19072)
         );
  OAI21_X1 U22072 ( .B1(n19073), .B2(n19072), .A(n19071), .ZN(P3_U3299) );
  INV_X1 U22073 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19076) );
  NAND2_X1 U22074 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20011), .ZN(n20000) );
  NAND2_X1 U22075 ( .A1(n19076), .A2(n19074), .ZN(n19997) );
  OAI21_X1 U22076 ( .B1(n19076), .B2(n20000), .A(n19997), .ZN(n20068) );
  AOI21_X1 U22077 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n20068), .ZN(n19075) );
  INV_X1 U22078 ( .A(n19075), .ZN(P2_U2815) );
  NAND2_X1 U22079 ( .A1(n19076), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20109) );
  INV_X2 U22080 ( .A(n20109), .ZN(n20108) );
  AOI21_X1 U22081 ( .B1(n19076), .B2(n20011), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19077) );
  AOI22_X1 U22082 ( .A1(n20108), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n19077), 
        .B2(n20109), .ZN(P2_U2817) );
  OAI21_X1 U22083 ( .B1(n20004), .B2(BS16), .A(n20068), .ZN(n20066) );
  OAI21_X1 U22084 ( .B1(n20068), .B2(n19541), .A(n20066), .ZN(P2_U2818) );
  NOR4_X1 U22085 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19081) );
  NOR4_X1 U22086 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19080) );
  NOR4_X1 U22087 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19079) );
  NOR4_X1 U22088 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19078) );
  NAND4_X1 U22089 ( .A1(n19081), .A2(n19080), .A3(n19079), .A4(n19078), .ZN(
        n19087) );
  NOR4_X1 U22090 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19085) );
  AOI211_X1 U22091 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19084) );
  NOR4_X1 U22092 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19083) );
  NOR4_X1 U22093 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19082) );
  NAND4_X1 U22094 ( .A1(n19085), .A2(n19084), .A3(n19083), .A4(n19082), .ZN(
        n19086) );
  NOR2_X1 U22095 ( .A1(n19087), .A2(n19086), .ZN(n19098) );
  INV_X1 U22096 ( .A(n19098), .ZN(n19096) );
  NOR2_X1 U22097 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19096), .ZN(n19090) );
  INV_X1 U22098 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19088) );
  AOI22_X1 U22099 ( .A1(n19090), .A2(n19091), .B1(n19096), .B2(n19088), .ZN(
        P2_U2820) );
  OR3_X1 U22100 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19095) );
  INV_X1 U22101 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19089) );
  AOI22_X1 U22102 ( .A1(n19090), .A2(n19095), .B1(n19096), .B2(n19089), .ZN(
        P2_U2821) );
  INV_X1 U22103 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20067) );
  NAND2_X1 U22104 ( .A1(n19090), .A2(n20067), .ZN(n19094) );
  OAI21_X1 U22105 ( .B1(n19091), .B2(n20013), .A(n19098), .ZN(n19092) );
  OAI21_X1 U22106 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19098), .A(n19092), 
        .ZN(n19093) );
  OAI221_X1 U22107 ( .B1(n19094), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19094), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19093), .ZN(P2_U2822) );
  INV_X1 U22108 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19097) );
  OAI221_X1 U22109 ( .B1(n19098), .B2(n19097), .C1(n19096), .C2(n19095), .A(
        n19094), .ZN(P2_U2823) );
  NAND2_X1 U22110 ( .A1(n13426), .A2(n19099), .ZN(n19101) );
  OAI211_X1 U22111 ( .C1(n9749), .C2(n19101), .A(n19100), .B(n19227), .ZN(
        n19111) );
  OAI22_X1 U22112 ( .A1(n19102), .A2(n19216), .B1(n20041), .B2(n19215), .ZN(
        n19103) );
  INV_X1 U22113 ( .A(n19103), .ZN(n19110) );
  AOI22_X1 U22114 ( .A1(n19183), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n19221), .ZN(n19109) );
  INV_X1 U22115 ( .A(n19104), .ZN(n19105) );
  OAI22_X1 U22116 ( .A1(n19106), .A2(n19129), .B1(n19105), .B2(n19231), .ZN(
        n19107) );
  INV_X1 U22117 ( .A(n19107), .ZN(n19108) );
  NAND4_X1 U22118 ( .A1(n19111), .A2(n19110), .A3(n19109), .A4(n19108), .ZN(
        P2_U2834) );
  INV_X1 U22119 ( .A(n19112), .ZN(n19133) );
  OAI21_X1 U22120 ( .B1(n19133), .B2(n19113), .A(n19227), .ZN(n19114) );
  AOI21_X1 U22121 ( .B1(n19151), .B2(n19114), .A(n9749), .ZN(n19122) );
  AOI22_X1 U22122 ( .A1(n19221), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n19199), .B2(P2_REIP_REG_20__SCAN_IN), .ZN(n19116) );
  NAND2_X1 U22123 ( .A1(n19183), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n19115) );
  OAI211_X1 U22124 ( .C1(n19117), .C2(n19129), .A(n19116), .B(n19115), .ZN(
        n19118) );
  AOI21_X1 U22125 ( .B1(n19119), .B2(n19189), .A(n19118), .ZN(n19120) );
  INV_X1 U22126 ( .A(n19120), .ZN(n19121) );
  AOI211_X1 U22127 ( .C1(n19209), .C2(n19123), .A(n19122), .B(n19121), .ZN(
        n19124) );
  INV_X1 U22128 ( .A(n19124), .ZN(P2_U2835) );
  INV_X1 U22129 ( .A(n19125), .ZN(n19137) );
  NAND2_X1 U22130 ( .A1(n19221), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n19126) );
  OAI211_X1 U22131 ( .C1(n20038), .C2(n19215), .A(n19126), .B(n19214), .ZN(
        n19127) );
  AOI21_X1 U22132 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n19183), .A(n19127), .ZN(
        n19128) );
  OAI21_X1 U22133 ( .B1(n19130), .B2(n19129), .A(n19128), .ZN(n19136) );
  OAI21_X1 U22134 ( .B1(n19132), .B2(n19131), .A(n19227), .ZN(n19134) );
  AOI21_X1 U22135 ( .B1(n19151), .B2(n19134), .A(n19133), .ZN(n19135) );
  AOI211_X1 U22136 ( .C1(n19189), .C2(n19137), .A(n19136), .B(n19135), .ZN(
        n19138) );
  OAI21_X1 U22137 ( .B1(n19139), .B2(n19231), .A(n19138), .ZN(P2_U2836) );
  AOI21_X1 U22138 ( .B1(n19199), .B2(P2_REIP_REG_17__SCAN_IN), .A(n19198), 
        .ZN(n19140) );
  OAI21_X1 U22139 ( .B1(n19186), .B2(n19141), .A(n19140), .ZN(n19142) );
  AOI21_X1 U22140 ( .B1(n19143), .B2(n19226), .A(n19142), .ZN(n19144) );
  OAI21_X1 U22141 ( .B1(n19218), .B2(n19145), .A(n19144), .ZN(n19153) );
  OAI21_X1 U22142 ( .B1(n19147), .B2(n19146), .A(n19227), .ZN(n19150) );
  INV_X1 U22143 ( .A(n19148), .ZN(n19149) );
  AOI21_X1 U22144 ( .B1(n19151), .B2(n19150), .A(n19149), .ZN(n19152) );
  AOI211_X1 U22145 ( .C1(n19189), .C2(n19154), .A(n19153), .B(n19152), .ZN(
        n19155) );
  OAI21_X1 U22146 ( .B1(n19156), .B2(n19231), .A(n19155), .ZN(P2_U2838) );
  OAI21_X1 U22147 ( .B1(n19215), .B2(n16401), .A(n19214), .ZN(n19157) );
  AOI21_X1 U22148 ( .B1(n19221), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n19157), .ZN(n19158) );
  OAI21_X1 U22149 ( .B1(n19218), .B2(n19159), .A(n19158), .ZN(n19163) );
  AOI21_X1 U22150 ( .B1(n19166), .B2(n19161), .A(n19160), .ZN(n19162) );
  AOI211_X1 U22151 ( .C1(n19189), .C2(n19164), .A(n19163), .B(n19162), .ZN(
        n19169) );
  AOI22_X1 U22152 ( .A1(n19167), .A2(n19166), .B1(n19226), .B2(n19165), .ZN(
        n19168) );
  OAI211_X1 U22153 ( .C1(n19231), .C2(n19279), .A(n19169), .B(n19168), .ZN(
        P2_U2842) );
  OAI21_X1 U22154 ( .B1(n19215), .B2(n19170), .A(n19214), .ZN(n19171) );
  AOI21_X1 U22155 ( .B1(n19221), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n19171), .ZN(n19173) );
  NAND2_X1 U22156 ( .A1(n19183), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n19172) );
  OAI211_X1 U22157 ( .C1(n19174), .C2(n19216), .A(n19173), .B(n19172), .ZN(
        n19175) );
  INV_X1 U22158 ( .A(n19175), .ZN(n19182) );
  NOR2_X1 U22159 ( .A1(n10085), .A2(n19176), .ZN(n19178) );
  XNOR2_X1 U22160 ( .A(n19178), .B(n19177), .ZN(n19180) );
  INV_X1 U22161 ( .A(n19245), .ZN(n19179) );
  AOI22_X1 U22162 ( .A1(n19180), .A2(n19227), .B1(n19226), .B2(n19179), .ZN(
        n19181) );
  OAI211_X1 U22163 ( .C1(n19231), .C2(n19281), .A(n19182), .B(n19181), .ZN(
        P2_U2843) );
  NAND2_X1 U22164 ( .A1(n19183), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n19185) );
  AOI21_X1 U22165 ( .B1(n19199), .B2(P2_REIP_REG_11__SCAN_IN), .A(n19198), 
        .ZN(n19184) );
  OAI211_X1 U22166 ( .C1(n19187), .C2(n19186), .A(n19185), .B(n19184), .ZN(
        n19188) );
  AOI21_X1 U22167 ( .B1(n19190), .B2(n19189), .A(n19188), .ZN(n19197) );
  NAND2_X1 U22168 ( .A1(n13426), .A2(n19191), .ZN(n19193) );
  XNOR2_X1 U22169 ( .A(n19193), .B(n19192), .ZN(n19195) );
  AOI22_X1 U22170 ( .A1(n19195), .A2(n19227), .B1(n19226), .B2(n19194), .ZN(
        n19196) );
  OAI211_X1 U22171 ( .C1(n19231), .C2(n19283), .A(n19197), .B(n19196), .ZN(
        P2_U2844) );
  AOI21_X1 U22172 ( .B1(n19199), .B2(P2_REIP_REG_6__SCAN_IN), .A(n19198), .ZN(
        n19201) );
  NAND2_X1 U22173 ( .A1(n19221), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n19200) );
  OAI211_X1 U22174 ( .C1(n19202), .C2(n19216), .A(n19201), .B(n19200), .ZN(
        n19203) );
  INV_X1 U22175 ( .A(n19203), .ZN(n19212) );
  NOR2_X1 U22176 ( .A1(n10085), .A2(n19204), .ZN(n19206) );
  XNOR2_X1 U22177 ( .A(n19206), .B(n19205), .ZN(n19210) );
  AOI222_X1 U22178 ( .A1(n19210), .A2(n19227), .B1(n19209), .B2(n19208), .C1(
        n19226), .C2(n19207), .ZN(n19211) );
  OAI211_X1 U22179 ( .C1(n19218), .C2(n19213), .A(n19212), .B(n19211), .ZN(
        P2_U2849) );
  OAI21_X1 U22180 ( .B1(n19215), .B2(n16460), .A(n19214), .ZN(n19220) );
  OAI22_X1 U22181 ( .A1(n19218), .A2(n10673), .B1(n19217), .B2(n19216), .ZN(
        n19219) );
  AOI211_X1 U22182 ( .C1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n19221), .A(
        n19220), .B(n19219), .ZN(n19230) );
  NAND2_X1 U22183 ( .A1(n13426), .A2(n19222), .ZN(n19224) );
  XNOR2_X1 U22184 ( .A(n19224), .B(n19223), .ZN(n19228) );
  AOI22_X1 U22185 ( .A1(n19228), .A2(n19227), .B1(n19226), .B2(n19225), .ZN(
        n19229) );
  OAI211_X1 U22186 ( .C1(n19231), .C2(n19303), .A(n19230), .B(n19229), .ZN(
        P2_U2850) );
  AOI21_X1 U22187 ( .B1(n19233), .B2(n19232), .A(n14347), .ZN(n19267) );
  AOI22_X1 U22188 ( .A1(n19267), .A2(n19260), .B1(P2_EBX_REG_16__SCAN_IN), 
        .B2(n19259), .ZN(n19234) );
  OAI21_X1 U22189 ( .B1(n19259), .B2(n19235), .A(n19234), .ZN(P2_U2871) );
  AOI211_X1 U22190 ( .C1(n19236), .C2(n13910), .A(n19254), .B(n14028), .ZN(
        n19237) );
  AOI21_X1 U22191 ( .B1(P2_EBX_REG_14__SCAN_IN), .B2(n19259), .A(n19237), .ZN(
        n19238) );
  OAI21_X1 U22192 ( .B1(n19239), .B2(n19259), .A(n19238), .ZN(P2_U2873) );
  AOI21_X1 U22193 ( .B1(n19246), .B2(n19241), .A(n19240), .ZN(n19242) );
  NOR3_X1 U22194 ( .A1(n19242), .A2(n9771), .A3(n19254), .ZN(n19243) );
  AOI21_X1 U22195 ( .B1(P2_EBX_REG_12__SCAN_IN), .B2(n19259), .A(n19243), .ZN(
        n19244) );
  OAI21_X1 U22196 ( .B1(n19245), .B2(n19259), .A(n19244), .ZN(P2_U2875) );
  AOI211_X1 U22197 ( .C1(n19248), .C2(n19247), .A(n19254), .B(n19246), .ZN(
        n19249) );
  AOI21_X1 U22198 ( .B1(n19250), .B2(n19252), .A(n19249), .ZN(n19251) );
  OAI21_X1 U22199 ( .B1(n19252), .B2(n9991), .A(n19251), .ZN(P2_U2877) );
  INV_X1 U22200 ( .A(n19253), .ZN(n19255) );
  AOI211_X1 U22201 ( .C1(n19255), .C2(n9780), .A(n19254), .B(n9697), .ZN(
        n19256) );
  AOI21_X1 U22202 ( .B1(P2_EBX_REG_8__SCAN_IN), .B2(n19259), .A(n19256), .ZN(
        n19257) );
  OAI21_X1 U22203 ( .B1(n19258), .B2(n19259), .A(n19257), .ZN(P2_U2879) );
  INV_X1 U22204 ( .A(n19307), .ZN(n19261) );
  AOI22_X1 U22205 ( .A1(n19261), .A2(n19260), .B1(P2_EBX_REG_4__SCAN_IN), .B2(
        n19259), .ZN(n19262) );
  OAI21_X1 U22206 ( .B1(n19259), .B2(n19263), .A(n19262), .ZN(P2_U2883) );
  AOI22_X1 U22207 ( .A1(n19264), .A2(n19360), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n19320), .ZN(n19271) );
  AOI22_X1 U22208 ( .A1(n19266), .A2(BUF2_REG_16__SCAN_IN), .B1(n19265), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n19270) );
  AOI22_X1 U22209 ( .A1(n19268), .A2(n19321), .B1(n19308), .B2(n19267), .ZN(
        n19269) );
  NAND3_X1 U22210 ( .A1(n19271), .A2(n19270), .A3(n19269), .ZN(P2_U2903) );
  OAI222_X1 U22211 ( .A1(n19273), .A2(n19304), .B1(n13598), .B2(n19293), .C1(
        n19272), .C2(n19329), .ZN(P2_U2904) );
  INV_X1 U22212 ( .A(n19274), .ZN(n19277) );
  AOI22_X1 U22213 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19320), .B1(n19275), 
        .B2(n19295), .ZN(n19276) );
  OAI21_X1 U22214 ( .B1(n19304), .B2(n19277), .A(n19276), .ZN(P2_U2905) );
  OAI222_X1 U22215 ( .A1(n19279), .A2(n19304), .B1(n13519), .B2(n19293), .C1(
        n19329), .C2(n19278), .ZN(P2_U2906) );
  AOI22_X1 U22216 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19320), .B1(n19371), 
        .B2(n19295), .ZN(n19280) );
  OAI21_X1 U22217 ( .B1(n19304), .B2(n19281), .A(n19280), .ZN(P2_U2907) );
  OAI222_X1 U22218 ( .A1(n19283), .A2(n19304), .B1(n13530), .B2(n19293), .C1(
        n19329), .C2(n19282), .ZN(P2_U2908) );
  INV_X1 U22219 ( .A(n19284), .ZN(n19286) );
  AOI22_X1 U22220 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19320), .B1(n19367), 
        .B2(n19295), .ZN(n19285) );
  OAI21_X1 U22221 ( .B1(n19304), .B2(n19286), .A(n19285), .ZN(P2_U2909) );
  OAI222_X1 U22222 ( .A1(n19288), .A2(n19304), .B1(n13527), .B2(n19293), .C1(
        n19329), .C2(n19287), .ZN(P2_U2910) );
  INV_X1 U22223 ( .A(n19289), .ZN(n19291) );
  AOI22_X1 U22224 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19320), .B1(n19363), .B2(
        n19295), .ZN(n19290) );
  OAI21_X1 U22225 ( .B1(n19304), .B2(n19291), .A(n19290), .ZN(P2_U2911) );
  INV_X1 U22226 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19342) );
  OAI222_X1 U22227 ( .A1(n19292), .A2(n19304), .B1(n19342), .B2(n19293), .C1(
        n19329), .C2(n19441), .ZN(P2_U2912) );
  INV_X1 U22228 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19344) );
  OAI222_X1 U22229 ( .A1(n19294), .A2(n19304), .B1(n19344), .B2(n19293), .C1(
        n19329), .C2(n19431), .ZN(P2_U2913) );
  INV_X1 U22230 ( .A(n19424), .ZN(n19296) );
  AOI22_X1 U22231 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19320), .B1(n19296), .B2(
        n19295), .ZN(n19302) );
  AOI21_X1 U22232 ( .B1(n19298), .B2(n20084), .A(n19297), .ZN(n19314) );
  XOR2_X1 U22233 ( .A(n20078), .B(n20074), .Z(n19315) );
  NOR2_X1 U22234 ( .A1(n19314), .A2(n19315), .ZN(n19313) );
  AOI21_X1 U22235 ( .B1(n20078), .B2(n19299), .A(n19313), .ZN(n19300) );
  NOR2_X1 U22236 ( .A1(n19300), .A2(n19305), .ZN(n19306) );
  OR3_X1 U22237 ( .A1(n19306), .A2(n19307), .A3(n19325), .ZN(n19301) );
  OAI211_X1 U22238 ( .C1(n19304), .C2(n19303), .A(n19302), .B(n19301), .ZN(
        P2_U2914) );
  AOI22_X1 U22239 ( .A1(n19321), .A2(n19305), .B1(n19320), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n19311) );
  XOR2_X1 U22240 ( .A(n19307), .B(n19306), .Z(n19309) );
  NAND2_X1 U22241 ( .A1(n19309), .A2(n19308), .ZN(n19310) );
  OAI211_X1 U22242 ( .C1(n19418), .C2(n19329), .A(n19311), .B(n19310), .ZN(
        P2_U2915) );
  INV_X1 U22243 ( .A(n20078), .ZN(n19312) );
  AOI22_X1 U22244 ( .A1(n19312), .A2(n19321), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19320), .ZN(n19318) );
  AOI21_X1 U22245 ( .B1(n19315), .B2(n19314), .A(n19313), .ZN(n19316) );
  OR2_X1 U22246 ( .A1(n19316), .A2(n19325), .ZN(n19317) );
  OAI211_X1 U22247 ( .C1(n19319), .C2(n19329), .A(n19318), .B(n19317), .ZN(
        P2_U2916) );
  AOI22_X1 U22248 ( .A1(n19321), .A2(n20096), .B1(n19320), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19328) );
  AOI21_X1 U22249 ( .B1(n19324), .B2(n19323), .A(n19322), .ZN(n19326) );
  OR2_X1 U22250 ( .A1(n19326), .A2(n19325), .ZN(n19327) );
  OAI211_X1 U22251 ( .C1(n19330), .C2(n19329), .A(n19328), .B(n19327), .ZN(
        P2_U2918) );
  AND2_X1 U22252 ( .A1(n19339), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  AOI22_X1 U22253 ( .A1(n19356), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19355), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19332) );
  OAI21_X1 U22254 ( .B1(n13598), .B2(n19358), .A(n19332), .ZN(P2_U2936) );
  INV_X1 U22255 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19391) );
  AOI22_X1 U22256 ( .A1(n19356), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19355), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19333) );
  OAI21_X1 U22257 ( .B1(n19391), .B2(n19358), .A(n19333), .ZN(P2_U2937) );
  AOI22_X1 U22258 ( .A1(n19356), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19355), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19334) );
  OAI21_X1 U22259 ( .B1(n13519), .B2(n19358), .A(n19334), .ZN(P2_U2938) );
  INV_X1 U22260 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19386) );
  AOI22_X1 U22261 ( .A1(n19356), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19355), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19335) );
  OAI21_X1 U22262 ( .B1(n19386), .B2(n19358), .A(n19335), .ZN(P2_U2939) );
  AOI22_X1 U22263 ( .A1(n19356), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19336) );
  OAI21_X1 U22264 ( .B1(n13530), .B2(n19358), .A(n19336), .ZN(P2_U2940) );
  INV_X1 U22265 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19383) );
  AOI22_X1 U22266 ( .A1(n19356), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19337) );
  OAI21_X1 U22267 ( .B1(n19383), .B2(n19358), .A(n19337), .ZN(P2_U2941) );
  AOI22_X1 U22268 ( .A1(n19356), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19338) );
  OAI21_X1 U22269 ( .B1(n13527), .B2(n19358), .A(n19338), .ZN(P2_U2942) );
  INV_X1 U22270 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19380) );
  AOI22_X1 U22271 ( .A1(n19356), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19339), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19340) );
  OAI21_X1 U22272 ( .B1(n19380), .B2(n19358), .A(n19340), .ZN(P2_U2943) );
  AOI22_X1 U22273 ( .A1(n19356), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19355), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19341) );
  OAI21_X1 U22274 ( .B1(n19342), .B2(n19358), .A(n19341), .ZN(P2_U2944) );
  AOI22_X1 U22275 ( .A1(n19356), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19355), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19343) );
  OAI21_X1 U22276 ( .B1(n19344), .B2(n19358), .A(n19343), .ZN(P2_U2945) );
  INV_X1 U22277 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19346) );
  AOI22_X1 U22278 ( .A1(n19356), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19355), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19345) );
  OAI21_X1 U22279 ( .B1(n19346), .B2(n19358), .A(n19345), .ZN(P2_U2946) );
  INV_X1 U22280 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19348) );
  AOI22_X1 U22281 ( .A1(n19356), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19355), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19347) );
  OAI21_X1 U22282 ( .B1(n19348), .B2(n19358), .A(n19347), .ZN(P2_U2947) );
  INV_X1 U22283 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19350) );
  AOI22_X1 U22284 ( .A1(n19356), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19355), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19349) );
  OAI21_X1 U22285 ( .B1(n19350), .B2(n19358), .A(n19349), .ZN(P2_U2948) );
  INV_X1 U22286 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19352) );
  AOI22_X1 U22287 ( .A1(n19356), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19355), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19351) );
  OAI21_X1 U22288 ( .B1(n19352), .B2(n19358), .A(n19351), .ZN(P2_U2949) );
  AOI22_X1 U22289 ( .A1(n19356), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19355), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19353) );
  OAI21_X1 U22290 ( .B1(n19354), .B2(n19358), .A(n19353), .ZN(P2_U2950) );
  AOI22_X1 U22291 ( .A1(n19356), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19355), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19357) );
  OAI21_X1 U22292 ( .B1(n13596), .B2(n19358), .A(n19357), .ZN(P2_U2951) );
  AOI22_X1 U22293 ( .A1(n19388), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19360), 
        .B2(n19359), .ZN(n19361) );
  OAI21_X1 U22294 ( .B1(n19362), .B2(n19390), .A(n19361), .ZN(P2_U2952) );
  INV_X1 U22295 ( .A(n19363), .ZN(n19364) );
  NOR2_X1 U22296 ( .A1(n19376), .A2(n19364), .ZN(n19378) );
  AOI21_X1 U22297 ( .B1(n19388), .B2(P2_UWORD_REG_8__SCAN_IN), .A(n19378), 
        .ZN(n19365) );
  OAI21_X1 U22298 ( .B1(n19366), .B2(n19390), .A(n19365), .ZN(P2_U2960) );
  INV_X1 U22299 ( .A(n19367), .ZN(n19368) );
  NOR2_X1 U22300 ( .A1(n19376), .A2(n19368), .ZN(n19381) );
  AOI21_X1 U22301 ( .B1(n19388), .B2(P2_UWORD_REG_10__SCAN_IN), .A(n19381), 
        .ZN(n19369) );
  OAI21_X1 U22302 ( .B1(n19370), .B2(n19390), .A(n19369), .ZN(P2_U2962) );
  INV_X1 U22303 ( .A(n19371), .ZN(n19372) );
  NOR2_X1 U22304 ( .A1(n19376), .A2(n19372), .ZN(n19384) );
  AOI21_X1 U22305 ( .B1(n19388), .B2(P2_UWORD_REG_12__SCAN_IN), .A(n19384), 
        .ZN(n19373) );
  OAI21_X1 U22306 ( .B1(n19374), .B2(n19390), .A(n19373), .ZN(P2_U2964) );
  NOR2_X1 U22307 ( .A1(n19376), .A2(n19375), .ZN(n19387) );
  AOI21_X1 U22308 ( .B1(n19388), .B2(P2_UWORD_REG_14__SCAN_IN), .A(n19387), 
        .ZN(n19377) );
  OAI21_X1 U22309 ( .B1(n13277), .B2(n19390), .A(n19377), .ZN(P2_U2966) );
  AOI21_X1 U22310 ( .B1(n19388), .B2(P2_LWORD_REG_8__SCAN_IN), .A(n19378), 
        .ZN(n19379) );
  OAI21_X1 U22311 ( .B1(n19380), .B2(n19390), .A(n19379), .ZN(P2_U2975) );
  AOI21_X1 U22312 ( .B1(n19388), .B2(P2_LWORD_REG_10__SCAN_IN), .A(n19381), 
        .ZN(n19382) );
  OAI21_X1 U22313 ( .B1(n19383), .B2(n19390), .A(n19382), .ZN(P2_U2977) );
  AOI21_X1 U22314 ( .B1(n19388), .B2(P2_LWORD_REG_12__SCAN_IN), .A(n19384), 
        .ZN(n19385) );
  OAI21_X1 U22315 ( .B1(n19386), .B2(n19390), .A(n19385), .ZN(P2_U2979) );
  AOI21_X1 U22316 ( .B1(n19388), .B2(P2_LWORD_REG_14__SCAN_IN), .A(n19387), 
        .ZN(n19389) );
  OAI21_X1 U22317 ( .B1(n19391), .B2(n19390), .A(n19389), .ZN(P2_U2981) );
  INV_X1 U22318 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19393) );
  OAI22_X1 U22319 ( .A1(n19394), .A2(n19393), .B1(n19214), .B2(n19392), .ZN(
        n19395) );
  INV_X1 U22320 ( .A(n19395), .ZN(n19403) );
  AOI222_X1 U22321 ( .A1(n19401), .A2(n19400), .B1(n19399), .B2(n19398), .C1(
        n19397), .C2(n19396), .ZN(n19402) );
  OAI211_X1 U22322 ( .C1(n19405), .C2(n19404), .A(n19403), .B(n19402), .ZN(
        P2_U3010) );
  AOI22_X1 U22323 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19437), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19436), .ZN(n19941) );
  OR2_X1 U22324 ( .A1(n19438), .A2(n10353), .ZN(n19869) );
  OAI22_X1 U22325 ( .A1(n19989), .A2(n19941), .B1(n19439), .B2(n19869), .ZN(
        n19406) );
  INV_X1 U22326 ( .A(n19406), .ZN(n19409) );
  NOR2_X2 U22327 ( .A1(n19865), .A2(n19407), .ZN(n19929) );
  AOI22_X1 U22328 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19437), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19436), .ZN(n19779) );
  AOI22_X1 U22329 ( .A1(n19929), .A2(n19442), .B1(n19465), .B2(n19938), .ZN(
        n19408) );
  OAI211_X1 U22330 ( .C1(n19435), .C2(n19410), .A(n19409), .B(n19408), .ZN(
        P2_U3048) );
  AOI22_X1 U22331 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19437), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19436), .ZN(n19953) );
  AOI22_X1 U22332 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19437), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19436), .ZN(n19883) );
  OR2_X1 U22333 ( .A1(n19438), .A2(n19411), .ZN(n19882) );
  OAI22_X1 U22334 ( .A1(n19989), .A2(n19883), .B1(n19439), .B2(n19882), .ZN(
        n19412) );
  INV_X1 U22335 ( .A(n19412), .ZN(n19415) );
  NOR2_X2 U22336 ( .A1(n19865), .A2(n19413), .ZN(n19949) );
  AOI22_X1 U22337 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19443), .B1(
        n19949), .B2(n19442), .ZN(n19414) );
  OAI211_X1 U22338 ( .C1(n19953), .C2(n19473), .A(n19415), .B(n19414), .ZN(
        P2_U3050) );
  INV_X1 U22339 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19421) );
  AOI22_X2 U22340 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19437), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19436), .ZN(n19896) );
  OR2_X1 U22341 ( .A1(n19438), .A2(n19416), .ZN(n19895) );
  OAI22_X1 U22342 ( .A1(n19989), .A2(n19896), .B1(n19439), .B2(n19895), .ZN(
        n19417) );
  INV_X1 U22343 ( .A(n19417), .ZN(n19420) );
  NOR2_X2 U22344 ( .A1(n19865), .A2(n19418), .ZN(n19961) );
  AOI22_X1 U22345 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19437), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19436), .ZN(n19965) );
  AOI22_X1 U22346 ( .A1(n19961), .A2(n19442), .B1(n19465), .B2(n19898), .ZN(
        n19419) );
  OAI211_X1 U22347 ( .C1(n19435), .C2(n19421), .A(n19420), .B(n19419), .ZN(
        P2_U3052) );
  AOI22_X1 U22348 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19436), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19437), .ZN(n19903) );
  OR2_X1 U22349 ( .A1(n19438), .A2(n19422), .ZN(n19902) );
  OAI22_X1 U22350 ( .A1(n19989), .A2(n19903), .B1(n19439), .B2(n19902), .ZN(
        n19423) );
  INV_X1 U22351 ( .A(n19423), .ZN(n19426) );
  NOR2_X2 U22352 ( .A1(n19865), .A2(n19424), .ZN(n19967) );
  AOI22_X1 U22353 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19443), .B1(
        n19967), .B2(n19442), .ZN(n19425) );
  OAI211_X1 U22354 ( .C1(n19971), .C2(n19473), .A(n19426), .B(n19425), .ZN(
        P2_U3053) );
  OAI22_X2 U22355 ( .A1(n19429), .A2(n19428), .B1(n20360), .B2(n19427), .ZN(
        n19909) );
  OR2_X1 U22356 ( .A1(n19438), .A2(n10357), .ZN(n19688) );
  AOI22_X1 U22357 ( .A1(n19975), .A2(n19909), .B1(n19430), .B2(n19972), .ZN(
        n19433) );
  NOR2_X2 U22358 ( .A1(n19865), .A2(n19431), .ZN(n19973) );
  INV_X1 U22359 ( .A(n19913), .ZN(n19974) );
  AOI22_X1 U22360 ( .A1(n19973), .A2(n19442), .B1(n19465), .B2(n19974), .ZN(
        n19432) );
  OAI211_X1 U22361 ( .C1(n19435), .C2(n19434), .A(n19433), .B(n19432), .ZN(
        P2_U3054) );
  AOI22_X2 U22362 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19436), .B1(
        BUF1_REG_23__SCAN_IN), .B2(n19437), .ZN(n19990) );
  AOI22_X1 U22363 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19437), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19436), .ZN(n19916) );
  OR2_X1 U22364 ( .A1(n19438), .A2(n9658), .ZN(n19915) );
  OAI22_X1 U22365 ( .A1(n19989), .A2(n19916), .B1(n19439), .B2(n19915), .ZN(
        n19440) );
  INV_X1 U22366 ( .A(n19440), .ZN(n19445) );
  NOR2_X2 U22367 ( .A1(n19865), .A2(n19441), .ZN(n19982) );
  AOI22_X1 U22368 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19443), .B1(
        n19982), .B2(n19442), .ZN(n19444) );
  OAI211_X1 U22369 ( .C1(n19990), .C2(n19473), .A(n19445), .B(n19444), .ZN(
        P2_U3055) );
  NOR2_X1 U22370 ( .A1(n19699), .A2(n19504), .ZN(n19468) );
  INV_X1 U22371 ( .A(n19451), .ZN(n19447) );
  AOI211_X2 U22372 ( .C1(n19448), .C2(n19926), .A(n19632), .B(n19447), .ZN(
        n19469) );
  AOI22_X1 U22373 ( .A1(n19469), .A2(n19929), .B1(n19928), .B2(n19468), .ZN(
        n19454) );
  OAI21_X1 U22374 ( .B1(n19634), .B2(n19700), .A(n19448), .ZN(n19452) );
  INV_X1 U22375 ( .A(n19468), .ZN(n19449) );
  NAND2_X1 U22376 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19449), .ZN(n19450) );
  NAND4_X1 U22377 ( .A1(n19452), .A2(n19936), .A3(n19451), .A4(n19450), .ZN(
        n19470) );
  INV_X1 U22378 ( .A(n19941), .ZN(n19776) );
  AOI22_X1 U22379 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19470), .B1(
        n19465), .B2(n19776), .ZN(n19453) );
  OAI211_X1 U22380 ( .C1(n19779), .C2(n19492), .A(n19454), .B(n19453), .ZN(
        P2_U3056) );
  AOI22_X1 U22381 ( .A1(n19469), .A2(n19943), .B1(n19942), .B2(n19468), .ZN(
        n19456) );
  AOI22_X1 U22382 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19470), .B1(
        n19465), .B2(n19944), .ZN(n19455) );
  OAI211_X1 U22383 ( .C1(n19947), .C2(n19492), .A(n19456), .B(n19455), .ZN(
        P2_U3057) );
  AOI22_X1 U22384 ( .A1(n19469), .A2(n19949), .B1(n19948), .B2(n19468), .ZN(
        n19458) );
  INV_X1 U22385 ( .A(n19953), .ZN(n19885) );
  AOI22_X1 U22386 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19470), .B1(
        n19499), .B2(n19885), .ZN(n19457) );
  OAI211_X1 U22387 ( .C1(n19883), .C2(n19473), .A(n19458), .B(n19457), .ZN(
        P2_U3058) );
  AOI22_X1 U22388 ( .A1(n19469), .A2(n19955), .B1(n19954), .B2(n19468), .ZN(
        n19460) );
  AOI22_X1 U22389 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19470), .B1(
        n19465), .B2(n19892), .ZN(n19459) );
  OAI211_X1 U22390 ( .C1(n19890), .C2(n19492), .A(n19460), .B(n19459), .ZN(
        P2_U3059) );
  AOI22_X1 U22391 ( .A1(n19469), .A2(n19961), .B1(n19960), .B2(n19468), .ZN(
        n19462) );
  AOI22_X1 U22392 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19470), .B1(
        n19499), .B2(n19898), .ZN(n19461) );
  OAI211_X1 U22393 ( .C1(n19896), .C2(n19473), .A(n19462), .B(n19461), .ZN(
        P2_U3060) );
  AOI22_X1 U22394 ( .A1(n19469), .A2(n19967), .B1(n19966), .B2(n19468), .ZN(
        n19464) );
  INV_X1 U22395 ( .A(n19903), .ZN(n19968) );
  AOI22_X1 U22396 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19470), .B1(
        n19465), .B2(n19968), .ZN(n19463) );
  OAI211_X1 U22397 ( .C1(n19971), .C2(n19492), .A(n19464), .B(n19463), .ZN(
        P2_U3061) );
  AOI22_X1 U22398 ( .A1(n19469), .A2(n19973), .B1(n19972), .B2(n19468), .ZN(
        n19467) );
  AOI22_X1 U22399 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19470), .B1(
        n19465), .B2(n19909), .ZN(n19466) );
  OAI211_X1 U22400 ( .C1(n19913), .C2(n19492), .A(n19467), .B(n19466), .ZN(
        P2_U3062) );
  INV_X1 U22401 ( .A(n19915), .ZN(n19980) );
  AOI22_X1 U22402 ( .A1(n19469), .A2(n19982), .B1(n19980), .B2(n19468), .ZN(
        n19472) );
  INV_X1 U22403 ( .A(n19990), .ZN(n19655) );
  AOI22_X1 U22404 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19470), .B1(
        n19499), .B2(n19655), .ZN(n19471) );
  OAI211_X1 U22405 ( .C1(n19916), .C2(n19473), .A(n19472), .B(n19471), .ZN(
        P2_U3063) );
  NOR2_X1 U22406 ( .A1(n19734), .A2(n19504), .ZN(n19497) );
  OAI21_X1 U22407 ( .B1(n10502), .B2(n19497), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19475) );
  NAND2_X1 U22408 ( .A1(n19598), .A2(n19474), .ZN(n19476) );
  NAND2_X1 U22409 ( .A1(n19475), .A2(n19476), .ZN(n19498) );
  AOI22_X1 U22410 ( .A1(n19498), .A2(n19929), .B1(n19928), .B2(n19497), .ZN(
        n19483) );
  OAI21_X1 U22411 ( .B1(n19518), .B2(n19499), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19477) );
  NAND3_X1 U22412 ( .A1(n19477), .A2(n20069), .A3(n19476), .ZN(n19481) );
  INV_X1 U22413 ( .A(n19497), .ZN(n19478) );
  OAI211_X1 U22414 ( .C1(n19479), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19860), 
        .B(n19478), .ZN(n19480) );
  NAND3_X1 U22415 ( .A1(n19481), .A2(n19936), .A3(n19480), .ZN(n19500) );
  AOI22_X1 U22416 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19500), .B1(
        n19518), .B2(n19938), .ZN(n19482) );
  OAI211_X1 U22417 ( .C1(n19941), .C2(n19492), .A(n19483), .B(n19482), .ZN(
        P2_U3064) );
  AOI22_X1 U22418 ( .A1(n19498), .A2(n19943), .B1(n19942), .B2(n19497), .ZN(
        n19485) );
  AOI22_X1 U22419 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19500), .B1(
        n19499), .B2(n19944), .ZN(n19484) );
  OAI211_X1 U22420 ( .C1(n19947), .C2(n19534), .A(n19485), .B(n19484), .ZN(
        P2_U3065) );
  AOI22_X1 U22421 ( .A1(n19498), .A2(n19949), .B1(n19948), .B2(n19497), .ZN(
        n19487) );
  INV_X1 U22422 ( .A(n19883), .ZN(n19950) );
  AOI22_X1 U22423 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19500), .B1(
        n19499), .B2(n19950), .ZN(n19486) );
  OAI211_X1 U22424 ( .C1(n19953), .C2(n19534), .A(n19487), .B(n19486), .ZN(
        P2_U3066) );
  INV_X1 U22425 ( .A(n19892), .ZN(n19959) );
  AOI22_X1 U22426 ( .A1(n19498), .A2(n19955), .B1(n19954), .B2(n19497), .ZN(
        n19489) );
  INV_X1 U22427 ( .A(n19890), .ZN(n19956) );
  AOI22_X1 U22428 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19500), .B1(
        n19518), .B2(n19956), .ZN(n19488) );
  OAI211_X1 U22429 ( .C1(n19959), .C2(n19492), .A(n19489), .B(n19488), .ZN(
        P2_U3067) );
  AOI22_X1 U22430 ( .A1(n19498), .A2(n19961), .B1(n19960), .B2(n19497), .ZN(
        n19491) );
  AOI22_X1 U22431 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19500), .B1(
        n19518), .B2(n19898), .ZN(n19490) );
  OAI211_X1 U22432 ( .C1(n19896), .C2(n19492), .A(n19491), .B(n19490), .ZN(
        P2_U3068) );
  AOI22_X1 U22433 ( .A1(n19498), .A2(n19967), .B1(n19966), .B2(n19497), .ZN(
        n19494) );
  AOI22_X1 U22434 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19500), .B1(
        n19499), .B2(n19968), .ZN(n19493) );
  OAI211_X1 U22435 ( .C1(n19971), .C2(n19534), .A(n19494), .B(n19493), .ZN(
        P2_U3069) );
  AOI22_X1 U22436 ( .A1(n19498), .A2(n19973), .B1(n19972), .B2(n19497), .ZN(
        n19496) );
  AOI22_X1 U22437 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19500), .B1(
        n19499), .B2(n19909), .ZN(n19495) );
  OAI211_X1 U22438 ( .C1(n19913), .C2(n19534), .A(n19496), .B(n19495), .ZN(
        P2_U3070) );
  AOI22_X1 U22439 ( .A1(n19498), .A2(n19982), .B1(n19980), .B2(n19497), .ZN(
        n19502) );
  INV_X1 U22440 ( .A(n19916), .ZN(n19984) );
  AOI22_X1 U22441 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19500), .B1(
        n19499), .B2(n19984), .ZN(n19501) );
  OAI211_X1 U22442 ( .C1(n19990), .C2(n19534), .A(n19502), .B(n19501), .ZN(
        P2_U3071) );
  NOR2_X1 U22443 ( .A1(n19765), .A2(n19504), .ZN(n19525) );
  INV_X1 U22444 ( .A(n19525), .ZN(n19528) );
  NOR2_X1 U22445 ( .A1(n19869), .A2(n19528), .ZN(n19503) );
  AOI21_X1 U22446 ( .B1(n19518), .B2(n19776), .A(n19503), .ZN(n19512) );
  OAI21_X1 U22447 ( .B1(n19634), .B2(n20071), .A(n20069), .ZN(n19510) );
  NOR2_X1 U22448 ( .A1(n20098), .A2(n19504), .ZN(n19507) );
  INV_X1 U22449 ( .A(n10648), .ZN(n19505) );
  OAI211_X1 U22450 ( .C1(n19505), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19860), 
        .B(n19528), .ZN(n19506) );
  OAI211_X1 U22451 ( .C1(n19510), .C2(n19507), .A(n19936), .B(n19506), .ZN(
        n19531) );
  INV_X1 U22452 ( .A(n19507), .ZN(n19509) );
  OAI21_X1 U22453 ( .B1(n10648), .B2(n19525), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19508) );
  OAI21_X1 U22454 ( .B1(n19510), .B2(n19509), .A(n19508), .ZN(n19530) );
  AOI22_X1 U22455 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19531), .B1(
        n19929), .B2(n19530), .ZN(n19511) );
  OAI211_X1 U22456 ( .C1(n19779), .C2(n19557), .A(n19512), .B(n19511), .ZN(
        P2_U3072) );
  AOI22_X1 U22457 ( .A1(n19518), .A2(n19944), .B1(n19942), .B2(n19525), .ZN(
        n19514) );
  AOI22_X1 U22458 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19531), .B1(
        n19943), .B2(n19530), .ZN(n19513) );
  OAI211_X1 U22459 ( .C1(n19947), .C2(n19557), .A(n19514), .B(n19513), .ZN(
        P2_U3073) );
  NOR2_X1 U22460 ( .A1(n19882), .A2(n19528), .ZN(n19515) );
  AOI21_X1 U22461 ( .B1(n19518), .B2(n19950), .A(n19515), .ZN(n19517) );
  AOI22_X1 U22462 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19531), .B1(
        n19949), .B2(n19530), .ZN(n19516) );
  OAI211_X1 U22463 ( .C1(n19953), .C2(n19557), .A(n19517), .B(n19516), .ZN(
        P2_U3074) );
  AOI22_X1 U22464 ( .A1(n19518), .A2(n19892), .B1(n19954), .B2(n19525), .ZN(
        n19520) );
  AOI22_X1 U22465 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19531), .B1(
        n19955), .B2(n19530), .ZN(n19519) );
  OAI211_X1 U22466 ( .C1(n19890), .C2(n19557), .A(n19520), .B(n19519), .ZN(
        P2_U3075) );
  AOI22_X1 U22467 ( .A1(n19898), .A2(n19564), .B1(n19525), .B2(n19960), .ZN(
        n19522) );
  AOI22_X1 U22468 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19531), .B1(
        n19961), .B2(n19530), .ZN(n19521) );
  OAI211_X1 U22469 ( .C1(n19896), .C2(n19534), .A(n19522), .B(n19521), .ZN(
        P2_U3076) );
  INV_X1 U22470 ( .A(n19971), .ZN(n19848) );
  AOI22_X1 U22471 ( .A1(n19564), .A2(n19848), .B1(n19525), .B2(n19966), .ZN(
        n19524) );
  AOI22_X1 U22472 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19531), .B1(
        n19967), .B2(n19530), .ZN(n19523) );
  OAI211_X1 U22473 ( .C1(n19903), .C2(n19534), .A(n19524), .B(n19523), .ZN(
        P2_U3077) );
  INV_X1 U22474 ( .A(n19909), .ZN(n19979) );
  AOI22_X1 U22475 ( .A1(n19974), .A2(n19564), .B1(n19525), .B2(n19972), .ZN(
        n19527) );
  AOI22_X1 U22476 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19531), .B1(
        n19973), .B2(n19530), .ZN(n19526) );
  OAI211_X1 U22477 ( .C1(n19979), .C2(n19534), .A(n19527), .B(n19526), .ZN(
        P2_U3078) );
  NOR2_X1 U22478 ( .A1(n19915), .A2(n19528), .ZN(n19529) );
  AOI21_X1 U22479 ( .B1(n19564), .B2(n19655), .A(n19529), .ZN(n19533) );
  AOI22_X1 U22480 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19531), .B1(
        n19982), .B2(n19530), .ZN(n19532) );
  OAI211_X1 U22481 ( .C1(n19916), .C2(n19534), .A(n19533), .B(n19532), .ZN(
        P2_U3079) );
  INV_X1 U22482 ( .A(n19535), .ZN(n19536) );
  OR2_X1 U22483 ( .A1(n19537), .A2(n19536), .ZN(n19805) );
  NOR2_X1 U22484 ( .A1(n19805), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19546) );
  INV_X1 U22485 ( .A(n19546), .ZN(n19539) );
  NAND2_X1 U22486 ( .A1(n20081), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19630) );
  OR2_X1 U22487 ( .A1(n19630), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19575) );
  NOR2_X1 U22488 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19575), .ZN(
        n19562) );
  OAI21_X1 U22489 ( .B1(n10637), .B2(n19562), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19538) );
  OAI21_X1 U22490 ( .B1(n19860), .B2(n19539), .A(n19538), .ZN(n19563) );
  AOI22_X1 U22491 ( .A1(n19563), .A2(n19929), .B1(n19928), .B2(n19562), .ZN(
        n19548) );
  AOI21_X1 U22492 ( .B1(n19557), .B2(n19589), .A(n19541), .ZN(n19545) );
  INV_X1 U22493 ( .A(n19562), .ZN(n19542) );
  OAI211_X1 U22494 ( .C1(n19543), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19860), 
        .B(n19542), .ZN(n19544) );
  OAI211_X1 U22495 ( .C1(n19546), .C2(n19545), .A(n19544), .B(n19936), .ZN(
        n19565) );
  AOI22_X1 U22496 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19565), .B1(
        n19592), .B2(n19938), .ZN(n19547) );
  OAI211_X1 U22497 ( .C1(n19941), .C2(n19557), .A(n19548), .B(n19547), .ZN(
        P2_U3080) );
  AOI22_X1 U22498 ( .A1(n19563), .A2(n19943), .B1(n19942), .B2(n19562), .ZN(
        n19550) );
  AOI22_X1 U22499 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19565), .B1(
        n19564), .B2(n19944), .ZN(n19549) );
  OAI211_X1 U22500 ( .C1(n19947), .C2(n19589), .A(n19550), .B(n19549), .ZN(
        P2_U3081) );
  AOI22_X1 U22501 ( .A1(n19563), .A2(n19949), .B1(n19948), .B2(n19562), .ZN(
        n19552) );
  AOI22_X1 U22502 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19565), .B1(
        n19564), .B2(n19950), .ZN(n19551) );
  OAI211_X1 U22503 ( .C1(n19953), .C2(n19589), .A(n19552), .B(n19551), .ZN(
        P2_U3082) );
  AOI22_X1 U22504 ( .A1(n19563), .A2(n19955), .B1(n19954), .B2(n19562), .ZN(
        n19554) );
  AOI22_X1 U22505 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19565), .B1(
        n19592), .B2(n19956), .ZN(n19553) );
  OAI211_X1 U22506 ( .C1(n19959), .C2(n19557), .A(n19554), .B(n19553), .ZN(
        P2_U3083) );
  AOI22_X1 U22507 ( .A1(n19563), .A2(n19961), .B1(n19960), .B2(n19562), .ZN(
        n19556) );
  AOI22_X1 U22508 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19565), .B1(
        n19592), .B2(n19898), .ZN(n19555) );
  OAI211_X1 U22509 ( .C1(n19896), .C2(n19557), .A(n19556), .B(n19555), .ZN(
        P2_U3084) );
  AOI22_X1 U22510 ( .A1(n19563), .A2(n19967), .B1(n19966), .B2(n19562), .ZN(
        n19559) );
  AOI22_X1 U22511 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19565), .B1(
        n19564), .B2(n19968), .ZN(n19558) );
  OAI211_X1 U22512 ( .C1(n19971), .C2(n19589), .A(n19559), .B(n19558), .ZN(
        P2_U3085) );
  AOI22_X1 U22513 ( .A1(n19563), .A2(n19973), .B1(n19972), .B2(n19562), .ZN(
        n19561) );
  AOI22_X1 U22514 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19565), .B1(
        n19564), .B2(n19909), .ZN(n19560) );
  OAI211_X1 U22515 ( .C1(n19913), .C2(n19589), .A(n19561), .B(n19560), .ZN(
        P2_U3086) );
  AOI22_X1 U22516 ( .A1(n19563), .A2(n19982), .B1(n19980), .B2(n19562), .ZN(
        n19567) );
  AOI22_X1 U22517 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19565), .B1(
        n19564), .B2(n19984), .ZN(n19566) );
  OAI211_X1 U22518 ( .C1(n19990), .C2(n19589), .A(n19567), .B(n19566), .ZN(
        P2_U3087) );
  NOR2_X1 U22519 ( .A1(n19699), .A2(n19630), .ZN(n19600) );
  AOI22_X1 U22520 ( .A1(n19938), .A2(n19618), .B1(n19928), .B2(n19600), .ZN(
        n19578) );
  INV_X1 U22521 ( .A(n10649), .ZN(n19568) );
  AOI21_X1 U22522 ( .B1(n19568), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19572) );
  INV_X1 U22523 ( .A(n19634), .ZN(n19570) );
  INV_X1 U22524 ( .A(n19836), .ZN(n19569) );
  AOI21_X1 U22525 ( .B1(n19570), .B2(n19569), .A(n19860), .ZN(n19573) );
  NAND2_X1 U22526 ( .A1(n19573), .A2(n19575), .ZN(n19571) );
  OAI211_X1 U22527 ( .C1(n19600), .C2(n19572), .A(n19571), .B(n19936), .ZN(
        n19594) );
  INV_X1 U22528 ( .A(n19573), .ZN(n19576) );
  OAI21_X1 U22529 ( .B1(n10649), .B2(n19600), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19574) );
  OAI21_X1 U22530 ( .B1(n19576), .B2(n19575), .A(n19574), .ZN(n19593) );
  AOI22_X1 U22531 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19594), .B1(
        n19929), .B2(n19593), .ZN(n19577) );
  OAI211_X1 U22532 ( .C1(n19941), .C2(n19589), .A(n19578), .B(n19577), .ZN(
        P2_U3088) );
  AOI22_X1 U22533 ( .A1(n19592), .A2(n19944), .B1(n19942), .B2(n19600), .ZN(
        n19580) );
  AOI22_X1 U22534 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19594), .B1(
        n19943), .B2(n19593), .ZN(n19579) );
  OAI211_X1 U22535 ( .C1(n19947), .C2(n19626), .A(n19580), .B(n19579), .ZN(
        P2_U3089) );
  AOI22_X1 U22536 ( .A1(n19592), .A2(n19950), .B1(n19600), .B2(n19948), .ZN(
        n19582) );
  AOI22_X1 U22537 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19594), .B1(
        n19949), .B2(n19593), .ZN(n19581) );
  OAI211_X1 U22538 ( .C1(n19953), .C2(n19626), .A(n19582), .B(n19581), .ZN(
        P2_U3090) );
  AOI22_X1 U22539 ( .A1(n19618), .A2(n19956), .B1(n19600), .B2(n19954), .ZN(
        n19584) );
  AOI22_X1 U22540 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19594), .B1(
        n19955), .B2(n19593), .ZN(n19583) );
  OAI211_X1 U22541 ( .C1(n19959), .C2(n19589), .A(n19584), .B(n19583), .ZN(
        P2_U3091) );
  AOI22_X1 U22542 ( .A1(n19898), .A2(n19618), .B1(n19600), .B2(n19960), .ZN(
        n19586) );
  AOI22_X1 U22543 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19594), .B1(
        n19961), .B2(n19593), .ZN(n19585) );
  OAI211_X1 U22544 ( .C1(n19896), .C2(n19589), .A(n19586), .B(n19585), .ZN(
        P2_U3092) );
  AOI22_X1 U22545 ( .A1(n19618), .A2(n19848), .B1(n19600), .B2(n19966), .ZN(
        n19588) );
  AOI22_X1 U22546 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19594), .B1(
        n19967), .B2(n19593), .ZN(n19587) );
  OAI211_X1 U22547 ( .C1(n19903), .C2(n19589), .A(n19588), .B(n19587), .ZN(
        P2_U3093) );
  AOI22_X1 U22548 ( .A1(n19592), .A2(n19909), .B1(n19600), .B2(n19972), .ZN(
        n19591) );
  AOI22_X1 U22549 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19594), .B1(
        n19973), .B2(n19593), .ZN(n19590) );
  OAI211_X1 U22550 ( .C1(n19913), .C2(n19626), .A(n19591), .B(n19590), .ZN(
        P2_U3094) );
  AOI22_X1 U22551 ( .A1(n19592), .A2(n19984), .B1(n19600), .B2(n19980), .ZN(
        n19596) );
  AOI22_X1 U22552 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19594), .B1(
        n19982), .B2(n19593), .ZN(n19595) );
  OAI211_X1 U22553 ( .C1(n19990), .C2(n19626), .A(n19596), .B(n19595), .ZN(
        P2_U3095) );
  INV_X1 U22554 ( .A(n19598), .ZN(n19741) );
  NOR2_X1 U22555 ( .A1(n19734), .A2(n19630), .ZN(n19621) );
  OAI21_X1 U22556 ( .B1(n10516), .B2(n19621), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19599) );
  OAI21_X1 U22557 ( .B1(n19630), .B2(n19741), .A(n19599), .ZN(n19622) );
  AOI22_X1 U22558 ( .A1(n19622), .A2(n19929), .B1(n19928), .B2(n19621), .ZN(
        n19607) );
  AOI221_X1 U22559 ( .B1(n19618), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19649), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19600), .ZN(n19601) );
  INV_X1 U22560 ( .A(n19621), .ZN(n19602) );
  OAI21_X1 U22561 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19601), .A(n19602), 
        .ZN(n19605) );
  NAND3_X1 U22562 ( .A1(n19603), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19602), 
        .ZN(n19604) );
  NAND3_X1 U22563 ( .A1(n19605), .A2(n19936), .A3(n19604), .ZN(n19623) );
  AOI22_X1 U22564 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19623), .B1(
        n19618), .B2(n19776), .ZN(n19606) );
  OAI211_X1 U22565 ( .C1(n19779), .C2(n19659), .A(n19607), .B(n19606), .ZN(
        P2_U3096) );
  AOI22_X1 U22566 ( .A1(n19622), .A2(n19943), .B1(n19942), .B2(n19621), .ZN(
        n19609) );
  AOI22_X1 U22567 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19623), .B1(
        n19618), .B2(n19944), .ZN(n19608) );
  OAI211_X1 U22568 ( .C1(n19947), .C2(n19659), .A(n19609), .B(n19608), .ZN(
        P2_U3097) );
  AOI22_X1 U22569 ( .A1(n19622), .A2(n19949), .B1(n19948), .B2(n19621), .ZN(
        n19611) );
  AOI22_X1 U22570 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19623), .B1(
        n19618), .B2(n19950), .ZN(n19610) );
  OAI211_X1 U22571 ( .C1(n19953), .C2(n19659), .A(n19611), .B(n19610), .ZN(
        P2_U3098) );
  AOI22_X1 U22572 ( .A1(n19622), .A2(n19955), .B1(n19954), .B2(n19621), .ZN(
        n19613) );
  AOI22_X1 U22573 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19623), .B1(
        n19649), .B2(n19956), .ZN(n19612) );
  OAI211_X1 U22574 ( .C1(n19959), .C2(n19626), .A(n19613), .B(n19612), .ZN(
        P2_U3099) );
  AOI22_X1 U22575 ( .A1(n19622), .A2(n19961), .B1(n19960), .B2(n19621), .ZN(
        n19615) );
  AOI22_X1 U22576 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19623), .B1(
        n19649), .B2(n19898), .ZN(n19614) );
  OAI211_X1 U22577 ( .C1(n19896), .C2(n19626), .A(n19615), .B(n19614), .ZN(
        P2_U3100) );
  AOI22_X1 U22578 ( .A1(n19622), .A2(n19967), .B1(n19966), .B2(n19621), .ZN(
        n19617) );
  AOI22_X1 U22579 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19623), .B1(
        n19649), .B2(n19848), .ZN(n19616) );
  OAI211_X1 U22580 ( .C1(n19903), .C2(n19626), .A(n19617), .B(n19616), .ZN(
        P2_U3101) );
  AOI22_X1 U22581 ( .A1(n19622), .A2(n19973), .B1(n19972), .B2(n19621), .ZN(
        n19620) );
  AOI22_X1 U22582 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19623), .B1(
        n19618), .B2(n19909), .ZN(n19619) );
  OAI211_X1 U22583 ( .C1(n19913), .C2(n19659), .A(n19620), .B(n19619), .ZN(
        P2_U3102) );
  AOI22_X1 U22584 ( .A1(n19622), .A2(n19982), .B1(n19980), .B2(n19621), .ZN(
        n19625) );
  AOI22_X1 U22585 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19623), .B1(
        n19649), .B2(n19655), .ZN(n19624) );
  OAI211_X1 U22586 ( .C1(n19916), .C2(n19626), .A(n19625), .B(n19624), .ZN(
        P2_U3103) );
  INV_X1 U22587 ( .A(n19627), .ZN(n19629) );
  INV_X1 U22588 ( .A(n19931), .ZN(n19628) );
  NOR2_X1 U22589 ( .A1(n19925), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19638) );
  INV_X1 U22590 ( .A(n19638), .ZN(n19633) );
  NOR2_X1 U22591 ( .A1(n19765), .A2(n19630), .ZN(n19665) );
  OR3_X1 U22592 ( .A1(n9708), .A2(n19665), .A3(n19926), .ZN(n19635) );
  INV_X1 U22593 ( .A(n19635), .ZN(n19631) );
  AOI211_X2 U22594 ( .C1(n19633), .C2(n19926), .A(n19632), .B(n19631), .ZN(
        n19654) );
  AOI22_X1 U22595 ( .A1(n19654), .A2(n19929), .B1(n19665), .B2(n19928), .ZN(
        n19640) );
  NOR2_X1 U22596 ( .A1(n19634), .A2(n19931), .ZN(n20070) );
  OAI211_X1 U22597 ( .C1(n19665), .C2(n13484), .A(n19635), .B(n19936), .ZN(
        n19636) );
  INV_X1 U22598 ( .A(n19636), .ZN(n19637) );
  OAI21_X1 U22599 ( .B1(n20070), .B2(n19638), .A(n19637), .ZN(n19656) );
  AOI22_X1 U22600 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19656), .B1(
        n19649), .B2(n19776), .ZN(n19639) );
  OAI211_X1 U22601 ( .C1(n19779), .C2(n19693), .A(n19640), .B(n19639), .ZN(
        P2_U3104) );
  AOI22_X1 U22602 ( .A1(n19654), .A2(n19943), .B1(n19942), .B2(n19665), .ZN(
        n19642) );
  AOI22_X1 U22603 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19656), .B1(
        n19649), .B2(n19944), .ZN(n19641) );
  OAI211_X1 U22604 ( .C1(n19947), .C2(n19693), .A(n19642), .B(n19641), .ZN(
        P2_U3105) );
  AOI22_X1 U22605 ( .A1(n19654), .A2(n19949), .B1(n19665), .B2(n19948), .ZN(
        n19644) );
  AOI22_X1 U22606 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19656), .B1(
        n19673), .B2(n19885), .ZN(n19643) );
  OAI211_X1 U22607 ( .C1(n19883), .C2(n19659), .A(n19644), .B(n19643), .ZN(
        P2_U3106) );
  AOI22_X1 U22608 ( .A1(n19654), .A2(n19955), .B1(n19954), .B2(n19665), .ZN(
        n19646) );
  AOI22_X1 U22609 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19656), .B1(
        n19673), .B2(n19956), .ZN(n19645) );
  OAI211_X1 U22610 ( .C1(n19959), .C2(n19659), .A(n19646), .B(n19645), .ZN(
        P2_U3107) );
  AOI22_X1 U22611 ( .A1(n19654), .A2(n19961), .B1(n19665), .B2(n19960), .ZN(
        n19648) );
  INV_X1 U22612 ( .A(n19896), .ZN(n19962) );
  AOI22_X1 U22613 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19656), .B1(
        n19649), .B2(n19962), .ZN(n19647) );
  OAI211_X1 U22614 ( .C1(n19965), .C2(n19693), .A(n19648), .B(n19647), .ZN(
        P2_U3108) );
  AOI22_X1 U22615 ( .A1(n19654), .A2(n19967), .B1(n19665), .B2(n19966), .ZN(
        n19651) );
  AOI22_X1 U22616 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19656), .B1(
        n19649), .B2(n19968), .ZN(n19650) );
  OAI211_X1 U22617 ( .C1(n19971), .C2(n19693), .A(n19651), .B(n19650), .ZN(
        P2_U3109) );
  AOI22_X1 U22618 ( .A1(n19654), .A2(n19973), .B1(n19665), .B2(n19972), .ZN(
        n19653) );
  AOI22_X1 U22619 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19656), .B1(
        n19673), .B2(n19974), .ZN(n19652) );
  OAI211_X1 U22620 ( .C1(n19979), .C2(n19659), .A(n19653), .B(n19652), .ZN(
        P2_U3110) );
  AOI22_X1 U22621 ( .A1(n19654), .A2(n19982), .B1(n19665), .B2(n19980), .ZN(
        n19658) );
  AOI22_X1 U22622 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19656), .B1(
        n19673), .B2(n19655), .ZN(n19657) );
  OAI211_X1 U22623 ( .C1(n19916), .C2(n19659), .A(n19658), .B(n19657), .ZN(
        P2_U3111) );
  NAND2_X1 U22624 ( .A1(n20088), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19769) );
  NOR2_X1 U22625 ( .A1(n19769), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19703) );
  INV_X1 U22626 ( .A(n19703), .ZN(n19706) );
  NOR2_X1 U22627 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19706), .ZN(
        n19672) );
  INV_X1 U22628 ( .A(n19672), .ZN(n19692) );
  OAI22_X1 U22629 ( .A1(n19779), .A2(n19726), .B1(n19869), .B2(n19692), .ZN(
        n19660) );
  INV_X1 U22630 ( .A(n19660), .ZN(n19671) );
  OAI21_X1 U22631 ( .B1(n19673), .B2(n19722), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19661) );
  NAND2_X1 U22632 ( .A1(n19661), .A2(n20069), .ZN(n19669) );
  NOR2_X1 U22633 ( .A1(n19669), .A2(n19665), .ZN(n19662) );
  AOI211_X1 U22634 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19663), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19662), .ZN(n19664) );
  NOR2_X1 U22635 ( .A1(n19665), .A2(n19672), .ZN(n19668) );
  OAI21_X1 U22636 ( .B1(n19666), .B2(n19672), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19667) );
  AOI22_X1 U22637 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19696), .B1(
        n19929), .B2(n19695), .ZN(n19670) );
  OAI211_X1 U22638 ( .C1(n19941), .C2(n19693), .A(n19671), .B(n19670), .ZN(
        P2_U3112) );
  AOI22_X1 U22639 ( .A1(n19673), .A2(n19944), .B1(n19942), .B2(n19672), .ZN(
        n19675) );
  AOI22_X1 U22640 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19696), .B1(
        n19695), .B2(n19943), .ZN(n19674) );
  OAI211_X1 U22641 ( .C1(n19947), .C2(n19726), .A(n19675), .B(n19674), .ZN(
        P2_U3113) );
  OAI22_X1 U22642 ( .A1(n19693), .A2(n19883), .B1(n19882), .B2(n19692), .ZN(
        n19676) );
  INV_X1 U22643 ( .A(n19676), .ZN(n19678) );
  AOI22_X1 U22644 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19696), .B1(
        n19695), .B2(n19949), .ZN(n19677) );
  OAI211_X1 U22645 ( .C1(n19953), .C2(n19726), .A(n19678), .B(n19677), .ZN(
        P2_U3114) );
  OAI22_X1 U22646 ( .A1(n19726), .A2(n19890), .B1(n19692), .B2(n19889), .ZN(
        n19679) );
  INV_X1 U22647 ( .A(n19679), .ZN(n19681) );
  AOI22_X1 U22648 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19696), .B1(
        n19695), .B2(n19955), .ZN(n19680) );
  OAI211_X1 U22649 ( .C1(n19959), .C2(n19693), .A(n19681), .B(n19680), .ZN(
        P2_U3115) );
  OAI22_X1 U22650 ( .A1(n19965), .A2(n19726), .B1(n19895), .B2(n19692), .ZN(
        n19682) );
  INV_X1 U22651 ( .A(n19682), .ZN(n19684) );
  AOI22_X1 U22652 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19696), .B1(
        n19695), .B2(n19961), .ZN(n19683) );
  OAI211_X1 U22653 ( .C1(n19896), .C2(n19693), .A(n19684), .B(n19683), .ZN(
        P2_U3116) );
  OAI22_X1 U22654 ( .A1(n19693), .A2(n19903), .B1(n19902), .B2(n19692), .ZN(
        n19685) );
  INV_X1 U22655 ( .A(n19685), .ZN(n19687) );
  AOI22_X1 U22656 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19696), .B1(
        n19695), .B2(n19967), .ZN(n19686) );
  OAI211_X1 U22657 ( .C1(n19971), .C2(n19726), .A(n19687), .B(n19686), .ZN(
        P2_U3117) );
  OAI22_X1 U22658 ( .A1(n19913), .A2(n19726), .B1(n19688), .B2(n19692), .ZN(
        n19689) );
  INV_X1 U22659 ( .A(n19689), .ZN(n19691) );
  AOI22_X1 U22660 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19696), .B1(
        n19695), .B2(n19973), .ZN(n19690) );
  OAI211_X1 U22661 ( .C1(n19979), .C2(n19693), .A(n19691), .B(n19690), .ZN(
        P2_U3118) );
  OAI22_X1 U22662 ( .A1(n19693), .A2(n19916), .B1(n19915), .B2(n19692), .ZN(
        n19694) );
  INV_X1 U22663 ( .A(n19694), .ZN(n19698) );
  AOI22_X1 U22664 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19696), .B1(
        n19695), .B2(n19982), .ZN(n19697) );
  OAI211_X1 U22665 ( .C1(n19990), .C2(n19726), .A(n19698), .B(n19697), .ZN(
        P2_U3119) );
  NOR2_X1 U22666 ( .A1(n19699), .A2(n19769), .ZN(n19732) );
  AOI22_X1 U22667 ( .A1(n19938), .A2(n19761), .B1(n19732), .B2(n19928), .ZN(
        n19709) );
  NAND2_X1 U22668 ( .A1(n20074), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19932) );
  OAI21_X1 U22669 ( .B1(n19932), .B2(n19700), .A(n20069), .ZN(n19707) );
  INV_X1 U22670 ( .A(n19732), .ZN(n19725) );
  OAI211_X1 U22671 ( .C1(n19701), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19860), 
        .B(n19725), .ZN(n19702) );
  OAI211_X1 U22672 ( .C1(n19707), .C2(n19703), .A(n19936), .B(n19702), .ZN(
        n19729) );
  OAI21_X1 U22673 ( .B1(n19704), .B2(n19732), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19705) );
  OAI21_X1 U22674 ( .B1(n19707), .B2(n19706), .A(n19705), .ZN(n19728) );
  AOI22_X1 U22675 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19729), .B1(
        n19929), .B2(n19728), .ZN(n19708) );
  OAI211_X1 U22676 ( .C1(n19941), .C2(n19726), .A(n19709), .B(n19708), .ZN(
        P2_U3120) );
  AOI22_X1 U22677 ( .A1(n19722), .A2(n19944), .B1(n19942), .B2(n19732), .ZN(
        n19711) );
  AOI22_X1 U22678 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19729), .B1(
        n19943), .B2(n19728), .ZN(n19710) );
  OAI211_X1 U22679 ( .C1(n19947), .C2(n19758), .A(n19711), .B(n19710), .ZN(
        P2_U3121) );
  AOI22_X1 U22680 ( .A1(n19885), .A2(n19761), .B1(n19948), .B2(n19732), .ZN(
        n19713) );
  AOI22_X1 U22681 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19729), .B1(
        n19949), .B2(n19728), .ZN(n19712) );
  OAI211_X1 U22682 ( .C1(n19883), .C2(n19726), .A(n19713), .B(n19712), .ZN(
        P2_U3122) );
  AOI22_X1 U22683 ( .A1(n19722), .A2(n19892), .B1(n19954), .B2(n19732), .ZN(
        n19715) );
  AOI22_X1 U22684 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19729), .B1(
        n19955), .B2(n19728), .ZN(n19714) );
  OAI211_X1 U22685 ( .C1(n19890), .C2(n19758), .A(n19715), .B(n19714), .ZN(
        P2_U3123) );
  OAI22_X1 U22686 ( .A1(n19726), .A2(n19896), .B1(n19895), .B2(n19725), .ZN(
        n19716) );
  INV_X1 U22687 ( .A(n19716), .ZN(n19718) );
  AOI22_X1 U22688 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19729), .B1(
        n19961), .B2(n19728), .ZN(n19717) );
  OAI211_X1 U22689 ( .C1(n19965), .C2(n19758), .A(n19718), .B(n19717), .ZN(
        P2_U3124) );
  OAI22_X1 U22690 ( .A1(n19726), .A2(n19903), .B1(n19902), .B2(n19725), .ZN(
        n19719) );
  INV_X1 U22691 ( .A(n19719), .ZN(n19721) );
  AOI22_X1 U22692 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19729), .B1(
        n19967), .B2(n19728), .ZN(n19720) );
  OAI211_X1 U22693 ( .C1(n19971), .C2(n19758), .A(n19721), .B(n19720), .ZN(
        P2_U3125) );
  AOI22_X1 U22694 ( .A1(n19722), .A2(n19909), .B1(n19972), .B2(n19732), .ZN(
        n19724) );
  AOI22_X1 U22695 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19729), .B1(
        n19973), .B2(n19728), .ZN(n19723) );
  OAI211_X1 U22696 ( .C1(n19913), .C2(n19758), .A(n19724), .B(n19723), .ZN(
        P2_U3126) );
  OAI22_X1 U22697 ( .A1(n19726), .A2(n19916), .B1(n19915), .B2(n19725), .ZN(
        n19727) );
  INV_X1 U22698 ( .A(n19727), .ZN(n19731) );
  AOI22_X1 U22699 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19729), .B1(
        n19982), .B2(n19728), .ZN(n19730) );
  OAI211_X1 U22700 ( .C1(n19990), .C2(n19758), .A(n19731), .B(n19730), .ZN(
        P2_U3127) );
  AOI221_X1 U22701 ( .B1(n19795), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19761), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19732), .ZN(n19733) );
  OR2_X1 U22702 ( .A1(n19733), .A2(n19860), .ZN(n19737) );
  NOR2_X1 U22703 ( .A1(n19926), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19735) );
  NOR2_X1 U22704 ( .A1(n19734), .A2(n19769), .ZN(n19759) );
  AOI21_X1 U22705 ( .B1(n19739), .B2(n19735), .A(n19759), .ZN(n19736) );
  NAND2_X1 U22706 ( .A1(n19737), .A2(n19736), .ZN(n19738) );
  AND2_X1 U22707 ( .A1(n19738), .A2(n19936), .ZN(n19747) );
  OAI21_X1 U22708 ( .B1(n19739), .B2(n19759), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19740) );
  OAI21_X1 U22709 ( .B1(n19769), .B2(n19741), .A(n19740), .ZN(n19760) );
  AOI22_X1 U22710 ( .A1(n19760), .A2(n19929), .B1(n19928), .B2(n19759), .ZN(
        n19743) );
  AOI22_X1 U22711 ( .A1(n19795), .A2(n19938), .B1(n19761), .B2(n19776), .ZN(
        n19742) );
  OAI211_X1 U22712 ( .C1(n19747), .C2(n19744), .A(n19743), .B(n19742), .ZN(
        P2_U3128) );
  AOI22_X1 U22713 ( .A1(n19760), .A2(n19943), .B1(n19942), .B2(n19759), .ZN(
        n19746) );
  AOI22_X1 U22714 ( .A1(n19761), .A2(n19944), .B1(n19795), .B2(n19878), .ZN(
        n19745) );
  OAI211_X1 U22715 ( .C1(n19747), .C2(n12451), .A(n19746), .B(n19745), .ZN(
        P2_U3129) );
  AOI22_X1 U22716 ( .A1(n19760), .A2(n19949), .B1(n19948), .B2(n19759), .ZN(
        n19749) );
  AOI22_X1 U22717 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19762), .B1(
        n19761), .B2(n19950), .ZN(n19748) );
  OAI211_X1 U22718 ( .C1(n19953), .C2(n19790), .A(n19749), .B(n19748), .ZN(
        P2_U3130) );
  AOI22_X1 U22719 ( .A1(n19760), .A2(n19955), .B1(n19954), .B2(n19759), .ZN(
        n19751) );
  AOI22_X1 U22720 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19762), .B1(
        n19795), .B2(n19956), .ZN(n19750) );
  OAI211_X1 U22721 ( .C1(n19959), .C2(n19758), .A(n19751), .B(n19750), .ZN(
        P2_U3131) );
  AOI22_X1 U22722 ( .A1(n19760), .A2(n19961), .B1(n19960), .B2(n19759), .ZN(
        n19753) );
  AOI22_X1 U22723 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19762), .B1(
        n19795), .B2(n19898), .ZN(n19752) );
  OAI211_X1 U22724 ( .C1(n19896), .C2(n19758), .A(n19753), .B(n19752), .ZN(
        P2_U3132) );
  AOI22_X1 U22725 ( .A1(n19760), .A2(n19967), .B1(n19966), .B2(n19759), .ZN(
        n19755) );
  AOI22_X1 U22726 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19762), .B1(
        n19761), .B2(n19968), .ZN(n19754) );
  OAI211_X1 U22727 ( .C1(n19971), .C2(n19790), .A(n19755), .B(n19754), .ZN(
        P2_U3133) );
  AOI22_X1 U22728 ( .A1(n19760), .A2(n19973), .B1(n19972), .B2(n19759), .ZN(
        n19757) );
  AOI22_X1 U22729 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19762), .B1(
        n19795), .B2(n19974), .ZN(n19756) );
  OAI211_X1 U22730 ( .C1(n19979), .C2(n19758), .A(n19757), .B(n19756), .ZN(
        P2_U3134) );
  AOI22_X1 U22731 ( .A1(n19760), .A2(n19982), .B1(n19980), .B2(n19759), .ZN(
        n19764) );
  AOI22_X1 U22732 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19762), .B1(
        n19761), .B2(n19984), .ZN(n19763) );
  OAI211_X1 U22733 ( .C1(n19990), .C2(n19790), .A(n19764), .B(n19763), .ZN(
        P2_U3135) );
  INV_X1 U22734 ( .A(n19765), .ZN(n19767) );
  INV_X1 U22735 ( .A(n19769), .ZN(n19766) );
  NAND2_X1 U22736 ( .A1(n19767), .A2(n19766), .ZN(n19772) );
  AND2_X1 U22737 ( .A1(n19772), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19768) );
  NAND2_X1 U22738 ( .A1(n10650), .A2(n19768), .ZN(n19774) );
  OR2_X1 U22739 ( .A1(n20098), .A2(n19769), .ZN(n19771) );
  OAI21_X1 U22740 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19771), .A(n19926), 
        .ZN(n19770) );
  INV_X1 U22741 ( .A(n19772), .ZN(n19793) );
  AOI22_X1 U22742 ( .A1(n19794), .A2(n19929), .B1(n19928), .B2(n19793), .ZN(
        n19778) );
  OAI21_X1 U22743 ( .B1(n19932), .B2(n20071), .A(n19771), .ZN(n19775) );
  NAND2_X1 U22744 ( .A1(n19772), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19773) );
  NAND4_X1 U22745 ( .A1(n19775), .A2(n19936), .A3(n19774), .A4(n19773), .ZN(
        n19796) );
  AOI22_X1 U22746 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19796), .B1(
        n19795), .B2(n19776), .ZN(n19777) );
  OAI211_X1 U22747 ( .C1(n19779), .C2(n19818), .A(n19778), .B(n19777), .ZN(
        P2_U3136) );
  AOI22_X1 U22748 ( .A1(n19794), .A2(n19943), .B1(n19942), .B2(n19793), .ZN(
        n19781) );
  AOI22_X1 U22749 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19796), .B1(
        n19795), .B2(n19944), .ZN(n19780) );
  OAI211_X1 U22750 ( .C1(n19947), .C2(n19818), .A(n19781), .B(n19780), .ZN(
        P2_U3137) );
  AOI22_X1 U22751 ( .A1(n19794), .A2(n19949), .B1(n19948), .B2(n19793), .ZN(
        n19783) );
  AOI22_X1 U22752 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19796), .B1(
        n19825), .B2(n19885), .ZN(n19782) );
  OAI211_X1 U22753 ( .C1(n19883), .C2(n19790), .A(n19783), .B(n19782), .ZN(
        P2_U3138) );
  AOI22_X1 U22754 ( .A1(n19794), .A2(n19955), .B1(n19954), .B2(n19793), .ZN(
        n19785) );
  AOI22_X1 U22755 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19796), .B1(
        n19795), .B2(n19892), .ZN(n19784) );
  OAI211_X1 U22756 ( .C1(n19890), .C2(n19818), .A(n19785), .B(n19784), .ZN(
        P2_U3139) );
  AOI22_X1 U22757 ( .A1(n19794), .A2(n19961), .B1(n19960), .B2(n19793), .ZN(
        n19787) );
  AOI22_X1 U22758 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19796), .B1(
        n19825), .B2(n19898), .ZN(n19786) );
  OAI211_X1 U22759 ( .C1(n19896), .C2(n19790), .A(n19787), .B(n19786), .ZN(
        P2_U3140) );
  AOI22_X1 U22760 ( .A1(n19794), .A2(n19967), .B1(n19966), .B2(n19793), .ZN(
        n19789) );
  AOI22_X1 U22761 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19796), .B1(
        n19825), .B2(n19848), .ZN(n19788) );
  OAI211_X1 U22762 ( .C1(n19903), .C2(n19790), .A(n19789), .B(n19788), .ZN(
        P2_U3141) );
  AOI22_X1 U22763 ( .A1(n19794), .A2(n19973), .B1(n19972), .B2(n19793), .ZN(
        n19792) );
  AOI22_X1 U22764 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19796), .B1(
        n19795), .B2(n19909), .ZN(n19791) );
  OAI211_X1 U22765 ( .C1(n19913), .C2(n19818), .A(n19792), .B(n19791), .ZN(
        P2_U3142) );
  AOI22_X1 U22766 ( .A1(n19794), .A2(n19982), .B1(n19980), .B2(n19793), .ZN(
        n19798) );
  AOI22_X1 U22767 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19796), .B1(
        n19795), .B2(n19984), .ZN(n19797) );
  OAI211_X1 U22768 ( .C1(n19990), .C2(n19818), .A(n19798), .B(n19797), .ZN(
        P2_U3143) );
  INV_X1 U22769 ( .A(n19799), .ZN(n19802) );
  NAND3_X1 U22770 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20098), .ZN(n19831) );
  NOR2_X1 U22771 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19831), .ZN(
        n19823) );
  OAI21_X1 U22772 ( .B1(n19800), .B2(n19823), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19801) );
  OAI21_X1 U22773 ( .B1(n19802), .B2(n19805), .A(n19801), .ZN(n19824) );
  AOI22_X1 U22774 ( .A1(n19824), .A2(n19929), .B1(n19928), .B2(n19823), .ZN(
        n19809) );
  AOI21_X1 U22775 ( .B1(n19803), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19807) );
  OAI21_X1 U22776 ( .B1(n19825), .B2(n19855), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19804) );
  OAI21_X1 U22777 ( .B1(n19805), .B2(n20081), .A(n19804), .ZN(n19806) );
  OAI211_X1 U22778 ( .C1(n19823), .C2(n19807), .A(n19806), .B(n19936), .ZN(
        n19826) );
  AOI22_X1 U22779 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19826), .B1(
        n19855), .B2(n19938), .ZN(n19808) );
  OAI211_X1 U22780 ( .C1(n19941), .C2(n19818), .A(n19809), .B(n19808), .ZN(
        P2_U3144) );
  AOI22_X1 U22781 ( .A1(n19824), .A2(n19943), .B1(n19942), .B2(n19823), .ZN(
        n19811) );
  AOI22_X1 U22782 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19826), .B1(
        n19825), .B2(n19944), .ZN(n19810) );
  OAI211_X1 U22783 ( .C1(n19947), .C2(n19851), .A(n19811), .B(n19810), .ZN(
        P2_U3145) );
  AOI22_X1 U22784 ( .A1(n19824), .A2(n19949), .B1(n19948), .B2(n19823), .ZN(
        n19813) );
  AOI22_X1 U22785 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19826), .B1(
        n19855), .B2(n19885), .ZN(n19812) );
  OAI211_X1 U22786 ( .C1(n19883), .C2(n19818), .A(n19813), .B(n19812), .ZN(
        P2_U3146) );
  AOI22_X1 U22787 ( .A1(n19824), .A2(n19955), .B1(n19954), .B2(n19823), .ZN(
        n19815) );
  AOI22_X1 U22788 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19826), .B1(
        n19825), .B2(n19892), .ZN(n19814) );
  OAI211_X1 U22789 ( .C1(n19890), .C2(n19851), .A(n19815), .B(n19814), .ZN(
        P2_U3147) );
  AOI22_X1 U22790 ( .A1(n19824), .A2(n19961), .B1(n19960), .B2(n19823), .ZN(
        n19817) );
  AOI22_X1 U22791 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19826), .B1(
        n19855), .B2(n19898), .ZN(n19816) );
  OAI211_X1 U22792 ( .C1(n19896), .C2(n19818), .A(n19817), .B(n19816), .ZN(
        P2_U3148) );
  AOI22_X1 U22793 ( .A1(n19824), .A2(n19967), .B1(n19966), .B2(n19823), .ZN(
        n19820) );
  AOI22_X1 U22794 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19826), .B1(
        n19825), .B2(n19968), .ZN(n19819) );
  OAI211_X1 U22795 ( .C1(n19971), .C2(n19851), .A(n19820), .B(n19819), .ZN(
        P2_U3149) );
  AOI22_X1 U22796 ( .A1(n19824), .A2(n19973), .B1(n19972), .B2(n19823), .ZN(
        n19822) );
  AOI22_X1 U22797 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19826), .B1(
        n19825), .B2(n19909), .ZN(n19821) );
  OAI211_X1 U22798 ( .C1(n19913), .C2(n19851), .A(n19822), .B(n19821), .ZN(
        P2_U3150) );
  AOI22_X1 U22799 ( .A1(n19824), .A2(n19982), .B1(n19980), .B2(n19823), .ZN(
        n19828) );
  AOI22_X1 U22800 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19826), .B1(
        n19825), .B2(n19984), .ZN(n19827) );
  OAI211_X1 U22801 ( .C1(n19990), .C2(n19851), .A(n19828), .B(n19827), .ZN(
        P2_U3151) );
  NOR2_X1 U22802 ( .A1(n20106), .A2(n19831), .ZN(n19862) );
  OAI21_X1 U22803 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19831), .A(n19926), 
        .ZN(n19830) );
  AND2_X1 U22804 ( .A1(n19834), .A2(n19830), .ZN(n19854) );
  AOI22_X1 U22805 ( .A1(n19854), .A2(n19929), .B1(n19928), .B2(n19862), .ZN(
        n19839) );
  OAI21_X1 U22806 ( .B1(n19932), .B2(n19836), .A(n19831), .ZN(n19835) );
  INV_X1 U22807 ( .A(n19862), .ZN(n19832) );
  NAND2_X1 U22808 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19832), .ZN(n19833) );
  NAND4_X1 U22809 ( .A1(n19835), .A2(n19936), .A3(n19834), .A4(n19833), .ZN(
        n19856) );
  AOI22_X1 U22810 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19856), .B1(
        n19910), .B2(n19938), .ZN(n19838) );
  OAI211_X1 U22811 ( .C1(n19941), .C2(n19851), .A(n19839), .B(n19838), .ZN(
        P2_U3152) );
  AOI22_X1 U22812 ( .A1(n19854), .A2(n19943), .B1(n19942), .B2(n19862), .ZN(
        n19841) );
  AOI22_X1 U22813 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19856), .B1(
        n19855), .B2(n19944), .ZN(n19840) );
  OAI211_X1 U22814 ( .C1(n19947), .C2(n19917), .A(n19841), .B(n19840), .ZN(
        P2_U3153) );
  AOI22_X1 U22815 ( .A1(n19854), .A2(n19949), .B1(n19948), .B2(n19862), .ZN(
        n19843) );
  AOI22_X1 U22816 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19856), .B1(
        n19910), .B2(n19885), .ZN(n19842) );
  OAI211_X1 U22817 ( .C1(n19883), .C2(n19851), .A(n19843), .B(n19842), .ZN(
        P2_U3154) );
  AOI22_X1 U22818 ( .A1(n19854), .A2(n19955), .B1(n19954), .B2(n19862), .ZN(
        n19845) );
  AOI22_X1 U22819 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19856), .B1(
        n19855), .B2(n19892), .ZN(n19844) );
  OAI211_X1 U22820 ( .C1(n19890), .C2(n19917), .A(n19845), .B(n19844), .ZN(
        P2_U3155) );
  AOI22_X1 U22821 ( .A1(n19854), .A2(n19961), .B1(n19960), .B2(n19862), .ZN(
        n19847) );
  AOI22_X1 U22822 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19856), .B1(
        n19855), .B2(n19962), .ZN(n19846) );
  OAI211_X1 U22823 ( .C1(n19965), .C2(n19917), .A(n19847), .B(n19846), .ZN(
        P2_U3156) );
  AOI22_X1 U22824 ( .A1(n19854), .A2(n19967), .B1(n19966), .B2(n19862), .ZN(
        n19850) );
  AOI22_X1 U22825 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19856), .B1(
        n19910), .B2(n19848), .ZN(n19849) );
  OAI211_X1 U22826 ( .C1(n19903), .C2(n19851), .A(n19850), .B(n19849), .ZN(
        P2_U3157) );
  AOI22_X1 U22827 ( .A1(n19854), .A2(n19973), .B1(n19972), .B2(n19862), .ZN(
        n19853) );
  AOI22_X1 U22828 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19856), .B1(
        n19855), .B2(n19909), .ZN(n19852) );
  OAI211_X1 U22829 ( .C1(n19913), .C2(n19917), .A(n19853), .B(n19852), .ZN(
        P2_U3158) );
  AOI22_X1 U22830 ( .A1(n19854), .A2(n19982), .B1(n19980), .B2(n19862), .ZN(
        n19858) );
  AOI22_X1 U22831 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19856), .B1(
        n19855), .B2(n19984), .ZN(n19857) );
  OAI211_X1 U22832 ( .C1(n19990), .C2(n19917), .A(n19858), .B(n19857), .ZN(
        P2_U3159) );
  NAND2_X1 U22833 ( .A1(n19978), .A2(n19917), .ZN(n19861) );
  AOI21_X1 U22834 ( .B1(n19861), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19860), 
        .ZN(n19871) );
  NOR3_X1 U22835 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20081), .A3(
        n19925), .ZN(n19908) );
  NOR2_X1 U22836 ( .A1(n19908), .A2(n19862), .ZN(n19873) );
  NAND2_X1 U22837 ( .A1(n19871), .A2(n19873), .ZN(n19868) );
  NAND2_X1 U22838 ( .A1(n19863), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19864) );
  NAND2_X1 U22839 ( .A1(n19864), .A2(n13484), .ZN(n19866) );
  INV_X1 U22840 ( .A(n19908), .ZN(n19914) );
  AOI21_X1 U22841 ( .B1(n19866), .B2(n19914), .A(n19865), .ZN(n19867) );
  INV_X1 U22842 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n19877) );
  OAI22_X1 U22843 ( .A1(n19917), .A2(n19941), .B1(n19869), .B2(n19914), .ZN(
        n19870) );
  INV_X1 U22844 ( .A(n19870), .ZN(n19876) );
  INV_X1 U22845 ( .A(n19871), .ZN(n19874) );
  OAI21_X1 U22846 ( .B1(n10511), .B2(n19908), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19872) );
  AOI22_X1 U22847 ( .A1(n19929), .A2(n19919), .B1(n19985), .B2(n19938), .ZN(
        n19875) );
  OAI211_X1 U22848 ( .C1(n19905), .C2(n19877), .A(n19876), .B(n19875), .ZN(
        P2_U3160) );
  INV_X1 U22849 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n19881) );
  AOI22_X1 U22850 ( .A1(n19910), .A2(n19944), .B1(n19942), .B2(n19908), .ZN(
        n19880) );
  AOI22_X1 U22851 ( .A1(n19943), .A2(n19919), .B1(n19985), .B2(n19878), .ZN(
        n19879) );
  OAI211_X1 U22852 ( .C1(n19905), .C2(n19881), .A(n19880), .B(n19879), .ZN(
        P2_U3161) );
  OAI22_X1 U22853 ( .A1(n19917), .A2(n19883), .B1(n19882), .B2(n19914), .ZN(
        n19884) );
  INV_X1 U22854 ( .A(n19884), .ZN(n19887) );
  AOI22_X1 U22855 ( .A1(n19949), .A2(n19919), .B1(n19985), .B2(n19885), .ZN(
        n19886) );
  OAI211_X1 U22856 ( .C1(n19905), .C2(n19888), .A(n19887), .B(n19886), .ZN(
        P2_U3162) );
  OAI22_X1 U22857 ( .A1(n19978), .A2(n19890), .B1(n19914), .B2(n19889), .ZN(
        n19891) );
  INV_X1 U22858 ( .A(n19891), .ZN(n19894) );
  AOI22_X1 U22859 ( .A1(n19955), .A2(n19919), .B1(n19910), .B2(n19892), .ZN(
        n19893) );
  OAI211_X1 U22860 ( .C1(n19905), .C2(n10471), .A(n19894), .B(n19893), .ZN(
        P2_U3163) );
  INV_X1 U22861 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n19901) );
  OAI22_X1 U22862 ( .A1(n19917), .A2(n19896), .B1(n19895), .B2(n19914), .ZN(
        n19897) );
  INV_X1 U22863 ( .A(n19897), .ZN(n19900) );
  AOI22_X1 U22864 ( .A1(n19961), .A2(n19919), .B1(n19985), .B2(n19898), .ZN(
        n19899) );
  OAI211_X1 U22865 ( .C1(n19905), .C2(n19901), .A(n19900), .B(n19899), .ZN(
        P2_U3164) );
  OAI22_X1 U22866 ( .A1(n19917), .A2(n19903), .B1(n19902), .B2(n19914), .ZN(
        n19904) );
  INV_X1 U22867 ( .A(n19904), .ZN(n19907) );
  INV_X1 U22868 ( .A(n19905), .ZN(n19920) );
  AOI22_X1 U22869 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19920), .B1(
        n19967), .B2(n19919), .ZN(n19906) );
  OAI211_X1 U22870 ( .C1(n19971), .C2(n19978), .A(n19907), .B(n19906), .ZN(
        P2_U3165) );
  AOI22_X1 U22871 ( .A1(n19910), .A2(n19909), .B1(n19972), .B2(n19908), .ZN(
        n19912) );
  AOI22_X1 U22872 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19920), .B1(
        n19973), .B2(n19919), .ZN(n19911) );
  OAI211_X1 U22873 ( .C1(n19913), .C2(n19978), .A(n19912), .B(n19911), .ZN(
        P2_U3166) );
  OAI22_X1 U22874 ( .A1(n19917), .A2(n19916), .B1(n19915), .B2(n19914), .ZN(
        n19918) );
  INV_X1 U22875 ( .A(n19918), .ZN(n19922) );
  AOI22_X1 U22876 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19920), .B1(
        n19982), .B2(n19919), .ZN(n19921) );
  OAI211_X1 U22877 ( .C1(n19990), .C2(n19978), .A(n19922), .B(n19921), .ZN(
        P2_U3167) );
  AND2_X1 U22878 ( .A1(n19933), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19923) );
  NAND2_X1 U22879 ( .A1(n19924), .A2(n19923), .ZN(n19935) );
  OR2_X1 U22880 ( .A1(n20081), .A2(n19925), .ZN(n19930) );
  OAI21_X1 U22881 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19930), .A(n19926), 
        .ZN(n19927) );
  AND2_X1 U22882 ( .A1(n19935), .A2(n19927), .ZN(n19983) );
  INV_X1 U22883 ( .A(n19933), .ZN(n19981) );
  AOI22_X1 U22884 ( .A1(n19983), .A2(n19929), .B1(n19981), .B2(n19928), .ZN(
        n19940) );
  OAI21_X1 U22885 ( .B1(n19932), .B2(n19931), .A(n19930), .ZN(n19937) );
  NAND2_X1 U22886 ( .A1(n19933), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19934) );
  NAND4_X1 U22887 ( .A1(n19937), .A2(n19936), .A3(n19935), .A4(n19934), .ZN(
        n19986) );
  AOI22_X1 U22888 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19986), .B1(
        n19975), .B2(n19938), .ZN(n19939) );
  OAI211_X1 U22889 ( .C1(n19941), .C2(n19978), .A(n19940), .B(n19939), .ZN(
        P2_U3168) );
  AOI22_X1 U22890 ( .A1(n19983), .A2(n19943), .B1(n19981), .B2(n19942), .ZN(
        n19946) );
  AOI22_X1 U22891 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19986), .B1(
        n19985), .B2(n19944), .ZN(n19945) );
  OAI211_X1 U22892 ( .C1(n19947), .C2(n19989), .A(n19946), .B(n19945), .ZN(
        P2_U3169) );
  AOI22_X1 U22893 ( .A1(n19983), .A2(n19949), .B1(n19981), .B2(n19948), .ZN(
        n19952) );
  AOI22_X1 U22894 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19986), .B1(
        n19985), .B2(n19950), .ZN(n19951) );
  OAI211_X1 U22895 ( .C1(n19953), .C2(n19989), .A(n19952), .B(n19951), .ZN(
        P2_U3170) );
  AOI22_X1 U22896 ( .A1(n19983), .A2(n19955), .B1(n19981), .B2(n19954), .ZN(
        n19958) );
  AOI22_X1 U22897 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19986), .B1(
        n19975), .B2(n19956), .ZN(n19957) );
  OAI211_X1 U22898 ( .C1(n19959), .C2(n19978), .A(n19958), .B(n19957), .ZN(
        P2_U3171) );
  AOI22_X1 U22899 ( .A1(n19983), .A2(n19961), .B1(n19981), .B2(n19960), .ZN(
        n19964) );
  AOI22_X1 U22900 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19986), .B1(
        n19985), .B2(n19962), .ZN(n19963) );
  OAI211_X1 U22901 ( .C1(n19965), .C2(n19989), .A(n19964), .B(n19963), .ZN(
        P2_U3172) );
  AOI22_X1 U22902 ( .A1(n19983), .A2(n19967), .B1(n19981), .B2(n19966), .ZN(
        n19970) );
  AOI22_X1 U22903 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19986), .B1(
        n19985), .B2(n19968), .ZN(n19969) );
  OAI211_X1 U22904 ( .C1(n19971), .C2(n19989), .A(n19970), .B(n19969), .ZN(
        P2_U3173) );
  AOI22_X1 U22905 ( .A1(n19983), .A2(n19973), .B1(n19981), .B2(n19972), .ZN(
        n19977) );
  AOI22_X1 U22906 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19986), .B1(
        n19975), .B2(n19974), .ZN(n19976) );
  OAI211_X1 U22907 ( .C1(n19979), .C2(n19978), .A(n19977), .B(n19976), .ZN(
        P2_U3174) );
  AOI22_X1 U22908 ( .A1(n19983), .A2(n19982), .B1(n19981), .B2(n19980), .ZN(
        n19988) );
  AOI22_X1 U22909 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19986), .B1(
        n19985), .B2(n19984), .ZN(n19987) );
  OAI211_X1 U22910 ( .C1(n19990), .C2(n19989), .A(n19988), .B(n19987), .ZN(
        P2_U3175) );
  AND2_X1 U22911 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19991), .ZN(
        P2_U3179) );
  AND2_X1 U22912 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19991), .ZN(
        P2_U3180) );
  AND2_X1 U22913 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19991), .ZN(
        P2_U3181) );
  AND2_X1 U22914 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19991), .ZN(
        P2_U3182) );
  AND2_X1 U22915 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19991), .ZN(
        P2_U3183) );
  AND2_X1 U22916 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19991), .ZN(
        P2_U3184) );
  AND2_X1 U22917 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19991), .ZN(
        P2_U3185) );
  AND2_X1 U22918 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19991), .ZN(
        P2_U3186) );
  AND2_X1 U22919 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19991), .ZN(
        P2_U3187) );
  AND2_X1 U22920 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19991), .ZN(
        P2_U3188) );
  AND2_X1 U22921 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19991), .ZN(
        P2_U3189) );
  AND2_X1 U22922 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19991), .ZN(
        P2_U3190) );
  AND2_X1 U22923 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19991), .ZN(
        P2_U3191) );
  AND2_X1 U22924 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19991), .ZN(
        P2_U3192) );
  AND2_X1 U22925 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19991), .ZN(
        P2_U3193) );
  AND2_X1 U22926 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19991), .ZN(
        P2_U3194) );
  AND2_X1 U22927 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19991), .ZN(
        P2_U3195) );
  AND2_X1 U22928 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19991), .ZN(
        P2_U3196) );
  AND2_X1 U22929 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19991), .ZN(
        P2_U3197) );
  AND2_X1 U22930 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19991), .ZN(
        P2_U3198) );
  AND2_X1 U22931 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19991), .ZN(
        P2_U3199) );
  AND2_X1 U22932 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19991), .ZN(
        P2_U3200) );
  AND2_X1 U22933 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19991), .ZN(P2_U3201) );
  AND2_X1 U22934 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19991), .ZN(P2_U3202) );
  AND2_X1 U22935 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19991), .ZN(P2_U3203) );
  AND2_X1 U22936 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19991), .ZN(P2_U3204) );
  AND2_X1 U22937 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19991), .ZN(P2_U3205) );
  AND2_X1 U22938 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19991), .ZN(P2_U3206) );
  AND2_X1 U22939 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19991), .ZN(P2_U3207) );
  AND2_X1 U22940 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19991), .ZN(P2_U3208) );
  NAND2_X1 U22941 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20003), .ZN(n20005) );
  NAND3_X1 U22942 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n20005), .ZN(n19993) );
  AOI211_X1 U22943 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n21115), .A(
        n20004), .B(n20108), .ZN(n19992) );
  NOR2_X1 U22944 ( .A1(n20898), .A2(n19997), .ZN(n20010) );
  AOI211_X1 U22945 ( .C1(n20011), .C2(n19993), .A(n19992), .B(n20010), .ZN(
        n19994) );
  INV_X1 U22946 ( .A(n19994), .ZN(P2_U3209) );
  INV_X1 U22947 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19995) );
  AOI21_X1 U22948 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21115), .A(n20011), 
        .ZN(n20001) );
  NOR2_X1 U22949 ( .A1(n19995), .A2(n20001), .ZN(n19998) );
  AOI21_X1 U22950 ( .B1(n19998), .B2(n19997), .A(n19996), .ZN(n19999) );
  OAI211_X1 U22951 ( .C1(n21115), .C2(n20000), .A(n19999), .B(n20005), .ZN(
        P2_U3210) );
  AOI21_X1 U22952 ( .B1(n20003), .B2(n20002), .A(n20001), .ZN(n20009) );
  INV_X1 U22953 ( .A(n20004), .ZN(n20006) );
  OAI22_X1 U22954 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n20006), .B1(NA), 
        .B2(n20005), .ZN(n20007) );
  OAI211_X1 U22955 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n20007), .ZN(n20008) );
  OAI21_X1 U22956 ( .B1(n20010), .B2(n20009), .A(n20008), .ZN(P2_U3211) );
  OAI222_X1 U22957 ( .A1(n20058), .A2(n20013), .B1(n20012), .B2(n20108), .C1(
        n20014), .C2(n20061), .ZN(P2_U3212) );
  OAI222_X1 U22958 ( .A1(n20061), .A2(n16471), .B1(n20015), .B2(n20108), .C1(
        n20014), .C2(n20058), .ZN(P2_U3213) );
  OAI222_X1 U22959 ( .A1(n20061), .A2(n19392), .B1(n20016), .B2(n20108), .C1(
        n16471), .C2(n20058), .ZN(P2_U3214) );
  OAI222_X1 U22960 ( .A1(n20061), .A2(n16460), .B1(n20017), .B2(n20108), .C1(
        n19392), .C2(n20058), .ZN(P2_U3215) );
  OAI222_X1 U22961 ( .A1(n20061), .A2(n20019), .B1(n20018), .B2(n20108), .C1(
        n16460), .C2(n20058), .ZN(P2_U3216) );
  OAI222_X1 U22962 ( .A1(n20061), .A2(n20021), .B1(n20020), .B2(n20108), .C1(
        n20019), .C2(n20058), .ZN(P2_U3217) );
  OAI222_X1 U22963 ( .A1(n20061), .A2(n11032), .B1(n20022), .B2(n20108), .C1(
        n20021), .C2(n20058), .ZN(P2_U3218) );
  OAI222_X1 U22964 ( .A1(n20061), .A2(n16436), .B1(n20023), .B2(n20108), .C1(
        n11032), .C2(n20058), .ZN(P2_U3219) );
  OAI222_X1 U22965 ( .A1(n20061), .A2(n15053), .B1(n20024), .B2(n20108), .C1(
        n16436), .C2(n20058), .ZN(P2_U3220) );
  INV_X1 U22966 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n20026) );
  OAI222_X1 U22967 ( .A1(n20061), .A2(n20026), .B1(n20025), .B2(n20108), .C1(
        n15053), .C2(n20058), .ZN(P2_U3221) );
  OAI222_X1 U22968 ( .A1(n20061), .A2(n19170), .B1(n20027), .B2(n20108), .C1(
        n20026), .C2(n20058), .ZN(P2_U3222) );
  OAI222_X1 U22969 ( .A1(n20061), .A2(n16401), .B1(n20028), .B2(n20108), .C1(
        n19170), .C2(n20058), .ZN(P2_U3223) );
  OAI222_X1 U22970 ( .A1(n20061), .A2(n11131), .B1(n20029), .B2(n20108), .C1(
        n16401), .C2(n20058), .ZN(P2_U3224) );
  OAI222_X1 U22971 ( .A1(n20061), .A2(n20031), .B1(n20030), .B2(n20108), .C1(
        n11131), .C2(n20058), .ZN(P2_U3225) );
  OAI222_X1 U22972 ( .A1(n20061), .A2(n20033), .B1(n20032), .B2(n20108), .C1(
        n20031), .C2(n20058), .ZN(P2_U3226) );
  OAI222_X1 U22973 ( .A1(n20061), .A2(n20035), .B1(n20034), .B2(n20108), .C1(
        n20033), .C2(n20058), .ZN(P2_U3227) );
  OAI222_X1 U22974 ( .A1(n20061), .A2(n15355), .B1(n20036), .B2(n20108), .C1(
        n20035), .C2(n20058), .ZN(P2_U3228) );
  OAI222_X1 U22975 ( .A1(n20061), .A2(n20038), .B1(n20037), .B2(n20108), .C1(
        n15355), .C2(n20058), .ZN(P2_U3229) );
  OAI222_X1 U22976 ( .A1(n20061), .A2(n11256), .B1(n20039), .B2(n20108), .C1(
        n20038), .C2(n20058), .ZN(P2_U3230) );
  OAI222_X1 U22977 ( .A1(n20061), .A2(n20041), .B1(n20040), .B2(n20108), .C1(
        n11256), .C2(n20058), .ZN(P2_U3231) );
  OAI222_X1 U22978 ( .A1(n20061), .A2(n11263), .B1(n20042), .B2(n20108), .C1(
        n20041), .C2(n20058), .ZN(P2_U3232) );
  OAI222_X1 U22979 ( .A1(n20061), .A2(n20044), .B1(n20043), .B2(n20108), .C1(
        n11263), .C2(n20058), .ZN(P2_U3233) );
  INV_X1 U22980 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20046) );
  OAI222_X1 U22981 ( .A1(n20061), .A2(n20046), .B1(n20045), .B2(n20108), .C1(
        n20044), .C2(n20058), .ZN(P2_U3234) );
  OAI222_X1 U22982 ( .A1(n20061), .A2(n20048), .B1(n20047), .B2(n20108), .C1(
        n20046), .C2(n20058), .ZN(P2_U3235) );
  OAI222_X1 U22983 ( .A1(n20061), .A2(n20050), .B1(n20049), .B2(n20108), .C1(
        n20048), .C2(n20058), .ZN(P2_U3236) );
  OAI222_X1 U22984 ( .A1(n20061), .A2(n20053), .B1(n20051), .B2(n20108), .C1(
        n20050), .C2(n20058), .ZN(P2_U3237) );
  INV_X1 U22985 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20054) );
  OAI222_X1 U22986 ( .A1(n20058), .A2(n20053), .B1(n20052), .B2(n20108), .C1(
        n20054), .C2(n20061), .ZN(P2_U3238) );
  OAI222_X1 U22987 ( .A1(n20061), .A2(n20056), .B1(n20055), .B2(n20108), .C1(
        n20054), .C2(n20058), .ZN(P2_U3239) );
  OAI222_X1 U22988 ( .A1(n20061), .A2(n14925), .B1(n20057), .B2(n20108), .C1(
        n20056), .C2(n20058), .ZN(P2_U3240) );
  INV_X1 U22989 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20059) );
  OAI222_X1 U22990 ( .A1(n20061), .A2(n20060), .B1(n20059), .B2(n20108), .C1(
        n14925), .C2(n20058), .ZN(P2_U3241) );
  OAI22_X1 U22991 ( .A1(n20109), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20108), .ZN(n20062) );
  INV_X1 U22992 ( .A(n20062), .ZN(P2_U3585) );
  MUX2_X1 U22993 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20109), .Z(P2_U3586) );
  OAI22_X1 U22994 ( .A1(n20109), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n20108), .ZN(n20063) );
  INV_X1 U22995 ( .A(n20063), .ZN(P2_U3587) );
  OAI22_X1 U22996 ( .A1(n20109), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20108), .ZN(n20064) );
  INV_X1 U22997 ( .A(n20064), .ZN(P2_U3588) );
  OAI21_X1 U22998 ( .B1(n20068), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20066), 
        .ZN(n20065) );
  INV_X1 U22999 ( .A(n20065), .ZN(P2_U3591) );
  OAI21_X1 U23000 ( .B1(n20068), .B2(n20067), .A(n20066), .ZN(P2_U3592) );
  INV_X1 U23001 ( .A(n20105), .ZN(n20104) );
  NAND2_X1 U23002 ( .A1(n20070), .A2(n20069), .ZN(n20077) );
  OR2_X1 U23003 ( .A1(n20071), .A2(n20093), .ZN(n20082) );
  NAND3_X1 U23004 ( .A1(n20094), .A2(n20072), .A3(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20073) );
  NAND2_X1 U23005 ( .A1(n20073), .A2(n20089), .ZN(n20083) );
  NAND2_X1 U23006 ( .A1(n20082), .A2(n20083), .ZN(n20075) );
  NAND2_X1 U23007 ( .A1(n20075), .A2(n20074), .ZN(n20076) );
  OAI211_X1 U23008 ( .C1(n20078), .C2(n13484), .A(n20077), .B(n20076), .ZN(
        n20079) );
  INV_X1 U23009 ( .A(n20079), .ZN(n20080) );
  AOI22_X1 U23010 ( .A1(n20104), .A2(n20081), .B1(n20080), .B2(n20105), .ZN(
        P2_U3602) );
  OAI21_X1 U23011 ( .B1(n20084), .B2(n20083), .A(n20082), .ZN(n20085) );
  AOI21_X1 U23012 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20086), .A(n20085), 
        .ZN(n20087) );
  AOI22_X1 U23013 ( .A1(n20104), .A2(n20088), .B1(n20087), .B2(n20105), .ZN(
        P2_U3603) );
  INV_X1 U23014 ( .A(n20089), .ZN(n20100) );
  AND2_X1 U23015 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20090) );
  OR3_X1 U23016 ( .A1(n20091), .A2(n20100), .A3(n20090), .ZN(n20092) );
  OAI21_X1 U23017 ( .B1(n20094), .B2(n20093), .A(n20092), .ZN(n20095) );
  AOI21_X1 U23018 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20096), .A(n20095), 
        .ZN(n20097) );
  AOI22_X1 U23019 ( .A1(n20104), .A2(n20098), .B1(n20097), .B2(n20105), .ZN(
        P2_U3604) );
  OAI22_X1 U23020 ( .A1(n20101), .A2(n20100), .B1(n19926), .B2(n20099), .ZN(
        n20102) );
  AOI21_X1 U23021 ( .B1(n20106), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20102), 
        .ZN(n20103) );
  OAI22_X1 U23022 ( .A1(n20106), .A2(n20105), .B1(n20104), .B2(n20103), .ZN(
        P2_U3605) );
  INV_X1 U23023 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20107) );
  AOI22_X1 U23024 ( .A1(n20108), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20107), 
        .B2(n20109), .ZN(P2_U3608) );
  OAI22_X1 U23025 ( .A1(n20109), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20108), .ZN(n20110) );
  INV_X1 U23026 ( .A(n20110), .ZN(P2_U3611) );
  AOI21_X1 U23027 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20885), .A(n12713), 
        .ZN(n20894) );
  INV_X1 U23028 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20111) );
  NAND2_X1 U23029 ( .A1(n12713), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20945) );
  AOI21_X1 U23030 ( .B1(n20894), .B2(n20111), .A(n20980), .ZN(P1_U2802) );
  NAND2_X1 U23031 ( .A1(n20885), .A2(n12713), .ZN(n20890) );
  INV_X1 U23032 ( .A(n20890), .ZN(n20112) );
  OAI21_X1 U23033 ( .B1(n20112), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20945), .ZN(
        n20113) );
  OAI21_X1 U23034 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20979), .A(n20113), 
        .ZN(P1_U2804) );
  INV_X1 U23035 ( .A(BS16), .ZN(n21102) );
  AOI21_X1 U23036 ( .B1(n21102), .B2(n20890), .A(n20884), .ZN(n20947) );
  AOI21_X1 U23037 ( .B1(n20884), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20947), 
        .ZN(n20114) );
  INV_X1 U23038 ( .A(n20114), .ZN(P1_U2805) );
  OAI21_X1 U23039 ( .B1(n20116), .B2(n21100), .A(n20115), .ZN(P1_U2806) );
  NOR4_X1 U23040 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20120) );
  NOR4_X1 U23041 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20119) );
  NOR4_X1 U23042 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20118) );
  NOR4_X1 U23043 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20117) );
  NAND4_X1 U23044 ( .A1(n20120), .A2(n20119), .A3(n20118), .A4(n20117), .ZN(
        n20126) );
  NOR4_X1 U23045 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20124) );
  AOI211_X1 U23046 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20123) );
  NOR4_X1 U23047 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20122) );
  NOR4_X1 U23048 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20121) );
  NAND4_X1 U23049 ( .A1(n20124), .A2(n20123), .A3(n20122), .A4(n20121), .ZN(
        n20125) );
  NOR2_X1 U23050 ( .A1(n20126), .A2(n20125), .ZN(n20965) );
  INV_X1 U23051 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21077) );
  NOR3_X1 U23052 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20128) );
  OAI21_X1 U23053 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20128), .A(n20965), .ZN(
        n20127) );
  OAI21_X1 U23054 ( .B1(n20965), .B2(n21077), .A(n20127), .ZN(P1_U2807) );
  INV_X1 U23055 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21093) );
  NOR2_X1 U23056 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20961) );
  OAI21_X1 U23057 ( .B1(n20128), .B2(n20961), .A(n20965), .ZN(n20129) );
  OAI21_X1 U23058 ( .B1(n20965), .B2(n21093), .A(n20129), .ZN(P1_U2808) );
  AOI22_X1 U23059 ( .A1(n20131), .A2(n20171), .B1(n20196), .B2(n20130), .ZN(
        n20140) );
  AOI22_X1 U23060 ( .A1(n20173), .A2(P1_EBX_REG_9__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n20186), .ZN(n20139) );
  INV_X1 U23061 ( .A(n20132), .ZN(n20137) );
  INV_X1 U23062 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20133) );
  OAI21_X1 U23063 ( .B1(n20175), .B2(n20134), .A(n20133), .ZN(n20135) );
  AOI22_X1 U23064 ( .A1(n20137), .A2(n20165), .B1(n20136), .B2(n20135), .ZN(
        n20138) );
  NAND4_X1 U23065 ( .A1(n20140), .A2(n20139), .A3(n20138), .A4(n20187), .ZN(
        P1_U2831) );
  NOR4_X1 U23066 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20175), .A3(n20174), .A4(
        n20145), .ZN(n20152) );
  OAI22_X1 U23067 ( .A1(n20190), .A2(n20143), .B1(n20142), .B2(n20141), .ZN(
        n20151) );
  NAND2_X1 U23068 ( .A1(n20146), .A2(n20174), .ZN(n20193) );
  NAND2_X1 U23069 ( .A1(n20193), .A2(n20144), .ZN(n20197) );
  AOI21_X1 U23070 ( .B1(n20146), .B2(n20145), .A(n20197), .ZN(n20169) );
  OAI22_X1 U23071 ( .A1(n20149), .A2(n20148), .B1(n20147), .B2(n20169), .ZN(
        n20150) );
  NOR4_X1 U23072 ( .A1(n20177), .A2(n20152), .A3(n20151), .A4(n20150), .ZN(
        n20155) );
  NAND2_X1 U23073 ( .A1(n20196), .A2(n20153), .ZN(n20154) );
  OAI211_X1 U23074 ( .C1(n20189), .C2(n20156), .A(n20155), .B(n20154), .ZN(
        P1_U2833) );
  INV_X1 U23075 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20168) );
  AOI21_X1 U23076 ( .B1(n20186), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20177), .ZN(n20157) );
  OAI21_X1 U23077 ( .B1(n20189), .B2(n20158), .A(n20157), .ZN(n20159) );
  AOI21_X1 U23078 ( .B1(n20173), .B2(P1_EBX_REG_6__SCAN_IN), .A(n20159), .ZN(
        n20160) );
  OAI21_X1 U23079 ( .B1(n20162), .B2(n20161), .A(n20160), .ZN(n20164) );
  NOR4_X1 U23080 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20174), .A3(n20175), .A4(
        n20908), .ZN(n20163) );
  AOI211_X1 U23081 ( .C1(n20166), .C2(n20165), .A(n20164), .B(n20163), .ZN(
        n20167) );
  OAI21_X1 U23082 ( .B1(n20169), .B2(n20168), .A(n20167), .ZN(P1_U2834) );
  INV_X1 U23083 ( .A(n20170), .ZN(n20172) );
  AOI22_X1 U23084 ( .A1(n20173), .A2(P1_EBX_REG_5__SCAN_IN), .B1(n20172), .B2(
        n20171), .ZN(n20183) );
  NOR2_X1 U23085 ( .A1(n20175), .A2(n20174), .ZN(n20176) );
  AOI22_X1 U23086 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n20186), .B1(
        n20176), .B2(n20908), .ZN(n20182) );
  AOI21_X1 U23087 ( .B1(n20196), .B2(n20178), .A(n20177), .ZN(n20181) );
  AOI22_X1 U23088 ( .A1(n20179), .A2(n20198), .B1(P1_REIP_REG_5__SCAN_IN), 
        .B2(n20197), .ZN(n20180) );
  NAND4_X1 U23089 ( .A1(n20183), .A2(n20182), .A3(n20181), .A4(n20180), .ZN(
        P1_U2835) );
  AOI22_X1 U23090 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n20186), .B1(
        n20185), .B2(n20184), .ZN(n20188) );
  OAI211_X1 U23091 ( .C1(n20189), .C2(n20242), .A(n20188), .B(n20187), .ZN(
        n20195) );
  NAND3_X1 U23092 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n20192) );
  OAI22_X1 U23093 ( .A1(n20193), .A2(n20192), .B1(n20191), .B2(n20190), .ZN(
        n20194) );
  AOI211_X1 U23094 ( .C1(n20196), .C2(n20257), .A(n20195), .B(n20194), .ZN(
        n20200) );
  AOI22_X1 U23095 ( .A1(n20239), .A2(n20198), .B1(P1_REIP_REG_4__SCAN_IN), 
        .B2(n20197), .ZN(n20199) );
  NAND2_X1 U23096 ( .A1(n20200), .A2(n20199), .ZN(P1_U2836) );
  AOI22_X1 U23097 ( .A1(n20231), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20230), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20202) );
  OAI21_X1 U23098 ( .B1(n14712), .B2(n20233), .A(n20202), .ZN(P1_U2921) );
  AOI22_X1 U23099 ( .A1(n20231), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20230), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20203) );
  OAI21_X1 U23100 ( .B1(n20204), .B2(n20233), .A(n20203), .ZN(P1_U2922) );
  AOI22_X1 U23101 ( .A1(n20231), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20230), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20205) );
  OAI21_X1 U23102 ( .B1(n20206), .B2(n20233), .A(n20205), .ZN(P1_U2923) );
  AOI22_X1 U23103 ( .A1(n20231), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20230), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20207) );
  OAI21_X1 U23104 ( .B1(n20208), .B2(n20233), .A(n20207), .ZN(P1_U2924) );
  AOI22_X1 U23105 ( .A1(n20231), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20218), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20209) );
  OAI21_X1 U23106 ( .B1(n20210), .B2(n20233), .A(n20209), .ZN(P1_U2925) );
  AOI22_X1 U23107 ( .A1(n20231), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20218), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20211) );
  OAI21_X1 U23108 ( .B1(n20212), .B2(n20233), .A(n20211), .ZN(P1_U2926) );
  AOI22_X1 U23109 ( .A1(n20231), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20218), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20213) );
  OAI21_X1 U23110 ( .B1(n20214), .B2(n20233), .A(n20213), .ZN(P1_U2927) );
  AOI22_X1 U23111 ( .A1(n20231), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20218), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20215) );
  OAI21_X1 U23112 ( .B1(n20216), .B2(n20233), .A(n20215), .ZN(P1_U2928) );
  AOI22_X1 U23113 ( .A1(n20231), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20218), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20217) );
  OAI21_X1 U23114 ( .B1(n11892), .B2(n20233), .A(n20217), .ZN(P1_U2929) );
  AOI22_X1 U23115 ( .A1(n20231), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20218), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20219) );
  OAI21_X1 U23116 ( .B1(n20220), .B2(n20233), .A(n20219), .ZN(P1_U2930) );
  AOI22_X1 U23117 ( .A1(n20231), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20230), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20221) );
  OAI21_X1 U23118 ( .B1(n11873), .B2(n20233), .A(n20221), .ZN(P1_U2931) );
  AOI22_X1 U23119 ( .A1(n20231), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20230), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20222) );
  OAI21_X1 U23120 ( .B1(n20223), .B2(n20233), .A(n20222), .ZN(P1_U2932) );
  AOI22_X1 U23121 ( .A1(n20231), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20230), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20224) );
  OAI21_X1 U23122 ( .B1(n20225), .B2(n20233), .A(n20224), .ZN(P1_U2933) );
  AOI22_X1 U23123 ( .A1(n20231), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20230), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20226) );
  OAI21_X1 U23124 ( .B1(n20227), .B2(n20233), .A(n20226), .ZN(P1_U2934) );
  AOI22_X1 U23125 ( .A1(n20231), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20230), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20228) );
  OAI21_X1 U23126 ( .B1(n20229), .B2(n20233), .A(n20228), .ZN(P1_U2935) );
  AOI22_X1 U23127 ( .A1(n20231), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20230), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20232) );
  OAI21_X1 U23128 ( .B1(n20234), .B2(n20233), .A(n20232), .ZN(P1_U2936) );
  AOI22_X1 U23129 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20290), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20241) );
  OAI21_X1 U23130 ( .B1(n20237), .B2(n20236), .A(n20235), .ZN(n20238) );
  INV_X1 U23131 ( .A(n20238), .ZN(n20262) );
  AOI22_X1 U23132 ( .A1(n20262), .A2(n20250), .B1(n20313), .B2(n20239), .ZN(
        n20240) );
  OAI211_X1 U23133 ( .C1(n20243), .C2(n20242), .A(n20241), .B(n20240), .ZN(
        P1_U2995) );
  AOI22_X1 U23134 ( .A1(n20244), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20290), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n20252) );
  OAI21_X1 U23135 ( .B1(n20246), .B2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n20245), .ZN(n20247) );
  INV_X1 U23136 ( .A(n20247), .ZN(n20297) );
  AOI22_X1 U23137 ( .A1(n20297), .A2(n20250), .B1(n20249), .B2(n20248), .ZN(
        n20251) );
  OAI211_X1 U23138 ( .C1(n20254), .C2(n20253), .A(n20252), .B(n20251), .ZN(
        P1_U2998) );
  NOR2_X1 U23139 ( .A1(n20259), .A2(n20279), .ZN(n20255) );
  OAI21_X1 U23140 ( .B1(n20276), .B2(n20255), .A(n20273), .ZN(n20272) );
  OAI21_X1 U23141 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20256), .ZN(n20265) );
  AOI22_X1 U23142 ( .A1(n20290), .A2(P1_REIP_REG_4__SCAN_IN), .B1(n20292), 
        .B2(n20257), .ZN(n20264) );
  AOI21_X1 U23143 ( .B1(n20260), .B2(n20259), .A(n20258), .ZN(n20283) );
  OAI21_X1 U23144 ( .B1(n20273), .B2(n20261), .A(n20283), .ZN(n20268) );
  AOI22_X1 U23145 ( .A1(n20262), .A2(n20296), .B1(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n20268), .ZN(n20263) );
  OAI211_X1 U23146 ( .C1(n20272), .C2(n20265), .A(n20264), .B(n20263), .ZN(
        P1_U3027) );
  AOI22_X1 U23147 ( .A1(n20290), .A2(P1_REIP_REG_3__SCAN_IN), .B1(n20292), 
        .B2(n20266), .ZN(n20271) );
  INV_X1 U23148 ( .A(n20267), .ZN(n20269) );
  AOI22_X1 U23149 ( .A1(n20269), .A2(n20296), .B1(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n20268), .ZN(n20270) );
  OAI211_X1 U23150 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n20272), .A(
        n20271), .B(n20270), .ZN(P1_U3028) );
  NAND2_X1 U23151 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20274) );
  OAI21_X1 U23152 ( .B1(n20274), .B2(n20282), .A(n20273), .ZN(n20275) );
  AOI22_X1 U23153 ( .A1(n20290), .A2(P1_REIP_REG_2__SCAN_IN), .B1(n20276), 
        .B2(n20275), .ZN(n20286) );
  NAND3_X1 U23154 ( .A1(n13791), .A2(n20277), .A3(n20296), .ZN(n20281) );
  NAND2_X1 U23155 ( .A1(n20282), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20278) );
  OR2_X1 U23156 ( .A1(n20279), .A2(n20278), .ZN(n20280) );
  OAI211_X1 U23157 ( .C1(n20283), .C2(n20282), .A(n20281), .B(n20280), .ZN(
        n20284) );
  INV_X1 U23158 ( .A(n20284), .ZN(n20285) );
  OAI211_X1 U23159 ( .C1(n20288), .C2(n20287), .A(n20286), .B(n20285), .ZN(
        P1_U3029) );
  INV_X1 U23160 ( .A(n20289), .ZN(n20291) );
  AOI22_X1 U23161 ( .A1(n20292), .A2(n20291), .B1(n20290), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n20299) );
  NOR2_X1 U23162 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20293), .ZN(
        n20295) );
  AOI22_X1 U23163 ( .A1(n20297), .A2(n20296), .B1(n20295), .B2(n20294), .ZN(
        n20298) );
  OAI211_X1 U23164 ( .C1(n20301), .C2(n20300), .A(n20299), .B(n20298), .ZN(
        P1_U3030) );
  NOR2_X1 U23165 ( .A1(n20303), .A2(n20302), .ZN(P1_U3032) );
  INV_X1 U23166 ( .A(n20635), .ZN(n20580) );
  OR2_X1 U23167 ( .A1(n20580), .A2(n20579), .ZN(n20471) );
  INV_X1 U23168 ( .A(n20318), .ZN(n20304) );
  NOR2_X1 U23169 ( .A1(n20304), .A2(n20968), .ZN(n20709) );
  INV_X1 U23170 ( .A(n20640), .ZN(n20413) );
  INV_X1 U23171 ( .A(n11838), .ZN(n20306) );
  OAI21_X1 U23172 ( .B1(n20876), .B2(n20405), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20307) );
  NAND2_X1 U23173 ( .A1(n20307), .A2(n20823), .ZN(n20320) );
  OR2_X1 U23174 ( .A1(n20578), .A2(n20308), .ZN(n20439) );
  OR2_X1 U23175 ( .A1(n20439), .A2(n20783), .ZN(n20319) );
  INV_X1 U23176 ( .A(n20319), .ZN(n20309) );
  NOR3_X1 U23177 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20388) );
  INV_X1 U23178 ( .A(n20388), .ZN(n20384) );
  NOR2_X1 U23179 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20384), .ZN(
        n20374) );
  OAI22_X1 U23180 ( .A1(n20320), .A2(n20309), .B1(n20374), .B2(n11516), .ZN(
        n20310) );
  AOI211_X2 U23181 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20471), .A(n20413), 
        .B(n20310), .ZN(n20375) );
  INV_X1 U23182 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20324) );
  INV_X1 U23183 ( .A(DATAI_24_), .ZN(n21079) );
  OAI22_X2 U23184 ( .A1(n20314), .A2(n20370), .B1(n21079), .B2(n20368), .ZN(
        n20829) );
  NOR2_X2 U23185 ( .A1(n20373), .A2(n20316), .ZN(n20820) );
  AOI22_X1 U23186 ( .A1(n20876), .A2(n20829), .B1(n20820), .B2(n20374), .ZN(
        n20323) );
  NOR2_X1 U23187 ( .A1(n20318), .A2(n20968), .ZN(n20637) );
  INV_X1 U23188 ( .A(n20637), .ZN(n20582) );
  OAI22_X1 U23189 ( .A1(n20320), .A2(n20319), .B1(n20582), .B2(n20471), .ZN(
        n20378) );
  INV_X1 U23190 ( .A(DATAI_16_), .ZN(n21143) );
  OAI22_X1 U23191 ( .A1(n20321), .A2(n20370), .B1(n21143), .B2(n20368), .ZN(
        n20711) );
  AOI22_X1 U23192 ( .A1(n20821), .A2(n20378), .B1(n20405), .B2(n20711), .ZN(
        n20322) );
  OAI211_X1 U23193 ( .C1(n20375), .C2(n20324), .A(n20323), .B(n20322), .ZN(
        P1_U3033) );
  INV_X1 U23194 ( .A(DATAI_25_), .ZN(n21105) );
  OAI22_X2 U23195 ( .A1(n20325), .A2(n20370), .B1(n21105), .B2(n20368), .ZN(
        n20792) );
  NOR2_X2 U23196 ( .A1(n20373), .A2(n20326), .ZN(n20833) );
  AOI22_X1 U23197 ( .A1(n20876), .A2(n20792), .B1(n20833), .B2(n20374), .ZN(
        n20329) );
  INV_X1 U23198 ( .A(DATAI_17_), .ZN(n21027) );
  AOI22_X1 U23199 ( .A1(n20834), .A2(n20378), .B1(n20405), .B2(n20835), .ZN(
        n20328) );
  OAI211_X1 U23200 ( .C1(n20375), .C2(n20330), .A(n20329), .B(n20328), .ZN(
        P1_U3034) );
  INV_X1 U23201 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n20336) );
  INV_X1 U23202 ( .A(DATAI_26_), .ZN(n21121) );
  OAI22_X2 U23203 ( .A1(n20331), .A2(n20370), .B1(n21121), .B2(n20368), .ZN(
        n20796) );
  NOR2_X2 U23204 ( .A1(n20373), .A2(n11563), .ZN(n20839) );
  AOI22_X1 U23205 ( .A1(n20876), .A2(n20796), .B1(n20839), .B2(n20374), .ZN(
        n20335) );
  INV_X1 U23206 ( .A(DATAI_18_), .ZN(n21108) );
  AOI22_X1 U23207 ( .A1(n20840), .A2(n20378), .B1(n20405), .B2(n20841), .ZN(
        n20334) );
  OAI211_X1 U23208 ( .C1(n20375), .C2(n20336), .A(n20335), .B(n20334), .ZN(
        P1_U3035) );
  INV_X1 U23209 ( .A(DATAI_27_), .ZN(n20337) );
  OAI22_X2 U23210 ( .A1(n20338), .A2(n20370), .B1(n20337), .B2(n20368), .ZN(
        n20847) );
  NOR2_X2 U23211 ( .A1(n20373), .A2(n20339), .ZN(n20845) );
  AOI22_X1 U23212 ( .A1(n20876), .A2(n20847), .B1(n20845), .B2(n20374), .ZN(
        n20343) );
  OAI22_X1 U23213 ( .A1(n14693), .A2(n20368), .B1(n20341), .B2(n20370), .ZN(
        n20726) );
  AOI22_X1 U23214 ( .A1(n20846), .A2(n20378), .B1(n20405), .B2(n20726), .ZN(
        n20342) );
  OAI211_X1 U23215 ( .C1(n20375), .C2(n20344), .A(n20343), .B(n20342), .ZN(
        P1_U3036) );
  INV_X1 U23216 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n20352) );
  INV_X1 U23217 ( .A(DATAI_28_), .ZN(n20345) );
  OAI22_X2 U23218 ( .A1(n20346), .A2(n20370), .B1(n20345), .B2(n20368), .ZN(
        n20853) );
  NOR2_X2 U23219 ( .A1(n20373), .A2(n20347), .ZN(n20852) );
  AOI22_X1 U23220 ( .A1(n20876), .A2(n20853), .B1(n20852), .B2(n20374), .ZN(
        n20351) );
  NAND2_X1 U23221 ( .A1(n20377), .A2(n20348), .ZN(n20733) );
  INV_X1 U23222 ( .A(DATAI_20_), .ZN(n21091) );
  OAI22_X1 U23223 ( .A1(n20349), .A2(n20370), .B1(n21091), .B2(n20368), .ZN(
        n20730) );
  AOI22_X1 U23224 ( .A1(n20851), .A2(n20378), .B1(n20405), .B2(n20730), .ZN(
        n20350) );
  OAI211_X1 U23225 ( .C1(n20375), .C2(n20352), .A(n20351), .B(n20350), .ZN(
        P1_U3037) );
  INV_X1 U23226 ( .A(DATAI_29_), .ZN(n21030) );
  OAI22_X2 U23227 ( .A1(n20353), .A2(n20370), .B1(n21030), .B2(n20368), .ZN(
        n20859) );
  NOR2_X2 U23228 ( .A1(n20373), .A2(n11510), .ZN(n20858) );
  AOI22_X1 U23229 ( .A1(n20876), .A2(n20859), .B1(n20858), .B2(n20374), .ZN(
        n20357) );
  NAND2_X1 U23230 ( .A1(n20377), .A2(n20354), .ZN(n20737) );
  INV_X1 U23231 ( .A(DATAI_21_), .ZN(n21083) );
  OAI22_X1 U23232 ( .A1(n20355), .A2(n20370), .B1(n21083), .B2(n20368), .ZN(
        n20734) );
  AOI22_X1 U23233 ( .A1(n20857), .A2(n20378), .B1(n20405), .B2(n20734), .ZN(
        n20356) );
  OAI211_X1 U23234 ( .C1(n20375), .C2(n20358), .A(n20357), .B(n20356), .ZN(
        P1_U3038) );
  INV_X1 U23235 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20365) );
  INV_X1 U23236 ( .A(DATAI_30_), .ZN(n20359) );
  OAI22_X2 U23237 ( .A1(n20360), .A2(n20370), .B1(n20359), .B2(n20368), .ZN(
        n20865) );
  AOI22_X1 U23238 ( .A1(n20876), .A2(n20865), .B1(n20864), .B2(n20374), .ZN(
        n20364) );
  NAND2_X1 U23239 ( .A1(n20377), .A2(n20361), .ZN(n20741) );
  INV_X1 U23240 ( .A(DATAI_22_), .ZN(n21017) );
  OAI22_X1 U23241 ( .A1(n21017), .A2(n20368), .B1(n20362), .B2(n20370), .ZN(
        n20738) );
  AOI22_X1 U23242 ( .A1(n20863), .A2(n20378), .B1(n20405), .B2(n20738), .ZN(
        n20363) );
  OAI211_X1 U23243 ( .C1(n20375), .C2(n20365), .A(n20364), .B(n20363), .ZN(
        P1_U3039) );
  INV_X1 U23244 ( .A(DATAI_23_), .ZN(n20366) );
  OAI22_X1 U23245 ( .A1(n20367), .A2(n20370), .B1(n20366), .B2(n20368), .ZN(
        n20875) );
  INV_X1 U23246 ( .A(n20875), .ZN(n20815) );
  INV_X1 U23247 ( .A(DATAI_31_), .ZN(n20369) );
  OAI22_X2 U23248 ( .A1(n20371), .A2(n20370), .B1(n20369), .B2(n20368), .ZN(
        n20810) );
  NOR2_X2 U23249 ( .A1(n20373), .A2(n20372), .ZN(n20874) );
  AOI22_X1 U23250 ( .A1(n20876), .A2(n20810), .B1(n20874), .B2(n20374), .ZN(
        n20381) );
  INV_X1 U23251 ( .A(n20375), .ZN(n20379) );
  NAND2_X1 U23252 ( .A1(n20377), .A2(n20376), .ZN(n20747) );
  AOI22_X1 U23253 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20379), .B1(
        n20871), .B2(n20378), .ZN(n20380) );
  OAI211_X1 U23254 ( .C1(n20815), .C2(n20382), .A(n20381), .B(n20380), .ZN(
        P1_U3040) );
  INV_X1 U23255 ( .A(n20711), .ZN(n20832) );
  INV_X1 U23256 ( .A(n20439), .ZN(n20383) );
  INV_X1 U23257 ( .A(n20753), .ZN(n20608) );
  NOR2_X1 U23258 ( .A1(n20751), .A2(n20384), .ZN(n20404) );
  AOI21_X1 U23259 ( .B1(n20383), .B2(n20608), .A(n20404), .ZN(n20385) );
  OAI22_X1 U23260 ( .A1(n20385), .A2(n20817), .B1(n20384), .B2(n20968), .ZN(
        n20403) );
  AOI22_X1 U23261 ( .A1(n20821), .A2(n20403), .B1(n20820), .B2(n20404), .ZN(
        n20390) );
  NOR2_X1 U23262 ( .A1(n20448), .A2(n20386), .ZN(n20387) );
  OAI21_X1 U23263 ( .B1(n20388), .B2(n20387), .A(n20827), .ZN(n20406) );
  AOI22_X1 U23264 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20406), .B1(
        n20405), .B2(n20829), .ZN(n20389) );
  OAI211_X1 U23265 ( .C1(n20832), .C2(n20409), .A(n20390), .B(n20389), .ZN(
        P1_U3041) );
  INV_X1 U23266 ( .A(n20835), .ZN(n20795) );
  AOI22_X1 U23267 ( .A1(n20834), .A2(n20403), .B1(n20833), .B2(n20404), .ZN(
        n20392) );
  AOI22_X1 U23268 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20406), .B1(
        n20405), .B2(n20792), .ZN(n20391) );
  OAI211_X1 U23269 ( .C1(n20795), .C2(n20409), .A(n20392), .B(n20391), .ZN(
        P1_U3042) );
  INV_X1 U23270 ( .A(n20841), .ZN(n20799) );
  AOI22_X1 U23271 ( .A1(n20840), .A2(n20403), .B1(n20839), .B2(n20404), .ZN(
        n20394) );
  AOI22_X1 U23272 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20406), .B1(
        n20405), .B2(n20796), .ZN(n20393) );
  OAI211_X1 U23273 ( .C1(n20799), .C2(n20409), .A(n20394), .B(n20393), .ZN(
        P1_U3043) );
  INV_X1 U23274 ( .A(n20726), .ZN(n20850) );
  AOI22_X1 U23275 ( .A1(n20846), .A2(n20403), .B1(n20845), .B2(n20404), .ZN(
        n20396) );
  AOI22_X1 U23276 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20406), .B1(
        n20405), .B2(n20847), .ZN(n20395) );
  OAI211_X1 U23277 ( .C1(n20850), .C2(n20409), .A(n20396), .B(n20395), .ZN(
        P1_U3044) );
  INV_X1 U23278 ( .A(n20730), .ZN(n20856) );
  AOI22_X1 U23279 ( .A1(n20852), .A2(n20404), .B1(n20403), .B2(n20851), .ZN(
        n20398) );
  AOI22_X1 U23280 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20406), .B1(
        n20405), .B2(n20853), .ZN(n20397) );
  OAI211_X1 U23281 ( .C1(n20856), .C2(n20409), .A(n20398), .B(n20397), .ZN(
        P1_U3045) );
  INV_X1 U23282 ( .A(n20734), .ZN(n20862) );
  AOI22_X1 U23283 ( .A1(n20858), .A2(n20404), .B1(n20403), .B2(n20857), .ZN(
        n20400) );
  AOI22_X1 U23284 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20406), .B1(
        n20405), .B2(n20859), .ZN(n20399) );
  OAI211_X1 U23285 ( .C1(n20862), .C2(n20409), .A(n20400), .B(n20399), .ZN(
        P1_U3046) );
  INV_X1 U23286 ( .A(n20738), .ZN(n20870) );
  AOI22_X1 U23287 ( .A1(n20864), .A2(n20404), .B1(n20403), .B2(n20863), .ZN(
        n20402) );
  AOI22_X1 U23288 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20406), .B1(
        n20405), .B2(n20865), .ZN(n20401) );
  OAI211_X1 U23289 ( .C1(n20870), .C2(n20409), .A(n20402), .B(n20401), .ZN(
        P1_U3047) );
  AOI22_X1 U23290 ( .A1(n20874), .A2(n20404), .B1(n20403), .B2(n20871), .ZN(
        n20408) );
  AOI22_X1 U23291 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20406), .B1(
        n20405), .B2(n20810), .ZN(n20407) );
  OAI211_X1 U23292 ( .C1(n20815), .C2(n20409), .A(n20408), .B(n20407), .ZN(
        P1_U3048) );
  NOR2_X2 U23293 ( .A1(n20448), .A2(n20778), .ZN(n20464) );
  NOR3_X1 U23294 ( .A1(n20464), .A2(n20433), .A3(n20817), .ZN(n20411) );
  NOR2_X1 U23295 ( .A1(n20411), .A2(n20410), .ZN(n20417) );
  INV_X1 U23296 ( .A(n20417), .ZN(n20412) );
  NOR2_X1 U23297 ( .A1(n20439), .A2(n13673), .ZN(n20416) );
  INV_X1 U23298 ( .A(n20821), .ZN(n20719) );
  NOR3_X1 U23299 ( .A1(n20638), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20443) );
  NAND2_X1 U23300 ( .A1(n20751), .A2(n20443), .ZN(n20414) );
  INV_X1 U23301 ( .A(n20414), .ZN(n20432) );
  AOI22_X1 U23302 ( .A1(n20464), .A2(n20711), .B1(n20432), .B2(n20820), .ZN(
        n20419) );
  NOR2_X1 U23303 ( .A1(n10210), .A2(n20968), .ZN(n20524) );
  AOI211_X1 U23304 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20414), .A(n20524), 
        .B(n20413), .ZN(n20415) );
  OAI21_X1 U23305 ( .B1(n20417), .B2(n20416), .A(n20415), .ZN(n20434) );
  AOI22_X1 U23306 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20434), .B1(
        n20433), .B2(n20829), .ZN(n20418) );
  OAI211_X1 U23307 ( .C1(n20437), .C2(n20719), .A(n20419), .B(n20418), .ZN(
        P1_U3049) );
  INV_X1 U23308 ( .A(n20834), .ZN(n20722) );
  AOI22_X1 U23309 ( .A1(n20433), .A2(n20792), .B1(n20833), .B2(n20432), .ZN(
        n20421) );
  AOI22_X1 U23310 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20434), .B1(
        n20464), .B2(n20835), .ZN(n20420) );
  OAI211_X1 U23311 ( .C1(n20437), .C2(n20722), .A(n20421), .B(n20420), .ZN(
        P1_U3050) );
  INV_X1 U23312 ( .A(n20840), .ZN(n20725) );
  AOI22_X1 U23313 ( .A1(n20433), .A2(n20796), .B1(n20839), .B2(n20432), .ZN(
        n20423) );
  AOI22_X1 U23314 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20434), .B1(
        n20464), .B2(n20841), .ZN(n20422) );
  OAI211_X1 U23315 ( .C1(n20437), .C2(n20725), .A(n20423), .B(n20422), .ZN(
        P1_U3051) );
  INV_X1 U23316 ( .A(n20846), .ZN(n20729) );
  AOI22_X1 U23317 ( .A1(n20433), .A2(n20847), .B1(n20432), .B2(n20845), .ZN(
        n20425) );
  AOI22_X1 U23318 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20434), .B1(
        n20464), .B2(n20726), .ZN(n20424) );
  OAI211_X1 U23319 ( .C1(n20437), .C2(n20729), .A(n20425), .B(n20424), .ZN(
        P1_U3052) );
  AOI22_X1 U23320 ( .A1(n20433), .A2(n20853), .B1(n20432), .B2(n20852), .ZN(
        n20427) );
  AOI22_X1 U23321 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20434), .B1(
        n20464), .B2(n20730), .ZN(n20426) );
  OAI211_X1 U23322 ( .C1(n20437), .C2(n20733), .A(n20427), .B(n20426), .ZN(
        P1_U3053) );
  AOI22_X1 U23323 ( .A1(n20433), .A2(n20859), .B1(n20858), .B2(n20432), .ZN(
        n20429) );
  AOI22_X1 U23324 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20434), .B1(
        n20464), .B2(n20734), .ZN(n20428) );
  OAI211_X1 U23325 ( .C1(n20437), .C2(n20737), .A(n20429), .B(n20428), .ZN(
        P1_U3054) );
  AOI22_X1 U23326 ( .A1(n20464), .A2(n20738), .B1(n20864), .B2(n20432), .ZN(
        n20431) );
  AOI22_X1 U23327 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20434), .B1(
        n20433), .B2(n20865), .ZN(n20430) );
  OAI211_X1 U23328 ( .C1(n20437), .C2(n20741), .A(n20431), .B(n20430), .ZN(
        P1_U3055) );
  AOI22_X1 U23329 ( .A1(n20433), .A2(n20810), .B1(n20874), .B2(n20432), .ZN(
        n20436) );
  AOI22_X1 U23330 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20434), .B1(
        n20464), .B2(n20875), .ZN(n20435) );
  OAI211_X1 U23331 ( .C1(n20437), .C2(n20747), .A(n20436), .B(n20435), .ZN(
        P1_U3056) );
  INV_X1 U23332 ( .A(n20448), .ZN(n20438) );
  INV_X1 U23333 ( .A(n20671), .ZN(n20822) );
  AOI21_X1 U23334 ( .B1(n20438), .B2(n20822), .A(n20817), .ZN(n20445) );
  AND2_X1 U23335 ( .A1(n9955), .A2(n11841), .ZN(n20667) );
  INV_X1 U23336 ( .A(n20667), .ZN(n20818) );
  OR2_X1 U23337 ( .A1(n20439), .A2(n20818), .ZN(n20441) );
  NOR2_X1 U23338 ( .A1(n20666), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20463) );
  INV_X1 U23339 ( .A(n20463), .ZN(n20440) );
  AND2_X1 U23340 ( .A1(n20441), .A2(n20440), .ZN(n20446) );
  INV_X1 U23341 ( .A(n20446), .ZN(n20442) );
  AOI22_X1 U23342 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20443), .B1(n20445), 
        .B2(n20442), .ZN(n20468) );
  AOI22_X1 U23343 ( .A1(n20464), .A2(n20829), .B1(n20463), .B2(n20820), .ZN(
        n20450) );
  OAI21_X1 U23344 ( .B1(n20823), .B2(n20443), .A(n20827), .ZN(n20444) );
  AOI21_X1 U23345 ( .B1(n20446), .B2(n20445), .A(n20444), .ZN(n20447) );
  NOR2_X2 U23346 ( .A1(n20448), .A2(n20674), .ZN(n20493) );
  AOI22_X1 U23347 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20465), .B1(
        n20493), .B2(n20711), .ZN(n20449) );
  OAI211_X1 U23348 ( .C1(n20468), .C2(n20719), .A(n20450), .B(n20449), .ZN(
        P1_U3057) );
  AOI22_X1 U23349 ( .A1(n20464), .A2(n20792), .B1(n20463), .B2(n20833), .ZN(
        n20452) );
  AOI22_X1 U23350 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20465), .B1(
        n20493), .B2(n20835), .ZN(n20451) );
  OAI211_X1 U23351 ( .C1(n20468), .C2(n20722), .A(n20452), .B(n20451), .ZN(
        P1_U3058) );
  AOI22_X1 U23352 ( .A1(n20493), .A2(n20841), .B1(n20839), .B2(n20463), .ZN(
        n20454) );
  AOI22_X1 U23353 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20465), .B1(
        n20464), .B2(n20796), .ZN(n20453) );
  OAI211_X1 U23354 ( .C1(n20468), .C2(n20725), .A(n20454), .B(n20453), .ZN(
        P1_U3059) );
  AOI22_X1 U23355 ( .A1(n20464), .A2(n20847), .B1(n20463), .B2(n20845), .ZN(
        n20456) );
  AOI22_X1 U23356 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20465), .B1(
        n20493), .B2(n20726), .ZN(n20455) );
  OAI211_X1 U23357 ( .C1(n20468), .C2(n20729), .A(n20456), .B(n20455), .ZN(
        P1_U3060) );
  AOI22_X1 U23358 ( .A1(n20464), .A2(n20853), .B1(n20463), .B2(n20852), .ZN(
        n20458) );
  AOI22_X1 U23359 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20465), .B1(
        n20493), .B2(n20730), .ZN(n20457) );
  OAI211_X1 U23360 ( .C1(n20468), .C2(n20733), .A(n20458), .B(n20457), .ZN(
        P1_U3061) );
  AOI22_X1 U23361 ( .A1(n20493), .A2(n20734), .B1(n20463), .B2(n20858), .ZN(
        n20460) );
  AOI22_X1 U23362 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20465), .B1(
        n20464), .B2(n20859), .ZN(n20459) );
  OAI211_X1 U23363 ( .C1(n20468), .C2(n20737), .A(n20460), .B(n20459), .ZN(
        P1_U3062) );
  AOI22_X1 U23364 ( .A1(n20493), .A2(n20738), .B1(n20463), .B2(n20864), .ZN(
        n20462) );
  AOI22_X1 U23365 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20465), .B1(
        n20464), .B2(n20865), .ZN(n20461) );
  OAI211_X1 U23366 ( .C1(n20468), .C2(n20741), .A(n20462), .B(n20461), .ZN(
        P1_U3063) );
  AOI22_X1 U23367 ( .A1(n20493), .A2(n20875), .B1(n20463), .B2(n20874), .ZN(
        n20467) );
  AOI22_X1 U23368 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20465), .B1(
        n20464), .B2(n20810), .ZN(n20466) );
  OAI211_X1 U23369 ( .C1(n20468), .C2(n20747), .A(n20467), .B(n20466), .ZN(
        P1_U3064) );
  INV_X1 U23370 ( .A(n20709), .ZN(n20780) );
  NOR2_X1 U23371 ( .A1(n13690), .A2(n20469), .ZN(n20550) );
  NAND3_X1 U23372 ( .A1(n20550), .A2(n20823), .A3(n13673), .ZN(n20470) );
  OAI21_X1 U23373 ( .B1(n20780), .B2(n20471), .A(n20470), .ZN(n20491) );
  NOR3_X1 U23374 ( .A1(n11776), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20500) );
  INV_X1 U23375 ( .A(n20500), .ZN(n20497) );
  NOR2_X1 U23376 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20497), .ZN(
        n20492) );
  AOI22_X1 U23377 ( .A1(n20821), .A2(n20491), .B1(n20820), .B2(n20492), .ZN(
        n20478) );
  INV_X1 U23378 ( .A(n20493), .ZN(n20472) );
  AOI21_X1 U23379 ( .B1(n20472), .B2(n20520), .A(n21106), .ZN(n20473) );
  AOI21_X1 U23380 ( .B1(n20550), .B2(n13673), .A(n20473), .ZN(n20474) );
  NOR2_X1 U23381 ( .A1(n20474), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20476) );
  AOI22_X1 U23382 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20494), .B1(
        n20493), .B2(n20829), .ZN(n20477) );
  OAI211_X1 U23383 ( .C1(n20832), .C2(n20520), .A(n20478), .B(n20477), .ZN(
        P1_U3065) );
  AOI22_X1 U23384 ( .A1(n20834), .A2(n20491), .B1(n20833), .B2(n20492), .ZN(
        n20480) );
  AOI22_X1 U23385 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20494), .B1(
        n20493), .B2(n20792), .ZN(n20479) );
  OAI211_X1 U23386 ( .C1(n20795), .C2(n20520), .A(n20480), .B(n20479), .ZN(
        P1_U3066) );
  AOI22_X1 U23387 ( .A1(n20840), .A2(n20491), .B1(n20839), .B2(n20492), .ZN(
        n20482) );
  AOI22_X1 U23388 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20494), .B1(
        n20493), .B2(n20796), .ZN(n20481) );
  OAI211_X1 U23389 ( .C1(n20799), .C2(n20520), .A(n20482), .B(n20481), .ZN(
        P1_U3067) );
  AOI22_X1 U23390 ( .A1(n20846), .A2(n20491), .B1(n20845), .B2(n20492), .ZN(
        n20484) );
  AOI22_X1 U23391 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20494), .B1(
        n20493), .B2(n20847), .ZN(n20483) );
  OAI211_X1 U23392 ( .C1(n20850), .C2(n20520), .A(n20484), .B(n20483), .ZN(
        P1_U3068) );
  AOI22_X1 U23393 ( .A1(n20852), .A2(n20492), .B1(n20491), .B2(n20851), .ZN(
        n20486) );
  AOI22_X1 U23394 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20494), .B1(
        n20493), .B2(n20853), .ZN(n20485) );
  OAI211_X1 U23395 ( .C1(n20856), .C2(n20520), .A(n20486), .B(n20485), .ZN(
        P1_U3069) );
  AOI22_X1 U23396 ( .A1(n20858), .A2(n20492), .B1(n20491), .B2(n20857), .ZN(
        n20488) );
  AOI22_X1 U23397 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20494), .B1(
        n20493), .B2(n20859), .ZN(n20487) );
  OAI211_X1 U23398 ( .C1(n20862), .C2(n20520), .A(n20488), .B(n20487), .ZN(
        P1_U3070) );
  AOI22_X1 U23399 ( .A1(n20864), .A2(n20492), .B1(n20491), .B2(n20863), .ZN(
        n20490) );
  AOI22_X1 U23400 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20494), .B1(
        n20493), .B2(n20865), .ZN(n20489) );
  OAI211_X1 U23401 ( .C1(n20870), .C2(n20520), .A(n20490), .B(n20489), .ZN(
        P1_U3071) );
  AOI22_X1 U23402 ( .A1(n20874), .A2(n20492), .B1(n20491), .B2(n20871), .ZN(
        n20496) );
  AOI22_X1 U23403 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20494), .B1(
        n20493), .B2(n20810), .ZN(n20495) );
  OAI211_X1 U23404 ( .C1(n20815), .C2(n20520), .A(n20496), .B(n20495), .ZN(
        P1_U3072) );
  INV_X1 U23405 ( .A(n20829), .ZN(n20678) );
  NOR2_X1 U23406 ( .A1(n20751), .A2(n20497), .ZN(n20516) );
  AOI21_X1 U23407 ( .B1(n20550), .B2(n20608), .A(n20516), .ZN(n20498) );
  OAI22_X1 U23408 ( .A1(n20498), .A2(n20817), .B1(n20497), .B2(n20968), .ZN(
        n20515) );
  AOI22_X1 U23409 ( .A1(n20821), .A2(n20515), .B1(n20820), .B2(n20516), .ZN(
        n20502) );
  OAI21_X1 U23410 ( .B1(n20553), .B2(n21106), .A(n20498), .ZN(n20499) );
  OAI221_X1 U23411 ( .B1(n20823), .B2(n20500), .C1(n20817), .C2(n20499), .A(
        n20827), .ZN(n20517) );
  AOI22_X1 U23412 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20517), .B1(
        n20543), .B2(n20711), .ZN(n20501) );
  OAI211_X1 U23413 ( .C1(n20678), .C2(n20520), .A(n20502), .B(n20501), .ZN(
        P1_U3073) );
  INV_X1 U23414 ( .A(n20792), .ZN(n20838) );
  AOI22_X1 U23415 ( .A1(n20834), .A2(n20515), .B1(n20833), .B2(n20516), .ZN(
        n20504) );
  AOI22_X1 U23416 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20517), .B1(
        n20543), .B2(n20835), .ZN(n20503) );
  OAI211_X1 U23417 ( .C1(n20838), .C2(n20520), .A(n20504), .B(n20503), .ZN(
        P1_U3074) );
  INV_X1 U23418 ( .A(n20796), .ZN(n20844) );
  AOI22_X1 U23419 ( .A1(n20840), .A2(n20515), .B1(n20839), .B2(n20516), .ZN(
        n20506) );
  AOI22_X1 U23420 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20517), .B1(
        n20543), .B2(n20841), .ZN(n20505) );
  OAI211_X1 U23421 ( .C1(n20844), .C2(n20520), .A(n20506), .B(n20505), .ZN(
        P1_U3075) );
  INV_X1 U23422 ( .A(n20847), .ZN(n20685) );
  AOI22_X1 U23423 ( .A1(n20846), .A2(n20515), .B1(n20845), .B2(n20516), .ZN(
        n20508) );
  AOI22_X1 U23424 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20517), .B1(
        n20543), .B2(n20726), .ZN(n20507) );
  OAI211_X1 U23425 ( .C1(n20685), .C2(n20520), .A(n20508), .B(n20507), .ZN(
        P1_U3076) );
  INV_X1 U23426 ( .A(n20853), .ZN(n20688) );
  AOI22_X1 U23427 ( .A1(n20852), .A2(n20516), .B1(n20515), .B2(n20851), .ZN(
        n20510) );
  AOI22_X1 U23428 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20517), .B1(
        n20543), .B2(n20730), .ZN(n20509) );
  OAI211_X1 U23429 ( .C1(n20688), .C2(n20520), .A(n20510), .B(n20509), .ZN(
        P1_U3077) );
  INV_X1 U23430 ( .A(n20859), .ZN(n20691) );
  AOI22_X1 U23431 ( .A1(n20858), .A2(n20516), .B1(n20515), .B2(n20857), .ZN(
        n20512) );
  AOI22_X1 U23432 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20517), .B1(
        n20543), .B2(n20734), .ZN(n20511) );
  OAI211_X1 U23433 ( .C1(n20691), .C2(n20520), .A(n20512), .B(n20511), .ZN(
        P1_U3078) );
  INV_X1 U23434 ( .A(n20865), .ZN(n20694) );
  AOI22_X1 U23435 ( .A1(n20864), .A2(n20516), .B1(n20515), .B2(n20863), .ZN(
        n20514) );
  AOI22_X1 U23436 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20517), .B1(
        n20543), .B2(n20738), .ZN(n20513) );
  OAI211_X1 U23437 ( .C1(n20694), .C2(n20520), .A(n20514), .B(n20513), .ZN(
        P1_U3079) );
  INV_X1 U23438 ( .A(n20810), .ZN(n20881) );
  AOI22_X1 U23439 ( .A1(n20874), .A2(n20516), .B1(n20515), .B2(n20871), .ZN(
        n20519) );
  AOI22_X1 U23440 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20517), .B1(
        n20543), .B2(n20875), .ZN(n20518) );
  OAI211_X1 U23441 ( .C1(n20881), .C2(n20520), .A(n20519), .B(n20518), .ZN(
        P1_U3080) );
  INV_X1 U23442 ( .A(n20543), .ZN(n20521) );
  NAND2_X1 U23443 ( .A1(n20521), .A2(n20823), .ZN(n20522) );
  NOR2_X2 U23444 ( .A1(n20553), .A2(n20778), .ZN(n20572) );
  OAI21_X1 U23445 ( .B1(n20522), .B2(n20572), .A(n20705), .ZN(n20526) );
  AND2_X1 U23446 ( .A1(n20550), .A2(n20783), .ZN(n20523) );
  NOR2_X1 U23447 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20551), .ZN(
        n20542) );
  AOI22_X1 U23448 ( .A1(n20572), .A2(n20711), .B1(n20820), .B2(n20542), .ZN(
        n20529) );
  INV_X1 U23449 ( .A(n20523), .ZN(n20525) );
  AOI21_X1 U23450 ( .B1(n20526), .B2(n20525), .A(n20524), .ZN(n20527) );
  OAI211_X1 U23451 ( .C1(n20542), .C2(n11516), .A(n20787), .B(n20527), .ZN(
        n20544) );
  AOI22_X1 U23452 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20829), .ZN(n20528) );
  OAI211_X1 U23453 ( .C1(n20547), .C2(n20719), .A(n20529), .B(n20528), .ZN(
        P1_U3081) );
  AOI22_X1 U23454 ( .A1(n20572), .A2(n20835), .B1(n20833), .B2(n20542), .ZN(
        n20531) );
  AOI22_X1 U23455 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20792), .ZN(n20530) );
  OAI211_X1 U23456 ( .C1(n20547), .C2(n20722), .A(n20531), .B(n20530), .ZN(
        P1_U3082) );
  AOI22_X1 U23457 ( .A1(n20572), .A2(n20841), .B1(n20839), .B2(n20542), .ZN(
        n20533) );
  AOI22_X1 U23458 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20796), .ZN(n20532) );
  OAI211_X1 U23459 ( .C1(n20547), .C2(n20725), .A(n20533), .B(n20532), .ZN(
        P1_U3083) );
  AOI22_X1 U23460 ( .A1(n20572), .A2(n20726), .B1(n20845), .B2(n20542), .ZN(
        n20535) );
  AOI22_X1 U23461 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20847), .ZN(n20534) );
  OAI211_X1 U23462 ( .C1(n20547), .C2(n20729), .A(n20535), .B(n20534), .ZN(
        P1_U3084) );
  AOI22_X1 U23463 ( .A1(n20572), .A2(n20730), .B1(n20852), .B2(n20542), .ZN(
        n20537) );
  AOI22_X1 U23464 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20853), .ZN(n20536) );
  OAI211_X1 U23465 ( .C1(n20547), .C2(n20733), .A(n20537), .B(n20536), .ZN(
        P1_U3085) );
  AOI22_X1 U23466 ( .A1(n20572), .A2(n20734), .B1(n20858), .B2(n20542), .ZN(
        n20539) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20859), .ZN(n20538) );
  OAI211_X1 U23468 ( .C1(n20547), .C2(n20737), .A(n20539), .B(n20538), .ZN(
        P1_U3086) );
  AOI22_X1 U23469 ( .A1(n20543), .A2(n20865), .B1(n20864), .B2(n20542), .ZN(
        n20541) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20544), .B1(
        n20572), .B2(n20738), .ZN(n20540) );
  OAI211_X1 U23471 ( .C1(n20547), .C2(n20741), .A(n20541), .B(n20540), .ZN(
        P1_U3087) );
  AOI22_X1 U23472 ( .A1(n20543), .A2(n20810), .B1(n20874), .B2(n20542), .ZN(
        n20546) );
  AOI22_X1 U23473 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20544), .B1(
        n20572), .B2(n20875), .ZN(n20545) );
  OAI211_X1 U23474 ( .C1(n20547), .C2(n20747), .A(n20546), .B(n20545), .ZN(
        P1_U3088) );
  AOI21_X1 U23475 ( .B1(n20550), .B2(n20667), .A(n20571), .ZN(n20552) );
  OAI22_X1 U23476 ( .A1(n20552), .A2(n20817), .B1(n20551), .B2(n20968), .ZN(
        n20570) );
  AOI22_X1 U23477 ( .A1(n20821), .A2(n20570), .B1(n20820), .B2(n20571), .ZN(
        n20557) );
  INV_X1 U23478 ( .A(n20551), .ZN(n20555) );
  OAI211_X1 U23479 ( .C1(n20553), .C2(n20671), .A(n20823), .B(n20552), .ZN(
        n20554) );
  OAI211_X1 U23480 ( .C1(n20823), .C2(n20555), .A(n20827), .B(n20554), .ZN(
        n20573) );
  AOI22_X1 U23481 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20573), .B1(
        n20572), .B2(n20829), .ZN(n20556) );
  OAI211_X1 U23482 ( .C1(n20832), .C2(n20583), .A(n20557), .B(n20556), .ZN(
        P1_U3089) );
  AOI22_X1 U23483 ( .A1(n20834), .A2(n20570), .B1(n20833), .B2(n20571), .ZN(
        n20559) );
  AOI22_X1 U23484 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20573), .B1(
        n20572), .B2(n20792), .ZN(n20558) );
  OAI211_X1 U23485 ( .C1(n20795), .C2(n20583), .A(n20559), .B(n20558), .ZN(
        P1_U3090) );
  AOI22_X1 U23486 ( .A1(n20840), .A2(n20570), .B1(n20839), .B2(n20571), .ZN(
        n20561) );
  AOI22_X1 U23487 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20573), .B1(
        n20572), .B2(n20796), .ZN(n20560) );
  OAI211_X1 U23488 ( .C1(n20799), .C2(n20583), .A(n20561), .B(n20560), .ZN(
        P1_U3091) );
  AOI22_X1 U23489 ( .A1(n20846), .A2(n20570), .B1(n20845), .B2(n20571), .ZN(
        n20563) );
  AOI22_X1 U23490 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20573), .B1(
        n20572), .B2(n20847), .ZN(n20562) );
  OAI211_X1 U23491 ( .C1(n20850), .C2(n20583), .A(n20563), .B(n20562), .ZN(
        P1_U3092) );
  AOI22_X1 U23492 ( .A1(n20852), .A2(n20571), .B1(n20570), .B2(n20851), .ZN(
        n20565) );
  AOI22_X1 U23493 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20573), .B1(
        n20572), .B2(n20853), .ZN(n20564) );
  OAI211_X1 U23494 ( .C1(n20856), .C2(n20583), .A(n20565), .B(n20564), .ZN(
        P1_U3093) );
  AOI22_X1 U23495 ( .A1(n20858), .A2(n20571), .B1(n20570), .B2(n20857), .ZN(
        n20567) );
  AOI22_X1 U23496 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20573), .B1(
        n20572), .B2(n20859), .ZN(n20566) );
  OAI211_X1 U23497 ( .C1(n20862), .C2(n20583), .A(n20567), .B(n20566), .ZN(
        P1_U3094) );
  AOI22_X1 U23498 ( .A1(n20864), .A2(n20571), .B1(n20570), .B2(n20863), .ZN(
        n20569) );
  AOI22_X1 U23499 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20573), .B1(
        n20572), .B2(n20865), .ZN(n20568) );
  OAI211_X1 U23500 ( .C1(n20870), .C2(n20583), .A(n20569), .B(n20568), .ZN(
        P1_U3095) );
  AOI22_X1 U23501 ( .A1(n20874), .A2(n20571), .B1(n20570), .B2(n20871), .ZN(
        n20575) );
  AOI22_X1 U23502 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20573), .B1(
        n20572), .B2(n20810), .ZN(n20574) );
  OAI211_X1 U23503 ( .C1(n20815), .C2(n20583), .A(n20575), .B(n20574), .ZN(
        P1_U3096) );
  INV_X1 U23504 ( .A(n20675), .ZN(n20577) );
  AND2_X1 U23505 ( .A1(n20578), .A2(n13690), .ZN(n20668) );
  NOR3_X1 U23506 ( .A1(n20710), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20612) );
  INV_X1 U23507 ( .A(n20612), .ZN(n20609) );
  NOR2_X1 U23508 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20609), .ZN(
        n20603) );
  AOI21_X1 U23509 ( .B1(n20668), .B2(n13673), .A(n20603), .ZN(n20585) );
  INV_X1 U23510 ( .A(n20579), .ZN(n20581) );
  NOR2_X1 U23511 ( .A1(n20581), .A2(n20580), .ZN(n20708) );
  INV_X1 U23512 ( .A(n20708), .ZN(n20713) );
  OAI22_X1 U23513 ( .A1(n20585), .A2(n20817), .B1(n20582), .B2(n20713), .ZN(
        n20602) );
  AOI22_X1 U23514 ( .A1(n20821), .A2(n20602), .B1(n20820), .B2(n20603), .ZN(
        n20589) );
  INV_X1 U23515 ( .A(n20632), .ZN(n20584) );
  OAI21_X1 U23516 ( .B1(n20584), .B2(n20604), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20586) );
  NAND2_X1 U23517 ( .A1(n20586), .A2(n20585), .ZN(n20587) );
  AOI22_X1 U23518 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20605), .B1(
        n20604), .B2(n20829), .ZN(n20588) );
  OAI211_X1 U23519 ( .C1(n20832), .C2(n20632), .A(n20589), .B(n20588), .ZN(
        P1_U3097) );
  AOI22_X1 U23520 ( .A1(n20834), .A2(n20602), .B1(n20833), .B2(n20603), .ZN(
        n20591) );
  AOI22_X1 U23521 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20605), .B1(
        n20604), .B2(n20792), .ZN(n20590) );
  OAI211_X1 U23522 ( .C1(n20795), .C2(n20632), .A(n20591), .B(n20590), .ZN(
        P1_U3098) );
  AOI22_X1 U23523 ( .A1(n20840), .A2(n20602), .B1(n20839), .B2(n20603), .ZN(
        n20593) );
  AOI22_X1 U23524 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20605), .B1(
        n20604), .B2(n20796), .ZN(n20592) );
  OAI211_X1 U23525 ( .C1(n20799), .C2(n20632), .A(n20593), .B(n20592), .ZN(
        P1_U3099) );
  AOI22_X1 U23526 ( .A1(n20846), .A2(n20602), .B1(n20845), .B2(n20603), .ZN(
        n20595) );
  AOI22_X1 U23527 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20605), .B1(
        n20604), .B2(n20847), .ZN(n20594) );
  OAI211_X1 U23528 ( .C1(n20850), .C2(n20632), .A(n20595), .B(n20594), .ZN(
        P1_U3100) );
  AOI22_X1 U23529 ( .A1(n20852), .A2(n20603), .B1(n20602), .B2(n20851), .ZN(
        n20597) );
  AOI22_X1 U23530 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20605), .B1(
        n20604), .B2(n20853), .ZN(n20596) );
  OAI211_X1 U23531 ( .C1(n20856), .C2(n20632), .A(n20597), .B(n20596), .ZN(
        P1_U3101) );
  AOI22_X1 U23532 ( .A1(n20858), .A2(n20603), .B1(n20602), .B2(n20857), .ZN(
        n20599) );
  AOI22_X1 U23533 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20605), .B1(
        n20604), .B2(n20859), .ZN(n20598) );
  OAI211_X1 U23534 ( .C1(n20862), .C2(n20632), .A(n20599), .B(n20598), .ZN(
        P1_U3102) );
  AOI22_X1 U23535 ( .A1(n20864), .A2(n20603), .B1(n20602), .B2(n20863), .ZN(
        n20601) );
  AOI22_X1 U23536 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20605), .B1(
        n20604), .B2(n20865), .ZN(n20600) );
  OAI211_X1 U23537 ( .C1(n20870), .C2(n20632), .A(n20601), .B(n20600), .ZN(
        P1_U3103) );
  AOI22_X1 U23538 ( .A1(n20874), .A2(n20603), .B1(n20602), .B2(n20871), .ZN(
        n20607) );
  AOI22_X1 U23539 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20605), .B1(
        n20604), .B2(n20810), .ZN(n20606) );
  OAI211_X1 U23540 ( .C1(n20815), .C2(n20632), .A(n20607), .B(n20606), .ZN(
        P1_U3104) );
  NOR2_X1 U23541 ( .A1(n20751), .A2(n20609), .ZN(n20628) );
  AOI21_X1 U23542 ( .B1(n20668), .B2(n20608), .A(n20628), .ZN(n20610) );
  OAI22_X1 U23543 ( .A1(n20610), .A2(n20817), .B1(n20609), .B2(n20968), .ZN(
        n20627) );
  AOI22_X1 U23544 ( .A1(n20821), .A2(n20627), .B1(n20820), .B2(n20628), .ZN(
        n20614) );
  OAI21_X1 U23545 ( .B1(n20675), .B2(n21106), .A(n20610), .ZN(n20611) );
  OAI221_X1 U23546 ( .B1(n20823), .B2(n20612), .C1(n20817), .C2(n20611), .A(
        n20827), .ZN(n20629) );
  AOI22_X1 U23547 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20629), .B1(
        n20661), .B2(n20711), .ZN(n20613) );
  OAI211_X1 U23548 ( .C1(n20678), .C2(n20632), .A(n20614), .B(n20613), .ZN(
        P1_U3105) );
  AOI22_X1 U23549 ( .A1(n20834), .A2(n20627), .B1(n20833), .B2(n20628), .ZN(
        n20616) );
  AOI22_X1 U23550 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20629), .B1(
        n20661), .B2(n20835), .ZN(n20615) );
  OAI211_X1 U23551 ( .C1(n20838), .C2(n20632), .A(n20616), .B(n20615), .ZN(
        P1_U3106) );
  AOI22_X1 U23552 ( .A1(n20840), .A2(n20627), .B1(n20839), .B2(n20628), .ZN(
        n20618) );
  AOI22_X1 U23553 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20629), .B1(
        n20661), .B2(n20841), .ZN(n20617) );
  OAI211_X1 U23554 ( .C1(n20844), .C2(n20632), .A(n20618), .B(n20617), .ZN(
        P1_U3107) );
  AOI22_X1 U23555 ( .A1(n20846), .A2(n20627), .B1(n20845), .B2(n20628), .ZN(
        n20620) );
  AOI22_X1 U23556 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20629), .B1(
        n20661), .B2(n20726), .ZN(n20619) );
  OAI211_X1 U23557 ( .C1(n20685), .C2(n20632), .A(n20620), .B(n20619), .ZN(
        P1_U3108) );
  AOI22_X1 U23558 ( .A1(n20852), .A2(n20628), .B1(n20627), .B2(n20851), .ZN(
        n20622) );
  AOI22_X1 U23559 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20629), .B1(
        n20661), .B2(n20730), .ZN(n20621) );
  OAI211_X1 U23560 ( .C1(n20688), .C2(n20632), .A(n20622), .B(n20621), .ZN(
        P1_U3109) );
  AOI22_X1 U23561 ( .A1(n20858), .A2(n20628), .B1(n20627), .B2(n20857), .ZN(
        n20624) );
  AOI22_X1 U23562 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20629), .B1(
        n20661), .B2(n20734), .ZN(n20623) );
  OAI211_X1 U23563 ( .C1(n20691), .C2(n20632), .A(n20624), .B(n20623), .ZN(
        P1_U3110) );
  AOI22_X1 U23564 ( .A1(n20864), .A2(n20628), .B1(n20627), .B2(n20863), .ZN(
        n20626) );
  AOI22_X1 U23565 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20629), .B1(
        n20661), .B2(n20738), .ZN(n20625) );
  OAI211_X1 U23566 ( .C1(n20694), .C2(n20632), .A(n20626), .B(n20625), .ZN(
        P1_U3111) );
  AOI22_X1 U23567 ( .A1(n20874), .A2(n20628), .B1(n20627), .B2(n20871), .ZN(
        n20631) );
  AOI22_X1 U23568 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20629), .B1(
        n20661), .B2(n20875), .ZN(n20630) );
  OAI211_X1 U23569 ( .C1(n20881), .C2(n20632), .A(n20631), .B(n20630), .ZN(
        P1_U3112) );
  NAND3_X1 U23570 ( .A1(n20700), .A2(n20633), .A3(n20823), .ZN(n20634) );
  NAND2_X1 U23571 ( .A1(n20634), .A2(n20705), .ZN(n20643) );
  AND2_X1 U23572 ( .A1(n20668), .A2(n20783), .ZN(n20639) );
  OR2_X1 U23573 ( .A1(n20635), .A2(n20710), .ZN(n20781) );
  INV_X1 U23574 ( .A(n20781), .ZN(n20636) );
  NOR3_X1 U23575 ( .A1(n20710), .A2(n20638), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20673) );
  INV_X1 U23576 ( .A(n20673), .ZN(n20669) );
  NOR2_X1 U23577 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20669), .ZN(
        n20659) );
  AOI22_X1 U23578 ( .A1(n20661), .A2(n20829), .B1(n20820), .B2(n20659), .ZN(
        n20646) );
  INV_X1 U23579 ( .A(n20639), .ZN(n20642) );
  NAND2_X1 U23580 ( .A1(n20781), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20786) );
  OAI211_X1 U23581 ( .C1(n11516), .C2(n20659), .A(n20786), .B(n20640), .ZN(
        n20641) );
  AOI21_X1 U23582 ( .B1(n20643), .B2(n20642), .A(n20641), .ZN(n20644) );
  AOI22_X1 U23583 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20662), .B1(
        n20660), .B2(n20711), .ZN(n20645) );
  OAI211_X1 U23584 ( .C1(n20665), .C2(n20719), .A(n20646), .B(n20645), .ZN(
        P1_U3113) );
  AOI22_X1 U23585 ( .A1(n20660), .A2(n20835), .B1(n20833), .B2(n20659), .ZN(
        n20648) );
  AOI22_X1 U23586 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20662), .B1(
        n20661), .B2(n20792), .ZN(n20647) );
  OAI211_X1 U23587 ( .C1(n20665), .C2(n20722), .A(n20648), .B(n20647), .ZN(
        P1_U3114) );
  AOI22_X1 U23588 ( .A1(n20660), .A2(n20841), .B1(n20839), .B2(n20659), .ZN(
        n20650) );
  AOI22_X1 U23589 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20662), .B1(
        n20661), .B2(n20796), .ZN(n20649) );
  OAI211_X1 U23590 ( .C1(n20665), .C2(n20725), .A(n20650), .B(n20649), .ZN(
        P1_U3115) );
  AOI22_X1 U23591 ( .A1(n20661), .A2(n20847), .B1(n20845), .B2(n20659), .ZN(
        n20652) );
  AOI22_X1 U23592 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20662), .B1(
        n20660), .B2(n20726), .ZN(n20651) );
  OAI211_X1 U23593 ( .C1(n20665), .C2(n20729), .A(n20652), .B(n20651), .ZN(
        P1_U3116) );
  AOI22_X1 U23594 ( .A1(n20661), .A2(n20853), .B1(n20852), .B2(n20659), .ZN(
        n20654) );
  AOI22_X1 U23595 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20662), .B1(
        n20660), .B2(n20730), .ZN(n20653) );
  OAI211_X1 U23596 ( .C1(n20665), .C2(n20733), .A(n20654), .B(n20653), .ZN(
        P1_U3117) );
  AOI22_X1 U23597 ( .A1(n20661), .A2(n20859), .B1(n20858), .B2(n20659), .ZN(
        n20656) );
  AOI22_X1 U23598 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20662), .B1(
        n20660), .B2(n20734), .ZN(n20655) );
  OAI211_X1 U23599 ( .C1(n20665), .C2(n20737), .A(n20656), .B(n20655), .ZN(
        P1_U3118) );
  AOI22_X1 U23600 ( .A1(n20661), .A2(n20865), .B1(n20864), .B2(n20659), .ZN(
        n20658) );
  AOI22_X1 U23601 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20662), .B1(
        n20660), .B2(n20738), .ZN(n20657) );
  OAI211_X1 U23602 ( .C1(n20665), .C2(n20741), .A(n20658), .B(n20657), .ZN(
        P1_U3119) );
  AOI22_X1 U23603 ( .A1(n20660), .A2(n20875), .B1(n20874), .B2(n20659), .ZN(
        n20664) );
  AOI22_X1 U23604 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20662), .B1(
        n20661), .B2(n20810), .ZN(n20663) );
  OAI211_X1 U23605 ( .C1(n20665), .C2(n20747), .A(n20664), .B(n20663), .ZN(
        P1_U3120) );
  NOR2_X1 U23606 ( .A1(n20666), .A2(n20710), .ZN(n20696) );
  AOI21_X1 U23607 ( .B1(n20668), .B2(n20667), .A(n20696), .ZN(n20670) );
  OAI22_X1 U23608 ( .A1(n20670), .A2(n20817), .B1(n20669), .B2(n20968), .ZN(
        n20695) );
  AOI22_X1 U23609 ( .A1(n20821), .A2(n20695), .B1(n20820), .B2(n20696), .ZN(
        n20677) );
  OAI21_X1 U23610 ( .B1(n20675), .B2(n20671), .A(n20670), .ZN(n20672) );
  OAI221_X1 U23611 ( .B1(n20823), .B2(n20673), .C1(n20817), .C2(n20672), .A(
        n20827), .ZN(n20697) );
  AOI22_X1 U23612 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20697), .B1(
        n20743), .B2(n20711), .ZN(n20676) );
  OAI211_X1 U23613 ( .C1(n20678), .C2(n20700), .A(n20677), .B(n20676), .ZN(
        P1_U3121) );
  AOI22_X1 U23614 ( .A1(n20834), .A2(n20695), .B1(n20833), .B2(n20696), .ZN(
        n20680) );
  AOI22_X1 U23615 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20697), .B1(
        n20743), .B2(n20835), .ZN(n20679) );
  OAI211_X1 U23616 ( .C1(n20838), .C2(n20700), .A(n20680), .B(n20679), .ZN(
        P1_U3122) );
  AOI22_X1 U23617 ( .A1(n20840), .A2(n20695), .B1(n20839), .B2(n20696), .ZN(
        n20682) );
  AOI22_X1 U23618 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20697), .B1(
        n20743), .B2(n20841), .ZN(n20681) );
  OAI211_X1 U23619 ( .C1(n20844), .C2(n20700), .A(n20682), .B(n20681), .ZN(
        P1_U3123) );
  AOI22_X1 U23620 ( .A1(n20846), .A2(n20695), .B1(n20845), .B2(n20696), .ZN(
        n20684) );
  AOI22_X1 U23621 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20697), .B1(
        n20743), .B2(n20726), .ZN(n20683) );
  OAI211_X1 U23622 ( .C1(n20685), .C2(n20700), .A(n20684), .B(n20683), .ZN(
        P1_U3124) );
  AOI22_X1 U23623 ( .A1(n20852), .A2(n20696), .B1(n20695), .B2(n20851), .ZN(
        n20687) );
  AOI22_X1 U23624 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20697), .B1(
        n20743), .B2(n20730), .ZN(n20686) );
  OAI211_X1 U23625 ( .C1(n20688), .C2(n20700), .A(n20687), .B(n20686), .ZN(
        P1_U3125) );
  AOI22_X1 U23626 ( .A1(n20858), .A2(n20696), .B1(n20695), .B2(n20857), .ZN(
        n20690) );
  AOI22_X1 U23627 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20697), .B1(
        n20743), .B2(n20734), .ZN(n20689) );
  OAI211_X1 U23628 ( .C1(n20691), .C2(n20700), .A(n20690), .B(n20689), .ZN(
        P1_U3126) );
  AOI22_X1 U23629 ( .A1(n20864), .A2(n20696), .B1(n20695), .B2(n20863), .ZN(
        n20693) );
  AOI22_X1 U23630 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20697), .B1(
        n20743), .B2(n20738), .ZN(n20692) );
  OAI211_X1 U23631 ( .C1(n20694), .C2(n20700), .A(n20693), .B(n20692), .ZN(
        P1_U3127) );
  AOI22_X1 U23632 ( .A1(n20874), .A2(n20696), .B1(n20695), .B2(n20871), .ZN(
        n20699) );
  AOI22_X1 U23633 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20697), .B1(
        n20743), .B2(n20875), .ZN(n20698) );
  OAI211_X1 U23634 ( .C1(n20881), .C2(n20700), .A(n20699), .B(n20698), .ZN(
        P1_U3128) );
  INV_X1 U23635 ( .A(n20774), .ZN(n20704) );
  NAND3_X1 U23636 ( .A1(n20704), .A2(n20823), .A3(n20703), .ZN(n20706) );
  NAND2_X1 U23637 ( .A1(n20706), .A2(n20705), .ZN(n20715) );
  OR2_X1 U23638 ( .A1(n13690), .A2(n20707), .ZN(n20752) );
  NOR2_X1 U23639 ( .A1(n20752), .A2(n20783), .ZN(n20712) );
  NOR3_X1 U23640 ( .A1(n11776), .A2(n20710), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20756) );
  INV_X1 U23641 ( .A(n20756), .ZN(n20754) );
  NOR2_X1 U23642 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20754), .ZN(
        n20742) );
  AOI22_X1 U23643 ( .A1(n20774), .A2(n20711), .B1(n20820), .B2(n20742), .ZN(
        n20718) );
  INV_X1 U23644 ( .A(n20712), .ZN(n20714) );
  AOI22_X1 U23645 ( .A1(n20715), .A2(n20714), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20713), .ZN(n20716) );
  OAI211_X1 U23646 ( .C1(n20742), .C2(n11516), .A(n20787), .B(n20716), .ZN(
        n20744) );
  AOI22_X1 U23647 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20744), .B1(
        n20743), .B2(n20829), .ZN(n20717) );
  OAI211_X1 U23648 ( .C1(n20748), .C2(n20719), .A(n20718), .B(n20717), .ZN(
        P1_U3129) );
  AOI22_X1 U23649 ( .A1(n20774), .A2(n20835), .B1(n20833), .B2(n20742), .ZN(
        n20721) );
  AOI22_X1 U23650 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20744), .B1(
        n20743), .B2(n20792), .ZN(n20720) );
  OAI211_X1 U23651 ( .C1(n20748), .C2(n20722), .A(n20721), .B(n20720), .ZN(
        P1_U3130) );
  AOI22_X1 U23652 ( .A1(n20774), .A2(n20841), .B1(n20839), .B2(n20742), .ZN(
        n20724) );
  AOI22_X1 U23653 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20744), .B1(
        n20743), .B2(n20796), .ZN(n20723) );
  OAI211_X1 U23654 ( .C1(n20748), .C2(n20725), .A(n20724), .B(n20723), .ZN(
        P1_U3131) );
  AOI22_X1 U23655 ( .A1(n20774), .A2(n20726), .B1(n20845), .B2(n20742), .ZN(
        n20728) );
  AOI22_X1 U23656 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20744), .B1(
        n20743), .B2(n20847), .ZN(n20727) );
  OAI211_X1 U23657 ( .C1(n20748), .C2(n20729), .A(n20728), .B(n20727), .ZN(
        P1_U3132) );
  AOI22_X1 U23658 ( .A1(n20774), .A2(n20730), .B1(n20852), .B2(n20742), .ZN(
        n20732) );
  AOI22_X1 U23659 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20744), .B1(
        n20743), .B2(n20853), .ZN(n20731) );
  OAI211_X1 U23660 ( .C1(n20748), .C2(n20733), .A(n20732), .B(n20731), .ZN(
        P1_U3133) );
  AOI22_X1 U23661 ( .A1(n20774), .A2(n20734), .B1(n20858), .B2(n20742), .ZN(
        n20736) );
  AOI22_X1 U23662 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20744), .B1(
        n20743), .B2(n20859), .ZN(n20735) );
  OAI211_X1 U23663 ( .C1(n20748), .C2(n20737), .A(n20736), .B(n20735), .ZN(
        P1_U3134) );
  AOI22_X1 U23664 ( .A1(n20774), .A2(n20738), .B1(n20864), .B2(n20742), .ZN(
        n20740) );
  AOI22_X1 U23665 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20744), .B1(
        n20743), .B2(n20865), .ZN(n20739) );
  OAI211_X1 U23666 ( .C1(n20748), .C2(n20741), .A(n20740), .B(n20739), .ZN(
        P1_U3135) );
  AOI22_X1 U23667 ( .A1(n20774), .A2(n20875), .B1(n20874), .B2(n20742), .ZN(
        n20746) );
  AOI22_X1 U23668 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20744), .B1(
        n20743), .B2(n20810), .ZN(n20745) );
  OAI211_X1 U23669 ( .C1(n20748), .C2(n20747), .A(n20746), .B(n20745), .ZN(
        P1_U3136) );
  INV_X1 U23670 ( .A(n20749), .ZN(n20750) );
  NOR2_X1 U23671 ( .A1(n20751), .A2(n20754), .ZN(n20773) );
  INV_X1 U23672 ( .A(n20773), .ZN(n20755) );
  INV_X1 U23673 ( .A(n20752), .ZN(n20784) );
  NAND2_X1 U23674 ( .A1(n20784), .A2(n20823), .ZN(n20819) );
  OAI222_X1 U23675 ( .A1(n20755), .A2(n20817), .B1(n20968), .B2(n20754), .C1(
        n20753), .C2(n20819), .ZN(n20772) );
  AOI22_X1 U23676 ( .A1(n20821), .A2(n20772), .B1(n20820), .B2(n20773), .ZN(
        n20759) );
  OAI21_X1 U23677 ( .B1(n20757), .B2(n20756), .A(n20827), .ZN(n20775) );
  AOI22_X1 U23678 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20775), .B1(
        n20774), .B2(n20829), .ZN(n20758) );
  OAI211_X1 U23679 ( .C1(n20832), .C2(n20789), .A(n20759), .B(n20758), .ZN(
        P1_U3137) );
  AOI22_X1 U23680 ( .A1(n20834), .A2(n20772), .B1(n20833), .B2(n20773), .ZN(
        n20761) );
  AOI22_X1 U23681 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20775), .B1(
        n20774), .B2(n20792), .ZN(n20760) );
  OAI211_X1 U23682 ( .C1(n20795), .C2(n20789), .A(n20761), .B(n20760), .ZN(
        P1_U3138) );
  AOI22_X1 U23683 ( .A1(n20840), .A2(n20772), .B1(n20839), .B2(n20773), .ZN(
        n20763) );
  AOI22_X1 U23684 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20775), .B1(
        n20774), .B2(n20796), .ZN(n20762) );
  OAI211_X1 U23685 ( .C1(n20799), .C2(n20789), .A(n20763), .B(n20762), .ZN(
        P1_U3139) );
  AOI22_X1 U23686 ( .A1(n20846), .A2(n20772), .B1(n20845), .B2(n20773), .ZN(
        n20765) );
  AOI22_X1 U23687 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20775), .B1(
        n20774), .B2(n20847), .ZN(n20764) );
  OAI211_X1 U23688 ( .C1(n20850), .C2(n20789), .A(n20765), .B(n20764), .ZN(
        P1_U3140) );
  AOI22_X1 U23689 ( .A1(n20852), .A2(n20773), .B1(n20772), .B2(n20851), .ZN(
        n20767) );
  AOI22_X1 U23690 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20775), .B1(
        n20774), .B2(n20853), .ZN(n20766) );
  OAI211_X1 U23691 ( .C1(n20856), .C2(n20789), .A(n20767), .B(n20766), .ZN(
        P1_U3141) );
  AOI22_X1 U23692 ( .A1(n20858), .A2(n20773), .B1(n20772), .B2(n20857), .ZN(
        n20769) );
  AOI22_X1 U23693 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20775), .B1(
        n20774), .B2(n20859), .ZN(n20768) );
  OAI211_X1 U23694 ( .C1(n20862), .C2(n20789), .A(n20769), .B(n20768), .ZN(
        P1_U3142) );
  AOI22_X1 U23695 ( .A1(n20864), .A2(n20773), .B1(n20772), .B2(n20863), .ZN(
        n20771) );
  AOI22_X1 U23696 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20775), .B1(
        n20774), .B2(n20865), .ZN(n20770) );
  OAI211_X1 U23697 ( .C1(n20870), .C2(n20789), .A(n20771), .B(n20770), .ZN(
        P1_U3143) );
  AOI22_X1 U23698 ( .A1(n20874), .A2(n20773), .B1(n20772), .B2(n20871), .ZN(
        n20777) );
  AOI22_X1 U23699 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20775), .B1(
        n20774), .B2(n20810), .ZN(n20776) );
  OAI211_X1 U23700 ( .C1(n20815), .C2(n20789), .A(n20777), .B(n20776), .ZN(
        P1_U3144) );
  INV_X1 U23701 ( .A(n20778), .ZN(n20779) );
  OAI22_X1 U23702 ( .A1(n20819), .A2(n13673), .B1(n20781), .B2(n20780), .ZN(
        n20808) );
  NOR2_X1 U23703 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20825), .ZN(
        n20809) );
  AOI22_X1 U23704 ( .A1(n20821), .A2(n20808), .B1(n20820), .B2(n20809), .ZN(
        n20791) );
  AOI21_X1 U23705 ( .B1(n20880), .B2(n20789), .A(n21106), .ZN(n20782) );
  AOI21_X1 U23706 ( .B1(n20784), .B2(n20783), .A(n20782), .ZN(n20785) );
  NOR2_X1 U23707 ( .A1(n20785), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20788) );
  AOI22_X1 U23708 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20812), .B1(
        n20811), .B2(n20829), .ZN(n20790) );
  OAI211_X1 U23709 ( .C1(n20832), .C2(n20880), .A(n20791), .B(n20790), .ZN(
        P1_U3145) );
  AOI22_X1 U23710 ( .A1(n20834), .A2(n20808), .B1(n20833), .B2(n20809), .ZN(
        n20794) );
  AOI22_X1 U23711 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20812), .B1(
        n20811), .B2(n20792), .ZN(n20793) );
  OAI211_X1 U23712 ( .C1(n20795), .C2(n20880), .A(n20794), .B(n20793), .ZN(
        P1_U3146) );
  AOI22_X1 U23713 ( .A1(n20840), .A2(n20808), .B1(n20839), .B2(n20809), .ZN(
        n20798) );
  AOI22_X1 U23714 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20812), .B1(
        n20811), .B2(n20796), .ZN(n20797) );
  OAI211_X1 U23715 ( .C1(n20799), .C2(n20880), .A(n20798), .B(n20797), .ZN(
        P1_U3147) );
  AOI22_X1 U23716 ( .A1(n20846), .A2(n20808), .B1(n20845), .B2(n20809), .ZN(
        n20801) );
  AOI22_X1 U23717 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20812), .B1(
        n20811), .B2(n20847), .ZN(n20800) );
  OAI211_X1 U23718 ( .C1(n20850), .C2(n20880), .A(n20801), .B(n20800), .ZN(
        P1_U3148) );
  AOI22_X1 U23719 ( .A1(n20852), .A2(n20809), .B1(n20808), .B2(n20851), .ZN(
        n20803) );
  AOI22_X1 U23720 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20812), .B1(
        n20811), .B2(n20853), .ZN(n20802) );
  OAI211_X1 U23721 ( .C1(n20856), .C2(n20880), .A(n20803), .B(n20802), .ZN(
        P1_U3149) );
  AOI22_X1 U23722 ( .A1(n20858), .A2(n20809), .B1(n20808), .B2(n20857), .ZN(
        n20805) );
  AOI22_X1 U23723 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20812), .B1(
        n20811), .B2(n20859), .ZN(n20804) );
  OAI211_X1 U23724 ( .C1(n20862), .C2(n20880), .A(n20805), .B(n20804), .ZN(
        P1_U3150) );
  AOI22_X1 U23725 ( .A1(n20864), .A2(n20809), .B1(n20808), .B2(n20863), .ZN(
        n20807) );
  AOI22_X1 U23726 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20812), .B1(
        n20811), .B2(n20865), .ZN(n20806) );
  OAI211_X1 U23727 ( .C1(n20870), .C2(n20880), .A(n20807), .B(n20806), .ZN(
        P1_U3151) );
  AOI22_X1 U23728 ( .A1(n20874), .A2(n20809), .B1(n20808), .B2(n20871), .ZN(
        n20814) );
  AOI22_X1 U23729 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20812), .B1(
        n20811), .B2(n20810), .ZN(n20813) );
  OAI211_X1 U23730 ( .C1(n20815), .C2(n20880), .A(n20814), .B(n20813), .ZN(
        P1_U3152) );
  INV_X1 U23731 ( .A(n20873), .ZN(n20816) );
  OAI222_X1 U23732 ( .A1(n20819), .A2(n20818), .B1(n20968), .B2(n20825), .C1(
        n20817), .C2(n20816), .ZN(n20872) );
  AOI22_X1 U23733 ( .A1(n20821), .A2(n20872), .B1(n20820), .B2(n20873), .ZN(
        n20831) );
  NAND3_X1 U23734 ( .A1(n20824), .A2(n20823), .A3(n20822), .ZN(n20826) );
  NAND2_X1 U23735 ( .A1(n20826), .A2(n20825), .ZN(n20828) );
  NAND2_X1 U23736 ( .A1(n20828), .A2(n20827), .ZN(n20877) );
  INV_X1 U23737 ( .A(n20880), .ZN(n20866) );
  AOI22_X1 U23738 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20877), .B1(
        n20866), .B2(n20829), .ZN(n20830) );
  OAI211_X1 U23739 ( .C1(n20832), .C2(n20869), .A(n20831), .B(n20830), .ZN(
        P1_U3153) );
  AOI22_X1 U23740 ( .A1(n20834), .A2(n20872), .B1(n20833), .B2(n20873), .ZN(
        n20837) );
  AOI22_X1 U23741 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20877), .B1(
        n20876), .B2(n20835), .ZN(n20836) );
  OAI211_X1 U23742 ( .C1(n20838), .C2(n20880), .A(n20837), .B(n20836), .ZN(
        P1_U3154) );
  AOI22_X1 U23743 ( .A1(n20840), .A2(n20872), .B1(n20839), .B2(n20873), .ZN(
        n20843) );
  AOI22_X1 U23744 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20877), .B1(
        n20876), .B2(n20841), .ZN(n20842) );
  OAI211_X1 U23745 ( .C1(n20844), .C2(n20880), .A(n20843), .B(n20842), .ZN(
        P1_U3155) );
  AOI22_X1 U23746 ( .A1(n20846), .A2(n20872), .B1(n20845), .B2(n20873), .ZN(
        n20849) );
  AOI22_X1 U23747 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20877), .B1(
        n20866), .B2(n20847), .ZN(n20848) );
  OAI211_X1 U23748 ( .C1(n20850), .C2(n20869), .A(n20849), .B(n20848), .ZN(
        P1_U3156) );
  AOI22_X1 U23749 ( .A1(n20852), .A2(n20873), .B1(n20872), .B2(n20851), .ZN(
        n20855) );
  AOI22_X1 U23750 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20877), .B1(
        n20866), .B2(n20853), .ZN(n20854) );
  OAI211_X1 U23751 ( .C1(n20856), .C2(n20869), .A(n20855), .B(n20854), .ZN(
        P1_U3157) );
  AOI22_X1 U23752 ( .A1(n20858), .A2(n20873), .B1(n20872), .B2(n20857), .ZN(
        n20861) );
  AOI22_X1 U23753 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20877), .B1(
        n20866), .B2(n20859), .ZN(n20860) );
  OAI211_X1 U23754 ( .C1(n20862), .C2(n20869), .A(n20861), .B(n20860), .ZN(
        P1_U3158) );
  AOI22_X1 U23755 ( .A1(n20864), .A2(n20873), .B1(n20872), .B2(n20863), .ZN(
        n20868) );
  AOI22_X1 U23756 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20877), .B1(
        n20866), .B2(n20865), .ZN(n20867) );
  OAI211_X1 U23757 ( .C1(n20870), .C2(n20869), .A(n20868), .B(n20867), .ZN(
        P1_U3159) );
  AOI22_X1 U23758 ( .A1(n20874), .A2(n20873), .B1(n20872), .B2(n20871), .ZN(
        n20879) );
  AOI22_X1 U23759 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20877), .B1(
        n20876), .B2(n20875), .ZN(n20878) );
  OAI211_X1 U23760 ( .C1(n20881), .C2(n20880), .A(n20879), .B(n20878), .ZN(
        P1_U3160) );
  NAND2_X1 U23761 ( .A1(n20883), .A2(n20882), .ZN(P1_U3163) );
  AND2_X1 U23762 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20884), .ZN(
        P1_U3164) );
  AND2_X1 U23763 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20884), .ZN(
        P1_U3165) );
  AND2_X1 U23764 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20884), .ZN(
        P1_U3166) );
  AND2_X1 U23765 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20884), .ZN(
        P1_U3167) );
  AND2_X1 U23766 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20884), .ZN(
        P1_U3168) );
  AND2_X1 U23767 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20884), .ZN(
        P1_U3169) );
  AND2_X1 U23768 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20884), .ZN(
        P1_U3170) );
  AND2_X1 U23769 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20884), .ZN(
        P1_U3171) );
  AND2_X1 U23770 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20884), .ZN(
        P1_U3172) );
  AND2_X1 U23771 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20884), .ZN(
        P1_U3173) );
  AND2_X1 U23772 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20884), .ZN(
        P1_U3174) );
  AND2_X1 U23773 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20884), .ZN(
        P1_U3175) );
  AND2_X1 U23774 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20884), .ZN(
        P1_U3176) );
  AND2_X1 U23775 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20884), .ZN(
        P1_U3177) );
  AND2_X1 U23776 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20884), .ZN(
        P1_U3178) );
  AND2_X1 U23777 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20884), .ZN(
        P1_U3179) );
  AND2_X1 U23778 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20884), .ZN(
        P1_U3180) );
  AND2_X1 U23779 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20884), .ZN(
        P1_U3181) );
  AND2_X1 U23780 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20884), .ZN(
        P1_U3182) );
  AND2_X1 U23781 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20884), .ZN(
        P1_U3183) );
  AND2_X1 U23782 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20884), .ZN(
        P1_U3184) );
  AND2_X1 U23783 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20884), .ZN(
        P1_U3185) );
  AND2_X1 U23784 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20884), .ZN(P1_U3186) );
  AND2_X1 U23785 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20884), .ZN(P1_U3187) );
  AND2_X1 U23786 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20884), .ZN(P1_U3188) );
  AND2_X1 U23787 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20884), .ZN(P1_U3189) );
  AND2_X1 U23788 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20884), .ZN(P1_U3190) );
  AND2_X1 U23789 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20884), .ZN(P1_U3191) );
  AND2_X1 U23790 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20884), .ZN(P1_U3192) );
  AND2_X1 U23791 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20884), .ZN(P1_U3193) );
  NAND2_X1 U23792 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20885), .ZN(n20891) );
  NAND2_X1 U23793 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n20886) );
  OAI211_X1 U23794 ( .C1(P1_STATE_REG_0__SCAN_IN), .C2(n20898), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .B(n20886), .ZN(n20887) );
  OAI21_X1 U23795 ( .B1(n20888), .B2(n20887), .A(n20945), .ZN(n20889) );
  OAI211_X1 U23796 ( .C1(n20892), .C2(n20891), .A(n20890), .B(n20889), .ZN(
        P1_U3194) );
  NOR3_X1 U23797 ( .A1(NA), .A2(n12713), .A3(n20892), .ZN(n20893) );
  INV_X1 U23798 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21028) );
  OAI22_X1 U23799 ( .A1(n20894), .A2(n20893), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n21028), .ZN(n20901) );
  NOR2_X1 U23800 ( .A1(n12713), .A2(n21028), .ZN(n20899) );
  INV_X1 U23801 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20896) );
  OAI221_X1 U23802 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(NA), .C1(
        P1_STATE_REG_0__SCAN_IN), .C2(n20896), .A(n20895), .ZN(n20897) );
  OAI221_X1 U23803 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n20899), .C1(
        P1_STATE_REG_2__SCAN_IN), .C2(n20898), .A(n20897), .ZN(n20900) );
  OAI21_X1 U23804 ( .B1(n21115), .B2(n20901), .A(n20900), .ZN(P1_U3196) );
  OR2_X1 U23805 ( .A1(n20979), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20928) );
  NAND2_X1 U23806 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20980), .ZN(n20926) );
  INV_X1 U23807 ( .A(n20926), .ZN(n20940) );
  AOI22_X1 U23808 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(n20945), .B1(
        P1_REIP_REG_1__SCAN_IN), .B2(n20940), .ZN(n20902) );
  OAI21_X1 U23809 ( .B1(n13786), .B2(n20928), .A(n20902), .ZN(P1_U3197) );
  AOI22_X1 U23810 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n20979), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20940), .ZN(n20903) );
  OAI21_X1 U23811 ( .B1(n20905), .B2(n20928), .A(n20903), .ZN(P1_U3198) );
  INV_X1 U23812 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20906) );
  OAI222_X1 U23813 ( .A1(n20926), .A2(n20905), .B1(n20904), .B2(n20980), .C1(
        n20906), .C2(n20928), .ZN(P1_U3199) );
  INV_X1 U23814 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20907) );
  OAI222_X1 U23815 ( .A1(n20928), .A2(n20908), .B1(n20907), .B2(n20980), .C1(
        n20906), .C2(n20926), .ZN(P1_U3200) );
  AOI222_X1 U23816 ( .A1(n20940), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20945), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20939), .ZN(n20909) );
  INV_X1 U23817 ( .A(n20909), .ZN(P1_U3201) );
  AOI222_X1 U23818 ( .A1(n20940), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20979), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20939), .ZN(n20910) );
  INV_X1 U23819 ( .A(n20910), .ZN(P1_U3202) );
  AOI222_X1 U23820 ( .A1(n20940), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20979), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20939), .ZN(n20911) );
  INV_X1 U23821 ( .A(n20911), .ZN(P1_U3203) );
  AOI222_X1 U23822 ( .A1(n20939), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20979), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20940), .ZN(n20912) );
  INV_X1 U23823 ( .A(n20912), .ZN(P1_U3204) );
  AOI222_X1 U23824 ( .A1(n20940), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20979), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20939), .ZN(n20913) );
  INV_X1 U23825 ( .A(n20913), .ZN(P1_U3205) );
  AOI222_X1 U23826 ( .A1(n20940), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20945), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n20939), .ZN(n20914) );
  INV_X1 U23827 ( .A(n20914), .ZN(P1_U3206) );
  AOI222_X1 U23828 ( .A1(n20940), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20945), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20939), .ZN(n20915) );
  INV_X1 U23829 ( .A(n20915), .ZN(P1_U3207) );
  AOI22_X1 U23830 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n20945), .B1(
        P1_REIP_REG_13__SCAN_IN), .B2(n20939), .ZN(n20916) );
  OAI21_X1 U23831 ( .B1(n20917), .B2(n20926), .A(n20916), .ZN(P1_U3208) );
  AOI22_X1 U23832 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20945), .B1(
        P1_REIP_REG_13__SCAN_IN), .B2(n20940), .ZN(n20918) );
  OAI21_X1 U23833 ( .B1(n20919), .B2(n20928), .A(n20918), .ZN(P1_U3209) );
  AOI222_X1 U23834 ( .A1(n20939), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20979), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20940), .ZN(n20920) );
  INV_X1 U23835 ( .A(n20920), .ZN(P1_U3210) );
  AOI222_X1 U23836 ( .A1(n20940), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20979), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20939), .ZN(n20921) );
  INV_X1 U23837 ( .A(n20921), .ZN(P1_U3211) );
  AOI22_X1 U23838 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20945), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20939), .ZN(n20922) );
  OAI21_X1 U23839 ( .B1(n20923), .B2(n20926), .A(n20922), .ZN(P1_U3212) );
  AOI22_X1 U23840 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20945), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20940), .ZN(n20924) );
  OAI21_X1 U23841 ( .B1(n14775), .B2(n20928), .A(n20924), .ZN(P1_U3213) );
  AOI22_X1 U23842 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n20945), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20939), .ZN(n20925) );
  OAI21_X1 U23843 ( .B1(n14775), .B2(n20926), .A(n20925), .ZN(P1_U3214) );
  AOI22_X1 U23844 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20945), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20940), .ZN(n20927) );
  OAI21_X1 U23845 ( .B1(n21073), .B2(n20928), .A(n20927), .ZN(P1_U3215) );
  AOI222_X1 U23846 ( .A1(n20939), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20945), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n20940), .ZN(n20929) );
  INV_X1 U23847 ( .A(n20929), .ZN(P1_U3216) );
  AOI222_X1 U23848 ( .A1(n20939), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20945), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20940), .ZN(n20930) );
  INV_X1 U23849 ( .A(n20930), .ZN(P1_U3217) );
  AOI222_X1 U23850 ( .A1(n20939), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20945), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n20940), .ZN(n20931) );
  INV_X1 U23851 ( .A(n20931), .ZN(P1_U3218) );
  AOI222_X1 U23852 ( .A1(n20940), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20945), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n20939), .ZN(n20932) );
  INV_X1 U23853 ( .A(n20932), .ZN(P1_U3219) );
  AOI222_X1 U23854 ( .A1(n20940), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20945), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20939), .ZN(n20933) );
  INV_X1 U23855 ( .A(n20933), .ZN(P1_U3220) );
  AOI222_X1 U23856 ( .A1(n20940), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20945), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20939), .ZN(n20934) );
  INV_X1 U23857 ( .A(n20934), .ZN(P1_U3221) );
  AOI222_X1 U23858 ( .A1(n20940), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20945), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20939), .ZN(n20935) );
  INV_X1 U23859 ( .A(n20935), .ZN(P1_U3222) );
  AOI222_X1 U23860 ( .A1(n20940), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20945), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20939), .ZN(n20936) );
  INV_X1 U23861 ( .A(n20936), .ZN(P1_U3223) );
  AOI222_X1 U23862 ( .A1(n20940), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20979), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20939), .ZN(n20937) );
  INV_X1 U23863 ( .A(n20937), .ZN(P1_U3224) );
  AOI222_X1 U23864 ( .A1(n20939), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20945), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20940), .ZN(n20938) );
  INV_X1 U23865 ( .A(n20938), .ZN(P1_U3225) );
  AOI222_X1 U23866 ( .A1(n20940), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20945), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20939), .ZN(n20941) );
  INV_X1 U23867 ( .A(n20941), .ZN(P1_U3226) );
  OAI22_X1 U23868 ( .A1(n20979), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20980), .ZN(n20942) );
  INV_X1 U23869 ( .A(n20942), .ZN(P1_U3458) );
  OAI22_X1 U23870 ( .A1(n20979), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20980), .ZN(n20943) );
  INV_X1 U23871 ( .A(n20943), .ZN(P1_U3459) );
  OAI22_X1 U23872 ( .A1(n20979), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20980), .ZN(n20944) );
  INV_X1 U23873 ( .A(n20944), .ZN(P1_U3460) );
  OAI22_X1 U23874 ( .A1(n20945), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20980), .ZN(n20946) );
  INV_X1 U23875 ( .A(n20946), .ZN(P1_U3461) );
  INV_X1 U23876 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20960) );
  AOI21_X1 U23877 ( .B1(n20960), .B2(n20884), .A(n20947), .ZN(P1_U3464) );
  AOI21_X1 U23878 ( .B1(n20884), .B2(P1_DATAWIDTH_REG_1__SCAN_IN), .A(n20947), 
        .ZN(n20948) );
  INV_X1 U23879 ( .A(n20948), .ZN(P1_U3465) );
  AOI21_X1 U23880 ( .B1(n20949), .B2(n11516), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n20951) );
  OAI22_X1 U23881 ( .A1(n20952), .A2(n20951), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20950), .ZN(n20954) );
  AOI22_X1 U23882 ( .A1(n20955), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20954), .B2(n20953), .ZN(n20956) );
  OAI21_X1 U23883 ( .B1(n20958), .B2(n20957), .A(n20956), .ZN(P1_U3474) );
  NOR3_X1 U23884 ( .A1(n20960), .A2(P1_REIP_REG_0__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .ZN(n20959) );
  AOI221_X1 U23885 ( .B1(n20961), .B2(n20960), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n20959), .ZN(n20962) );
  INV_X1 U23886 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21059) );
  INV_X1 U23887 ( .A(n20965), .ZN(n20963) );
  AOI22_X1 U23888 ( .A1(n20965), .A2(n20962), .B1(n21059), .B2(n20963), .ZN(
        P1_U3481) );
  NOR2_X1 U23889 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n20964) );
  INV_X1 U23890 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21109) );
  AOI22_X1 U23891 ( .A1(n20965), .A2(n20964), .B1(n21109), .B2(n20963), .ZN(
        P1_U3482) );
  INV_X1 U23892 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20966) );
  AOI22_X1 U23893 ( .A1(n20980), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20966), 
        .B2(n20979), .ZN(P1_U3483) );
  AOI211_X1 U23894 ( .C1(n20969), .C2(n21106), .A(n20968), .B(n20967), .ZN(
        n20972) );
  OAI21_X1 U23895 ( .B1(n20972), .B2(n20971), .A(n20970), .ZN(n20978) );
  AOI211_X1 U23896 ( .C1(n20976), .C2(n20975), .A(n20974), .B(n20973), .ZN(
        n20977) );
  MUX2_X1 U23897 ( .A(n20978), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n20977), 
        .Z(P1_U3485) );
  INV_X1 U23898 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n21122) );
  AOI22_X1 U23899 ( .A1(n20980), .A2(n21122), .B1(n21118), .B2(n20979), .ZN(
        P1_U3486) );
  INV_X1 U23900 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n21174) );
  AOI22_X1 U23901 ( .A1(DATAI_16_), .A2(keyinput_f16), .B1(
        P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_f44), .ZN(n20981) );
  OAI221_X1 U23902 ( .B1(DATAI_16_), .B2(keyinput_f16), .C1(
        P1_STATEBS16_REG_SCAN_IN), .C2(keyinput_f44), .A(n20981), .ZN(n20988)
         );
  AOI22_X1 U23903 ( .A1(DATAI_30_), .A2(keyinput_f2), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(keyinput_f62), .ZN(n20982) );
  OAI221_X1 U23904 ( .B1(DATAI_30_), .B2(keyinput_f2), .C1(
        P1_REIP_REG_21__SCAN_IN), .C2(keyinput_f62), .A(n20982), .ZN(n20987)
         );
  AOI22_X1 U23905 ( .A1(DATAI_0_), .A2(keyinput_f32), .B1(DATAI_11_), .B2(
        keyinput_f21), .ZN(n20983) );
  OAI221_X1 U23906 ( .B1(DATAI_0_), .B2(keyinput_f32), .C1(DATAI_11_), .C2(
        keyinput_f21), .A(n20983), .ZN(n20986) );
  AOI22_X1 U23907 ( .A1(DATAI_21_), .A2(keyinput_f11), .B1(DATAI_28_), .B2(
        keyinput_f4), .ZN(n20984) );
  OAI221_X1 U23908 ( .B1(DATAI_21_), .B2(keyinput_f11), .C1(DATAI_28_), .C2(
        keyinput_f4), .A(n20984), .ZN(n20985) );
  NOR4_X1 U23909 ( .A1(n20988), .A2(n20987), .A3(n20986), .A4(n20985), .ZN(
        n21015) );
  INV_X1 U23910 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21099) );
  XNOR2_X1 U23911 ( .A(n21099), .B(keyinput_f55), .ZN(n20995) );
  AOI22_X1 U23912 ( .A1(DATAI_23_), .A2(keyinput_f9), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(keyinput_f58), .ZN(n20989) );
  OAI221_X1 U23913 ( .B1(DATAI_23_), .B2(keyinput_f9), .C1(
        P1_REIP_REG_25__SCAN_IN), .C2(keyinput_f58), .A(n20989), .ZN(n20994)
         );
  AOI22_X1 U23914 ( .A1(keyinput_f51), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        DATAI_3_), .B2(keyinput_f29), .ZN(n20990) );
  OAI221_X1 U23915 ( .B1(keyinput_f51), .B2(P1_BYTEENABLE_REG_3__SCAN_IN), 
        .C1(DATAI_3_), .C2(keyinput_f29), .A(n20990), .ZN(n20993) );
  AOI22_X1 U23916 ( .A1(keyinput_f33), .A2(HOLD), .B1(P1_FLUSH_REG_SCAN_IN), 
        .B2(keyinput_f46), .ZN(n20991) );
  OAI221_X1 U23917 ( .B1(keyinput_f33), .B2(HOLD), .C1(P1_FLUSH_REG_SCAN_IN), 
        .C2(keyinput_f46), .A(n20991), .ZN(n20992) );
  NOR4_X1 U23918 ( .A1(n20995), .A2(n20994), .A3(n20993), .A4(n20992), .ZN(
        n21014) );
  AOI22_X1 U23919 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(keyinput_f40), .B1(
        DATAI_2_), .B2(keyinput_f30), .ZN(n20996) );
  OAI221_X1 U23920 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_f40), .C1(
        DATAI_2_), .C2(keyinput_f30), .A(n20996), .ZN(n21003) );
  AOI22_X1 U23921 ( .A1(keyinput_f34), .A2(NA), .B1(DATAI_20_), .B2(
        keyinput_f12), .ZN(n20997) );
  OAI221_X1 U23922 ( .B1(keyinput_f34), .B2(NA), .C1(DATAI_20_), .C2(
        keyinput_f12), .A(n20997), .ZN(n21002) );
  AOI22_X1 U23923 ( .A1(DATAI_18_), .A2(keyinput_f14), .B1(DATAI_6_), .B2(
        keyinput_f26), .ZN(n20998) );
  OAI221_X1 U23924 ( .B1(DATAI_18_), .B2(keyinput_f14), .C1(DATAI_6_), .C2(
        keyinput_f26), .A(n20998), .ZN(n21001) );
  AOI22_X1 U23925 ( .A1(DATAI_8_), .A2(keyinput_f24), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(keyinput_f60), .ZN(n20999) );
  OAI221_X1 U23926 ( .B1(DATAI_8_), .B2(keyinput_f24), .C1(
        P1_REIP_REG_23__SCAN_IN), .C2(keyinput_f60), .A(n20999), .ZN(n21000)
         );
  NOR4_X1 U23927 ( .A1(n21003), .A2(n21002), .A3(n21001), .A4(n21000), .ZN(
        n21013) );
  AOI22_X1 U23928 ( .A1(DATAI_24_), .A2(keyinput_f8), .B1(DATAI_25_), .B2(
        keyinput_f7), .ZN(n21004) );
  OAI221_X1 U23929 ( .B1(DATAI_24_), .B2(keyinput_f8), .C1(DATAI_25_), .C2(
        keyinput_f7), .A(n21004), .ZN(n21011) );
  AOI22_X1 U23930 ( .A1(DATAI_10_), .A2(keyinput_f22), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(keyinput_f61), .ZN(n21005) );
  OAI221_X1 U23931 ( .B1(DATAI_10_), .B2(keyinput_f22), .C1(
        P1_REIP_REG_22__SCAN_IN), .C2(keyinput_f61), .A(n21005), .ZN(n21010)
         );
  AOI22_X1 U23932 ( .A1(READY2), .A2(keyinput_f37), .B1(DATAI_27_), .B2(
        keyinput_f5), .ZN(n21006) );
  OAI221_X1 U23933 ( .B1(READY2), .B2(keyinput_f37), .C1(DATAI_27_), .C2(
        keyinput_f5), .A(n21006), .ZN(n21009) );
  AOI22_X1 U23934 ( .A1(keyinput_f39), .A2(P1_ADS_N_REG_SCAN_IN), .B1(DATAI_1_), .B2(keyinput_f31), .ZN(n21007) );
  OAI221_X1 U23935 ( .B1(keyinput_f39), .B2(P1_ADS_N_REG_SCAN_IN), .C1(
        DATAI_1_), .C2(keyinput_f31), .A(n21007), .ZN(n21008) );
  NOR4_X1 U23936 ( .A1(n21011), .A2(n21010), .A3(n21009), .A4(n21008), .ZN(
        n21012) );
  NAND4_X1 U23937 ( .A1(n21015), .A2(n21014), .A3(n21013), .A4(n21012), .ZN(
        n21070) );
  INV_X1 U23938 ( .A(READY1), .ZN(n21076) );
  AOI22_X1 U23939 ( .A1(n21076), .A2(keyinput_f36), .B1(keyinput_f10), .B2(
        n21017), .ZN(n21016) );
  OAI221_X1 U23940 ( .B1(n21076), .B2(keyinput_f36), .C1(n21017), .C2(
        keyinput_f10), .A(n21016), .ZN(n21025) );
  AOI22_X1 U23941 ( .A1(n21103), .A2(keyinput_f23), .B1(keyinput_f0), .B2(
        n21122), .ZN(n21018) );
  OAI221_X1 U23942 ( .B1(n21103), .B2(keyinput_f23), .C1(n21122), .C2(
        keyinput_f0), .A(n21018), .ZN(n21024) );
  AOI22_X1 U23943 ( .A1(n14543), .A2(keyinput_f57), .B1(keyinput_f49), .B2(
        n21077), .ZN(n21019) );
  OAI221_X1 U23944 ( .B1(n14543), .B2(keyinput_f57), .C1(n21077), .C2(
        keyinput_f49), .A(n21019), .ZN(n21023) );
  INV_X1 U23945 ( .A(DATAI_14_), .ZN(n21021) );
  INV_X1 U23946 ( .A(DATAI_13_), .ZN(n21124) );
  AOI22_X1 U23947 ( .A1(n21021), .A2(keyinput_f18), .B1(keyinput_f19), .B2(
        n21124), .ZN(n21020) );
  OAI221_X1 U23948 ( .B1(n21021), .B2(keyinput_f18), .C1(n21124), .C2(
        keyinput_f19), .A(n21020), .ZN(n21022) );
  NOR4_X1 U23949 ( .A1(n21025), .A2(n21024), .A3(n21023), .A4(n21022), .ZN(
        n21068) );
  AOI22_X1 U23950 ( .A1(n21028), .A2(keyinput_f43), .B1(n21027), .B2(
        keyinput_f15), .ZN(n21026) );
  OAI221_X1 U23951 ( .B1(n21028), .B2(keyinput_f43), .C1(n21027), .C2(
        keyinput_f15), .A(n21026), .ZN(n21039) );
  AOI22_X1 U23952 ( .A1(DATAI_31_), .A2(keyinput_f1), .B1(n21030), .B2(
        keyinput_f3), .ZN(n21029) );
  OAI221_X1 U23953 ( .B1(DATAI_31_), .B2(keyinput_f1), .C1(n21030), .C2(
        keyinput_f3), .A(n21029), .ZN(n21038) );
  INV_X1 U23954 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n21033) );
  INV_X1 U23955 ( .A(keyinput_f47), .ZN(n21032) );
  AOI22_X1 U23956 ( .A1(n21033), .A2(keyinput_f38), .B1(P1_W_R_N_REG_SCAN_IN), 
        .B2(n21032), .ZN(n21031) );
  OAI221_X1 U23957 ( .B1(n21033), .B2(keyinput_f38), .C1(n21032), .C2(
        P1_W_R_N_REG_SCAN_IN), .A(n21031), .ZN(n21037) );
  AOI22_X1 U23958 ( .A1(n21035), .A2(keyinput_f25), .B1(keyinput_f48), .B2(
        n21109), .ZN(n21034) );
  OAI221_X1 U23959 ( .B1(n21035), .B2(keyinput_f25), .C1(n21109), .C2(
        keyinput_f48), .A(n21034), .ZN(n21036) );
  NOR4_X1 U23960 ( .A1(n21039), .A2(n21038), .A3(n21037), .A4(n21036), .ZN(
        n21067) );
  AOI22_X1 U23961 ( .A1(n14693), .A2(keyinput_f13), .B1(n21041), .B2(
        keyinput_f27), .ZN(n21040) );
  OAI221_X1 U23962 ( .B1(n14693), .B2(keyinput_f13), .C1(n21041), .C2(
        keyinput_f27), .A(n21040), .ZN(n21051) );
  AOI22_X1 U23963 ( .A1(n21043), .A2(keyinput_f20), .B1(keyinput_f6), .B2(
        n21121), .ZN(n21042) );
  OAI221_X1 U23964 ( .B1(n21043), .B2(keyinput_f20), .C1(n21121), .C2(
        keyinput_f6), .A(n21042), .ZN(n21050) );
  INV_X1 U23965 ( .A(keyinput_f42), .ZN(n21045) );
  AOI22_X1 U23966 ( .A1(n21046), .A2(keyinput_f54), .B1(P1_D_C_N_REG_SCAN_IN), 
        .B2(n21045), .ZN(n21044) );
  OAI221_X1 U23967 ( .B1(n21046), .B2(keyinput_f54), .C1(n21045), .C2(
        P1_D_C_N_REG_SCAN_IN), .A(n21044), .ZN(n21049) );
  AOI22_X1 U23968 ( .A1(n21073), .A2(keyinput_f63), .B1(n21082), .B2(
        keyinput_f52), .ZN(n21047) );
  OAI221_X1 U23969 ( .B1(n21073), .B2(keyinput_f63), .C1(n21082), .C2(
        keyinput_f52), .A(n21047), .ZN(n21048) );
  NOR4_X1 U23970 ( .A1(n21051), .A2(n21050), .A3(n21049), .A4(n21048), .ZN(
        n21066) );
  AOI22_X1 U23971 ( .A1(n21118), .A2(keyinput_f41), .B1(n21053), .B2(
        keyinput_f56), .ZN(n21052) );
  OAI221_X1 U23972 ( .B1(n21118), .B2(keyinput_f41), .C1(n21053), .C2(
        keyinput_f56), .A(n21052), .ZN(n21064) );
  AOI22_X1 U23973 ( .A1(n21056), .A2(keyinput_f45), .B1(n21055), .B2(
        keyinput_f59), .ZN(n21054) );
  OAI221_X1 U23974 ( .B1(n21056), .B2(keyinput_f45), .C1(n21055), .C2(
        keyinput_f59), .A(n21054), .ZN(n21063) );
  INV_X1 U23975 ( .A(DATAI_4_), .ZN(n21080) );
  AOI22_X1 U23976 ( .A1(n21080), .A2(keyinput_f28), .B1(keyinput_f35), .B2(
        n21102), .ZN(n21057) );
  OAI221_X1 U23977 ( .B1(n21080), .B2(keyinput_f28), .C1(n21102), .C2(
        keyinput_f35), .A(n21057), .ZN(n21062) );
  AOI22_X1 U23978 ( .A1(n21060), .A2(keyinput_f17), .B1(keyinput_f50), .B2(
        n21059), .ZN(n21058) );
  OAI221_X1 U23979 ( .B1(n21060), .B2(keyinput_f17), .C1(n21059), .C2(
        keyinput_f50), .A(n21058), .ZN(n21061) );
  NOR4_X1 U23980 ( .A1(n21064), .A2(n21063), .A3(n21062), .A4(n21061), .ZN(
        n21065) );
  NAND4_X1 U23981 ( .A1(n21068), .A2(n21067), .A3(n21066), .A4(n21065), .ZN(
        n21069) );
  OAI22_X1 U23982 ( .A1(n21070), .A2(n21069), .B1(keyinput_f53), .B2(
        P1_REIP_REG_30__SCAN_IN), .ZN(n21071) );
  AOI21_X1 U23983 ( .B1(keyinput_f53), .B2(P1_REIP_REG_30__SCAN_IN), .A(n21071), .ZN(n21173) );
  INV_X1 U23984 ( .A(READY2), .ZN(n21074) );
  AOI22_X1 U23985 ( .A1(n21074), .A2(keyinput_g37), .B1(n21073), .B2(
        keyinput_g63), .ZN(n21072) );
  OAI221_X1 U23986 ( .B1(n21074), .B2(keyinput_g37), .C1(n21073), .C2(
        keyinput_g63), .A(n21072), .ZN(n21087) );
  AOI22_X1 U23987 ( .A1(n21077), .A2(keyinput_g49), .B1(n21076), .B2(
        keyinput_g36), .ZN(n21075) );
  OAI221_X1 U23988 ( .B1(n21077), .B2(keyinput_g49), .C1(n21076), .C2(
        keyinput_g36), .A(n21075), .ZN(n21086) );
  AOI22_X1 U23989 ( .A1(n21080), .A2(keyinput_g28), .B1(n21079), .B2(
        keyinput_g8), .ZN(n21078) );
  OAI221_X1 U23990 ( .B1(n21080), .B2(keyinput_g28), .C1(n21079), .C2(
        keyinput_g8), .A(n21078), .ZN(n21085) );
  AOI22_X1 U23991 ( .A1(n21083), .A2(keyinput_g11), .B1(n21082), .B2(
        keyinput_g52), .ZN(n21081) );
  OAI221_X1 U23992 ( .B1(n21083), .B2(keyinput_g11), .C1(n21082), .C2(
        keyinput_g52), .A(n21081), .ZN(n21084) );
  NOR4_X1 U23993 ( .A1(n21087), .A2(n21086), .A3(n21085), .A4(n21084), .ZN(
        n21133) );
  AOI22_X1 U23994 ( .A1(DATAI_23_), .A2(keyinput_g9), .B1(DATAI_12_), .B2(
        keyinput_g20), .ZN(n21088) );
  OAI221_X1 U23995 ( .B1(DATAI_23_), .B2(keyinput_g9), .C1(DATAI_12_), .C2(
        keyinput_g20), .A(n21088), .ZN(n21097) );
  AOI22_X1 U23996 ( .A1(DATAI_22_), .A2(keyinput_g10), .B1(DATAI_30_), .B2(
        keyinput_g2), .ZN(n21089) );
  OAI221_X1 U23997 ( .B1(DATAI_22_), .B2(keyinput_g10), .C1(DATAI_30_), .C2(
        keyinput_g2), .A(n21089), .ZN(n21096) );
  AOI22_X1 U23998 ( .A1(n21091), .A2(keyinput_g12), .B1(n14543), .B2(
        keyinput_g57), .ZN(n21090) );
  OAI221_X1 U23999 ( .B1(n21091), .B2(keyinput_g12), .C1(n14543), .C2(
        keyinput_g57), .A(n21090), .ZN(n21095) );
  AOI22_X1 U24000 ( .A1(P1_MORE_REG_SCAN_IN), .A2(keyinput_g45), .B1(n21093), 
        .B2(keyinput_g51), .ZN(n21092) );
  OAI221_X1 U24001 ( .B1(P1_MORE_REG_SCAN_IN), .B2(keyinput_g45), .C1(n21093), 
        .C2(keyinput_g51), .A(n21092), .ZN(n21094) );
  NOR4_X1 U24002 ( .A1(n21097), .A2(n21096), .A3(n21095), .A4(n21094), .ZN(
        n21132) );
  AOI22_X1 U24003 ( .A1(n21100), .A2(keyinput_g46), .B1(n21099), .B2(
        keyinput_g55), .ZN(n21098) );
  OAI221_X1 U24004 ( .B1(n21100), .B2(keyinput_g46), .C1(n21099), .C2(
        keyinput_g55), .A(n21098), .ZN(n21113) );
  AOI22_X1 U24005 ( .A1(n21103), .A2(keyinput_g23), .B1(keyinput_g35), .B2(
        n21102), .ZN(n21101) );
  OAI221_X1 U24006 ( .B1(n21103), .B2(keyinput_g23), .C1(n21102), .C2(
        keyinput_g35), .A(n21101), .ZN(n21112) );
  AOI22_X1 U24007 ( .A1(n21106), .A2(keyinput_g44), .B1(keyinput_g7), .B2(
        n21105), .ZN(n21104) );
  OAI221_X1 U24008 ( .B1(n21106), .B2(keyinput_g44), .C1(n21105), .C2(
        keyinput_g7), .A(n21104), .ZN(n21111) );
  AOI22_X1 U24009 ( .A1(n21109), .A2(keyinput_g48), .B1(n21108), .B2(
        keyinput_g14), .ZN(n21107) );
  OAI221_X1 U24010 ( .B1(n21109), .B2(keyinput_g48), .C1(n21108), .C2(
        keyinput_g14), .A(n21107), .ZN(n21110) );
  NOR4_X1 U24011 ( .A1(n21113), .A2(n21112), .A3(n21111), .A4(n21110), .ZN(
        n21131) );
  AOI22_X1 U24012 ( .A1(n21116), .A2(keyinput_g58), .B1(keyinput_g33), .B2(
        n21115), .ZN(n21114) );
  OAI221_X1 U24013 ( .B1(n21116), .B2(keyinput_g58), .C1(n21115), .C2(
        keyinput_g33), .A(n21114), .ZN(n21129) );
  INV_X1 U24014 ( .A(DATAI_6_), .ZN(n21119) );
  AOI22_X1 U24015 ( .A1(n21119), .A2(keyinput_g26), .B1(keyinput_g41), .B2(
        n21118), .ZN(n21117) );
  OAI221_X1 U24016 ( .B1(n21119), .B2(keyinput_g26), .C1(n21118), .C2(
        keyinput_g41), .A(n21117), .ZN(n21128) );
  AOI22_X1 U24017 ( .A1(n21122), .A2(keyinput_g0), .B1(n21121), .B2(
        keyinput_g6), .ZN(n21120) );
  OAI221_X1 U24018 ( .B1(n21122), .B2(keyinput_g0), .C1(n21121), .C2(
        keyinput_g6), .A(n21120), .ZN(n21127) );
  INV_X1 U24019 ( .A(DATAI_1_), .ZN(n21125) );
  AOI22_X1 U24020 ( .A1(n21125), .A2(keyinput_g31), .B1(n21124), .B2(
        keyinput_g19), .ZN(n21123) );
  OAI221_X1 U24021 ( .B1(n21125), .B2(keyinput_g31), .C1(n21124), .C2(
        keyinput_g19), .A(n21123), .ZN(n21126) );
  NOR4_X1 U24022 ( .A1(n21129), .A2(n21128), .A3(n21127), .A4(n21126), .ZN(
        n21130) );
  NAND4_X1 U24023 ( .A1(n21133), .A2(n21132), .A3(n21131), .A4(n21130), .ZN(
        n21171) );
  AOI22_X1 U24024 ( .A1(DATAI_5_), .A2(keyinput_g27), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(keyinput_g62), .ZN(n21134) );
  OAI221_X1 U24025 ( .B1(DATAI_5_), .B2(keyinput_g27), .C1(
        P1_REIP_REG_21__SCAN_IN), .C2(keyinput_g62), .A(n21134), .ZN(n21141)
         );
  AOI22_X1 U24026 ( .A1(DATAI_19_), .A2(keyinput_g13), .B1(DATAI_14_), .B2(
        keyinput_g18), .ZN(n21135) );
  OAI221_X1 U24027 ( .B1(DATAI_19_), .B2(keyinput_g13), .C1(DATAI_14_), .C2(
        keyinput_g18), .A(n21135), .ZN(n21140) );
  AOI22_X1 U24028 ( .A1(P1_READREQUEST_REG_SCAN_IN), .A2(keyinput_g38), .B1(
        DATAI_27_), .B2(keyinput_g5), .ZN(n21136) );
  OAI221_X1 U24029 ( .B1(P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_g38), .C1(
        DATAI_27_), .C2(keyinput_g5), .A(n21136), .ZN(n21139) );
  AOI22_X1 U24030 ( .A1(DATAI_31_), .A2(keyinput_g1), .B1(
        P1_REIP_REG_27__SCAN_IN), .B2(keyinput_g56), .ZN(n21137) );
  OAI221_X1 U24031 ( .B1(DATAI_31_), .B2(keyinput_g1), .C1(
        P1_REIP_REG_27__SCAN_IN), .C2(keyinput_g56), .A(n21137), .ZN(n21138)
         );
  NOR4_X1 U24032 ( .A1(n21141), .A2(n21140), .A3(n21139), .A4(n21138), .ZN(
        n21169) );
  XNOR2_X1 U24033 ( .A(P1_W_R_N_REG_SCAN_IN), .B(keyinput_g47), .ZN(n21149) );
  AOI22_X1 U24034 ( .A1(DATAI_11_), .A2(keyinput_g21), .B1(n21143), .B2(
        keyinput_g16), .ZN(n21142) );
  OAI221_X1 U24035 ( .B1(DATAI_11_), .B2(keyinput_g21), .C1(n21143), .C2(
        keyinput_g16), .A(n21142), .ZN(n21148) );
  AOI22_X1 U24036 ( .A1(P1_REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_g43), 
        .B1(DATAI_10_), .B2(keyinput_g22), .ZN(n21144) );
  OAI221_X1 U24037 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_g43), 
        .C1(DATAI_10_), .C2(keyinput_g22), .A(n21144), .ZN(n21147) );
  AOI22_X1 U24038 ( .A1(DATAI_15_), .A2(keyinput_g17), .B1(DATAI_0_), .B2(
        keyinput_g32), .ZN(n21145) );
  OAI221_X1 U24039 ( .B1(DATAI_15_), .B2(keyinput_g17), .C1(DATAI_0_), .C2(
        keyinput_g32), .A(n21145), .ZN(n21146) );
  NOR4_X1 U24040 ( .A1(n21149), .A2(n21148), .A3(n21147), .A4(n21146), .ZN(
        n21168) );
  AOI22_X1 U24041 ( .A1(P1_BYTEENABLE_REG_2__SCAN_IN), .A2(keyinput_g50), .B1(
        DATAI_29_), .B2(keyinput_g3), .ZN(n21150) );
  OAI221_X1 U24042 ( .B1(P1_BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_g50), 
        .C1(DATAI_29_), .C2(keyinput_g3), .A(n21150), .ZN(n21157) );
  AOI22_X1 U24043 ( .A1(DATAI_2_), .A2(keyinput_g30), .B1(DATAI_8_), .B2(
        keyinput_g24), .ZN(n21151) );
  OAI221_X1 U24044 ( .B1(DATAI_2_), .B2(keyinput_g30), .C1(DATAI_8_), .C2(
        keyinput_g24), .A(n21151), .ZN(n21156) );
  AOI22_X1 U24045 ( .A1(DATAI_3_), .A2(keyinput_g29), .B1(DATAI_28_), .B2(
        keyinput_g4), .ZN(n21152) );
  OAI221_X1 U24046 ( .B1(DATAI_3_), .B2(keyinput_g29), .C1(DATAI_28_), .C2(
        keyinput_g4), .A(n21152), .ZN(n21155) );
  AOI22_X1 U24047 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(keyinput_g39), .B1(
        DATAI_17_), .B2(keyinput_g15), .ZN(n21153) );
  OAI221_X1 U24048 ( .B1(P1_ADS_N_REG_SCAN_IN), .B2(keyinput_g39), .C1(
        DATAI_17_), .C2(keyinput_g15), .A(n21153), .ZN(n21154) );
  NOR4_X1 U24049 ( .A1(n21157), .A2(n21156), .A3(n21155), .A4(n21154), .ZN(
        n21167) );
  AOI22_X1 U24050 ( .A1(DATAI_7_), .A2(keyinput_g25), .B1(
        P1_REIP_REG_24__SCAN_IN), .B2(keyinput_g59), .ZN(n21158) );
  OAI221_X1 U24051 ( .B1(DATAI_7_), .B2(keyinput_g25), .C1(
        P1_REIP_REG_24__SCAN_IN), .C2(keyinput_g59), .A(n21158), .ZN(n21165)
         );
  AOI22_X1 U24052 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(keyinput_g40), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(keyinput_g61), .ZN(n21159) );
  OAI221_X1 U24053 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_g40), .C1(
        P1_REIP_REG_22__SCAN_IN), .C2(keyinput_g61), .A(n21159), .ZN(n21164)
         );
  AOI22_X1 U24054 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(keyinput_g60), .B1(
        P1_REIP_REG_29__SCAN_IN), .B2(keyinput_g54), .ZN(n21160) );
  OAI221_X1 U24055 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(keyinput_g60), .C1(
        P1_REIP_REG_29__SCAN_IN), .C2(keyinput_g54), .A(n21160), .ZN(n21163)
         );
  AOI22_X1 U24056 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(keyinput_g42), .B1(NA), 
        .B2(keyinput_g34), .ZN(n21161) );
  OAI221_X1 U24057 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(keyinput_g42), .C1(NA), 
        .C2(keyinput_g34), .A(n21161), .ZN(n21162) );
  NOR4_X1 U24058 ( .A1(n21165), .A2(n21164), .A3(n21163), .A4(n21162), .ZN(
        n21166) );
  NAND4_X1 U24059 ( .A1(n21169), .A2(n21168), .A3(n21167), .A4(n21166), .ZN(
        n21170) );
  OAI22_X1 U24060 ( .A1(keyinput_g53), .A2(n21174), .B1(n21171), .B2(n21170), 
        .ZN(n21172) );
  AOI211_X1 U24061 ( .C1(keyinput_g53), .C2(n21174), .A(n21173), .B(n21172), 
        .ZN(n21176) );
  AOI22_X1 U24062 ( .A1(n16686), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n16688), .ZN(n21175) );
  XNOR2_X1 U24063 ( .A(n21176), .B(n21175), .ZN(U355) );
  INV_X2 U11186 ( .A(n16086), .ZN(n16110) );
  AND2_X1 U11159 ( .A1(n9989), .A2(n9988), .ZN(n10046) );
  INV_X1 U19103 ( .A(n15942), .ZN(n17593) );
  INV_X4 U12511 ( .A(n12912), .ZN(n12945) );
  AOI21_X1 U11099 ( .B1(n12859), .B2(n15877), .A(n12855), .ZN(n11523) );
  CLKBUF_X1 U11103 ( .A(n11428), .Z(n12303) );
  CLKBUF_X1 U11120 ( .A(n12267), .Z(n12294) );
  CLKBUF_X1 U11122 ( .A(n11499), .Z(n13629) );
  NAND2_X1 U11124 ( .A1(n11494), .A2(n11504), .ZN(n12856) );
  INV_X1 U11132 ( .A(n11520), .ZN(n11597) );
  NAND2_X2 U11139 ( .A1(n11494), .A2(n11505), .ZN(n12849) );
  CLKBUF_X1 U11148 ( .A(n12742), .Z(n9674) );
  CLKBUF_X1 U11151 ( .A(n11437), .Z(n12845) );
  CLKBUF_X1 U11168 ( .A(n10437), .Z(n10438) );
  CLKBUF_X1 U11179 ( .A(n11504), .Z(n11531) );
  CLKBUF_X1 U11203 ( .A(n11840), .Z(n11841) );
  CLKBUF_X1 U11204 ( .A(n10366), .Z(n13279) );
  CLKBUF_X1 U11698 ( .A(n19339), .Z(n19355) );
  CLKBUF_X1 U12038 ( .A(n10983), .Z(n9676) );
  CLKBUF_X1 U12316 ( .A(n18996), .Z(n18990) );
endmodule

