

module b21_C_gen_AntiSAT_k_256_6 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2, 
        keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7, 
        keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12, 
        keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17, 
        keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22, 
        keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27, 
        keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32, 
        keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37, 
        keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42, 
        keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47, 
        keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52, 
        keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57, 
        keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62, 
        keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67, 
        keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72, 
        keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77, 
        keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82, 
        keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87, 
        keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92, 
        keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97, 
        keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524;

  NAND2_X1 U4986 ( .A1(n9320), .A2(n9215), .ZN(n9217) );
  NAND2_X1 U4987 ( .A1(n4779), .A2(n4778), .ZN(n8464) );
  AOI21_X1 U4988 ( .B1(n7073), .B2(n7072), .A(n7071), .ZN(n7228) );
  INV_X2 U4989 ( .A(n5946), .ZN(n6538) );
  NAND4_X1 U4990 ( .A1(n5310), .A2(n5309), .A3(n5308), .A4(n5307), .ZN(n7020)
         );
  INV_X1 U4991 ( .A(n5950), .ZN(n5973) );
  CLKBUF_X2 U4992 ( .A(n5311), .Z(n4484) );
  NAND2_X1 U4993 ( .A1(n5916), .A2(n5919), .ZN(n7912) );
  OAI21_X1 U4994 ( .B1(n5211), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5213) );
  AND2_X1 U4995 ( .A1(n7679), .A2(n8629), .ZN(n7735) );
  INV_X1 U4996 ( .A(n6043), .ZN(n7885) );
  INV_X1 U4997 ( .A(n7043), .ZN(n5749) );
  INV_X1 U4998 ( .A(n8151), .ZN(n5227) );
  BUF_X1 U4999 ( .A(n5311), .Z(n4485) );
  NAND2_X1 U5000 ( .A1(n7287), .A2(n8953), .ZN(n7554) );
  INV_X1 U5001 ( .A(n7853), .ZN(n7720) );
  OR2_X1 U5002 ( .A1(n8379), .A2(n8567), .ZN(n8363) );
  OR2_X1 U5003 ( .A1(n8427), .A2(n4768), .ZN(n8379) );
  NAND2_X2 U5004 ( .A1(n6351), .A2(n6350), .ZN(n5946) );
  INV_X1 U5005 ( .A(n9561), .ZN(n5223) );
  INV_X1 U5006 ( .A(n5086), .ZN(n5896) );
  NAND2_X1 U5007 ( .A1(n6007), .A2(n6006), .ZN(n10347) );
  OAI21_X1 U5008 ( .B1(n5773), .B2(n5772), .A(n8753), .ZN(n8738) );
  XNOR2_X1 U5009 ( .A(n5213), .B(n5212), .ZN(n7764) );
  CLKBUF_X3 U5010 ( .A(n5974), .Z(n4488) );
  NAND2_X1 U5011 ( .A1(n6468), .A2(n5850), .ZN(n4481) );
  NAND2_X1 U5012 ( .A1(n6468), .A2(n5850), .ZN(n4482) );
  NAND2_X1 U5013 ( .A1(n6468), .A2(n5850), .ZN(n5478) );
  OAI21_X2 U5014 ( .B1(n9217), .B2(n5035), .A(n5033), .ZN(n9271) );
  NOR2_X2 U5015 ( .A1(n7423), .A2(n7424), .ZN(n4764) );
  NAND2_X2 U5016 ( .A1(n5916), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5915) );
  XNOR2_X2 U5017 ( .A(n7975), .B(n8255), .ZN(n8108) );
  NAND2_X1 U5018 ( .A1(n6349), .A2(n8131), .ZN(n10431) );
  AND2_X1 U5019 ( .A1(n5863), .A2(n7080), .ZN(n5491) );
  NAND2_X1 U5020 ( .A1(n5921), .A2(n5922), .ZN(n4483) );
  NAND2_X1 U5021 ( .A1(n5921), .A2(n5922), .ZN(n6016) );
  NAND2_X1 U5022 ( .A1(n4481), .A2(n5896), .ZN(n5311) );
  NAND2_X1 U5023 ( .A1(n5302), .A2(n5303), .ZN(n6632) );
  OR2_X2 U5024 ( .A1(n10431), .A2(n8103), .ZN(n10462) );
  XNOR2_X1 U5025 ( .A(n4889), .B(P2_IR_REG_19__SCAN_IN), .ZN(n10367) );
  NOR2_X1 U5026 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9972) );
  OR2_X1 U5027 ( .A1(n8566), .A2(n10432), .ZN(n4614) );
  OR2_X1 U5028 ( .A1(n4815), .A2(n4673), .ZN(n9532) );
  AND2_X1 U5029 ( .A1(n9439), .A2(n10295), .ZN(n4815) );
  OR2_X1 U5030 ( .A1(n8165), .A2(n4698), .ZN(n4697) );
  OAI21_X1 U5031 ( .B1(n8426), .B2(n4792), .A(n4789), .ZN(n4788) );
  INV_X1 U5032 ( .A(n8159), .ZN(n8165) );
  NAND2_X1 U5033 ( .A1(n4816), .A2(n4674), .ZN(n4673) );
  NOR2_X1 U5034 ( .A1(n9442), .A2(n4675), .ZN(n4674) );
  NAND2_X1 U5035 ( .A1(n9214), .A2(n9213), .ZN(n9320) );
  NOR2_X1 U5036 ( .A1(n9321), .A2(n9238), .ZN(n9295) );
  INV_X1 U5037 ( .A(n4790), .ZN(n4789) );
  NAND2_X1 U5038 ( .A1(n4793), .A2(n8394), .ZN(n4792) );
  AOI21_X1 U5039 ( .B1(n9369), .B2(n9234), .A(n9233), .ZN(n9360) );
  OAI21_X1 U5040 ( .B1(n7706), .B2(n8853), .A(n8969), .ZN(n7746) );
  AOI21_X1 U5041 ( .B1(n5046), .B2(n5049), .A(n5045), .ZN(n7607) );
  NAND2_X1 U5042 ( .A1(n6183), .A2(n6182), .ZN(n8618) );
  OR2_X1 U5043 ( .A1(n7170), .A2(n4639), .ZN(n7287) );
  NAND2_X1 U5044 ( .A1(n6074), .A2(n6073), .ZN(n7274) );
  INV_X1 U5045 ( .A(n8108), .ZN(n4486) );
  NAND2_X2 U5046 ( .A1(n6360), .A2(n8468), .ZN(n10376) );
  AOI21_X1 U5047 ( .B1(n7944), .B2(n7943), .A(n7942), .ZN(n7948) );
  AND2_X1 U5048 ( .A1(n6626), .A2(n5288), .ZN(n5302) );
  AND2_X2 U5049 ( .A1(n7027), .A2(n10237), .ZN(n10215) );
  OR2_X1 U5050 ( .A1(n6382), .A2(n6381), .ZN(n6383) );
  AND4_X1 U5051 ( .A1(n6042), .A2(n6041), .A3(n6040), .A4(n6039), .ZN(n8225)
         );
  AND4_X1 U5052 ( .A1(n6014), .A2(n6013), .A3(n6012), .A4(n6011), .ZN(n7966)
         );
  NAND4_X1 U5053 ( .A1(n5994), .A2(n5993), .A3(n5992), .A4(n5991), .ZN(n8258)
         );
  NAND4_X1 U5054 ( .A1(n5966), .A2(n5965), .A3(n5964), .A4(n5963), .ZN(n5971)
         );
  NAND4_X1 U5055 ( .A1(n5957), .A2(n5956), .A3(n5955), .A4(n5954), .ZN(n8262)
         );
  INV_X1 U5056 ( .A(n6865), .ZN(n5984) );
  NAND2_X1 U5057 ( .A1(n5277), .A2(n5276), .ZN(n6932) );
  INV_X1 U5058 ( .A(n10257), .ZN(n7018) );
  AND3_X1 U5059 ( .A1(n6025), .A2(n6024), .A3(n6023), .ZN(n6824) );
  INV_X1 U5060 ( .A(n5285), .ZN(n5767) );
  AND3_X1 U5061 ( .A1(n5336), .A2(n5335), .A3(n5334), .ZN(n10264) );
  AND2_X2 U5062 ( .A1(n5285), .A2(n6923), .ZN(n5278) );
  AND3_X1 U5063 ( .A1(n5317), .A2(n5316), .A3(n5315), .ZN(n10257) );
  AND3_X1 U5064 ( .A1(n5983), .A2(n5982), .A3(n5981), .ZN(n6865) );
  NAND2_X2 U5065 ( .A1(n6922), .A2(n6936), .ZN(n7043) );
  INV_X1 U5066 ( .A(n7912), .ZN(n5922) );
  INV_X1 U5067 ( .A(n5491), .ZN(n4487) );
  OR2_X2 U5068 ( .A1(n8097), .A2(n8350), .ZN(n8093) );
  NAND2_X2 U5069 ( .A1(n5227), .A2(n9561), .ZN(n6526) );
  NAND2_X1 U5070 ( .A1(n8141), .A2(n10367), .ZN(n8128) );
  AND2_X2 U5071 ( .A1(n8151), .A2(n9561), .ZN(n5325) );
  XNOR2_X1 U5072 ( .A(n5204), .B(n5203), .ZN(n6468) );
  AND2_X1 U5073 ( .A1(n6323), .A2(n4504), .ZN(n8103) );
  OR2_X1 U5074 ( .A1(n5209), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5211) );
  XNOR2_X1 U5075 ( .A(n4891), .B(n6321), .ZN(n8131) );
  XNOR2_X1 U5076 ( .A(n5895), .B(n5891), .ZN(n6351) );
  NAND2_X1 U5077 ( .A1(n4504), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4891) );
  OR2_X1 U5078 ( .A1(n6307), .A2(n5917), .ZN(n4889) );
  INV_X1 U5079 ( .A(n5215), .ZN(n5196) );
  AND2_X1 U5080 ( .A1(n5057), .A2(n4805), .ZN(n4804) );
  NAND2_X2 U5081 ( .A1(n4677), .A2(n4676), .ZN(n5086) );
  AND2_X1 U5082 ( .A1(n5414), .A2(n5184), .ZN(n5463) );
  AND3_X1 U5083 ( .A1(n5187), .A2(n5186), .A3(n5185), .ZN(n5191) );
  AND4_X1 U5084 ( .A1(n5884), .A2(n6117), .A3(n6045), .A4(n6131), .ZN(n5885)
         );
  AND4_X1 U5085 ( .A1(n5562), .A2(n5189), .A3(n5565), .A4(n5188), .ZN(n5190)
         );
  NAND3_X1 U5086 ( .A1(n5192), .A2(n4647), .A3(n4648), .ZN(n5352) );
  NOR2_X1 U5087 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5884) );
  INV_X1 U5088 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5240) );
  INV_X4 U5089 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U5090 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5839) );
  INV_X4 U5091 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U5092 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5186) );
  NOR2_X1 U5093 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5185) );
  NOR2_X1 U5094 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5184) );
  NOR2_X1 U5095 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5414) );
  AND2_X1 U5096 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n9971) );
  NAND2_X2 U5097 ( .A1(n8450), .A2(n8449), .ZN(n8451) );
  NOR3_X2 U5098 ( .A1(n7997), .A2(n7996), .A3(n7995), .ZN(n8000) );
  OAI22_X2 U5099 ( .A1(n8378), .A2(n4636), .B1(n8572), .B2(n8244), .ZN(n8362)
         );
  AND2_X2 U5100 ( .A1(n5921), .A2(n7912), .ZN(n5950) );
  NAND2_X1 U5101 ( .A1(n5920), .A2(n5922), .ZN(n5974) );
  NAND2_X1 U5102 ( .A1(n6376), .A2(n8140), .ZN(n4489) );
  NAND2_X2 U5103 ( .A1(n6376), .A2(n8140), .ZN(n4490) );
  NAND2_X1 U5104 ( .A1(n6376), .A2(n8140), .ZN(n7853) );
  XNOR2_X2 U5105 ( .A(n4775), .B(n5893), .ZN(n6350) );
  XNOR2_X2 U5106 ( .A(n5915), .B(n5914), .ZN(n5921) );
  INV_X1 U5107 ( .A(n5894), .ZN(n5892) );
  NAND2_X1 U5108 ( .A1(n4841), .A2(n4840), .ZN(n5734) );
  AOI21_X1 U5109 ( .B1(n4496), .B2(n4846), .A(n4563), .ZN(n4840) );
  NAND2_X1 U5110 ( .A1(n4880), .A2(n4877), .ZN(n4876) );
  AND2_X1 U5111 ( .A1(n4879), .A2(n4875), .ZN(n4874) );
  NOR2_X1 U5112 ( .A1(n4852), .A2(n7873), .ZN(n4851) );
  INV_X1 U5113 ( .A(n4854), .ZN(n4852) );
  AND2_X1 U5114 ( .A1(n4680), .A2(n5466), .ZN(n4685) );
  NAND2_X1 U5115 ( .A1(n4864), .A2(n5103), .ZN(n4680) );
  NAND2_X1 U5116 ( .A1(n9972), .A2(n5073), .ZN(n4677) );
  INV_X1 U5117 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5073) );
  NAND2_X1 U5118 ( .A1(n9971), .A2(n5074), .ZN(n4676) );
  INV_X1 U5119 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5074) );
  NAND2_X1 U5120 ( .A1(n7910), .A2(n7848), .ZN(n7849) );
  OR2_X1 U5121 ( .A1(n8397), .A2(n8204), .ZN(n8071) );
  NOR2_X1 U5122 ( .A1(n8490), .A2(n4786), .ZN(n4785) );
  AND2_X1 U5123 ( .A1(n4787), .A2(n4508), .ZN(n4786) );
  NOR2_X1 U5124 ( .A1(n8521), .A2(n8618), .ZN(n4773) );
  OR2_X1 U5125 ( .A1(n8618), .A2(n8514), .ZN(n8507) );
  OR2_X1 U5126 ( .A1(n7683), .A2(n7729), .ZN(n8024) );
  INV_X1 U5127 ( .A(n4938), .ZN(n4937) );
  INV_X1 U5128 ( .A(n8712), .ZN(n4977) );
  OR2_X1 U5129 ( .A1(n9450), .A2(n9259), .ZN(n9043) );
  INV_X1 U5130 ( .A(n5039), .ZN(n5034) );
  OR2_X1 U5131 ( .A1(n9305), .A2(n9218), .ZN(n9031) );
  AOI21_X1 U5132 ( .B1(n4821), .B2(n4818), .A(n9230), .ZN(n4817) );
  INV_X1 U5133 ( .A(n4825), .ZN(n4818) );
  NAND2_X1 U5134 ( .A1(n9418), .A2(n7788), .ZN(n5027) );
  INV_X1 U5135 ( .A(n7746), .ZN(n7709) );
  OR2_X1 U5136 ( .A1(n10020), .A2(n7555), .ZN(n8962) );
  XNOR2_X1 U5137 ( .A(n6920), .B(n10251), .ZN(n7013) );
  OR2_X1 U5138 ( .A1(n9444), .A2(n9275), .ZN(n9242) );
  NAND2_X1 U5139 ( .A1(n4546), .A2(n5195), .ZN(n5012) );
  OAI21_X1 U5140 ( .B1(n5261), .B2(n5168), .A(n5170), .ZN(n5775) );
  NAND2_X1 U5141 ( .A1(n5146), .A2(n5145), .ZN(n5654) );
  OAI21_X1 U5142 ( .B1(n5125), .B2(n4691), .A(n4689), .ZN(n5600) );
  INV_X1 U5143 ( .A(n4690), .ZN(n4689) );
  OAI21_X1 U5144 ( .B1(n4693), .B2(n4691), .A(n5133), .ZN(n4690) );
  NAND2_X1 U5145 ( .A1(n4692), .A2(n5128), .ZN(n4691) );
  NAND2_X1 U5146 ( .A1(n5133), .A2(n5132), .ZN(n5582) );
  INV_X1 U5147 ( .A(n5520), .ZN(n4619) );
  AND2_X1 U5148 ( .A1(n5124), .A2(n5123), .ZN(n5542) );
  NAND2_X1 U5149 ( .A1(n5100), .A2(n9844), .ZN(n5103) );
  NOR2_X1 U5150 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5236) );
  INV_X1 U5151 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4648) );
  INV_X1 U5152 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4647) );
  NAND2_X1 U5153 ( .A1(n7336), .A2(n4893), .ZN(n7485) );
  NOR2_X1 U5154 ( .A1(n6441), .A2(n4894), .ZN(n4893) );
  INV_X1 U5155 ( .A(n6434), .ZN(n4894) );
  XNOR2_X1 U5156 ( .A(n7849), .B(n4507), .ZN(n8176) );
  NAND2_X1 U5157 ( .A1(n4904), .A2(n8184), .ZN(n4903) );
  NAND2_X1 U5158 ( .A1(n8163), .A2(n8164), .ZN(n4904) );
  INV_X1 U5159 ( .A(n4903), .ZN(n4900) );
  AND2_X1 U5160 ( .A1(n6443), .A2(n6438), .ZN(n6450) );
  NAND2_X1 U5161 ( .A1(n4607), .A2(n4606), .ZN(n8159) );
  INV_X1 U5162 ( .A(n7855), .ZN(n4606) );
  INV_X1 U5163 ( .A(n7854), .ZN(n4607) );
  INV_X1 U5164 ( .A(n6016), .ZN(n5923) );
  INV_X1 U5165 ( .A(n5962), .ZN(n6353) );
  NAND2_X1 U5166 ( .A1(n8384), .A2(n4769), .ZN(n4768) );
  INV_X1 U5167 ( .A(n4795), .ZN(n4794) );
  OAI21_X1 U5168 ( .B1(n4796), .B2(n4799), .A(n6242), .ZN(n4795) );
  OR2_X1 U5169 ( .A1(n8583), .A2(n8437), .ZN(n6242) );
  OR2_X1 U5170 ( .A1(n8583), .A2(n6241), .ZN(n8402) );
  NOR2_X1 U5171 ( .A1(n8427), .A2(n8583), .ZN(n6359) );
  NOR2_X2 U5172 ( .A1(n8593), .A2(n8465), .ZN(n8452) );
  OR2_X1 U5173 ( .A1(n8467), .A2(n8179), .ZN(n8444) );
  NOR2_X1 U5174 ( .A1(n8545), .A2(n8521), .ZN(n4787) );
  OR2_X1 U5175 ( .A1(n8618), .A2(n8247), .ZN(n6190) );
  OR2_X1 U5176 ( .A1(n8538), .A2(n8514), .ZN(n5058) );
  AND2_X1 U5177 ( .A1(n4557), .A2(n5891), .ZN(n4956) );
  OR2_X1 U5178 ( .A1(n5769), .A2(n4977), .ZN(n4976) );
  OR2_X1 U5179 ( .A1(n8832), .A2(n6590), .ZN(n5290) );
  NOR2_X1 U5180 ( .A1(n4560), .A2(n5042), .ZN(n5041) );
  AND2_X1 U5181 ( .A1(n9507), .A2(n9421), .ZN(n7786) );
  INV_X1 U5182 ( .A(n5047), .ZN(n5045) );
  INV_X1 U5183 ( .A(n7559), .ZN(n5046) );
  AOI21_X1 U5184 ( .B1(n5049), .B2(n5048), .A(n5052), .ZN(n5047) );
  INV_X1 U5185 ( .A(n4485), .ZN(n5673) );
  INV_X1 U5186 ( .A(n5439), .ZN(n8866) );
  OAI21_X1 U5187 ( .B1(n5032), .B2(n5029), .A(n5028), .ZN(n7073) );
  AOI21_X1 U5188 ( .B1(n5030), .B2(n10208), .A(n4538), .ZN(n5028) );
  INV_X1 U5189 ( .A(n5030), .ZN(n5029) );
  NAND2_X1 U5190 ( .A1(n4482), .A2(n7875), .ZN(n5439) );
  XNOR2_X1 U5191 ( .A(n7881), .B(n7880), .ZN(n8682) );
  OAI21_X1 U5192 ( .B1(n7884), .B2(n9845), .A(n7878), .ZN(n7881) );
  AND2_X1 U5193 ( .A1(n5056), .A2(n5203), .ZN(n5055) );
  OAI21_X1 U5194 ( .B1(n5734), .B2(n5733), .A(n5161), .ZN(n5756) );
  AND2_X1 U5195 ( .A1(n5165), .A2(n5164), .ZN(n5755) );
  XNOR2_X1 U5196 ( .A(n5094), .B(n5093), .ZN(n5369) );
  NAND2_X1 U5197 ( .A1(n10148), .A2(n10149), .ZN(n10146) );
  MUX2_X1 U5198 ( .A(n7991), .B(n7990), .S(n8093), .Z(n7992) );
  INV_X1 U5199 ( .A(n7982), .ZN(n4873) );
  OAI211_X1 U5200 ( .C1(n4871), .C2(n4869), .A(n4868), .B(n8003), .ZN(n8005)
         );
  NAND2_X1 U5201 ( .A1(n7992), .A2(n4866), .ZN(n4868) );
  INV_X1 U5202 ( .A(n4869), .ZN(n4866) );
  NAND2_X1 U5203 ( .A1(n8001), .A2(n4870), .ZN(n4869) );
  NAND2_X1 U5204 ( .A1(n8013), .A2(n8089), .ZN(n4888) );
  NOR2_X1 U5205 ( .A1(n8120), .A2(n8028), .ZN(n4887) );
  NAND2_X1 U5206 ( .A1(n4880), .A2(n8064), .ZN(n4875) );
  NAND2_X1 U5207 ( .A1(n4965), .A2(n4964), .ZN(n4963) );
  OAI21_X1 U5208 ( .B1(n4491), .B2(n4962), .A(n4965), .ZN(n4961) );
  INV_X1 U5209 ( .A(n4963), .ZN(n4960) );
  NAND2_X1 U5210 ( .A1(n4636), .A2(n8069), .ZN(n4635) );
  INV_X1 U5211 ( .A(n5005), .ZN(n5002) );
  NAND2_X1 U5212 ( .A1(n4685), .A2(n4683), .ZN(n4682) );
  INV_X1 U5213 ( .A(n5103), .ZN(n4683) );
  AND2_X1 U5214 ( .A1(n4836), .A2(n5498), .ZN(n4492) );
  NAND2_X1 U5215 ( .A1(n5109), .A2(n9669), .ZN(n5112) );
  INV_X1 U5216 ( .A(n6388), .ZN(n4923) );
  INV_X1 U5217 ( .A(n4927), .ZN(n4576) );
  INV_X1 U5218 ( .A(n7841), .ZN(n4598) );
  INV_X1 U5219 ( .A(n4601), .ZN(n4597) );
  INV_X1 U5220 ( .A(n7840), .ZN(n4595) );
  INV_X1 U5221 ( .A(n7839), .ZN(n4594) );
  OAI21_X1 U5222 ( .B1(n4794), .B2(n4791), .A(n4541), .ZN(n4790) );
  OR2_X1 U5223 ( .A1(n8587), .A2(n8210), .ZN(n8062) );
  AND2_X1 U5224 ( .A1(n8495), .A2(n4773), .ZN(n4772) );
  NOR2_X1 U5225 ( .A1(n8117), .A2(n8020), .ZN(n4626) );
  AND2_X1 U5226 ( .A1(n7927), .A2(n4628), .ZN(n4627) );
  AND2_X1 U5227 ( .A1(n8019), .A2(n7419), .ZN(n4628) );
  OR2_X1 U5228 ( .A1(n4946), .A2(n8020), .ZN(n4625) );
  INV_X1 U5229 ( .A(n6128), .ZN(n4811) );
  OR2_X1 U5230 ( .A1(n8003), .A2(n8004), .ZN(n7993) );
  NAND2_X1 U5231 ( .A1(n5900), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6052) );
  INV_X1 U5232 ( .A(n6037), .ZN(n5900) );
  INV_X1 U5233 ( .A(n4991), .ZN(n4988) );
  OR2_X1 U5234 ( .A1(n8747), .A2(n4982), .ZN(n4981) );
  NAND2_X1 U5235 ( .A1(n4518), .A2(n4982), .ZN(n4979) );
  NAND2_X1 U5236 ( .A1(n7314), .A2(n5475), .ZN(n5009) );
  AND2_X1 U5237 ( .A1(n5863), .A2(n6936), .ZN(n5285) );
  NOR2_X1 U5238 ( .A1(n5001), .A2(n4997), .ZN(n4996) );
  INV_X1 U5239 ( .A(n7636), .ZN(n4997) );
  INV_X1 U5240 ( .A(n4721), .ZN(n9166) );
  NOR2_X1 U5241 ( .A1(n5037), .A2(n9221), .ZN(n5036) );
  INV_X1 U5242 ( .A(n9219), .ZN(n5037) );
  NOR2_X1 U5243 ( .A1(n9474), .A2(n9481), .ZN(n4753) );
  AND2_X1 U5244 ( .A1(n9358), .A2(n9348), .ZN(n9236) );
  OR2_X1 U5245 ( .A1(n9481), .A2(n9385), .ZN(n8879) );
  NOR2_X1 U5246 ( .A1(n9229), .A2(n4826), .ZN(n4825) );
  OAI21_X1 U5247 ( .B1(n9227), .B2(n9228), .A(n4824), .ZN(n4823) );
  OR2_X1 U5248 ( .A1(n9229), .A2(n8992), .ZN(n4824) );
  AND2_X1 U5249 ( .A1(n10020), .A2(n9133), .ZN(n5052) );
  AND2_X1 U5250 ( .A1(n7022), .A2(n8908), .ZN(n9088) );
  AND2_X1 U5251 ( .A1(n10227), .A2(n8908), .ZN(n4649) );
  OR2_X1 U5252 ( .A1(n10225), .A2(n10264), .ZN(n9083) );
  NAND2_X1 U5253 ( .A1(n7018), .A2(n7019), .ZN(n9082) );
  NAND2_X1 U5254 ( .A1(n9082), .A2(n9080), .ZN(n7033) );
  INV_X1 U5255 ( .A(n9224), .ZN(n9244) );
  OR2_X1 U5256 ( .A1(n9397), .A2(n9486), .ZN(n9386) );
  AND2_X1 U5257 ( .A1(n6932), .A2(n6946), .ZN(n6921) );
  XNOR2_X1 U5258 ( .A(n7877), .B(n7876), .ZN(n7884) );
  AOI21_X1 U5259 ( .B1(n4855), .B2(n6275), .A(n4571), .ZN(n4854) );
  INV_X1 U5260 ( .A(n5798), .ZN(n4855) );
  INV_X1 U5261 ( .A(n6275), .ZN(n4856) );
  NAND2_X1 U5262 ( .A1(n5245), .A2(n5244), .ZN(n5180) );
  NAND2_X1 U5263 ( .A1(n5236), .A2(n5240), .ZN(n5193) );
  INV_X1 U5264 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5565) );
  INV_X1 U5265 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5562) );
  NOR2_X1 U5266 ( .A1(n5129), .A2(n4694), .ZN(n4693) );
  INV_X1 U5267 ( .A(n5124), .ZN(n4694) );
  INV_X1 U5268 ( .A(n5560), .ZN(n5129) );
  NAND2_X1 U5269 ( .A1(n5119), .A2(n5118), .ZN(n5520) );
  AOI21_X1 U5270 ( .B1(n5476), .B2(n4838), .A(n4837), .ZN(n4836) );
  INV_X1 U5271 ( .A(n5112), .ZN(n4837) );
  INV_X1 U5272 ( .A(n5107), .ZN(n4838) );
  INV_X1 U5273 ( .A(n5476), .ZN(n4839) );
  NAND2_X1 U5274 ( .A1(n4681), .A2(n4685), .ZN(n5108) );
  NAND2_X1 U5275 ( .A1(n5438), .A2(n5103), .ZN(n4681) );
  NAND2_X1 U5276 ( .A1(n5086), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4609) );
  NAND2_X1 U5277 ( .A1(n5907), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U5278 ( .A1(n6375), .A2(n8131), .ZN(n6376) );
  AND2_X1 U5279 ( .A1(n4516), .A2(n4604), .ZN(n4601) );
  OR2_X1 U5280 ( .A1(n4602), .A2(n4600), .ZN(n4599) );
  INV_X1 U5281 ( .A(n4604), .ZN(n4600) );
  AND2_X1 U5282 ( .A1(n7773), .A2(n4605), .ZN(n4602) );
  AND2_X1 U5283 ( .A1(n7865), .A2(n6413), .ZN(n6414) );
  NAND2_X1 U5284 ( .A1(n7155), .A2(n6430), .ZN(n7336) );
  OR2_X1 U5285 ( .A1(n6091), .A2(n6090), .ZN(n6109) );
  AND2_X1 U5286 ( .A1(n7049), .A2(n6418), .ZN(n4913) );
  NOR2_X1 U5287 ( .A1(n6414), .A2(n4910), .ZN(n4909) );
  INV_X1 U5288 ( .A(n6418), .ZN(n4910) );
  INV_X1 U5289 ( .A(n6423), .ZN(n4912) );
  AND2_X1 U5290 ( .A1(n7517), .A2(n4932), .ZN(n4929) );
  INV_X1 U5291 ( .A(n7821), .ZN(n4931) );
  XNOR2_X1 U5292 ( .A(n7737), .B(n7720), .ZN(n7823) );
  AND2_X1 U5293 ( .A1(n6240), .A2(n6239), .ZN(n6241) );
  OR3_X1 U5294 ( .A1(n7551), .A2(n7688), .A3(n7630), .ZN(n6650) );
  OR2_X1 U5295 ( .A1(n6717), .A2(n6716), .ZN(n4715) );
  NAND2_X1 U5296 ( .A1(n8298), .A2(n4711), .ZN(n4710) );
  AOI21_X1 U5297 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n8324), .A(n8323), .ZN(
        n8338) );
  NAND2_X1 U5298 ( .A1(n4798), .A2(n4797), .ZN(n4796) );
  NAND2_X1 U5299 ( .A1(n4799), .A2(n8434), .ZN(n4797) );
  AND2_X1 U5300 ( .A1(n8420), .A2(n6348), .ZN(n8404) );
  NOR2_X1 U5301 ( .A1(n8427), .A2(n4767), .ZN(n8396) );
  INV_X1 U5302 ( .A(n4769), .ZN(n4767) );
  NAND2_X1 U5303 ( .A1(n8417), .A2(n8098), .ZN(n8420) );
  NOR2_X1 U5304 ( .A1(n4801), .A2(n8587), .ZN(n4800) );
  OAI21_X1 U5305 ( .B1(n8459), .B2(n4498), .A(n4953), .ZN(n8435) );
  OR2_X1 U5306 ( .A1(n6345), .A2(n4954), .ZN(n4953) );
  INV_X1 U5307 ( .A(n8060), .ZN(n4954) );
  AND2_X1 U5308 ( .A1(n8062), .A2(n8059), .ZN(n8434) );
  NOR2_X1 U5309 ( .A1(n8426), .A2(n8434), .ZN(n8425) );
  INV_X1 U5310 ( .A(n8459), .ZN(n4955) );
  AOI21_X1 U5311 ( .B1(n4785), .B2(n4782), .A(n4547), .ZN(n4781) );
  INV_X1 U5312 ( .A(n4508), .ZN(n4782) );
  INV_X1 U5313 ( .A(n4785), .ZN(n4783) );
  NAND2_X1 U5314 ( .A1(n6341), .A2(n8490), .ZN(n8501) );
  INV_X1 U5315 ( .A(n8497), .ZN(n6341) );
  AND2_X1 U5316 ( .A1(n6210), .A2(n6209), .ZN(n8499) );
  NAND2_X1 U5317 ( .A1(n4612), .A2(n4942), .ZN(n8512) );
  AND2_X1 U5318 ( .A1(n6340), .A2(n4943), .ZN(n4942) );
  NAND2_X1 U5319 ( .A1(n8540), .A2(n8031), .ZN(n4943) );
  NAND2_X1 U5320 ( .A1(n7726), .A2(n8030), .ZN(n8541) );
  NAND2_X1 U5321 ( .A1(n8541), .A2(n8540), .ZN(n8539) );
  AOI21_X1 U5322 ( .B1(n4493), .B2(n8118), .A(n4537), .ZN(n4808) );
  NAND2_X1 U5323 ( .A1(n7728), .A2(n7727), .ZN(n7726) );
  OR2_X1 U5324 ( .A1(n7668), .A2(n8118), .ZN(n4809) );
  NAND2_X1 U5325 ( .A1(n7540), .A2(n6337), .ZN(n7538) );
  INV_X1 U5326 ( .A(n4947), .ZN(n6337) );
  OAI21_X1 U5327 ( .B1(n7360), .B2(n7359), .A(n6116), .ZN(n7416) );
  NAND2_X1 U5328 ( .A1(n4506), .A2(n7419), .ZN(n7540) );
  INV_X1 U5329 ( .A(n6059), .ZN(n4803) );
  NAND2_X1 U5330 ( .A1(n5902), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6075) );
  INV_X1 U5331 ( .A(n6064), .ZN(n5902) );
  NAND2_X1 U5332 ( .A1(n4940), .A2(n4939), .ZN(n4938) );
  INV_X1 U5333 ( .A(n8515), .ZN(n8544) );
  NAND2_X1 U5334 ( .A1(n6281), .A2(n6280), .ZN(n8562) );
  AND2_X1 U5335 ( .A1(n4615), .A2(n4565), .ZN(n8565) );
  NAND2_X1 U5336 ( .A1(n4616), .A2(n10369), .ZN(n4615) );
  NAND2_X1 U5337 ( .A1(n5930), .A2(n5929), .ZN(n8521) );
  NAND2_X1 U5338 ( .A1(n6148), .A2(n6147), .ZN(n8638) );
  NAND2_X1 U5339 ( .A1(n6120), .A2(n6119), .ZN(n7424) );
  INV_X1 U5340 ( .A(n10460), .ZN(n8644) );
  NOR2_X1 U5341 ( .A1(n7688), .A2(n6312), .ZN(n10391) );
  AND2_X1 U5342 ( .A1(n7630), .A2(n6311), .ZN(n6312) );
  OAI21_X1 U5343 ( .B1(n5912), .B2(P2_IR_REG_28__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n4777) );
  AND2_X1 U5344 ( .A1(n6303), .A2(n5890), .ZN(n4805) );
  INV_X1 U5345 ( .A(n5928), .ZN(n4941) );
  INV_X1 U5346 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6303) );
  OAI21_X2 U5347 ( .B1(n4504), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6320) );
  INV_X1 U5348 ( .A(n5541), .ZN(n5004) );
  NAND2_X1 U5349 ( .A1(n5323), .A2(n5324), .ZN(n4968) );
  NOR2_X1 U5350 ( .A1(n4988), .A2(n4985), .ZN(n4984) );
  INV_X1 U5351 ( .A(n8739), .ZN(n4985) );
  OR2_X1 U5352 ( .A1(n4989), .A2(n4988), .ZN(n4987) );
  NAND2_X1 U5353 ( .A1(n4969), .A2(n4972), .ZN(n8753) );
  INV_X1 U5354 ( .A(n4973), .ZN(n4972) );
  OAI21_X1 U5355 ( .B1(n4976), .B2(n4974), .A(n8755), .ZN(n4973) );
  AND2_X1 U5356 ( .A1(n8814), .A2(n4993), .ZN(n4989) );
  OR2_X1 U5357 ( .A1(n5856), .A2(n7203), .ZN(n5307) );
  OAI21_X1 U5358 ( .B1(n6505), .B2(n6476), .A(n9146), .ZN(n10072) );
  NAND2_X1 U5359 ( .A1(n9158), .A2(n6479), .ZN(n6579) );
  OR2_X1 U5360 ( .A1(n6579), .A2(n6578), .ZN(n4582) );
  AND2_X1 U5361 ( .A1(n4582), .A2(n4581), .ZN(n6565) );
  NAND2_X1 U5362 ( .A1(n6588), .A2(n6480), .ZN(n4581) );
  AND2_X1 U5363 ( .A1(n6467), .A2(n6583), .ZN(n6570) );
  NOR2_X1 U5364 ( .A1(n9178), .A2(n4568), .ZN(n9181) );
  AOI21_X1 U5365 ( .B1(n9177), .B2(P1_REG2_REG_17__SCAN_IN), .A(n10138), .ZN(
        n10153) );
  NOR2_X1 U5366 ( .A1(n9251), .A2(n4737), .ZN(n4736) );
  NAND2_X1 U5367 ( .A1(n4738), .A2(n9284), .ZN(n4737) );
  AND2_X1 U5368 ( .A1(n9058), .A2(n8928), .ZN(n9224) );
  NAND2_X1 U5369 ( .A1(n9046), .A2(n9241), .ZN(n4667) );
  NAND2_X1 U5370 ( .A1(n9046), .A2(n9222), .ZN(n4668) );
  OAI21_X1 U5371 ( .B1(n9324), .B2(n4829), .A(n4827), .ZN(n9273) );
  AOI21_X1 U5372 ( .B1(n4830), .B2(n9238), .A(n4828), .ZN(n4827) );
  INV_X1 U5373 ( .A(n4830), .ZN(n4829) );
  INV_X1 U5374 ( .A(n9239), .ZN(n4828) );
  AND4_X1 U5375 ( .A1(n5811), .A2(n5810), .A3(n5809), .A4(n5808), .ZN(n9275)
         );
  NOR2_X1 U5376 ( .A1(n9313), .A2(n5040), .ZN(n5039) );
  AND2_X1 U5377 ( .A1(n9031), .A2(n9030), .ZN(n9313) );
  OAI21_X1 U5378 ( .B1(n9360), .B2(n9236), .A(n9235), .ZN(n9346) );
  NAND2_X1 U5379 ( .A1(n9210), .A2(n4527), .ZN(n5043) );
  INV_X1 U5380 ( .A(n9209), .ZN(n5044) );
  NAND2_X1 U5381 ( .A1(n4661), .A2(n4660), .ZN(n9369) );
  NAND2_X1 U5382 ( .A1(n4665), .A2(n4655), .ZN(n4661) );
  AOI21_X1 U5383 ( .B1(n4817), .B2(n9232), .A(n9231), .ZN(n4658) );
  INV_X1 U5384 ( .A(n4821), .ZN(n4819) );
  NOR2_X1 U5385 ( .A1(n7707), .A2(n7708), .ZN(n4664) );
  OR2_X1 U5386 ( .A1(n7709), .A2(n7707), .ZN(n4665) );
  INV_X1 U5387 ( .A(n4817), .ZN(n4659) );
  OR2_X1 U5388 ( .A1(n9491), .A2(n9203), .ZN(n9202) );
  NOR2_X1 U5389 ( .A1(n4823), .A2(n9407), .ZN(n4821) );
  NAND2_X1 U5390 ( .A1(n7780), .A2(n4825), .ZN(n4822) );
  INV_X1 U5391 ( .A(n4823), .ZN(n4820) );
  NAND2_X1 U5392 ( .A1(n4549), .A2(n5027), .ZN(n5024) );
  AND2_X1 U5393 ( .A1(n8874), .A2(n8883), .ZN(n9419) );
  AOI21_X1 U5394 ( .B1(n7709), .B2(n7708), .A(n7707), .ZN(n7780) );
  OR2_X1 U5395 ( .A1(n7804), .A2(n9131), .ZN(n7704) );
  NAND2_X1 U5396 ( .A1(n7612), .A2(n8965), .ZN(n7706) );
  NOR2_X1 U5397 ( .A1(n10021), .A2(n9516), .ZN(n7608) );
  OR2_X1 U5398 ( .A1(n7563), .A2(n10020), .ZN(n10021) );
  INV_X1 U5399 ( .A(n7560), .ZN(n5050) );
  AND2_X1 U5400 ( .A1(n7165), .A2(n7164), .ZN(n5053) );
  NAND2_X1 U5401 ( .A1(n4747), .A2(n4745), .ZN(n7239) );
  AND2_X1 U5402 ( .A1(n4746), .A2(n10292), .ZN(n4745) );
  INV_X1 U5403 ( .A(n4748), .ZN(n4746) );
  AND3_X1 U5404 ( .A1(n5375), .A2(n5374), .A3(n5373), .ZN(n10189) );
  AND2_X1 U5405 ( .A1(n10178), .A2(n4515), .ZN(n5030) );
  NOR2_X1 U5406 ( .A1(n10218), .A2(n10200), .ZN(n10197) );
  INV_X1 U5407 ( .A(n9358), .ZN(n9474) );
  NAND2_X1 U5408 ( .A1(n5605), .A2(n5604), .ZN(n9507) );
  AND2_X1 U5409 ( .A1(n5482), .A2(n5481), .ZN(n10002) );
  AND2_X1 U5410 ( .A1(n5055), .A2(n4654), .ZN(n4653) );
  AND2_X1 U5411 ( .A1(n4551), .A2(n9885), .ZN(n4654) );
  NOR2_X1 U5412 ( .A1(n5220), .A2(n5464), .ZN(n5016) );
  NAND2_X1 U5413 ( .A1(n9552), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5015) );
  NAND3_X1 U5414 ( .A1(n5196), .A2(n9885), .A3(n5055), .ZN(n5219) );
  INV_X1 U5415 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5220) );
  INV_X1 U5416 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9885) );
  NOR2_X1 U5417 ( .A1(n5199), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n5056) );
  INV_X1 U5418 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5203) );
  NAND2_X1 U5419 ( .A1(n4842), .A2(n4843), .ZN(n5715) );
  OR2_X1 U5420 ( .A1(n5654), .A2(n4846), .ZN(n4842) );
  OAI21_X1 U5421 ( .B1(n5654), .B2(n5653), .A(n5151), .ZN(n5696) );
  XNOR2_X1 U5422 ( .A(n5633), .B(n5632), .ZN(n6885) );
  NAND2_X1 U5423 ( .A1(n5138), .A2(n5137), .ZN(n5633) );
  NAND2_X1 U5424 ( .A1(n5102), .A2(n5103), .ZN(n4864) );
  AND2_X1 U5425 ( .A1(n5237), .A2(n5236), .ZN(n5462) );
  XNOR2_X1 U5426 ( .A(n5091), .B(n9944), .ZN(n5389) );
  NAND2_X1 U5427 ( .A1(n5090), .A2(n5089), .ZN(n5390) );
  INV_X1 U5428 ( .A(n5082), .ZN(n4645) );
  XNOR2_X1 U5429 ( .A(n5314), .B(P1_IR_REG_2__SCAN_IN), .ZN(n10053) );
  NAND2_X1 U5430 ( .A1(n4648), .A2(n4647), .ZN(n4646) );
  NAND2_X1 U5431 ( .A1(n6221), .A2(n6220), .ZN(n8593) );
  NAND2_X1 U5432 ( .A1(n4900), .A2(n4896), .ZN(n4895) );
  INV_X1 U5433 ( .A(n8196), .ZN(n4896) );
  INV_X1 U5434 ( .A(n4902), .ZN(n4901) );
  OAI21_X1 U5435 ( .B1(n4903), .B2(n8163), .A(n8194), .ZN(n4902) );
  OR2_X1 U5436 ( .A1(n8193), .A2(n8192), .ZN(n8194) );
  AOI21_X1 U5437 ( .B1(n4900), .B2(n4899), .A(n4898), .ZN(n4897) );
  INV_X1 U5438 ( .A(n8195), .ZN(n4898) );
  NOR2_X1 U5439 ( .A1(n8196), .A2(n8163), .ZN(n4899) );
  NAND2_X1 U5440 ( .A1(n6231), .A2(n6230), .ZN(n8583) );
  NAND2_X1 U5441 ( .A1(n4930), .A2(n4929), .ZN(n7822) );
  INV_X1 U5442 ( .A(n8217), .ZN(n7859) );
  NAND2_X1 U5443 ( .A1(n6212), .A2(n6211), .ZN(n8467) );
  NAND2_X1 U5444 ( .A1(n4931), .A2(n7659), .ZN(n4928) );
  AND2_X1 U5445 ( .A1(n6770), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8229) );
  NAND2_X1 U5446 ( .A1(n6244), .A2(n6243), .ZN(n8397) );
  NAND2_X1 U5447 ( .A1(n6442), .A2(n8468), .ZN(n8230) );
  NAND2_X1 U5448 ( .A1(n4699), .A2(n8235), .ZN(n4698) );
  NAND2_X1 U5449 ( .A1(n7854), .A2(n7855), .ZN(n4699) );
  OR2_X1 U5450 ( .A1(n4483), .A2(n5989), .ZN(n5992) );
  OR2_X1 U5451 ( .A1(n4488), .A2(n7110), .ZN(n6018) );
  OR2_X1 U5452 ( .A1(n5962), .A2(n7101), .ZN(n5963) );
  NAND4_X2 U5453 ( .A1(n5941), .A2(n5062), .A3(n5939), .A4(n5940), .ZN(n8261)
         );
  OR2_X1 U5454 ( .A1(n5962), .A2(n5938), .ZN(n5939) );
  OR2_X1 U5455 ( .A1(n4483), .A2(n5952), .ZN(n5956) );
  AOI22_X1 U5456 ( .A1(n5996), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6538), .B2(
        n6694), .ZN(n6006) );
  OR2_X1 U5457 ( .A1(n10390), .A2(n6734), .ZN(n8468) );
  NAND2_X1 U5458 ( .A1(n7883), .A2(n7882), .ZN(n7922) );
  INV_X1 U5459 ( .A(n8558), .ZN(n4757) );
  NAND2_X1 U5460 ( .A1(n4762), .A2(n4760), .ZN(n4759) );
  OR2_X1 U5461 ( .A1(n10469), .A2(n4761), .ZN(n4760) );
  NAND2_X1 U5462 ( .A1(n7922), .A2(n8650), .ZN(n4762) );
  INV_X1 U5463 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n4761) );
  OR2_X1 U5464 ( .A1(n5946), .A2(n6516), .ZN(n5968) );
  AND4_X1 U5465 ( .A1(n5683), .A2(n5682), .A3(n5681), .A4(n5680), .ZN(n9411)
         );
  AND3_X1 U5466 ( .A1(n5357), .A2(n5356), .A3(n5355), .ZN(n10270) );
  INV_X1 U5467 ( .A(n9361), .ZN(n9385) );
  AND2_X1 U5468 ( .A1(n5505), .A2(n5504), .ZN(n7558) );
  AND4_X1 U5469 ( .A1(n5786), .A2(n5785), .A3(n5784), .A4(n5783), .ZN(n9218)
         );
  INV_X1 U5470 ( .A(n8773), .ZN(n8812) );
  OR2_X1 U5471 ( .A1(n5856), .A2(n6596), .ZN(n5293) );
  NAND2_X1 U5472 ( .A1(n9160), .A2(n9159), .ZN(n9158) );
  XNOR2_X1 U5473 ( .A(n9181), .B(n9180), .ZN(n10119) );
  NAND2_X1 U5474 ( .A1(n10119), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n10118) );
  NAND2_X1 U5475 ( .A1(n10130), .A2(n4574), .ZN(n10148) );
  NOR2_X1 U5476 ( .A1(n10166), .A2(n10167), .ZN(n10165) );
  NAND2_X1 U5477 ( .A1(n10079), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4731) );
  OAI21_X1 U5478 ( .B1(n9192), .B2(n10159), .A(n4728), .ZN(n4727) );
  OR2_X1 U5479 ( .A1(n9191), .A2(n10169), .ZN(n4728) );
  OAI21_X1 U5480 ( .B1(n9190), .B2(n9189), .A(n4733), .ZN(n4732) );
  AOI21_X1 U5481 ( .B1(n9191), .B2(n10147), .A(n10129), .ZN(n4733) );
  NOR2_X1 U5482 ( .A1(n7984), .A2(n7983), .ZN(n4867) );
  INV_X1 U5483 ( .A(n7992), .ZN(n4865) );
  AND2_X1 U5484 ( .A1(n4887), .A2(n4556), .ZN(n4883) );
  NAND2_X1 U5485 ( .A1(n4887), .A2(n4530), .ZN(n4885) );
  AND2_X1 U5486 ( .A1(n8098), .A2(n8065), .ZN(n4879) );
  OR2_X1 U5487 ( .A1(n8063), .A2(n8093), .ZN(n4880) );
  INV_X1 U5488 ( .A(n8061), .ZN(n4877) );
  OAI21_X1 U5489 ( .B1(n8058), .B2(n8093), .A(n8446), .ZN(n4882) );
  NOR2_X1 U5490 ( .A1(n8057), .A2(n8089), .ZN(n4878) );
  AOI21_X1 U5491 ( .B1(n8040), .B2(n8039), .A(n8038), .ZN(n8058) );
  NAND2_X1 U5492 ( .A1(n8092), .A2(n8080), .ZN(n8085) );
  NOR2_X1 U5493 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5880) );
  NOR2_X1 U5494 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5881) );
  NOR2_X1 U5495 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5882) );
  INV_X1 U5496 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U5497 ( .A1(n4850), .A2(n4849), .ZN(n7877) );
  AOI21_X1 U5498 ( .B1(n4851), .B2(n4856), .A(n4572), .ZN(n4849) );
  AND2_X1 U5499 ( .A1(n4848), .A2(n5695), .ZN(n4847) );
  NAND2_X1 U5500 ( .A1(n5653), .A2(n5151), .ZN(n4848) );
  NOR2_X1 U5501 ( .A1(n4860), .A2(n4859), .ZN(n4858) );
  INV_X1 U5502 ( .A(n5137), .ZN(n4859) );
  INV_X1 U5503 ( .A(n5632), .ZN(n4860) );
  INV_X1 U5504 ( .A(n5582), .ZN(n4692) );
  NAND2_X1 U5505 ( .A1(n5116), .A2(n9868), .ZN(n5119) );
  INV_X1 U5506 ( .A(SI_8_), .ZN(n9844) );
  INV_X1 U5507 ( .A(SI_10_), .ZN(n9669) );
  INV_X1 U5508 ( .A(n4959), .ZN(n4958) );
  OAI21_X1 U5509 ( .B1(n4963), .B2(n8073), .A(n4961), .ZN(n4959) );
  INV_X1 U5510 ( .A(n8085), .ZN(n8127) );
  NAND2_X1 U5511 ( .A1(n4861), .A2(n7919), .ZN(n8092) );
  INV_X1 U5512 ( .A(n7922), .ZN(n4861) );
  AND2_X1 U5513 ( .A1(n7922), .A2(n7921), .ZN(n8090) );
  NOR2_X1 U5514 ( .A1(n4635), .A2(n4798), .ZN(n4634) );
  NAND2_X1 U5515 ( .A1(n4633), .A2(n4632), .ZN(n4631) );
  INV_X1 U5516 ( .A(n6348), .ZN(n4632) );
  INV_X1 U5517 ( .A(n4635), .ZN(n4633) );
  INV_X1 U5518 ( .A(n4796), .ZN(n4793) );
  INV_X1 U5519 ( .A(n4800), .ZN(n4799) );
  NOR2_X1 U5520 ( .A1(n8397), .A2(n8583), .ZN(n4769) );
  NOR2_X1 U5521 ( .A1(n4944), .A2(n8120), .ZN(n4613) );
  NAND2_X1 U5522 ( .A1(n4812), .A2(n7539), .ZN(n4947) );
  NAND2_X1 U5523 ( .A1(n10454), .A2(n8253), .ZN(n7987) );
  AND2_X1 U5524 ( .A1(n10448), .A2(n6963), .ZN(n4766) );
  NOR2_X1 U5525 ( .A1(n4486), .A2(n7971), .ZN(n4950) );
  NAND2_X1 U5526 ( .A1(n4952), .A2(n6954), .ZN(n4951) );
  NAND2_X1 U5527 ( .A1(n5899), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6037) );
  OR2_X1 U5528 ( .A1(n10363), .A2(n8258), .ZN(n6026) );
  NAND2_X1 U5529 ( .A1(n8258), .A2(n10437), .ZN(n7960) );
  NAND2_X1 U5530 ( .A1(n5985), .A2(n5984), .ZN(n7931) );
  AND2_X1 U5531 ( .A1(n7959), .A2(n7931), .ZN(n8104) );
  XNOR2_X1 U5532 ( .A(n4520), .B(n8125), .ZN(n4616) );
  NAND2_X1 U5533 ( .A1(n4937), .A2(n6306), .ZN(n4933) );
  OR2_X1 U5534 ( .A1(n6047), .A2(n6046), .ZN(n6060) );
  AND2_X1 U5535 ( .A1(n8778), .A2(n4975), .ZN(n4970) );
  NAND2_X1 U5536 ( .A1(n8745), .A2(n5652), .ZN(n8721) );
  NAND2_X1 U5538 ( .A1(n10099), .A2(n4722), .ZN(n4721) );
  NAND2_X1 U5539 ( .A1(n7407), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4722) );
  OR2_X1 U5540 ( .A1(n9251), .A2(n9258), .ZN(n9058) );
  AOI21_X1 U5541 ( .B1(n4831), .B2(n9022), .A(n9240), .ZN(n4830) );
  NAND2_X1 U5542 ( .A1(n4832), .A2(n9237), .ZN(n4831) );
  INV_X1 U5543 ( .A(n9322), .ZN(n4832) );
  INV_X1 U5544 ( .A(n9211), .ZN(n5042) );
  NAND2_X1 U5545 ( .A1(n9345), .A2(n4753), .ZN(n4752) );
  NOR2_X1 U5546 ( .A1(n4819), .A2(n4656), .ZN(n4655) );
  NAND2_X1 U5547 ( .A1(n4662), .A2(n4657), .ZN(n4656) );
  INV_X1 U5548 ( .A(n4664), .ZN(n4657) );
  NOR2_X1 U5549 ( .A1(n9507), .A2(n7804), .ZN(n4743) );
  INV_X1 U5550 ( .A(n5068), .ZN(n5048) );
  NAND2_X1 U5551 ( .A1(n10189), .A2(n10278), .ZN(n4748) );
  NAND2_X1 U5552 ( .A1(n7753), .A2(n9510), .ZN(n7752) );
  AND2_X1 U5553 ( .A1(n7608), .A2(n10029), .ZN(n7753) );
  NAND2_X1 U5554 ( .A1(n7222), .A2(n9083), .ZN(n10230) );
  NOR2_X1 U5555 ( .A1(n7018), .A2(n7205), .ZN(n7216) );
  AND2_X1 U5556 ( .A1(n5798), .A2(n5183), .ZN(n5796) );
  OAI21_X1 U5557 ( .B1(n5775), .B2(n5774), .A(n5174), .ZN(n5245) );
  AND2_X1 U5558 ( .A1(n5179), .A2(n5178), .ZN(n5244) );
  AOI21_X1 U5559 ( .B1(n4847), .B2(n4845), .A(n4844), .ZN(n4843) );
  INV_X1 U5560 ( .A(n5156), .ZN(n4844) );
  INV_X1 U5561 ( .A(n5151), .ZN(n4845) );
  INV_X1 U5562 ( .A(n4847), .ZN(n4846) );
  NAND2_X1 U5563 ( .A1(n5121), .A2(n5120), .ZN(n5124) );
  AOI21_X1 U5564 ( .B1(n4492), .B2(n4839), .A(n4543), .ZN(n4834) );
  OR2_X1 U5565 ( .A1(n4620), .A2(n4678), .ZN(n4618) );
  NAND2_X1 U5566 ( .A1(n4682), .A2(n4492), .ZN(n4678) );
  NAND3_X1 U5567 ( .A1(n4682), .A2(n4492), .A3(n4684), .ZN(n4679) );
  INV_X1 U5568 ( .A(n4685), .ZN(n4684) );
  AND2_X1 U5569 ( .A1(n5107), .A2(n5106), .ZN(n5466) );
  OAI21_X1 U5570 ( .B1(n7875), .B2(P1_DATAO_REG_8__SCAN_IN), .A(n4637), .ZN(
        n5100) );
  NAND2_X1 U5571 ( .A1(n7875), .A2(n6522), .ZN(n4637) );
  INV_X1 U5572 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5440) );
  NOR2_X1 U5573 ( .A1(n4645), .A2(n4505), .ZN(n4644) );
  OR2_X1 U5574 ( .A1(n5330), .A2(n4505), .ZN(n4641) );
  NAND2_X1 U5575 ( .A1(n5282), .A2(n4833), .ZN(n5077) );
  NAND2_X1 U5576 ( .A1(n7485), .A2(n7484), .ZN(n7509) );
  AND2_X1 U5577 ( .A1(n8184), .A2(n8157), .ZN(n8163) );
  NOR2_X1 U5578 ( .A1(n4924), .A2(n4919), .ZN(n4918) );
  OR2_X1 U5579 ( .A1(n6788), .A2(n4914), .ZN(n4919) );
  INV_X1 U5580 ( .A(n6802), .ZN(n4914) );
  NAND2_X1 U5581 ( .A1(n5906), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6184) );
  INV_X1 U5582 ( .A(n6175), .ZN(n5906) );
  INV_X1 U5583 ( .A(n7514), .ZN(n4932) );
  OAI21_X1 U5584 ( .B1(n8176), .B2(n8174), .A(n7850), .ZN(n4687) );
  NAND2_X1 U5585 ( .A1(n4922), .A2(n6392), .ZN(n4921) );
  NAND2_X1 U5586 ( .A1(n6794), .A2(n4923), .ZN(n4922) );
  INV_X1 U5587 ( .A(n6794), .ZN(n4924) );
  NAND2_X1 U5588 ( .A1(n5908), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6213) );
  NAND2_X1 U5589 ( .A1(n4595), .A2(n4594), .ZN(n4593) );
  NAND2_X1 U5590 ( .A1(n4892), .A2(n4608), .ZN(n7854) );
  NAND2_X1 U5591 ( .A1(n8203), .A2(n8201), .ZN(n4892) );
  INV_X1 U5592 ( .A(n8131), .ZN(n7944) );
  OR2_X1 U5593 ( .A1(n6729), .A2(n6728), .ZN(n4707) );
  NAND2_X1 U5594 ( .A1(n4707), .A2(n4706), .ZN(n4705) );
  NAND2_X1 U5595 ( .A1(n6732), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4706) );
  AOI21_X1 U5596 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n6763), .A(n6762), .ZN(
        n6764) );
  AND2_X1 U5597 ( .A1(n6979), .A2(n4716), .ZN(n8265) );
  NAND2_X1 U5598 ( .A1(n6980), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4716) );
  NOR2_X1 U5599 ( .A1(n8265), .A2(n8264), .ZN(n8263) );
  OR2_X1 U5600 ( .A1(n6984), .A2(n6983), .ZN(n4702) );
  NAND2_X1 U5601 ( .A1(n7306), .A2(n4700), .ZN(n7308) );
  OR2_X1 U5602 ( .A1(n7307), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4700) );
  NAND2_X1 U5603 ( .A1(n7574), .A2(n4717), .ZN(n7576) );
  OR2_X1 U5604 ( .A1(n7575), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4717) );
  AND2_X1 U5605 ( .A1(n6274), .A2(n6273), .ZN(n8187) );
  AND2_X1 U5606 ( .A1(n8081), .A2(n4965), .ZN(n8125) );
  AND2_X1 U5607 ( .A1(n6287), .A2(n6286), .ZN(n8372) );
  AOI21_X1 U5608 ( .B1(n8382), .B2(n6262), .A(n6261), .ZN(n8371) );
  AND2_X1 U5609 ( .A1(n4629), .A2(n4630), .ZN(n8370) );
  AND2_X1 U5610 ( .A1(n4631), .A2(n8073), .ZN(n4629) );
  NOR2_X1 U5611 ( .A1(n8370), .A2(n8369), .ZN(n8368) );
  NAND2_X1 U5612 ( .A1(n4630), .A2(n4631), .ZN(n8385) );
  AOI21_X1 U5613 ( .B1(n4495), .B2(n4783), .A(n4542), .ZN(n4778) );
  NOR2_X1 U5614 ( .A1(n8603), .A2(n4771), .ZN(n4770) );
  INV_X1 U5615 ( .A(n4772), .ZN(n4771) );
  NAND2_X1 U5616 ( .A1(n8512), .A2(n8045), .ZN(n8497) );
  NAND2_X1 U5617 ( .A1(n8531), .A2(n4773), .ZN(n8519) );
  NAND2_X1 U5618 ( .A1(n8531), .A2(n8538), .ZN(n8532) );
  AND3_X1 U5619 ( .A1(n6189), .A2(n6188), .A3(n6187), .ZN(n8514) );
  NOR2_X1 U5620 ( .A1(n4626), .A2(n8026), .ZN(n4624) );
  OR2_X1 U5621 ( .A1(n6167), .A2(n9926), .ZN(n6175) );
  AND2_X1 U5622 ( .A1(n4623), .A2(n4622), .ZN(n4621) );
  INV_X1 U5623 ( .A(n4626), .ZN(n4622) );
  OR2_X1 U5624 ( .A1(n6137), .A2(n9929), .ZN(n6150) );
  NAND2_X1 U5625 ( .A1(n5905), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6167) );
  INV_X1 U5626 ( .A(n6150), .ZN(n5905) );
  NOR2_X1 U5627 ( .A1(n4812), .A2(n4811), .ZN(n4810) );
  NOR2_X1 U5628 ( .A1(n7533), .A2(n8638), .ZN(n7679) );
  AND4_X1 U5629 ( .A1(n6156), .A2(n6155), .A3(n6154), .A4(n6153), .ZN(n7672)
         );
  NAND2_X1 U5630 ( .A1(n4764), .A2(n4763), .ZN(n7533) );
  NAND2_X1 U5631 ( .A1(n5903), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6122) );
  INV_X1 U5632 ( .A(n6109), .ZN(n5903) );
  AND2_X1 U5633 ( .A1(n7379), .A2(n7441), .ZN(n7380) );
  INV_X1 U5634 ( .A(n7987), .ZN(n7984) );
  NAND3_X1 U5635 ( .A1(n4766), .A2(n4765), .A3(n10349), .ZN(n7352) );
  NOR2_X2 U5636 ( .A1(n7352), .A2(n7274), .ZN(n7379) );
  INV_X1 U5637 ( .A(n6052), .ZN(n5901) );
  AND4_X1 U5638 ( .A1(n6080), .A2(n6079), .A3(n6078), .A4(n6077), .ZN(n7346)
         );
  AND2_X1 U5639 ( .A1(n10349), .A2(n6963), .ZN(n7146) );
  NAND2_X1 U5640 ( .A1(n4766), .A2(n10349), .ZN(n7351) );
  AND2_X1 U5641 ( .A1(n4951), .A2(n7968), .ZN(n7140) );
  NAND2_X1 U5642 ( .A1(n4951), .A2(n4950), .ZN(n7139) );
  AND4_X1 U5643 ( .A1(n6069), .A2(n6068), .A3(n6067), .A4(n6066), .ZN(n7263)
         );
  OR2_X1 U5644 ( .A1(n6649), .A2(n8138), .ZN(n8515) );
  INV_X1 U5645 ( .A(n6332), .ZN(n10370) );
  INV_X1 U5646 ( .A(n8104), .ZN(n7953) );
  NOR2_X2 U5647 ( .A1(n6856), .A2(n5984), .ZN(n6855) );
  OR2_X1 U5648 ( .A1(n10462), .A2(n8350), .ZN(n6734) );
  NAND2_X1 U5649 ( .A1(n7888), .A2(n7887), .ZN(n8355) );
  NAND2_X1 U5650 ( .A1(n6264), .A2(n6263), .ZN(n8567) );
  NAND2_X1 U5651 ( .A1(n6255), .A2(n6254), .ZN(n8572) );
  INV_X1 U5652 ( .A(n6737), .ZN(n6750) );
  NAND2_X1 U5653 ( .A1(n5912), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4775) );
  AND2_X1 U5654 ( .A1(n5057), .A2(n6303), .ZN(n4806) );
  NAND2_X1 U5655 ( .A1(n4937), .A2(n4935), .ZN(n4934) );
  AND2_X1 U5656 ( .A1(n6306), .A2(n4936), .ZN(n4935) );
  INV_X1 U5657 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4936) );
  INV_X1 U5658 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6021) );
  NAND2_X1 U5659 ( .A1(n5381), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5406) );
  INV_X1 U5660 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U5661 ( .A1(n5794), .A2(n4992), .ZN(n4991) );
  OR2_X1 U5662 ( .A1(n7645), .A2(n7644), .ZN(n5005) );
  INV_X1 U5663 ( .A(n5738), .ZN(n5761) );
  OR2_X1 U5664 ( .A1(n5456), .A2(n5455), .ZN(n5483) );
  NAND2_X1 U5665 ( .A1(n6932), .A2(n5278), .ZN(n5284) );
  NAND2_X1 U5666 ( .A1(n6932), .A2(n5491), .ZN(n5287) );
  AND2_X1 U5667 ( .A1(n5699), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5718) );
  NAND2_X1 U5668 ( .A1(n4980), .A2(n4536), .ZN(n8764) );
  INV_X1 U5669 ( .A(n5007), .ZN(n5006) );
  OAI21_X1 U5670 ( .B1(n5008), .B2(n5475), .A(n7496), .ZN(n5007) );
  NAND2_X1 U5671 ( .A1(n5009), .A2(n7497), .ZN(n5008) );
  NAND2_X1 U5672 ( .A1(n5306), .A2(n6633), .ZN(n8787) );
  INV_X1 U5673 ( .A(n4968), .ZN(n8788) );
  NAND2_X1 U5674 ( .A1(n5793), .A2(n5792), .ZN(n4993) );
  NAND2_X1 U5675 ( .A1(n5589), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5607) );
  NAND2_X1 U5676 ( .A1(n4995), .A2(n4998), .ZN(n7809) );
  AOI21_X1 U5677 ( .B1(n5000), .B2(n4999), .A(n4544), .ZN(n4998) );
  INV_X1 U5678 ( .A(n4510), .ZN(n4999) );
  NAND2_X1 U5679 ( .A1(n5272), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5274) );
  NAND2_X1 U5680 ( .A1(n4580), .A2(n4579), .ZN(n10056) );
  INV_X1 U5681 ( .A(n6475), .ZN(n4579) );
  NOR2_X1 U5682 ( .A1(n9139), .A2(n4725), .ZN(n10067) );
  NOR2_X1 U5683 ( .A1(n6505), .A2(n7215), .ZN(n4725) );
  NAND2_X1 U5684 ( .A1(n10067), .A2(n4724), .ZN(n10066) );
  NAND2_X1 U5685 ( .A1(n10066), .A2(n4723), .ZN(n9154) );
  OR2_X1 U5686 ( .A1(n10069), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4723) );
  CLKBUF_X1 U5687 ( .A(n5414), .Z(n5415) );
  NAND2_X1 U5688 ( .A1(n10087), .A2(n6483), .ZN(n6485) );
  NOR2_X1 U5689 ( .A1(n6834), .A2(n4561), .ZN(n6838) );
  NOR2_X1 U5690 ( .A1(n6838), .A2(n6837), .ZN(n6872) );
  NOR2_X1 U5691 ( .A1(n6485), .A2(n6484), .ZN(n6829) );
  NOR2_X1 U5692 ( .A1(n6872), .A2(n4719), .ZN(n6874) );
  NOR2_X1 U5693 ( .A1(n4720), .A2(n7178), .ZN(n4719) );
  NAND2_X1 U5694 ( .A1(n6874), .A2(n6875), .ZN(n7062) );
  NAND2_X1 U5695 ( .A1(n10095), .A2(n10094), .ZN(n10099) );
  XNOR2_X1 U5696 ( .A(n4721), .B(n9179), .ZN(n7408) );
  NOR2_X1 U5697 ( .A1(n9170), .A2(n10113), .ZN(n10125) );
  XNOR2_X1 U5698 ( .A(n9188), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9191) );
  NAND2_X1 U5699 ( .A1(n8827), .A2(n8826), .ZN(n9197) );
  NAND2_X1 U5700 ( .A1(n9278), .A2(n9251), .ZN(n4734) );
  NAND2_X1 U5701 ( .A1(n9251), .A2(n9444), .ZN(n4739) );
  AND4_X1 U5702 ( .A1(n5231), .A2(n5230), .A3(n5229), .A4(n5228), .ZN(n9259)
         );
  NOR2_X1 U5703 ( .A1(n9273), .A2(n9274), .ZN(n9272) );
  AOI21_X1 U5704 ( .B1(n5034), .B2(n5036), .A(n4548), .ZN(n5033) );
  INV_X1 U5705 ( .A(n5036), .ZN(n5035) );
  AND2_X1 U5706 ( .A1(n9304), .A2(n9293), .ZN(n9289) );
  NAND2_X1 U5707 ( .A1(n5777), .A2(n5776), .ZN(n9305) );
  NOR2_X1 U5708 ( .A1(n9329), .A2(n9305), .ZN(n9304) );
  NAND2_X1 U5709 ( .A1(n5263), .A2(n5262), .ZN(n9330) );
  NOR2_X1 U5710 ( .A1(n9386), .A2(n4751), .ZN(n9355) );
  INV_X1 U5711 ( .A(n4753), .ZN(n4751) );
  AND2_X1 U5712 ( .A1(n7753), .A2(n4740), .ZN(n9396) );
  NOR2_X1 U5713 ( .A1(n4742), .A2(n8796), .ZN(n4740) );
  NAND2_X1 U5714 ( .A1(n5019), .A2(n5018), .ZN(n9395) );
  AOI21_X1 U5715 ( .B1(n5021), .B2(n5023), .A(n4545), .ZN(n5018) );
  OR2_X1 U5716 ( .A1(n5677), .A2(n5676), .ZN(n5679) );
  INV_X1 U5717 ( .A(n5024), .ZN(n5023) );
  INV_X1 U5718 ( .A(n5022), .ZN(n5021) );
  OAI21_X1 U5719 ( .B1(n4512), .B2(n5023), .A(n8856), .ZN(n5022) );
  AOI21_X1 U5720 ( .B1(n7780), .B2(n8993), .A(n7779), .ZN(n9420) );
  NAND2_X1 U5721 ( .A1(n7753), .A2(n4743), .ZN(n9414) );
  NOR2_X1 U5722 ( .A1(n7703), .A2(n7702), .ZN(n7745) );
  NOR2_X1 U5723 ( .A1(n8897), .A2(n9132), .ZN(n7702) );
  OR2_X1 U5724 ( .A1(n8986), .A2(n7707), .ZN(n8985) );
  OR2_X1 U5725 ( .A1(n5549), .A2(n5548), .ZN(n5571) );
  NOR2_X1 U5726 ( .A1(n5571), .A2(n7409), .ZN(n5589) );
  AOI21_X1 U5727 ( .B1(n7554), .B2(n8960), .A(n8890), .ZN(n10011) );
  NOR2_X1 U5728 ( .A1(n5508), .A2(n5507), .ZN(n5527) );
  NOR2_X1 U5729 ( .A1(n7176), .A2(n7503), .ZN(n7291) );
  AND2_X1 U5730 ( .A1(n8950), .A2(n8953), .ZN(n8848) );
  INV_X1 U5731 ( .A(n7239), .ZN(n4744) );
  OR2_X1 U5732 ( .A1(n7241), .A2(n7322), .ZN(n7176) );
  NAND2_X1 U5733 ( .A1(n4651), .A2(n4650), .ZN(n7024) );
  NAND2_X1 U5734 ( .A1(n10232), .A2(n4535), .ZN(n4651) );
  NOR2_X1 U5735 ( .A1(n10218), .A2(n4748), .ZN(n10191) );
  AND2_X1 U5736 ( .A1(n6927), .A2(n9437), .ZN(n7080) );
  NAND2_X1 U5737 ( .A1(n7017), .A2(n7016), .ZN(n4638) );
  OR2_X1 U5738 ( .A1(n6920), .A2(n10251), .ZN(n7016) );
  INV_X1 U5739 ( .A(n7080), .ZN(n6936) );
  NAND2_X1 U5740 ( .A1(n10251), .A2(n6615), .ZN(n7205) );
  NOR2_X1 U5741 ( .A1(n6932), .A2(n6615), .ZN(n7014) );
  INV_X1 U5742 ( .A(n9249), .ZN(n4675) );
  NAND2_X1 U5743 ( .A1(n4494), .A2(n9424), .ZN(n4816) );
  NOR2_X1 U5744 ( .A1(n9257), .A2(n9243), .ZN(n9245) );
  AND3_X1 U5745 ( .A1(n5420), .A2(n5419), .A3(n5418), .ZN(n10292) );
  XNOR2_X1 U5746 ( .A(n7884), .B(SI_30_), .ZN(n8825) );
  XNOR2_X1 U5747 ( .A(n7874), .B(n6279), .ZN(n8833) );
  NAND2_X1 U5748 ( .A1(n4853), .A2(n4854), .ZN(n7874) );
  OR2_X1 U5749 ( .A1(n5799), .A2(n4856), .ZN(n4853) );
  XNOR2_X1 U5750 ( .A(n5245), .B(n5244), .ZN(n7686) );
  NOR2_X1 U5751 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5187) );
  NAND2_X1 U5752 ( .A1(n4688), .A2(n5128), .ZN(n5583) );
  NAND2_X1 U5753 ( .A1(n4836), .A2(n4835), .ZN(n5499) );
  OR2_X1 U5754 ( .A1(n5108), .A2(n4839), .ZN(n4835) );
  XNOR2_X1 U5755 ( .A(n5476), .B(n5477), .ZN(n6552) );
  XNOR2_X1 U5756 ( .A(n4611), .B(n5466), .ZN(n6533) );
  OAI21_X1 U5757 ( .B1(n5438), .B2(n4864), .A(n5103), .ZN(n4611) );
  XNOR2_X1 U5758 ( .A(n5096), .B(SI_7_), .ZN(n5412) );
  INV_X1 U5759 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5192) );
  OAI21_X1 U5760 ( .B1(n8165), .B2(n8164), .A(n8163), .ZN(n8185) );
  AND4_X1 U5761 ( .A1(n6127), .A2(n6126), .A3(n6125), .A4(n6124), .ZN(n7543)
         );
  INV_X1 U5762 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9692) );
  AND2_X1 U5763 ( .A1(n7870), .A2(n6418), .ZN(n7048) );
  NAND2_X1 U5764 ( .A1(n4925), .A2(n6388), .ZN(n6795) );
  NAND2_X1 U5765 ( .A1(n4920), .A2(n4926), .ZN(n4925) );
  AND2_X1 U5766 ( .A1(n4927), .A2(n4499), .ZN(n7719) );
  NAND2_X1 U5767 ( .A1(n4890), .A2(n6772), .ZN(n6771) );
  NAND2_X1 U5768 ( .A1(n4592), .A2(n4599), .ZN(n7842) );
  NAND2_X1 U5769 ( .A1(n4927), .A2(n4601), .ZN(n4592) );
  AND4_X1 U5770 ( .A1(n6096), .A2(n6095), .A3(n6094), .A4(n6093), .ZN(n7364)
         );
  NAND2_X1 U5771 ( .A1(n6106), .A2(n6105), .ZN(n8003) );
  AND2_X1 U5772 ( .A1(n4930), .A2(n4932), .ZN(n7518) );
  NAND2_X1 U5773 ( .A1(n4686), .A2(n6174), .ZN(n7737) );
  NAND2_X1 U5774 ( .A1(n6885), .A2(n7885), .ZN(n4686) );
  XNOR2_X1 U5775 ( .A(n4687), .B(n7851), .ZN(n8213) );
  INV_X1 U5776 ( .A(n7852), .ZN(n7851) );
  NAND2_X1 U5777 ( .A1(n4917), .A2(n4915), .ZN(n6804) );
  INV_X1 U5778 ( .A(n4921), .ZN(n4917) );
  NAND2_X1 U5779 ( .A1(n4920), .A2(n4916), .ZN(n4915) );
  NOR2_X1 U5780 ( .A1(n4924), .A2(n6788), .ZN(n4916) );
  NAND2_X1 U5781 ( .A1(n7864), .A2(n6414), .ZN(n7870) );
  AND2_X1 U5782 ( .A1(n8227), .A2(n8544), .ZN(n8216) );
  AND2_X1 U5783 ( .A1(n4603), .A2(n4605), .ZN(n7774) );
  NAND2_X1 U5784 ( .A1(n4927), .A2(n4516), .ZN(n4603) );
  INV_X1 U5785 ( .A(n8216), .ZN(n7827) );
  NAND2_X1 U5786 ( .A1(n7336), .A2(n6434), .ZN(n6440) );
  OAI21_X1 U5787 ( .B1(n7864), .B2(n4911), .A(n4908), .ZN(n6428) );
  OAI21_X1 U5788 ( .B1(n8134), .B2(n8133), .A(n4863), .ZN(n4862) );
  NAND2_X1 U5789 ( .A1(n8136), .A2(n8135), .ZN(n4863) );
  AND2_X1 U5790 ( .A1(n6253), .A2(n6252), .ZN(n8204) );
  INV_X1 U5791 ( .A(n8499), .ZN(n8246) );
  OR2_X1 U5792 ( .A1(n6650), .A2(n10425), .ZN(n8245) );
  NOR2_X1 U5793 ( .A1(n9989), .A2(n4514), .ZN(n6717) );
  NOR2_X1 U5794 ( .A1(n6704), .A2(n6703), .ZN(n6702) );
  AND2_X1 U5795 ( .A1(n4715), .A2(n4714), .ZN(n6704) );
  NAND2_X1 U5796 ( .A1(n6720), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4714) );
  INV_X1 U5797 ( .A(n4707), .ZN(n6727) );
  INV_X1 U5798 ( .A(n4705), .ZN(n6691) );
  AND2_X1 U5799 ( .A1(n4705), .A2(n4704), .ZN(n6689) );
  INV_X1 U5800 ( .A(n6690), .ZN(n4704) );
  AND2_X1 U5801 ( .A1(n6032), .A2(n6005), .ZN(n6694) );
  NOR2_X1 U5802 ( .A1(n6689), .A2(n4703), .ZN(n6656) );
  AND2_X1 U5803 ( .A1(n6694), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4703) );
  OR2_X1 U5804 ( .A1(n6764), .A2(n6765), .ZN(n6979) );
  INV_X1 U5805 ( .A(n4702), .ZN(n7184) );
  NAND2_X1 U5806 ( .A1(n7185), .A2(n7186), .ZN(n7306) );
  AND2_X1 U5807 ( .A1(n4702), .A2(n4701), .ZN(n7185) );
  NAND2_X1 U5808 ( .A1(n7188), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4701) );
  OR2_X1 U5809 ( .A1(n7309), .A2(n7308), .ZN(n7449) );
  NAND2_X1 U5810 ( .A1(n7451), .A2(n7452), .ZN(n7574) );
  AND2_X1 U5811 ( .A1(n7449), .A2(n4718), .ZN(n7451) );
  NAND2_X1 U5812 ( .A1(n7450), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4718) );
  INV_X1 U5813 ( .A(n4710), .ZN(n8310) );
  OAI22_X1 U5814 ( .A1(n4709), .A2(n4708), .B1(n4503), .B2(n8312), .ZN(n8323)
         );
  INV_X1 U5815 ( .A(n8298), .ZN(n4709) );
  NAND2_X1 U5816 ( .A1(n4711), .A2(n4713), .ZN(n4708) );
  INV_X1 U5817 ( .A(n8567), .ZN(n8367) );
  OAI21_X1 U5818 ( .B1(n8426), .B2(n4796), .A(n4794), .ZN(n8395) );
  OR2_X1 U5819 ( .A1(n8404), .A2(n8403), .ZN(n8405) );
  INV_X1 U5820 ( .A(n6359), .ZN(n8412) );
  NOR2_X1 U5821 ( .A1(n8425), .A2(n4800), .ZN(n8411) );
  AND2_X1 U5822 ( .A1(n8439), .A2(n8438), .ZN(n8590) );
  NAND2_X1 U5823 ( .A1(n8443), .A2(n6345), .ZN(n8445) );
  NAND2_X1 U5824 ( .A1(n8501), .A2(n8048), .ZN(n8484) );
  NAND2_X1 U5825 ( .A1(n4780), .A2(n4781), .ZN(n8476) );
  OR2_X1 U5826 ( .A1(n8506), .A2(n4783), .ZN(n4780) );
  AND2_X1 U5827 ( .A1(n4784), .A2(n4508), .ZN(n8491) );
  OR2_X1 U5828 ( .A1(n8506), .A2(n4787), .ZN(n4784) );
  AND2_X1 U5829 ( .A1(n8547), .A2(n8546), .ZN(n8621) );
  AND2_X1 U5830 ( .A1(n4809), .A2(n4550), .ZN(n7734) );
  NAND2_X1 U5831 ( .A1(n6166), .A2(n6165), .ZN(n7683) );
  NAND2_X1 U5832 ( .A1(n7538), .A2(n7927), .ZN(n7523) );
  NAND2_X1 U5833 ( .A1(n7418), .A2(n6128), .ZN(n7532) );
  NAND2_X1 U5834 ( .A1(n7137), .A2(n6059), .ZN(n7344) );
  INV_X1 U5835 ( .A(n10437), .ZN(n10363) );
  INV_X1 U5836 ( .A(n8537), .ZN(n10381) );
  AND2_X1 U5837 ( .A1(n10383), .A2(n10360), .ZN(n8551) );
  NAND2_X1 U5838 ( .A1(n8565), .A2(n4528), .ZN(n8654) );
  INV_X1 U5839 ( .A(n7737), .ZN(n6180) );
  INV_X1 U5840 ( .A(n10469), .ZN(n10468) );
  NAND2_X1 U5841 ( .A1(n4776), .A2(n5918), .ZN(n5919) );
  NAND2_X1 U5842 ( .A1(n5913), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5918) );
  NAND2_X1 U5843 ( .A1(n4777), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n4776) );
  NAND2_X1 U5844 ( .A1(n5894), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5895) );
  XNOR2_X1 U5845 ( .A(n6310), .B(n6309), .ZN(n7551) );
  INV_X1 U5846 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6557) );
  INV_X1 U5847 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6554) );
  INV_X1 U5848 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6536) );
  INV_X1 U5849 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6513) );
  INV_X1 U5850 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6499) );
  NAND2_X1 U5851 ( .A1(n5945), .A2(n5944), .ZN(n9981) );
  NAND2_X1 U5852 ( .A1(n8813), .A2(n4991), .ZN(n8704) );
  NAND2_X1 U5853 ( .A1(n5206), .A2(n5205), .ZN(n9450) );
  NAND2_X1 U5854 ( .A1(n5003), .A2(n5005), .ZN(n7692) );
  NAND2_X1 U5855 ( .A1(n7634), .A2(n4510), .ZN(n5003) );
  NOR2_X1 U5856 ( .A1(n4978), .A2(n5769), .ZN(n8711) );
  NAND2_X1 U5857 ( .A1(n5758), .A2(n5757), .ZN(n9469) );
  NAND2_X1 U5858 ( .A1(n7317), .A2(n5475), .ZN(n7499) );
  NAND2_X1 U5859 ( .A1(n5324), .A2(n4968), .ZN(n4966) );
  NAND2_X1 U5860 ( .A1(n5656), .A2(n5655), .ZN(n9491) );
  NAND2_X1 U5861 ( .A1(n4983), .A2(n4986), .ZN(n5879) );
  AND2_X1 U5862 ( .A1(n4990), .A2(n4987), .ZN(n4986) );
  OR2_X1 U5863 ( .A1(n8702), .A2(n5845), .ZN(n4990) );
  NAND2_X1 U5864 ( .A1(n8763), .A2(n8767), .ZN(n8732) );
  INV_X1 U5865 ( .A(n9362), .ZN(n8836) );
  NAND2_X1 U5866 ( .A1(n4971), .A2(n4975), .ZN(n8754) );
  NAND2_X1 U5867 ( .A1(n4978), .A2(n4976), .ZN(n4971) );
  NAND2_X1 U5868 ( .A1(n5011), .A2(n5010), .ZN(n7317) );
  INV_X1 U5869 ( .A(n7314), .ZN(n5010) );
  INV_X1 U5870 ( .A(n7315), .ZN(n5011) );
  NAND2_X1 U5871 ( .A1(n5698), .A2(n5697), .ZN(n9486) );
  NAND2_X1 U5872 ( .A1(n7634), .A2(n5541), .ZN(n7647) );
  NAND2_X1 U5873 ( .A1(n5547), .A2(n5546), .ZN(n9516) );
  OR2_X1 U5874 ( .A1(n5843), .A2(n5842), .ZN(n8773) );
  AND2_X1 U5875 ( .A1(n8795), .A2(n9524), .ZN(n8791) );
  XNOR2_X1 U5876 ( .A(n5235), .B(P1_IR_REG_22__SCAN_IN), .ZN(n9125) );
  OR2_X1 U5877 ( .A1(n6526), .A2(n7204), .ZN(n5308) );
  AND2_X1 U5878 ( .A1(n10042), .A2(n6465), .ZN(n10043) );
  NAND2_X1 U5879 ( .A1(n4578), .A2(n4577), .ZN(n9146) );
  INV_X1 U5880 ( .A(n9144), .ZN(n4577) );
  NAND2_X1 U5881 ( .A1(n10056), .A2(n9145), .ZN(n4578) );
  AND2_X1 U5882 ( .A1(n6478), .A2(n6477), .ZN(n9160) );
  INV_X1 U5883 ( .A(n4582), .ZN(n6577) );
  OR2_X1 U5884 ( .A1(n6582), .A2(n6466), .ZN(n6583) );
  NOR2_X1 U5885 ( .A1(n6564), .A2(n6482), .ZN(n10089) );
  NAND2_X1 U5886 ( .A1(n10089), .A2(n10088), .ZN(n10087) );
  NAND2_X1 U5887 ( .A1(n9182), .A2(n10118), .ZN(n10132) );
  OR2_X1 U5888 ( .A1(n10159), .A2(n10141), .ZN(n10143) );
  NAND2_X1 U5889 ( .A1(n10146), .A2(n4570), .ZN(n10166) );
  OR2_X1 U5890 ( .A1(n10159), .A2(n10158), .ZN(n10161) );
  AOI21_X1 U5891 ( .B1(n8682), .B2(n8866), .A(n8865), .ZN(n9431) );
  INV_X1 U5892 ( .A(n9197), .ZN(n9436) );
  NAND2_X1 U5893 ( .A1(n5038), .A2(n9219), .ZN(n9288) );
  NAND2_X1 U5894 ( .A1(n9217), .A2(n5039), .ZN(n5038) );
  NAND2_X1 U5895 ( .A1(n5043), .A2(n9211), .ZN(n9339) );
  AND2_X1 U5896 ( .A1(n5736), .A2(n5735), .ZN(n9358) );
  NAND2_X1 U5897 ( .A1(n9210), .A2(n9209), .ZN(n9354) );
  NAND2_X1 U5898 ( .A1(n5717), .A2(n5716), .ZN(n9481) );
  AOI21_X1 U5899 ( .B1(n4665), .B2(n4663), .A(n4659), .ZN(n9382) );
  NOR2_X1 U5900 ( .A1(n4819), .A2(n4664), .ZN(n4663) );
  NAND2_X1 U5901 ( .A1(n4822), .A2(n4820), .ZN(n9408) );
  NAND2_X1 U5902 ( .A1(n5020), .A2(n5024), .ZN(n7789) );
  NAND2_X1 U5903 ( .A1(n7787), .A2(n4512), .ZN(n5020) );
  OAI21_X1 U5904 ( .B1(n7787), .B2(n5023), .A(n5021), .ZN(n9494) );
  INV_X1 U5905 ( .A(n7786), .ZN(n5025) );
  NAND2_X1 U5906 ( .A1(n7787), .A2(n8988), .ZN(n5026) );
  INV_X1 U5907 ( .A(n10187), .ZN(n10239) );
  NAND2_X1 U5908 ( .A1(n5525), .A2(n5524), .ZN(n10020) );
  AND2_X1 U5909 ( .A1(n5051), .A2(n5049), .ZN(n10009) );
  NAND2_X1 U5910 ( .A1(n5051), .A2(n7560), .ZN(n10010) );
  NAND2_X1 U5911 ( .A1(n7559), .A2(n5068), .ZN(n5051) );
  INV_X1 U5912 ( .A(n10002), .ZN(n7503) );
  NAND2_X1 U5913 ( .A1(n5031), .A2(n5030), .ZN(n10173) );
  NAND2_X1 U5914 ( .A1(n5032), .A2(n7041), .ZN(n5031) );
  OR2_X1 U5915 ( .A1(n6502), .A2(n5439), .ZN(n4669) );
  NAND2_X1 U5916 ( .A1(n7032), .A2(n7031), .ZN(n7202) );
  INV_X1 U5917 ( .A(n10251), .ZN(n7030) );
  AND2_X1 U5918 ( .A1(n9403), .A2(n10201), .ZN(n10187) );
  AND2_X1 U5919 ( .A1(n9406), .A2(n10198), .ZN(n10221) );
  NAND2_X1 U5920 ( .A1(n5218), .A2(n5220), .ZN(n9555) );
  NAND2_X1 U5921 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n5017) );
  OAI21_X1 U5922 ( .B1(n5016), .B2(n9552), .A(n5015), .ZN(n5014) );
  NAND2_X1 U5923 ( .A1(n4653), .A2(n5196), .ZN(n5013) );
  XNOR2_X1 U5924 ( .A(n6276), .B(n6275), .ZN(n8149) );
  NAND2_X1 U5925 ( .A1(n5799), .A2(n5798), .ZN(n6276) );
  NAND2_X1 U5926 ( .A1(n5200), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5201) );
  NAND2_X1 U5927 ( .A1(n5196), .A2(n5055), .ZN(n5200) );
  XNOR2_X1 U5928 ( .A(n5756), .B(n5755), .ZN(n7435) );
  INV_X1 U5929 ( .A(n6927), .ZN(n9076) );
  INV_X1 U5930 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9703) );
  INV_X1 U5931 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9738) );
  INV_X1 U5932 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9728) );
  INV_X1 U5933 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9934) );
  INV_X1 U5934 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9680) );
  INV_X1 U5935 ( .A(n4864), .ZN(n5437) );
  INV_X1 U5936 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6522) );
  INV_X1 U5937 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6511) );
  NAND2_X1 U5938 ( .A1(n4589), .A2(n5092), .ZN(n5370) );
  NAND2_X1 U5939 ( .A1(n5390), .A2(n5389), .ZN(n4589) );
  OR2_X1 U5940 ( .A1(n5371), .A2(n5464), .ZN(n5372) );
  XNOR2_X1 U5941 ( .A(n5390), .B(n5389), .ZN(n6502) );
  INV_X1 U5942 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6496) );
  OAI21_X1 U5943 ( .B1(n5083), .B2(n4642), .A(n4640), .ZN(n5351) );
  AOI21_X1 U5944 ( .B1(n4645), .B2(n5330), .A(n4505), .ZN(n4640) );
  NAND2_X1 U5945 ( .A1(n5083), .A2(n5082), .ZN(n5331) );
  NAND2_X1 U5946 ( .A1(n4583), .A2(n4646), .ZN(n6602) );
  INV_X1 U5947 ( .A(n4584), .ZN(n4583) );
  OAI21_X1 U5948 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(P1_IR_REG_1__SCAN_IN), .A(
        n4585), .ZN(n4584) );
  NOR2_X1 U5949 ( .A1(n9588), .A2(n10506), .ZN(n10505) );
  AOI21_X1 U5950 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10503), .ZN(n10502) );
  NOR2_X1 U5951 ( .A1(n10502), .A2(n10501), .ZN(n10500) );
  AND2_X1 U5952 ( .A1(n8198), .A2(n8199), .ZN(n4905) );
  NAND2_X1 U5953 ( .A1(n4927), .A2(n4928), .ZN(n7832) );
  NAND2_X1 U5954 ( .A1(n4697), .A2(n4695), .ZN(P2_U3242) );
  NOR2_X1 U5955 ( .A1(n7856), .A2(n4696), .ZN(n4695) );
  AND2_X1 U5956 ( .A1(n8397), .A2(n8230), .ZN(n4696) );
  NOR2_X1 U5957 ( .A1(n6368), .A2(n6367), .ZN(n6369) );
  NAND2_X1 U5958 ( .A1(n10469), .A2(n10360), .ZN(n4758) );
  NOR2_X1 U5959 ( .A1(n4759), .A2(n4567), .ZN(n4756) );
  NAND2_X1 U5960 ( .A1(n4729), .A2(n4726), .ZN(P1_U3260) );
  AOI21_X1 U5961 ( .B1(n4732), .B2(n10206), .A(n4730), .ZN(n4729) );
  NAND2_X1 U5962 ( .A1(n4731), .A2(n9165), .ZN(n4730) );
  OR2_X1 U5963 ( .A1(n10326), .A2(n4671), .ZN(n4670) );
  NAND2_X1 U5964 ( .A1(n9532), .A2(n10326), .ZN(n4672) );
  INV_X1 U5965 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n4671) );
  OR2_X1 U5966 ( .A1(n10315), .A2(n5854), .ZN(n4813) );
  NAND2_X1 U5967 ( .A1(n9532), .A2(n10315), .ZN(n4814) );
  AND2_X1 U5968 ( .A1(n8367), .A2(n8243), .ZN(n4491) );
  INV_X1 U5969 ( .A(n10462), .ZN(n10360) );
  AND2_X1 U5970 ( .A1(n8120), .A2(n4550), .ZN(n4493) );
  AND2_X1 U5971 ( .A1(n5937), .A2(n5936), .ZN(n8498) );
  XOR2_X1 U5972 ( .A(n9245), .B(n9244), .Z(n4494) );
  NAND2_X1 U5973 ( .A1(n4955), .A2(n6344), .ZN(n8443) );
  AND2_X1 U5974 ( .A1(n9043), .A2(n9044), .ZN(n9222) );
  AND2_X1 U5975 ( .A1(n4781), .A2(n4529), .ZN(n4495) );
  AND2_X1 U5976 ( .A1(n4843), .A2(n5714), .ZN(n4496) );
  NAND2_X1 U5977 ( .A1(n8010), .A2(n7927), .ZN(n8014) );
  AND2_X1 U5978 ( .A1(n8562), .A2(n8372), .ZN(n8082) );
  INV_X1 U5979 ( .A(n8082), .ZN(n4965) );
  NAND2_X1 U5980 ( .A1(n8071), .A2(n8069), .ZN(n8394) );
  INV_X1 U5981 ( .A(n8394), .ZN(n4791) );
  INV_X1 U5982 ( .A(n8897), .ZN(n10029) );
  NAND2_X1 U5983 ( .A1(n5569), .A2(n5568), .ZN(n8897) );
  NAND2_X1 U5984 ( .A1(n5898), .A2(n5897), .ZN(n8587) );
  AND2_X1 U5985 ( .A1(n8030), .A2(n8029), .ZN(n7727) );
  INV_X1 U5986 ( .A(n7727), .ZN(n8120) );
  AND2_X1 U5987 ( .A1(n4739), .A2(n10198), .ZN(n4497) );
  INV_X1 U5988 ( .A(n4742), .ZN(n4741) );
  NAND2_X1 U5989 ( .A1(n4743), .A2(n9418), .ZN(n4742) );
  NAND2_X1 U5990 ( .A1(n6344), .A2(n8060), .ZN(n4498) );
  AND2_X1 U5991 ( .A1(n4928), .A2(n4533), .ZN(n4499) );
  INV_X1 U5992 ( .A(n9220), .ZN(n9317) );
  AND2_X1 U5993 ( .A1(n8133), .A2(n6375), .ZN(n4500) );
  AND2_X1 U5994 ( .A1(n8940), .A2(n8936), .ZN(n4501) );
  AND2_X1 U5995 ( .A1(n4948), .A2(n4558), .ZN(n4502) );
  INV_X1 U5996 ( .A(n7717), .ZN(n4605) );
  INV_X1 U5997 ( .A(n6788), .ZN(n4926) );
  NAND2_X1 U5998 ( .A1(n8313), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4503) );
  OR2_X1 U5999 ( .A1(n6158), .A2(n4934), .ZN(n4504) );
  AND2_X1 U6000 ( .A1(n5085), .A2(SI_3_), .ZN(n4505) );
  AND2_X1 U6001 ( .A1(n6336), .A2(n7993), .ZN(n4506) );
  XOR2_X1 U6002 ( .A(n8593), .B(n7853), .Z(n4507) );
  OAI211_X1 U6003 ( .C1(n5478), .C2(n6503), .A(n5391), .B(n4669), .ZN(n10200)
         );
  INV_X1 U6004 ( .A(n10200), .ZN(n10278) );
  NAND2_X1 U6005 ( .A1(n8521), .A2(n8545), .ZN(n4508) );
  NAND2_X1 U6006 ( .A1(n10444), .A2(n7966), .ZN(n4509) );
  NOR2_X1 U6007 ( .A1(n5559), .A2(n5004), .ZN(n4510) );
  OR2_X1 U6008 ( .A1(n9510), .A2(n7815), .ZN(n4511) );
  AND2_X1 U6009 ( .A1(n5027), .A2(n8988), .ZN(n4512) );
  AND2_X1 U6010 ( .A1(n4687), .A2(n7852), .ZN(n4513) );
  AND2_X1 U6011 ( .A1(n5943), .A2(n5883), .ZN(n5995) );
  INV_X1 U6012 ( .A(n9237), .ZN(n9323) );
  OR2_X1 U6013 ( .A1(n9469), .A2(n8836), .ZN(n9237) );
  XNOR2_X1 U6014 ( .A(n8567), .B(n8187), .ZN(n8369) );
  INV_X1 U6015 ( .A(n8369), .ZN(n4964) );
  AND2_X1 U6016 ( .A1(n9993), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4514) );
  NAND2_X1 U6017 ( .A1(n10224), .A2(n10200), .ZN(n4515) );
  AND2_X1 U6018 ( .A1(n4499), .A2(n7718), .ZN(n4516) );
  OR4_X2 U6019 ( .A1(n8016), .A2(n8015), .A3(n8014), .A4(n8093), .ZN(n4517) );
  AND2_X1 U6020 ( .A1(n5069), .A2(n4981), .ZN(n4518) );
  NAND2_X1 U6021 ( .A1(n5801), .A2(n5800), .ZN(n9444) );
  INV_X1 U6022 ( .A(n9444), .ZN(n4738) );
  AND2_X1 U6023 ( .A1(n6398), .A2(n6403), .ZN(n4519) );
  NAND2_X1 U6024 ( .A1(n5637), .A2(n5636), .ZN(n9500) );
  NOR2_X1 U6025 ( .A1(n8368), .A2(n4491), .ZN(n4520) );
  AND2_X1 U6026 ( .A1(n4978), .A2(n5769), .ZN(n4521) );
  OR3_X1 U6027 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4522) );
  NOR2_X1 U6028 ( .A1(n10012), .A2(n5050), .ZN(n5049) );
  NOR2_X1 U6029 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n6044) );
  AND4_X1 U6030 ( .A1(n6044), .A2(n5882), .A3(n5881), .A4(n5880), .ZN(n4523)
         );
  AND2_X1 U6031 ( .A1(n9500), .A2(n9130), .ZN(n4524) );
  AND2_X1 U6032 ( .A1(n8002), .A2(n8001), .ZN(n4525) );
  NAND2_X1 U6033 ( .A1(n9242), .A2(n9048), .ZN(n9267) );
  NOR2_X1 U6034 ( .A1(n9272), .A2(n9241), .ZN(n4526) );
  INV_X1 U6035 ( .A(n8603), .ZN(n8482) );
  NAND2_X1 U6036 ( .A1(n6201), .A2(n6200), .ZN(n8603) );
  AND2_X1 U6037 ( .A1(n8507), .A2(n8041), .ZN(n8540) );
  INV_X1 U6038 ( .A(n8540), .ZN(n4944) );
  NOR2_X1 U6039 ( .A1(n9212), .A2(n5044), .ZN(n4527) );
  AND2_X1 U6040 ( .A1(n4614), .A2(n8564), .ZN(n4528) );
  OR2_X1 U6041 ( .A1(n8482), .A2(n8499), .ZN(n4529) );
  INV_X1 U6042 ( .A(n7804), .ZN(n9510) );
  NAND2_X1 U6043 ( .A1(n5587), .A2(n5586), .ZN(n7804) );
  NAND2_X1 U6044 ( .A1(n8835), .A2(n8834), .ZN(n9251) );
  OR2_X1 U6045 ( .A1(n8023), .A2(n8022), .ZN(n4530) );
  XNOR2_X1 U6046 ( .A(n5113), .B(SI_11_), .ZN(n5498) );
  AND2_X1 U6047 ( .A1(n4834), .A2(n4619), .ZN(n4531) );
  AND2_X1 U6048 ( .A1(n4822), .A2(n4821), .ZN(n4532) );
  NAND2_X1 U6049 ( .A1(n7661), .A2(n7660), .ZN(n4533) );
  AND2_X1 U6050 ( .A1(n8907), .A2(n9083), .ZN(n4534) );
  AND2_X1 U6051 ( .A1(n4649), .A2(n7022), .ZN(n4535) );
  AND2_X1 U6052 ( .A1(n4979), .A2(n5694), .ZN(n4536) );
  AND2_X1 U6053 ( .A1(n6180), .A2(n7828), .ZN(n4537) );
  NOR2_X1 U6054 ( .A1(n10204), .A2(n10188), .ZN(n4538) );
  OR2_X1 U6055 ( .A1(n8165), .A2(n4895), .ZN(n4539) );
  NOR2_X1 U6056 ( .A1(n9278), .A2(n9444), .ZN(n4540) );
  INV_X1 U6057 ( .A(n5001), .ZN(n5000) );
  OR2_X1 U6058 ( .A1(n5623), .A2(n5002), .ZN(n5001) );
  INV_X1 U6059 ( .A(n4735), .ZN(n9250) );
  NAND2_X1 U6060 ( .A1(n8660), .A2(n8204), .ZN(n4541) );
  NOR2_X1 U6061 ( .A1(n8603), .A2(n8246), .ZN(n4542) );
  NAND2_X1 U6062 ( .A1(n8073), .A2(n8072), .ZN(n8386) );
  INV_X1 U6063 ( .A(n8386), .ZN(n4636) );
  AND2_X1 U6064 ( .A1(n8402), .A2(n8067), .ZN(n8098) );
  INV_X1 U6065 ( .A(n8098), .ZN(n4798) );
  AND2_X1 U6066 ( .A1(n9392), .A2(n9206), .ZN(n9231) );
  INV_X1 U6067 ( .A(n9231), .ZN(n4662) );
  INV_X1 U6068 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5917) );
  AND2_X1 U6069 ( .A1(n5114), .A2(SI_11_), .ZN(n4543) );
  NAND2_X1 U6070 ( .A1(n5622), .A2(n5621), .ZN(n4544) );
  INV_X1 U6071 ( .A(n9454), .ZN(n9293) );
  NAND2_X1 U6072 ( .A1(n5247), .A2(n5246), .ZN(n9454) );
  NOR2_X1 U6073 ( .A1(n9201), .A2(n9411), .ZN(n4545) );
  AND2_X1 U6074 ( .A1(n5207), .A2(n5232), .ZN(n4546) );
  NOR2_X1 U6075 ( .A1(n8495), .A2(n8516), .ZN(n4547) );
  AND2_X1 U6076 ( .A1(n9454), .A2(n9220), .ZN(n4548) );
  INV_X1 U6077 ( .A(n8117), .ZN(n8017) );
  AND2_X1 U6078 ( .A1(n8019), .A2(n8018), .ZN(n8117) );
  OR2_X1 U6079 ( .A1(n4524), .A2(n7786), .ZN(n4549) );
  NAND2_X1 U6080 ( .A1(n6193), .A2(n6192), .ZN(n8608) );
  OR2_X1 U6081 ( .A1(n7737), .A2(n7828), .ZN(n8030) );
  NAND2_X1 U6082 ( .A1(n7683), .A2(n8248), .ZN(n4550) );
  OR2_X1 U6083 ( .A1(n8638), .A2(n7672), .ZN(n8019) );
  AND2_X1 U6084 ( .A1(n9552), .A2(n5220), .ZN(n4551) );
  OR2_X1 U6085 ( .A1(n8562), .A2(n8372), .ZN(n8081) );
  INV_X1 U6086 ( .A(n8081), .ZN(n4962) );
  OR2_X1 U6087 ( .A1(n9134), .A2(n10002), .ZN(n8950) );
  INV_X1 U6088 ( .A(n8950), .ZN(n4639) );
  OR2_X1 U6089 ( .A1(n8608), .A2(n8516), .ZN(n8048) );
  INV_X1 U6090 ( .A(n8048), .ZN(n4945) );
  OR2_X1 U6091 ( .A1(n6158), .A2(n4933), .ZN(n4552) );
  AND3_X1 U6092 ( .A1(n5446), .A2(n5445), .A3(n5444), .ZN(n7128) );
  NOR2_X1 U6093 ( .A1(n8483), .A2(n4945), .ZN(n4553) );
  OR2_X1 U6094 ( .A1(n4738), .A2(n9275), .ZN(n4554) );
  OR2_X1 U6095 ( .A1(n8643), .A2(n7591), .ZN(n7927) );
  OR2_X1 U6096 ( .A1(n9507), .A2(n7747), .ZN(n8992) );
  INV_X1 U6097 ( .A(n4975), .ZN(n4974) );
  NAND2_X1 U6098 ( .A1(n5769), .A2(n4977), .ZN(n4975) );
  AND2_X1 U6099 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4555) );
  AND2_X1 U6100 ( .A1(n8117), .A2(n4888), .ZN(n4556) );
  AND2_X1 U6101 ( .A1(n5913), .A2(n5893), .ZN(n4557) );
  AND2_X1 U6102 ( .A1(n7988), .A2(n7981), .ZN(n8110) );
  OR2_X1 U6103 ( .A1(n8572), .A2(n8371), .ZN(n8073) );
  NAND2_X1 U6104 ( .A1(n7975), .A2(n7858), .ZN(n4558) );
  OAI21_X1 U6105 ( .B1(n8554), .B2(n4758), .A(n4756), .ZN(P2_U3519) );
  INV_X1 U6106 ( .A(n6873), .ZN(n4720) );
  NAND2_X1 U6107 ( .A1(n7586), .A2(n7515), .ZN(n4930) );
  INV_X1 U6108 ( .A(n9132), .ZN(n8976) );
  AND2_X1 U6109 ( .A1(n7753), .A2(n4741), .ZN(n4559) );
  NOR2_X1 U6110 ( .A1(n9469), .A2(n9362), .ZN(n4560) );
  INV_X1 U6111 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4610) );
  AND2_X1 U6112 ( .A1(n4621), .A2(n4625), .ZN(n7671) );
  AND2_X1 U6113 ( .A1(n6835), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4561) );
  INV_X1 U6114 ( .A(n8993), .ZN(n4826) );
  NAND2_X1 U6115 ( .A1(n4809), .A2(n4493), .ZN(n7733) );
  NOR3_X1 U6116 ( .A1(n9386), .A2(n9330), .A3(n4752), .ZN(n4749) );
  AND4_X1 U6117 ( .A1(n6115), .A2(n6114), .A3(n6113), .A4(n6112), .ZN(n8004)
         );
  INV_X1 U6118 ( .A(n8004), .ZN(n4870) );
  AND2_X1 U6119 ( .A1(n4710), .A2(n4503), .ZN(n4562) );
  NAND2_X1 U6120 ( .A1(n8531), .A2(n4772), .ZN(n4774) );
  INV_X1 U6121 ( .A(n4754), .ZN(n9372) );
  NOR2_X1 U6122 ( .A1(n9386), .A2(n9481), .ZN(n4754) );
  NAND2_X1 U6123 ( .A1(n5675), .A2(n5674), .ZN(n8796) );
  INV_X1 U6124 ( .A(n4750), .ZN(n9340) );
  NOR2_X1 U6125 ( .A1(n9386), .A2(n4752), .ZN(n4750) );
  AND2_X1 U6126 ( .A1(n5157), .A2(SI_21_), .ZN(n4563) );
  AND2_X1 U6127 ( .A1(n5026), .A2(n5025), .ZN(n4564) );
  AND2_X1 U6128 ( .A1(n6358), .A2(n6357), .ZN(n4565) );
  OR2_X1 U6129 ( .A1(n6158), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n4566) );
  NAND2_X1 U6130 ( .A1(n6450), .A2(n6439), .ZN(n8211) );
  NAND2_X1 U6131 ( .A1(n6428), .A2(n7152), .ZN(n7155) );
  NAND2_X1 U6132 ( .A1(n7870), .A2(n4913), .ZN(n7047) );
  NAND2_X1 U6133 ( .A1(n4806), .A2(n4941), .ZN(n6299) );
  AND2_X1 U6134 ( .A1(n10469), .A2(n4757), .ZN(n4567) );
  NAND2_X1 U6135 ( .A1(n10232), .A2(n10227), .ZN(n10207) );
  INV_X1 U6136 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4939) );
  NAND2_X1 U6137 ( .A1(n6135), .A2(n6134), .ZN(n8643) );
  INV_X1 U6138 ( .A(n8643), .ZN(n4763) );
  NAND2_X1 U6139 ( .A1(n7137), .A2(n4802), .ZN(n7342) );
  NAND2_X1 U6140 ( .A1(n5054), .A2(n7164), .ZN(n7166) );
  AND2_X1 U6141 ( .A1(n9179), .A2(n5570), .ZN(n4568) );
  NOR2_X1 U6142 ( .A1(n6819), .A2(n8101), .ZN(n4569) );
  NAND2_X1 U6143 ( .A1(n4941), .A2(n5057), .ZN(n6302) );
  INV_X1 U6144 ( .A(n4764), .ZN(n7535) );
  OR2_X1 U6145 ( .A1(n10144), .A2(n9185), .ZN(n4570) );
  AND2_X1 U6146 ( .A1(n6278), .A2(n9681), .ZN(n4571) );
  AND2_X1 U6147 ( .A1(n7872), .A2(SI_29_), .ZN(n4572) );
  AND2_X1 U6148 ( .A1(n5031), .A2(n4515), .ZN(n4573) );
  INV_X1 U6149 ( .A(n7356), .ZN(n4765) );
  OR2_X1 U6150 ( .A1(n6614), .A2(n6926), .ZN(n10306) );
  INV_X1 U6151 ( .A(n10306), .ZN(n10198) );
  XNOR2_X1 U6152 ( .A(n5201), .B(n9885), .ZN(n5850) );
  INV_X1 U6153 ( .A(n10227), .ZN(n4652) );
  NAND4_X1 U6154 ( .A1(n5979), .A2(n5978), .A3(n5977), .A4(n5976), .ZN(n8260)
         );
  INV_X1 U6155 ( .A(n8260), .ZN(n5985) );
  OR2_X1 U6156 ( .A1(n10217), .A2(n7038), .ZN(n10218) );
  INV_X1 U6157 ( .A(n10218), .ZN(n4747) );
  OR2_X1 U6158 ( .A1(n9184), .A2(n9183), .ZN(n4574) );
  INV_X1 U6159 ( .A(n10367), .ZN(n8350) );
  INV_X1 U6160 ( .A(n10055), .ZN(n4580) );
  INV_X1 U6161 ( .A(n10065), .ZN(n4724) );
  NAND2_X1 U6162 ( .A1(n10431), .A2(n8128), .ZN(n8097) );
  NAND2_X1 U6163 ( .A1(n4727), .A2(n9332), .ZN(n4726) );
  AND2_X1 U6164 ( .A1(n9403), .A2(n9332), .ZN(n9406) );
  OR2_X1 U6165 ( .A1(n10306), .A2(n9332), .ZN(n6918) );
  NAND2_X1 U6166 ( .A1(n7163), .A2(n7162), .ZN(n5054) );
  NAND2_X1 U6167 ( .A1(n7200), .A2(n7034), .ZN(n7214) );
  AOI21_X2 U6168 ( .B1(n9223), .B2(n9274), .A(n5060), .ZN(n9268) );
  NAND2_X1 U6169 ( .A1(n4672), .A2(n4670), .ZN(P1_U3552) );
  NAND2_X2 U6170 ( .A1(n7705), .A2(n4511), .ZN(n7787) );
  XNOR2_X2 U6171 ( .A(n5221), .B(n5220), .ZN(n9561) );
  NAND2_X1 U6172 ( .A1(n5600), .A2(n5599), .ZN(n5138) );
  OAI21_X1 U6173 ( .B1(n8203), .B2(n8201), .A(n8200), .ZN(n4608) );
  NAND2_X1 U6174 ( .A1(n4857), .A2(n5142), .ZN(n5669) );
  NAND3_X1 U6175 ( .A1(n4596), .A2(n4593), .A3(n4575), .ZN(n7847) );
  NAND3_X1 U6176 ( .A1(n4599), .A2(n4598), .A3(n4576), .ZN(n4575) );
  NAND2_X1 U6177 ( .A1(n4871), .A2(n4865), .ZN(n8002) );
  OAI21_X2 U6178 ( .B1(n4590), .B2(n4588), .A(n5095), .ZN(n5413) );
  NAND2_X1 U6179 ( .A1(n4886), .A2(n4885), .ZN(n8034) );
  NOR2_X1 U6180 ( .A1(n4862), .A2(n4500), .ZN(n8146) );
  OAI21_X1 U6181 ( .B1(n4881), .B2(n4876), .A(n4874), .ZN(n8066) );
  NAND3_X1 U6182 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n4585) );
  NOR2_X1 U6183 ( .A1(n5390), .A2(n4591), .ZN(n4588) );
  NAND2_X1 U6184 ( .A1(n5369), .A2(n4586), .ZN(n4590) );
  NAND2_X1 U6185 ( .A1(n4587), .A2(n5092), .ZN(n4586) );
  INV_X1 U6186 ( .A(n5389), .ZN(n4587) );
  INV_X1 U6187 ( .A(n5092), .ZN(n4591) );
  NAND3_X1 U6188 ( .A1(n4597), .A2(n4599), .A3(n4598), .ZN(n4596) );
  NAND2_X1 U6189 ( .A1(n7771), .A2(n7772), .ZN(n4604) );
  OAI21_X1 U6190 ( .B1(n5086), .B2(n4610), .A(n4609), .ZN(n5085) );
  NAND2_X2 U6191 ( .A1(n5099), .A2(n5098), .ZN(n5438) );
  NAND2_X1 U6192 ( .A1(n7728), .A2(n4613), .ZN(n4612) );
  INV_X1 U6193 ( .A(n5438), .ZN(n4620) );
  NAND2_X1 U6194 ( .A1(n4617), .A2(n5119), .ZN(n5543) );
  NAND3_X1 U6195 ( .A1(n4618), .A2(n4531), .A3(n4679), .ZN(n4617) );
  NAND3_X1 U6196 ( .A1(n4618), .A2(n4679), .A3(n4834), .ZN(n5521) );
  NAND2_X1 U6197 ( .A1(n4506), .A2(n4627), .ZN(n4623) );
  NAND3_X1 U6198 ( .A1(n4625), .A2(n4624), .A3(n4623), .ZN(n6338) );
  NAND2_X1 U6199 ( .A1(n8417), .A2(n4634), .ZN(n4630) );
  NAND2_X1 U6200 ( .A1(n4638), .A2(n8838), .ZN(n7021) );
  OAI21_X1 U6201 ( .B1(n9081), .B2(n4638), .A(n9080), .ZN(n9084) );
  XNOR2_X1 U6202 ( .A(n4638), .B(n8838), .ZN(n7209) );
  NAND2_X1 U6203 ( .A1(n5083), .A2(n4644), .ZN(n4643) );
  INV_X1 U6204 ( .A(n5330), .ZN(n4642) );
  NAND3_X1 U6205 ( .A1(n4643), .A2(n5350), .A3(n4641), .ZN(n5090) );
  NAND2_X1 U6206 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n4646), .ZN(n5314) );
  NAND2_X1 U6207 ( .A1(n9089), .A2(n9088), .ZN(n4650) );
  NAND2_X1 U6208 ( .A1(n7222), .A2(n4534), .ZN(n10232) );
  NAND2_X1 U6209 ( .A1(n7024), .A2(n7023), .ZN(n7075) );
  INV_X1 U6210 ( .A(n5219), .ZN(n5218) );
  INV_X1 U6211 ( .A(n4658), .ZN(n4660) );
  OAI21_X1 U6212 ( .B1(n5086), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n4666), .ZN(
        n5080) );
  NAND2_X1 U6213 ( .A1(n5086), .A2(n6495), .ZN(n4666) );
  OAI21_X1 U6214 ( .B1(n9273), .B2(n4668), .A(n4667), .ZN(n9257) );
  NAND2_X1 U6215 ( .A1(n5413), .A2(n5412), .ZN(n5099) );
  NAND3_X1 U6216 ( .A1(n4677), .A2(n4676), .A3(n4555), .ZN(n4833) );
  NAND2_X1 U6217 ( .A1(n5125), .A2(n4693), .ZN(n4688) );
  NAND2_X1 U6218 ( .A1(n5125), .A2(n5124), .ZN(n5561) );
  NAND3_X1 U6219 ( .A1(n4930), .A2(n4931), .A3(n4929), .ZN(n4927) );
  NAND2_X1 U6220 ( .A1(n8298), .A2(n8299), .ZN(n8301) );
  NOR2_X1 U6221 ( .A1(n8300), .A2(n4712), .ZN(n4711) );
  INV_X1 U6222 ( .A(n8299), .ZN(n4712) );
  INV_X1 U6223 ( .A(n8312), .ZN(n4713) );
  INV_X1 U6224 ( .A(n4715), .ZN(n6715) );
  MUX2_X1 U6225 ( .A(n5289), .B(P1_REG2_REG_1__SCAN_IN), .S(n6602), .Z(n6599)
         );
  NAND2_X1 U6226 ( .A1(n4814), .A2(n4813), .ZN(P1_U3520) );
  NAND2_X1 U6227 ( .A1(n9289), .A2(n4736), .ZN(n4735) );
  NAND2_X1 U6228 ( .A1(n9289), .A2(n9284), .ZN(n9278) );
  NAND3_X1 U6229 ( .A1(n4735), .A2(n4734), .A3(n4497), .ZN(n9441) );
  NAND2_X1 U6230 ( .A1(n4744), .A2(n7128), .ZN(n7241) );
  INV_X1 U6231 ( .A(n4749), .ZN(n9329) );
  AND3_X2 U6232 ( .A1(n5298), .A2(n5296), .A3(n5297), .ZN(n10251) );
  OAI21_X1 U6233 ( .B1(n8554), .B2(n10462), .A(n8558), .ZN(n8649) );
  NAND2_X1 U6234 ( .A1(n4770), .A2(n8531), .ZN(n8477) );
  INV_X1 U6235 ( .A(n4774), .ZN(n8492) );
  NAND2_X1 U6236 ( .A1(n7938), .A2(n7945), .ZN(n7087) );
  NAND2_X1 U6237 ( .A1(n8261), .A2(n7903), .ZN(n7945) );
  NAND2_X1 U6238 ( .A1(n8506), .A2(n4495), .ZN(n4779) );
  INV_X1 U6239 ( .A(n4788), .ZN(n8378) );
  INV_X1 U6240 ( .A(n8210), .ZN(n4801) );
  NOR2_X1 U6241 ( .A1(n8110), .A2(n4803), .ZN(n4802) );
  NAND2_X1 U6242 ( .A1(n4941), .A2(n4804), .ZN(n5894) );
  NAND2_X1 U6243 ( .A1(n7668), .A2(n4493), .ZN(n4807) );
  NAND2_X1 U6244 ( .A1(n4807), .A2(n4808), .ZN(n8530) );
  INV_X1 U6245 ( .A(n4809), .ZN(n7669) );
  NAND2_X1 U6246 ( .A1(n7418), .A2(n4810), .ZN(n6144) );
  OR2_X2 U6247 ( .A1(n7416), .A2(n7419), .ZN(n7418) );
  INV_X1 U6248 ( .A(n8014), .ZN(n4812) );
  INV_X1 U6249 ( .A(n7033), .ZN(n8838) );
  NAND2_X1 U6250 ( .A1(n4816), .A2(n9249), .ZN(n9443) );
  NOR2_X1 U6251 ( .A1(n9324), .A2(n4831), .ZN(n9321) );
  NAND2_X1 U6252 ( .A1(n7221), .A2(n8839), .ZN(n7222) );
  NAND2_X1 U6253 ( .A1(n7075), .A2(n4501), .ZN(n7168) );
  NAND2_X1 U6254 ( .A1(n7168), .A2(n8884), .ZN(n7169) );
  AND2_X1 U6255 ( .A1(n7075), .A2(n8936), .ZN(n7232) );
  OR2_X1 U6256 ( .A1(n5439), .A2(n6517), .ZN(n5316) );
  NAND2_X1 U6257 ( .A1(n5196), .A2(n5056), .ZN(n5202) );
  NAND2_X1 U6258 ( .A1(n7342), .A2(n6070), .ZN(n7269) );
  XNOR2_X2 U6259 ( .A(n7922), .B(n8356), .ZN(n8554) );
  AND3_X4 U6260 ( .A1(n5949), .A2(n5948), .A3(n5947), .ZN(n7903) );
  OR2_X2 U6261 ( .A1(n7093), .A2(n7106), .ZN(n6856) );
  NAND2_X1 U6262 ( .A1(n5086), .A2(n5075), .ZN(n5282) );
  NAND2_X1 U6263 ( .A1(n5108), .A2(n5107), .ZN(n5477) );
  NAND2_X1 U6264 ( .A1(n5654), .A2(n4496), .ZN(n4841) );
  NAND2_X1 U6265 ( .A1(n5799), .A2(n4851), .ZN(n4850) );
  NAND2_X1 U6266 ( .A1(n5138), .A2(n4858), .ZN(n4857) );
  AOI21_X2 U6267 ( .B1(n8096), .B2(n8095), .A(n8103), .ZN(n8133) );
  OR2_X2 U6268 ( .A1(n7985), .A2(n4872), .ZN(n4871) );
  NAND2_X1 U6269 ( .A1(n4873), .A2(n4867), .ZN(n4872) );
  NOR2_X1 U6270 ( .A1(n4882), .A2(n4878), .ZN(n4881) );
  NAND2_X1 U6271 ( .A1(n8012), .A2(n8093), .ZN(n4884) );
  NAND3_X1 U6272 ( .A1(n4517), .A2(n4884), .A3(n4883), .ZN(n4886) );
  OAI21_X1 U6273 ( .B1(n6772), .B2(n4890), .A(n6771), .ZN(n6775) );
  AND2_X1 U6274 ( .A1(n6383), .A2(n6385), .ZN(n4890) );
  XNOR2_X2 U6275 ( .A(n6320), .B(n6319), .ZN(n6349) );
  AOI21_X2 U6276 ( .B1(n8213), .B2(n8212), .A(n4513), .ZN(n8203) );
  NAND3_X1 U6277 ( .A1(n4907), .A2(n4897), .A3(n4539), .ZN(n4906) );
  OAI21_X1 U6278 ( .B1(n8165), .B2(n4903), .A(n4901), .ZN(n4907) );
  NAND2_X1 U6279 ( .A1(n4906), .A2(n4905), .ZN(P2_U3222) );
  AOI21_X1 U6280 ( .B1(n7049), .B2(n4909), .A(n4912), .ZN(n4908) );
  INV_X1 U6281 ( .A(n4913), .ZN(n4911) );
  INV_X1 U6282 ( .A(n6789), .ZN(n4920) );
  AOI22_X1 U6283 ( .A1(n4921), .A2(n6802), .B1(n4920), .B2(n4918), .ZN(n6393)
         );
  NOR2_X1 U6284 ( .A1(n6158), .A2(n4938), .ZN(n6307) );
  INV_X1 U6285 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4940) );
  NAND2_X1 U6286 ( .A1(n8501), .A2(n4553), .ZN(n6343) );
  NAND2_X1 U6287 ( .A1(n4947), .A2(n7927), .ZN(n4946) );
  NAND2_X1 U6288 ( .A1(n4949), .A2(n4502), .ZN(n7345) );
  NAND3_X1 U6289 ( .A1(n8108), .A2(n7968), .A3(n8107), .ZN(n4948) );
  NAND2_X1 U6290 ( .A1(n6955), .A2(n4950), .ZN(n4949) );
  INV_X1 U6291 ( .A(n6955), .ZN(n4952) );
  NAND2_X1 U6292 ( .A1(n5892), .A2(n5891), .ZN(n5912) );
  NAND2_X1 U6293 ( .A1(n5892), .A2(n4956), .ZN(n5916) );
  NAND2_X1 U6294 ( .A1(n8385), .A2(n4960), .ZN(n4957) );
  NAND2_X1 U6295 ( .A1(n4957), .A2(n4958), .ZN(n7916) );
  NAND3_X1 U6296 ( .A1(n4967), .A2(n4966), .A3(n6780), .ZN(n6778) );
  NAND3_X1 U6297 ( .A1(n5324), .A2(n5306), .A3(n6633), .ZN(n4967) );
  NAND2_X1 U6298 ( .A1(n8786), .A2(n5324), .ZN(n6779) );
  NAND2_X1 U6299 ( .A1(n8787), .A2(n8788), .ZN(n8786) );
  NAND2_X1 U6300 ( .A1(n8776), .A2(n8778), .ZN(n4978) );
  NAND2_X1 U6301 ( .A1(n4970), .A2(n8776), .ZN(n4969) );
  NAND2_X1 U6302 ( .A1(n8746), .A2(n4518), .ZN(n4980) );
  INV_X1 U6303 ( .A(n5652), .ZN(n4982) );
  NAND2_X1 U6304 ( .A1(n8746), .A2(n8747), .ZN(n8745) );
  NAND2_X1 U6305 ( .A1(n8738), .A2(n8739), .ZN(n4994) );
  NAND2_X1 U6306 ( .A1(n8738), .A2(n4984), .ZN(n4983) );
  NAND2_X1 U6307 ( .A1(n4994), .A2(n4989), .ZN(n8813) );
  AND2_X1 U6308 ( .A1(n4994), .A2(n4993), .ZN(n8815) );
  INV_X1 U6309 ( .A(n5795), .ZN(n4992) );
  NAND2_X1 U6310 ( .A1(n7635), .A2(n7636), .ZN(n7634) );
  NAND2_X1 U6311 ( .A1(n7635), .A2(n4996), .ZN(n4995) );
  OAI21_X1 U6312 ( .B1(n7315), .B2(n5008), .A(n5006), .ZN(n7465) );
  OAI21_X2 U6313 ( .B1(n7001), .B2(n5398), .A(n5404), .ZN(n8692) );
  NAND2_X2 U6314 ( .A1(n6849), .A2(n6844), .ZN(n7001) );
  NAND2_X1 U6315 ( .A1(n5362), .A2(n5361), .ZN(n6849) );
  NOR2_X2 U6316 ( .A1(n5215), .A2(n5012), .ZN(n5837) );
  OAI211_X2 U6317 ( .C1(n5218), .C2(n5017), .A(n5014), .B(n5013), .ZN(n8151)
         );
  NAND2_X1 U6318 ( .A1(n7787), .A2(n5021), .ZN(n5019) );
  INV_X1 U6319 ( .A(n10196), .ZN(n5032) );
  NAND2_X1 U6320 ( .A1(n9217), .A2(n9216), .ZN(n9303) );
  INV_X1 U6321 ( .A(n9216), .ZN(n5040) );
  INV_X1 U6322 ( .A(n9271), .ZN(n9223) );
  NAND2_X1 U6323 ( .A1(n5043), .A2(n5041), .ZN(n9214) );
  NAND2_X1 U6324 ( .A1(n5054), .A2(n5053), .ZN(n7285) );
  NAND3_X1 U6325 ( .A1(n7032), .A2(n7031), .A3(n7033), .ZN(n7200) );
  INV_X1 U6326 ( .A(n7020), .ZN(n7019) );
  AND2_X1 U6327 ( .A1(n5284), .A2(n5283), .ZN(n6628) );
  INV_X1 U6328 ( .A(n6845), .ZN(n5362) );
  NAND2_X1 U6329 ( .A1(n5430), .A2(n5429), .ZN(n7127) );
  CLKBUF_X1 U6330 ( .A(n7013), .Z(n8843) );
  OAI22_X2 U6331 ( .A1(n7607), .A2(n7561), .B1(n7693), .B2(n7611), .ZN(n7701)
         );
  AND2_X1 U6332 ( .A1(n6219), .A2(n6218), .ZN(n8179) );
  INV_X1 U6333 ( .A(n8179), .ZN(n7844) );
  AND4_X1 U6334 ( .A1(n5889), .A2(n5888), .A3(n5887), .A4(n5886), .ZN(n5057)
         );
  AND2_X1 U6335 ( .A1(n8367), .A2(n8187), .ZN(n5059) );
  AND2_X1 U6336 ( .A1(n9284), .A2(n9259), .ZN(n5060) );
  OR2_X1 U6337 ( .A1(n9440), .A2(n10304), .ZN(n5061) );
  OR2_X1 U6338 ( .A1(n4483), .A2(n6662), .ZN(n5062) );
  NAND2_X1 U6339 ( .A1(n10342), .A2(n4509), .ZN(n5063) );
  AND4_X1 U6340 ( .A1(n9053), .A2(n9440), .A3(n9057), .A4(n9258), .ZN(n5064)
         );
  AND2_X1 U6341 ( .A1(n5872), .A2(n8812), .ZN(n5065) );
  INV_X1 U6342 ( .A(n8986), .ZN(n7708) );
  AND4_X1 U6343 ( .A1(n8127), .A2(n8126), .A3(n4964), .A4(n5067), .ZN(n5066)
         );
  AOI21_X1 U6344 ( .B1(n6406), .B2(n5071), .A(n5070), .ZN(n6892) );
  AND4_X1 U6345 ( .A1(n5513), .A2(n5512), .A3(n5511), .A4(n5510), .ZN(n7639)
         );
  AND3_X1 U6346 ( .A1(n6179), .A2(n6178), .A3(n6177), .ZN(n7828) );
  AND4_X1 U6347 ( .A1(n8125), .A2(n4636), .A3(n4791), .A4(n8124), .ZN(n5067)
         );
  OR2_X1 U6348 ( .A1(n7558), .A2(n7639), .ZN(n5068) );
  INV_X1 U6349 ( .A(n7558), .ZN(n9523) );
  AND2_X1 U6350 ( .A1(n8723), .A2(n5688), .ZN(n5069) );
  NOR2_X1 U6351 ( .A1(n6894), .A2(n6890), .ZN(n5070) );
  NOR2_X1 U6352 ( .A1(n6889), .A2(n6894), .ZN(n5071) );
  OR2_X1 U6353 ( .A1(n8256), .A2(n7252), .ZN(n5072) );
  INV_X1 U6354 ( .A(n10344), .ZN(n6015) );
  INV_X1 U6355 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5195) );
  OR2_X1 U6356 ( .A1(n8720), .A2(n8719), .ZN(n5688) );
  INV_X1 U6357 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5207) );
  NOR2_X1 U6358 ( .A1(n8090), .A2(n8088), .ZN(n8126) );
  INV_X1 U6359 ( .A(n8111), .ZN(n6081) );
  INV_X1 U6360 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6045) );
  OR2_X1 U6361 ( .A1(n6627), .A2(n5749), .ZN(n5288) );
  INV_X1 U6362 ( .A(n6203), .ZN(n5908) );
  INV_X1 U6363 ( .A(n6233), .ZN(n6232) );
  XNOR2_X1 U6364 ( .A(n4489), .B(n7903), .ZN(n6382) );
  INV_X1 U6365 ( .A(n6186), .ZN(n5907) );
  INV_X1 U6366 ( .A(n8463), .ZN(n6344) );
  OR2_X1 U6367 ( .A1(n6184), .A2(n9871), .ZN(n6186) );
  NAND2_X1 U6368 ( .A1(n8243), .A2(n8543), .ZN(n6358) );
  INV_X1 U6369 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6131) );
  OR2_X1 U6370 ( .A1(n5856), .A2(n6947), .ZN(n5273) );
  INV_X1 U6371 ( .A(n8898), .ZN(n7707) );
  INV_X1 U6372 ( .A(n8848), .ZN(n7165) );
  NOR2_X1 U6373 ( .A1(n5193), .A2(n5352), .ZN(n5194) );
  INV_X1 U6374 ( .A(SI_12_), .ZN(n9868) );
  INV_X1 U6375 ( .A(SI_9_), .ZN(n9905) );
  OR2_X1 U6376 ( .A1(n6075), .A2(n9692), .ZN(n6091) );
  NAND2_X1 U6377 ( .A1(n6232), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6247) );
  OR2_X1 U6378 ( .A1(n7849), .A2(n4507), .ZN(n7850) );
  INV_X1 U6379 ( .A(n6122), .ZN(n5904) );
  OR2_X1 U6380 ( .A1(n6222), .A2(n5909), .ZN(n6233) );
  AND2_X1 U6381 ( .A1(n7455), .A2(n7454), .ZN(n7457) );
  OR2_X1 U6382 ( .A1(n8003), .A2(n4870), .ZN(n6116) );
  NAND2_X1 U6383 ( .A1(n5901), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6064) );
  NOR2_X1 U6384 ( .A1(n5607), .A2(n7813), .ZN(n5638) );
  INV_X1 U6385 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5455) );
  NAND2_X1 U6386 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(n5761), .ZN(n5760) );
  AND2_X1 U6387 ( .A1(n5718), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5737) );
  OR2_X1 U6388 ( .A1(n5483), .A2(n6840), .ZN(n5508) );
  NAND2_X1 U6389 ( .A1(n5226), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5804) );
  NOR2_X1 U6390 ( .A1(n5679), .A2(n5657), .ZN(n5699) );
  INV_X1 U6391 ( .A(n7072), .ZN(n7023) );
  NAND2_X1 U6392 ( .A1(n5130), .A2(n9941), .ZN(n5133) );
  OR3_X1 U6393 ( .A1(n5522), .A2(P1_IR_REG_11__SCAN_IN), .A3(
        P1_IR_REG_10__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U6394 ( .A1(n5104), .A2(n9905), .ZN(n5107) );
  OR2_X1 U6395 ( .A1(n6256), .A2(n8168), .ZN(n6267) );
  OR2_X1 U6396 ( .A1(n6213), .A2(n7904), .ZN(n6222) );
  OR2_X1 U6397 ( .A1(n6387), .A2(n6386), .ZN(n6388) );
  NAND2_X1 U6398 ( .A1(n7509), .A2(n7508), .ZN(n7586) );
  AND2_X1 U6399 ( .A1(n7654), .A2(n7656), .ZN(n7717) );
  NAND2_X1 U6400 ( .A1(n5904), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6137) );
  INV_X1 U6401 ( .A(n8248), .ZN(n7729) );
  OR2_X1 U6402 ( .A1(n8197), .A2(n4488), .ZN(n6274) );
  OR2_X1 U6403 ( .A1(n6194), .A2(n9900), .ZN(n6203) );
  INV_X1 U6404 ( .A(n8355), .ZN(n7889) );
  OAI21_X1 U6405 ( .B1(n6953), .B2(n6954), .A(n5072), .ZN(n7135) );
  NAND2_X1 U6406 ( .A1(n7937), .A2(n7940), .ZN(n8099) );
  NAND2_X1 U6407 ( .A1(n10376), .A2(n10364), .ZN(n8537) );
  OR2_X1 U6408 ( .A1(n6649), .A2(n6350), .ZN(n8513) );
  AND2_X1 U6409 ( .A1(n7987), .A2(n7986), .ZN(n8111) );
  NOR2_X1 U6410 ( .A1(n5406), .A2(n5405), .ZN(n5431) );
  AND3_X1 U6411 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5381) );
  INV_X1 U6412 ( .A(n6846), .ZN(n5361) );
  NAND2_X1 U6413 ( .A1(n5737), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5738) );
  INV_X1 U6414 ( .A(n7464), .ZN(n5515) );
  OR2_X1 U6415 ( .A1(n5856), .A2(n9282), .ZN(n5229) );
  INV_X1 U6416 ( .A(n5325), .ZN(n5855) );
  INV_X1 U6417 ( .A(n8832), .ZN(n5853) );
  INV_X1 U6418 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6840) );
  INV_X1 U6419 ( .A(n9450), .ZN(n9284) );
  INV_X1 U6420 ( .A(n9469), .ZN(n9345) );
  NAND2_X1 U6421 ( .A1(n9441), .A2(n5061), .ZN(n9442) );
  AND2_X1 U6422 ( .A1(n8962), .A2(n8961), .ZN(n10012) );
  AND2_X1 U6423 ( .A1(n6929), .A2(n6928), .ZN(n10228) );
  NAND2_X1 U6424 ( .A1(n5166), .A2(n5165), .ZN(n5261) );
  AND2_X1 U6425 ( .A1(n5156), .A2(n5155), .ZN(n5695) );
  AND2_X1 U6426 ( .A1(n5137), .A2(n5136), .ZN(n5599) );
  XNOR2_X1 U6427 ( .A(n5126), .B(SI_14_), .ZN(n5560) );
  AND2_X1 U6428 ( .A1(n5112), .A2(n5111), .ZN(n5476) );
  AND2_X1 U6429 ( .A1(n6267), .A2(n6257), .ZN(n8382) );
  AND2_X1 U6430 ( .A1(n8227), .A2(n8543), .ZN(n8217) );
  INV_X1 U6431 ( .A(n8587), .ZN(n8432) );
  NAND2_X1 U6432 ( .A1(n6412), .A2(n6903), .ZN(n7864) );
  INV_X1 U6433 ( .A(n8229), .ZN(n8206) );
  NOR2_X1 U6434 ( .A1(n6453), .A2(n6452), .ZN(n8227) );
  NAND2_X1 U6435 ( .A1(n7926), .A2(n7925), .ZN(n8135) );
  AND4_X1 U6436 ( .A1(n6142), .A2(n6141), .A3(n6140), .A4(n6139), .ZN(n7591)
         );
  OR2_X1 U6437 ( .A1(P2_U3966), .A2(n6672), .ZN(n6657) );
  INV_X1 U6438 ( .A(n9988), .ZN(n10331) );
  NAND2_X1 U6439 ( .A1(n8357), .A2(n7889), .ZN(n8356) );
  INV_X1 U6440 ( .A(n8513), .ZN(n8543) );
  INV_X1 U6441 ( .A(n8553), .ZN(n10352) );
  AND2_X1 U6442 ( .A1(n10423), .A2(n6326), .ZN(n6737) );
  AND2_X1 U6443 ( .A1(n7676), .A2(n8633), .ZN(n10432) );
  INV_X1 U6444 ( .A(n10432), .ZN(n10466) );
  AND3_X1 U6445 ( .A1(n6736), .A2(n6735), .A3(n6734), .ZN(n6751) );
  NAND2_X1 U6446 ( .A1(n6650), .A2(n6318), .ZN(n10390) );
  AND2_X1 U6447 ( .A1(n6145), .A2(n6133), .ZN(n8278) );
  INV_X1 U6448 ( .A(n5478), .ZN(n6545) );
  INV_X1 U6449 ( .A(n10304), .ZN(n9524) );
  AND2_X1 U6450 ( .A1(n9115), .A2(n9114), .ZN(n9120) );
  AND4_X1 U6451 ( .A1(n5861), .A2(n5860), .A3(n5859), .A4(n5858), .ZN(n9258)
         );
  AND2_X1 U6452 ( .A1(n5746), .A2(n5745), .ZN(n9371) );
  AND4_X1 U6453 ( .A1(n5613), .A2(n5612), .A3(n5611), .A4(n5610), .ZN(n7747)
         );
  AND4_X1 U6454 ( .A1(n5533), .A2(n5532), .A3(n5531), .A4(n5530), .ZN(n7555)
         );
  NAND2_X1 U6455 ( .A1(n5325), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5386) );
  INV_X1 U6456 ( .A(n10163), .ZN(n10129) );
  INV_X1 U6457 ( .A(n9222), .ZN(n9274) );
  OR2_X1 U6458 ( .A1(n9231), .A2(n8878), .ZN(n9381) );
  AND2_X1 U6459 ( .A1(n8894), .A2(n8965), .ZN(n8850) );
  AND2_X1 U6460 ( .A1(n6931), .A2(n10049), .ZN(n10226) );
  INV_X1 U6461 ( .A(n10183), .ZN(n10223) );
  NAND2_X1 U6462 ( .A1(n9122), .A2(n6919), .ZN(n10237) );
  OR2_X1 U6463 ( .A1(n6614), .A2(n9116), .ZN(n10304) );
  INV_X1 U6464 ( .A(n10295), .ZN(n9520) );
  AND2_X1 U6465 ( .A1(n6939), .A2(n6918), .ZN(n6620) );
  INV_X4 U6466 ( .A(n5896), .ZN(n7875) );
  OR2_X1 U6467 ( .A1(n8211), .A2(n8186), .ZN(n8224) );
  INV_X1 U6468 ( .A(n8230), .ZN(n8220) );
  INV_X1 U6469 ( .A(n8187), .ZN(n8243) );
  INV_X1 U6470 ( .A(n6241), .ZN(n8437) );
  OR2_X1 U6471 ( .A1(n6172), .A2(n6171), .ZN(n8248) );
  INV_X1 U6472 ( .A(n10376), .ZN(n8548) );
  INV_X1 U6473 ( .A(n10376), .ZN(n10389) );
  INV_X1 U6474 ( .A(n10477), .ZN(n10475) );
  INV_X1 U6475 ( .A(n8397), .ZN(n8660) );
  INV_X1 U6476 ( .A(n8521), .ZN(n8673) );
  CLKBUF_X1 U6477 ( .A(n10406), .Z(n10427) );
  INV_X1 U6478 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6641) );
  INV_X1 U6479 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6524) );
  AND2_X1 U6480 ( .A1(n5868), .A2(n5867), .ZN(n8804) );
  INV_X1 U6481 ( .A(n8791), .ZN(n8824) );
  OR2_X1 U6482 ( .A1(n5724), .A2(n5723), .ZN(n9361) );
  AND2_X1 U6483 ( .A1(n7785), .A2(n7784), .ZN(n9498) );
  INV_X1 U6484 ( .A(n10326), .ZN(n10324) );
  INV_X1 U6485 ( .A(n10315), .ZN(n10313) );
  AND2_X1 U6486 ( .A1(n5863), .A2(n5841), .ZN(n9122) );
  INV_X1 U6487 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9726) );
  INV_X1 U6488 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9899) );
  INV_X1 U6489 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9750) );
  NOR2_X1 U6490 ( .A1(n10508), .A2(n10507), .ZN(n10506) );
  NOR2_X1 U6491 ( .A1(n10505), .A2(n10504), .ZN(n10503) );
  INV_X1 U6492 ( .A(n9138), .ZN(P1_U4006) );
  AND2_X1 U6493 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5075) );
  INV_X1 U6494 ( .A(SI_1_), .ZN(n5076) );
  XNOR2_X1 U6495 ( .A(n5077), .B(n5076), .ZN(n5295) );
  MUX2_X1 U6496 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5086), .Z(n5294) );
  NAND2_X1 U6497 ( .A1(n5295), .A2(n5294), .ZN(n5079) );
  NAND2_X1 U6498 ( .A1(n5077), .A2(SI_1_), .ZN(n5078) );
  NAND2_X1 U6499 ( .A1(n5079), .A2(n5078), .ZN(n5313) );
  INV_X1 U6500 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6518) );
  INV_X1 U6501 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6495) );
  XNOR2_X1 U6502 ( .A(n5080), .B(SI_2_), .ZN(n5312) );
  NAND2_X1 U6503 ( .A1(n5313), .A2(n5312), .ZN(n5083) );
  INV_X1 U6504 ( .A(n5080), .ZN(n5081) );
  NAND2_X1 U6505 ( .A1(n5081), .A2(SI_2_), .ZN(n5082) );
  INV_X1 U6506 ( .A(SI_3_), .ZN(n5084) );
  XNOR2_X1 U6507 ( .A(n5085), .B(n5084), .ZN(n5330) );
  MUX2_X1 U6508 ( .A(n6499), .B(n6496), .S(n5086), .Z(n5087) );
  XNOR2_X1 U6509 ( .A(n5087), .B(SI_4_), .ZN(n5350) );
  INV_X1 U6510 ( .A(n5087), .ZN(n5088) );
  NAND2_X1 U6511 ( .A1(n5088), .A2(SI_4_), .ZN(n5089) );
  MUX2_X1 U6512 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5086), .Z(n5091) );
  INV_X1 U6513 ( .A(SI_5_), .ZN(n9944) );
  NAND2_X1 U6514 ( .A1(n5091), .A2(SI_5_), .ZN(n5092) );
  MUX2_X1 U6515 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7875), .Z(n5094) );
  INV_X1 U6516 ( .A(SI_6_), .ZN(n5093) );
  NAND2_X1 U6517 ( .A1(n5094), .A2(SI_6_), .ZN(n5095) );
  MUX2_X1 U6518 ( .A(n6513), .B(n6511), .S(n7875), .Z(n5096) );
  INV_X1 U6519 ( .A(n5096), .ZN(n5097) );
  NAND2_X1 U6520 ( .A1(n5097), .A2(SI_7_), .ZN(n5098) );
  INV_X1 U6521 ( .A(n5100), .ZN(n5101) );
  NAND2_X1 U6522 ( .A1(n5101), .A2(SI_8_), .ZN(n5102) );
  MUX2_X1 U6523 ( .A(n6536), .B(n9680), .S(n7875), .Z(n5104) );
  INV_X1 U6524 ( .A(n5104), .ZN(n5105) );
  NAND2_X1 U6525 ( .A1(n5105), .A2(SI_9_), .ZN(n5106) );
  MUX2_X1 U6526 ( .A(n6554), .B(n9750), .S(n7875), .Z(n5109) );
  INV_X1 U6527 ( .A(n5109), .ZN(n5110) );
  NAND2_X1 U6528 ( .A1(n5110), .A2(SI_10_), .ZN(n5111) );
  MUX2_X1 U6529 ( .A(n6557), .B(n9934), .S(n7875), .Z(n5113) );
  INV_X1 U6530 ( .A(n5113), .ZN(n5114) );
  INV_X1 U6531 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5115) );
  MUX2_X1 U6532 ( .A(n5115), .B(n9728), .S(n7875), .Z(n5116) );
  INV_X1 U6533 ( .A(n5116), .ZN(n5117) );
  NAND2_X1 U6534 ( .A1(n5117), .A2(SI_12_), .ZN(n5118) );
  MUX2_X1 U6535 ( .A(n6641), .B(n9738), .S(n7875), .Z(n5121) );
  INV_X1 U6536 ( .A(SI_13_), .ZN(n5120) );
  INV_X1 U6537 ( .A(n5121), .ZN(n5122) );
  NAND2_X1 U6538 ( .A1(n5122), .A2(SI_13_), .ZN(n5123) );
  NAND2_X1 U6539 ( .A1(n5543), .A2(n5542), .ZN(n5125) );
  INV_X1 U6540 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6682) );
  MUX2_X1 U6541 ( .A(n6682), .B(n9703), .S(n7875), .Z(n5126) );
  INV_X1 U6542 ( .A(n5126), .ZN(n5127) );
  NAND2_X1 U6543 ( .A1(n5127), .A2(SI_14_), .ZN(n5128) );
  INV_X1 U6544 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6815) );
  MUX2_X1 U6545 ( .A(n6815), .B(n9899), .S(n7875), .Z(n5130) );
  INV_X1 U6546 ( .A(SI_15_), .ZN(n9941) );
  INV_X1 U6547 ( .A(n5130), .ZN(n5131) );
  NAND2_X1 U6548 ( .A1(n5131), .A2(SI_15_), .ZN(n5132) );
  INV_X1 U6549 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6883) );
  MUX2_X1 U6550 ( .A(n6883), .B(n9726), .S(n7875), .Z(n5134) );
  INV_X1 U6551 ( .A(SI_16_), .ZN(n9875) );
  NAND2_X1 U6552 ( .A1(n5134), .A2(n9875), .ZN(n5137) );
  INV_X1 U6553 ( .A(n5134), .ZN(n5135) );
  NAND2_X1 U6554 ( .A1(n5135), .A2(SI_16_), .ZN(n5136) );
  INV_X1 U6555 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6945) );
  INV_X1 U6556 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5139) );
  MUX2_X1 U6557 ( .A(n6945), .B(n5139), .S(n7875), .Z(n5140) );
  XNOR2_X1 U6558 ( .A(n5140), .B(SI_17_), .ZN(n5632) );
  INV_X1 U6559 ( .A(n5140), .ZN(n5141) );
  NAND2_X1 U6560 ( .A1(n5141), .A2(SI_17_), .ZN(n5142) );
  MUX2_X1 U6561 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7875), .Z(n5144) );
  XNOR2_X1 U6562 ( .A(n5144), .B(SI_18_), .ZN(n5668) );
  INV_X1 U6563 ( .A(n5668), .ZN(n5143) );
  NAND2_X1 U6564 ( .A1(n5669), .A2(n5143), .ZN(n5146) );
  NAND2_X1 U6565 ( .A1(n5144), .A2(SI_18_), .ZN(n5145) );
  INV_X1 U6566 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7055) );
  INV_X1 U6567 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n9748) );
  MUX2_X1 U6568 ( .A(n7055), .B(n9748), .S(n7875), .Z(n5148) );
  INV_X1 U6569 ( .A(SI_19_), .ZN(n5147) );
  NAND2_X1 U6570 ( .A1(n5148), .A2(n5147), .ZN(n5151) );
  INV_X1 U6571 ( .A(n5148), .ZN(n5149) );
  NAND2_X1 U6572 ( .A1(n5149), .A2(SI_19_), .ZN(n5150) );
  NAND2_X1 U6573 ( .A1(n5151), .A2(n5150), .ZN(n5653) );
  INV_X1 U6574 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7260) );
  INV_X1 U6575 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7280) );
  MUX2_X1 U6576 ( .A(n7260), .B(n7280), .S(n7875), .Z(n5153) );
  INV_X1 U6577 ( .A(SI_20_), .ZN(n5152) );
  NAND2_X1 U6578 ( .A1(n5153), .A2(n5152), .ZN(n5156) );
  INV_X1 U6579 ( .A(n5153), .ZN(n5154) );
  NAND2_X1 U6580 ( .A1(n5154), .A2(SI_20_), .ZN(n5155) );
  MUX2_X1 U6581 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n7875), .Z(n5157) );
  INV_X1 U6582 ( .A(SI_21_), .ZN(n9877) );
  XNOR2_X1 U6583 ( .A(n5157), .B(n9877), .ZN(n5714) );
  INV_X1 U6584 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7915) );
  INV_X1 U6585 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7373) );
  MUX2_X1 U6586 ( .A(n7915), .B(n7373), .S(n7875), .Z(n5158) );
  INV_X1 U6587 ( .A(SI_22_), .ZN(n9915) );
  NAND2_X1 U6588 ( .A1(n5158), .A2(n9915), .ZN(n5161) );
  INV_X1 U6589 ( .A(n5158), .ZN(n5159) );
  NAND2_X1 U6590 ( .A1(n5159), .A2(SI_22_), .ZN(n5160) );
  NAND2_X1 U6591 ( .A1(n5161), .A2(n5160), .ZN(n5733) );
  INV_X1 U6592 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7437) );
  INV_X1 U6593 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7434) );
  MUX2_X1 U6594 ( .A(n7437), .B(n7434), .S(n7875), .Z(n5162) );
  INV_X1 U6595 ( .A(SI_23_), .ZN(n9884) );
  NAND2_X1 U6596 ( .A1(n5162), .A2(n9884), .ZN(n5165) );
  INV_X1 U6597 ( .A(n5162), .ZN(n5163) );
  NAND2_X1 U6598 ( .A1(n5163), .A2(SI_23_), .ZN(n5164) );
  NAND2_X1 U6599 ( .A1(n5756), .A2(n5755), .ZN(n5166) );
  MUX2_X1 U6600 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n7875), .Z(n5169) );
  INV_X1 U6601 ( .A(SI_24_), .ZN(n5167) );
  XNOR2_X1 U6602 ( .A(n5169), .B(n5167), .ZN(n5260) );
  INV_X1 U6603 ( .A(n5260), .ZN(n5168) );
  NAND2_X1 U6604 ( .A1(n5169), .A2(SI_24_), .ZN(n5170) );
  INV_X1 U6605 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7631) );
  INV_X1 U6606 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9859) );
  MUX2_X1 U6607 ( .A(n7631), .B(n9859), .S(n7875), .Z(n5171) );
  INV_X1 U6608 ( .A(SI_25_), .ZN(n9857) );
  NAND2_X1 U6609 ( .A1(n5171), .A2(n9857), .ZN(n5174) );
  INV_X1 U6610 ( .A(n5171), .ZN(n5172) );
  NAND2_X1 U6611 ( .A1(n5172), .A2(SI_25_), .ZN(n5173) );
  NAND2_X1 U6612 ( .A1(n5174), .A2(n5173), .ZN(n5774) );
  INV_X1 U6613 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7687) );
  INV_X1 U6614 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9940) );
  MUX2_X1 U6615 ( .A(n7687), .B(n9940), .S(n7875), .Z(n5176) );
  INV_X1 U6616 ( .A(SI_26_), .ZN(n5175) );
  NAND2_X1 U6617 ( .A1(n5176), .A2(n5175), .ZN(n5179) );
  INV_X1 U6618 ( .A(n5176), .ZN(n5177) );
  NAND2_X1 U6619 ( .A1(n5177), .A2(SI_26_), .ZN(n5178) );
  NAND2_X1 U6620 ( .A1(n5180), .A2(n5179), .ZN(n5797) );
  INV_X1 U6621 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7762) );
  INV_X1 U6622 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9946) );
  MUX2_X1 U6623 ( .A(n7762), .B(n9946), .S(n7875), .Z(n5181) );
  INV_X1 U6624 ( .A(SI_27_), .ZN(n9753) );
  NAND2_X1 U6625 ( .A1(n5181), .A2(n9753), .ZN(n5798) );
  INV_X1 U6626 ( .A(n5181), .ZN(n5182) );
  NAND2_X1 U6627 ( .A1(n5182), .A2(SI_27_), .ZN(n5183) );
  XNOR2_X1 U6628 ( .A(n5797), .B(n5796), .ZN(n7761) );
  INV_X1 U6629 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5189) );
  INV_X1 U6630 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5188) );
  AND3_X2 U6631 ( .A1(n5463), .A2(n5191), .A3(n5190), .ZN(n5238) );
  NAND2_X1 U6632 ( .A1(n5238), .A2(n5194), .ZN(n5215) );
  NOR2_X1 U6633 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n5198) );
  NOR2_X1 U6634 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5197) );
  NAND4_X1 U6635 ( .A1(n5198), .A2(n5197), .A3(n5207), .A4(n5839), .ZN(n5199)
         );
  NAND2_X1 U6636 ( .A1(n5202), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5204) );
  NAND2_X1 U6637 ( .A1(n7761), .A2(n8866), .ZN(n5206) );
  OR2_X1 U6638 ( .A1(n4484), .A2(n9946), .ZN(n5205) );
  INV_X1 U6639 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5232) );
  NAND2_X1 U6640 ( .A1(n5837), .A2(n5839), .ZN(n5209) );
  NAND2_X1 U6641 ( .A1(n5211), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5208) );
  XNOR2_X1 U6642 ( .A(n5208), .B(P1_IR_REG_25__SCAN_IN), .ZN(n5821) );
  NAND2_X1 U6643 ( .A1(n5209), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5210) );
  XNOR2_X1 U6644 ( .A(n5210), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5820) );
  NAND2_X1 U6645 ( .A1(n5821), .A2(n5820), .ZN(n5214) );
  INV_X1 U6646 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5212) );
  OR2_X2 U6647 ( .A1(n5214), .A2(n7764), .ZN(n5863) );
  NAND2_X1 U6648 ( .A1(n5215), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5217) );
  NAND2_X1 U6649 ( .A1(n5217), .A2(n5195), .ZN(n5216) );
  NAND2_X1 U6650 ( .A1(n5216), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5233) );
  XNOR2_X1 U6651 ( .A(n5233), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6927) );
  XNOR2_X1 U6652 ( .A(n5217), .B(n5195), .ZN(n9437) );
  INV_X2 U6653 ( .A(n4487), .ZN(n5816) );
  INV_X1 U6654 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9552) );
  NAND2_X1 U6655 ( .A1(n5219), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5221) );
  NAND2_X4 U6656 ( .A1(n8151), .A2(n5223), .ZN(n8832) );
  NAND2_X1 U6657 ( .A1(n5853), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5231) );
  INV_X1 U6658 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n5222) );
  OR2_X1 U6659 ( .A1(n5855), .A2(n5222), .ZN(n5230) );
  NAND2_X4 U6660 ( .A1(n5227), .A2(n5223), .ZN(n5856) );
  NAND2_X1 U6661 ( .A1(n5431), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5456) );
  INV_X1 U6662 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U6663 ( .A1(n5527), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5549) );
  INV_X1 U6664 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5548) );
  INV_X1 U6665 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7409) );
  INV_X1 U6666 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7813) );
  NAND2_X1 U6667 ( .A1(n5638), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5677) );
  INV_X1 U6668 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5676) );
  INV_X1 U6669 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5657) );
  INV_X1 U6670 ( .A(n5760), .ZN(n5224) );
  NAND2_X1 U6671 ( .A1(n5224), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5779) );
  INV_X1 U6672 ( .A(n5779), .ZN(n5225) );
  NAND2_X1 U6673 ( .A1(n5225), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5781) );
  INV_X1 U6674 ( .A(n5781), .ZN(n5226) );
  INV_X1 U6675 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8705) );
  XNOR2_X1 U6676 ( .A(n5804), .B(n8705), .ZN(n9282) );
  INV_X1 U6677 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9283) );
  OR2_X1 U6678 ( .A1(n6526), .A2(n9283), .ZN(n5228) );
  NAND2_X1 U6679 ( .A1(n5233), .A2(n5232), .ZN(n5234) );
  NAND2_X1 U6680 ( .A1(n5234), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5235) );
  INV_X1 U6681 ( .A(n9125), .ZN(n8938) );
  INV_X1 U6682 ( .A(n5352), .ZN(n5237) );
  NAND2_X1 U6683 ( .A1(n5462), .A2(n5238), .ZN(n5239) );
  NAND2_X1 U6684 ( .A1(n5239), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5241) );
  XNOR2_X1 U6685 ( .A(n5241), .B(n5240), .ZN(n9332) );
  AND2_X1 U6686 ( .A1(n9437), .A2(n9332), .ZN(n9116) );
  NAND2_X1 U6687 ( .A1(n8938), .A2(n9116), .ZN(n6923) );
  INV_X1 U6688 ( .A(n5278), .ZN(n5812) );
  NOR2_X1 U6689 ( .A1(n9259), .A2(n5812), .ZN(n5242) );
  AOI21_X1 U6690 ( .B1(n9450), .B2(n5816), .A(n5242), .ZN(n8701) );
  INV_X1 U6691 ( .A(n8701), .ZN(n5845) );
  OAI22_X1 U6692 ( .A1(n9284), .A2(n5767), .B1(n9259), .B2(n4487), .ZN(n5243)
         );
  NAND2_X1 U6693 ( .A1(n9125), .A2(n9332), .ZN(n6922) );
  XNOR2_X1 U6694 ( .A(n5243), .B(n7043), .ZN(n8702) );
  NAND2_X1 U6695 ( .A1(n7686), .A2(n8866), .ZN(n5247) );
  OR2_X1 U6696 ( .A1(n4485), .A2(n9940), .ZN(n5246) );
  NAND2_X1 U6697 ( .A1(n5853), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5255) );
  INV_X1 U6698 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n5248) );
  OR2_X1 U6699 ( .A1(n5855), .A2(n5248), .ZN(n5254) );
  INV_X1 U6700 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U6701 ( .A1(n5781), .A2(n5249), .ZN(n5250) );
  NAND2_X1 U6702 ( .A1(n5804), .A2(n5250), .ZN(n8816) );
  OR2_X1 U6703 ( .A1(n5856), .A2(n8816), .ZN(n5253) );
  INV_X1 U6704 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n5251) );
  OR2_X1 U6705 ( .A1(n6526), .A2(n5251), .ZN(n5252) );
  NAND4_X1 U6706 ( .A1(n5255), .A2(n5254), .A3(n5253), .A4(n5252), .ZN(n9220)
         );
  AND2_X1 U6707 ( .A1(n9220), .A2(n5278), .ZN(n5256) );
  AOI21_X1 U6708 ( .B1(n9454), .B2(n5816), .A(n5256), .ZN(n5795) );
  NAND2_X1 U6709 ( .A1(n9454), .A2(n5817), .ZN(n5258) );
  NAND2_X1 U6710 ( .A1(n9220), .A2(n5816), .ZN(n5257) );
  NAND2_X1 U6711 ( .A1(n5258), .A2(n5257), .ZN(n5259) );
  XNOR2_X1 U6712 ( .A(n5259), .B(n7043), .ZN(n5794) );
  XNOR2_X1 U6713 ( .A(n5261), .B(n5260), .ZN(n7549) );
  NAND2_X1 U6714 ( .A1(n7549), .A2(n8866), .ZN(n5263) );
  INV_X1 U6715 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n9928) );
  OR2_X1 U6716 ( .A1(n4484), .A2(n9928), .ZN(n5262) );
  NAND2_X1 U6717 ( .A1(n5325), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5270) );
  INV_X1 U6718 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9334) );
  OR2_X1 U6719 ( .A1(n6526), .A2(n9334), .ZN(n5269) );
  INV_X1 U6720 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5264) );
  NAND2_X1 U6721 ( .A1(n5760), .A2(n5264), .ZN(n5265) );
  NAND2_X1 U6722 ( .A1(n5779), .A2(n5265), .ZN(n8757) );
  OR2_X1 U6723 ( .A1(n5856), .A2(n8757), .ZN(n5268) );
  INV_X1 U6724 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5266) );
  OR2_X1 U6725 ( .A1(n8832), .A2(n5266), .ZN(n5267) );
  NAND4_X1 U6726 ( .A1(n5270), .A2(n5269), .A3(n5268), .A4(n5267), .ZN(n9349)
         );
  AOI22_X1 U6727 ( .A1(n9330), .A2(n5816), .B1(n5278), .B2(n9349), .ZN(n5771)
         );
  INV_X1 U6728 ( .A(n5771), .ZN(n5773) );
  AOI22_X1 U6729 ( .A1(n9330), .A2(n5817), .B1(n5816), .B2(n9349), .ZN(n5271)
         );
  XNOR2_X1 U6730 ( .A(n5271), .B(n7043), .ZN(n5770) );
  INV_X1 U6731 ( .A(n5770), .ZN(n5772) );
  NAND2_X1 U6732 ( .A1(n5325), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5275) );
  INV_X1 U6733 ( .A(n8832), .ZN(n5272) );
  INV_X1 U6734 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6947) );
  AND3_X1 U6735 ( .A1(n5275), .A2(n5274), .A3(n5273), .ZN(n5277) );
  INV_X1 U6736 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6542) );
  OR2_X1 U6737 ( .A1(n6526), .A2(n6542), .ZN(n5276) );
  NAND2_X1 U6738 ( .A1(n7875), .A2(SI_0_), .ZN(n5280) );
  INV_X1 U6739 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5279) );
  NAND2_X1 U6740 ( .A1(n5280), .A2(n5279), .ZN(n5281) );
  AND2_X1 U6741 ( .A1(n5282), .A2(n5281), .ZN(n9563) );
  MUX2_X1 U6742 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9563), .S(n5478), .Z(n6946) );
  INV_X1 U6743 ( .A(n5863), .ZN(n6371) );
  AOI22_X1 U6744 ( .A1(n5491), .A2(n6946), .B1(n6371), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5283) );
  AOI22_X1 U6745 ( .A1(n5285), .A2(n6946), .B1(n6371), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U6746 ( .A1(n5287), .A2(n5286), .ZN(n6627) );
  NAND2_X1 U6747 ( .A1(n6628), .A2(n6627), .ZN(n6626) );
  INV_X1 U6748 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6596) );
  NAND2_X1 U6749 ( .A1(n5325), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5292) );
  INV_X1 U6750 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5289) );
  OR2_X1 U6751 ( .A1(n6526), .A2(n5289), .ZN(n5291) );
  INV_X1 U6752 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6590) );
  NAND4_X2 U6753 ( .A1(n5293), .A2(n5292), .A3(n5291), .A4(n5290), .ZN(n6920)
         );
  NAND2_X1 U6754 ( .A1(n6920), .A2(n5491), .ZN(n5300) );
  XNOR2_X1 U6755 ( .A(n5295), .B(n5294), .ZN(n6514) );
  OR2_X1 U6756 ( .A1(n5439), .A2(n6514), .ZN(n5298) );
  INV_X1 U6757 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6509) );
  OR2_X1 U6758 ( .A1(n4484), .A2(n6509), .ZN(n5297) );
  OR2_X1 U6759 ( .A1(n5478), .A2(n6602), .ZN(n5296) );
  OR2_X1 U6760 ( .A1(n5767), .A2(n10251), .ZN(n5299) );
  NAND2_X1 U6761 ( .A1(n5300), .A2(n5299), .ZN(n5301) );
  XNOR2_X1 U6762 ( .A(n5301), .B(n7043), .ZN(n5303) );
  AOI22_X1 U6763 ( .A1(n6920), .A2(n5278), .B1(n7030), .B2(n5491), .ZN(n6634)
         );
  NAND2_X1 U6764 ( .A1(n6632), .A2(n6634), .ZN(n5306) );
  INV_X1 U6765 ( .A(n5302), .ZN(n5305) );
  INV_X1 U6766 ( .A(n5303), .ZN(n5304) );
  NAND2_X1 U6767 ( .A1(n5305), .A2(n5304), .ZN(n6633) );
  NAND2_X1 U6768 ( .A1(n5325), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5310) );
  INV_X1 U6769 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10054) );
  OR2_X1 U6770 ( .A1(n8832), .A2(n10054), .ZN(n5309) );
  INV_X1 U6771 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7204) );
  INV_X1 U6772 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7203) );
  NAND2_X1 U6773 ( .A1(n7020), .A2(n5491), .ZN(n5319) );
  OR2_X1 U6774 ( .A1(n4485), .A2(n6495), .ZN(n5317) );
  XNOR2_X1 U6775 ( .A(n5313), .B(n5312), .ZN(n6517) );
  INV_X1 U6776 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5464) );
  INV_X1 U6777 ( .A(n10053), .ZN(n10059) );
  OR2_X1 U6778 ( .A1(n5478), .A2(n10059), .ZN(n5315) );
  OR2_X1 U6779 ( .A1(n5767), .A2(n10257), .ZN(n5318) );
  NAND2_X1 U6780 ( .A1(n5319), .A2(n5318), .ZN(n5320) );
  XNOR2_X1 U6781 ( .A(n5320), .B(n5749), .ZN(n5322) );
  AOI22_X1 U6782 ( .A1(n7020), .A2(n5278), .B1(n7018), .B2(n5491), .ZN(n5321)
         );
  NAND2_X1 U6783 ( .A1(n5322), .A2(n5321), .ZN(n5324) );
  OR2_X1 U6784 ( .A1(n5322), .A2(n5321), .ZN(n5323) );
  NAND2_X1 U6785 ( .A1(n5325), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5329) );
  INV_X1 U6786 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7215) );
  OR2_X1 U6787 ( .A1(n6526), .A2(n7215), .ZN(n5328) );
  INV_X1 U6788 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6476) );
  OR2_X1 U6789 ( .A1(n8832), .A2(n6476), .ZN(n5327) );
  OR2_X1 U6790 ( .A1(n5856), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5326) );
  NAND4_X1 U6791 ( .A1(n5329), .A2(n5328), .A3(n5327), .A4(n5326), .ZN(n10225)
         );
  NAND2_X1 U6792 ( .A1(n10225), .A2(n5491), .ZN(n5338) );
  XNOR2_X1 U6793 ( .A(n5331), .B(n5330), .ZN(n6506) );
  OR2_X1 U6794 ( .A1(n5439), .A2(n6506), .ZN(n5336) );
  INV_X1 U6795 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6507) );
  OR2_X1 U6796 ( .A1(n4484), .A2(n6507), .ZN(n5335) );
  NAND2_X1 U6797 ( .A1(n5352), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5333) );
  INV_X1 U6798 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5332) );
  XNOR2_X1 U6799 ( .A(n5333), .B(n5332), .ZN(n6505) );
  OR2_X1 U6800 ( .A1(n4482), .A2(n6505), .ZN(n5334) );
  OR2_X1 U6801 ( .A1(n5767), .A2(n10264), .ZN(n5337) );
  NAND2_X1 U6802 ( .A1(n5338), .A2(n5337), .ZN(n5339) );
  XNOR2_X1 U6803 ( .A(n5339), .B(n7043), .ZN(n5340) );
  INV_X1 U6804 ( .A(n10264), .ZN(n7220) );
  AOI22_X1 U6805 ( .A1(n10225), .A2(n5278), .B1(n7220), .B2(n5491), .ZN(n5341)
         );
  XNOR2_X1 U6806 ( .A(n5340), .B(n5341), .ZN(n6780) );
  INV_X1 U6807 ( .A(n5340), .ZN(n5342) );
  NAND2_X1 U6808 ( .A1(n5342), .A2(n5341), .ZN(n5343) );
  NAND2_X1 U6809 ( .A1(n6778), .A2(n5343), .ZN(n6845) );
  NAND2_X1 U6810 ( .A1(n5325), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5349) );
  INV_X1 U6811 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5344) );
  OR2_X1 U6812 ( .A1(n8832), .A2(n5344), .ZN(n5348) );
  XNOR2_X1 U6813 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n10238) );
  OR2_X1 U6814 ( .A1(n5856), .A2(n10238), .ZN(n5347) );
  INV_X1 U6815 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5345) );
  OR2_X1 U6816 ( .A1(n6526), .A2(n5345), .ZN(n5346) );
  NAND4_X1 U6817 ( .A1(n5349), .A2(n5348), .A3(n5347), .A4(n5346), .ZN(n9137)
         );
  NAND2_X1 U6818 ( .A1(n9137), .A2(n5491), .ZN(n5359) );
  OR2_X1 U6819 ( .A1(n4484), .A2(n6496), .ZN(n5357) );
  XNOR2_X1 U6820 ( .A(n5351), .B(n5350), .ZN(n6498) );
  OR2_X1 U6821 ( .A1(n5439), .A2(n6498), .ZN(n5356) );
  OR2_X1 U6822 ( .A1(n5352), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U6823 ( .A1(n5353), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5354) );
  XNOR2_X1 U6824 ( .A(n5354), .B(P1_IR_REG_4__SCAN_IN), .ZN(n10069) );
  INV_X1 U6825 ( .A(n10069), .ZN(n6497) );
  OR2_X1 U6826 ( .A1(n5478), .A2(n6497), .ZN(n5355) );
  OR2_X1 U6827 ( .A1(n5767), .A2(n10270), .ZN(n5358) );
  NAND2_X1 U6828 ( .A1(n5359), .A2(n5358), .ZN(n5360) );
  XNOR2_X1 U6829 ( .A(n5360), .B(n5749), .ZN(n5364) );
  INV_X1 U6830 ( .A(n10270), .ZN(n7038) );
  AOI22_X1 U6831 ( .A1(n9137), .A2(n5278), .B1(n7038), .B2(n5816), .ZN(n5363)
         );
  AND2_X1 U6832 ( .A1(n5364), .A2(n5363), .ZN(n6846) );
  OR2_X1 U6833 ( .A1(n5364), .A2(n5363), .ZN(n6844) );
  NAND2_X1 U6834 ( .A1(n5325), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5368) );
  INV_X1 U6835 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6480) );
  OR2_X1 U6836 ( .A1(n8832), .A2(n6480), .ZN(n5367) );
  OAI21_X1 U6837 ( .B1(n5381), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5406), .ZN(
        n10185) );
  OR2_X1 U6838 ( .A1(n5856), .A2(n10185), .ZN(n5366) );
  INV_X1 U6839 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6461) );
  OR2_X1 U6840 ( .A1(n6526), .A2(n6461), .ZN(n5365) );
  NAND4_X1 U6841 ( .A1(n5368), .A2(n5367), .A3(n5366), .A4(n5365), .ZN(n10204)
         );
  NAND2_X1 U6842 ( .A1(n10204), .A2(n5491), .ZN(n5377) );
  XNOR2_X1 U6843 ( .A(n5370), .B(n5369), .ZN(n6508) );
  OR2_X1 U6844 ( .A1(n5439), .A2(n6508), .ZN(n5375) );
  INV_X1 U6845 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9755) );
  OR2_X1 U6846 ( .A1(n4485), .A2(n9755), .ZN(n5374) );
  INV_X1 U6847 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9932) );
  AND2_X1 U6848 ( .A1(n5462), .A2(n9932), .ZN(n5371) );
  INV_X1 U6849 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9620) );
  XNOR2_X1 U6850 ( .A(n5372), .B(n9620), .ZN(n6588) );
  OR2_X1 U6851 ( .A1(n4482), .A2(n6588), .ZN(n5373) );
  OR2_X1 U6852 ( .A1(n5767), .A2(n10189), .ZN(n5376) );
  NAND2_X1 U6853 ( .A1(n5377), .A2(n5376), .ZN(n5378) );
  XNOR2_X1 U6854 ( .A(n5378), .B(n7043), .ZN(n7004) );
  NAND2_X1 U6855 ( .A1(n10204), .A2(n5278), .ZN(n5380) );
  OR2_X1 U6856 ( .A1(n4487), .A2(n10189), .ZN(n5379) );
  NAND2_X1 U6857 ( .A1(n5380), .A2(n5379), .ZN(n7003) );
  NAND2_X1 U6858 ( .A1(n7004), .A2(n7003), .ZN(n5402) );
  INV_X1 U6859 ( .A(n5856), .ZN(n5740) );
  AOI21_X1 U6860 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5382) );
  NOR2_X1 U6861 ( .A1(n5382), .A2(n5381), .ZN(n10202) );
  NAND2_X1 U6862 ( .A1(n5740), .A2(n10202), .ZN(n5387) );
  INV_X1 U6863 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6472) );
  OR2_X1 U6864 ( .A1(n8832), .A2(n6472), .ZN(n5385) );
  INV_X1 U6865 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5383) );
  OR2_X1 U6866 ( .A1(n6526), .A2(n5383), .ZN(n5384) );
  NAND4_X1 U6867 ( .A1(n5387), .A2(n5386), .A3(n5385), .A4(n5384), .ZN(n10224)
         );
  NAND2_X1 U6868 ( .A1(n10224), .A2(n5491), .ZN(n5393) );
  OR2_X1 U6869 ( .A1(n5462), .A2(n5464), .ZN(n5388) );
  XNOR2_X1 U6870 ( .A(n5388), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9156) );
  INV_X1 U6871 ( .A(n9156), .ZN(n6503) );
  INV_X1 U6872 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6501) );
  OR2_X1 U6873 ( .A1(n4484), .A2(n6501), .ZN(n5391) );
  NAND2_X1 U6874 ( .A1(n5817), .A2(n10200), .ZN(n5392) );
  NAND2_X1 U6875 ( .A1(n5393), .A2(n5392), .ZN(n5394) );
  XNOR2_X1 U6876 ( .A(n5394), .B(n7043), .ZN(n7002) );
  NAND2_X1 U6877 ( .A1(n10224), .A2(n5278), .ZN(n5396) );
  NAND2_X1 U6878 ( .A1(n5491), .A2(n10200), .ZN(n5395) );
  NAND2_X1 U6879 ( .A1(n5396), .A2(n5395), .ZN(n5399) );
  NAND2_X1 U6880 ( .A1(n7002), .A2(n5399), .ZN(n5397) );
  NAND2_X1 U6881 ( .A1(n5402), .A2(n5397), .ZN(n5398) );
  INV_X1 U6882 ( .A(n7002), .ZN(n6967) );
  INV_X1 U6883 ( .A(n5399), .ZN(n6969) );
  AND2_X1 U6884 ( .A1(n6967), .A2(n6969), .ZN(n5403) );
  INV_X1 U6885 ( .A(n7003), .ZN(n5401) );
  INV_X1 U6886 ( .A(n7004), .ZN(n5400) );
  AOI22_X1 U6887 ( .A1(n5403), .A2(n5402), .B1(n5401), .B2(n5400), .ZN(n5404)
         );
  NAND2_X1 U6888 ( .A1(n5325), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5411) );
  INV_X1 U6889 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6481) );
  OR2_X1 U6890 ( .A1(n8832), .A2(n6481), .ZN(n5410) );
  AND2_X1 U6891 ( .A1(n5406), .A2(n5405), .ZN(n5407) );
  OR2_X1 U6892 ( .A1(n5407), .A2(n5431), .ZN(n8696) );
  OR2_X1 U6893 ( .A1(n5856), .A2(n8696), .ZN(n5409) );
  INV_X1 U6894 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7026) );
  OR2_X1 U6895 ( .A1(n6526), .A2(n7026), .ZN(n5408) );
  NAND4_X1 U6896 ( .A1(n5411), .A2(n5410), .A3(n5409), .A4(n5408), .ZN(n10174)
         );
  NAND2_X1 U6897 ( .A1(n10174), .A2(n5278), .ZN(n5422) );
  XNOR2_X1 U6898 ( .A(n5413), .B(n5412), .ZN(n6512) );
  OR2_X1 U6899 ( .A1(n5439), .A2(n6512), .ZN(n5420) );
  OR2_X1 U6900 ( .A1(n4484), .A2(n6511), .ZN(n5419) );
  NAND2_X1 U6901 ( .A1(n5462), .A2(n5415), .ZN(n5416) );
  NAND2_X1 U6902 ( .A1(n5416), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5417) );
  XNOR2_X1 U6903 ( .A(n5417), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6573) );
  INV_X1 U6904 ( .A(n6573), .ZN(n6510) );
  OR2_X1 U6905 ( .A1(n4482), .A2(n6510), .ZN(n5418) );
  OR2_X1 U6906 ( .A1(n4487), .A2(n10292), .ZN(n5421) );
  AND2_X1 U6907 ( .A1(n5422), .A2(n5421), .ZN(n8689) );
  NAND2_X1 U6908 ( .A1(n8692), .A2(n8689), .ZN(n5426) );
  NAND2_X1 U6909 ( .A1(n10174), .A2(n5491), .ZN(n5424) );
  OR2_X1 U6910 ( .A1(n5767), .A2(n10292), .ZN(n5423) );
  NAND2_X1 U6911 ( .A1(n5424), .A2(n5423), .ZN(n5425) );
  XNOR2_X1 U6912 ( .A(n5425), .B(n7043), .ZN(n8690) );
  NAND2_X1 U6913 ( .A1(n5426), .A2(n8690), .ZN(n5430) );
  INV_X1 U6914 ( .A(n8692), .ZN(n5428) );
  INV_X1 U6915 ( .A(n8689), .ZN(n5427) );
  NAND2_X1 U6916 ( .A1(n5428), .A2(n5427), .ZN(n5429) );
  NAND2_X1 U6917 ( .A1(n5325), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5436) );
  INV_X1 U6918 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7238) );
  OR2_X1 U6919 ( .A1(n6526), .A2(n7238), .ZN(n5435) );
  OR2_X1 U6920 ( .A1(n5431), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5432) );
  NAND2_X1 U6921 ( .A1(n5456), .A2(n5432), .ZN(n7237) );
  OR2_X1 U6922 ( .A1(n5856), .A2(n7237), .ZN(n5434) );
  INV_X1 U6923 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6471) );
  OR2_X1 U6924 ( .A1(n8832), .A2(n6471), .ZN(n5433) );
  NAND4_X1 U6925 ( .A1(n5436), .A2(n5435), .A3(n5434), .A4(n5433), .ZN(n9136)
         );
  NAND2_X1 U6926 ( .A1(n9136), .A2(n5278), .ZN(n5448) );
  XNOR2_X1 U6927 ( .A(n5438), .B(n5437), .ZN(n6523) );
  OR2_X1 U6928 ( .A1(n5439), .A2(n6523), .ZN(n5446) );
  OR2_X1 U6929 ( .A1(n4484), .A2(n6522), .ZN(n5445) );
  AND2_X1 U6930 ( .A1(n5415), .A2(n5440), .ZN(n5441) );
  NAND2_X1 U6931 ( .A1(n5462), .A2(n5441), .ZN(n5442) );
  NAND2_X1 U6932 ( .A1(n5442), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5443) );
  XNOR2_X1 U6933 ( .A(n5443), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10080) );
  INV_X1 U6934 ( .A(n10080), .ZN(n6521) );
  OR2_X1 U6935 ( .A1(n5478), .A2(n6521), .ZN(n5444) );
  OR2_X1 U6936 ( .A1(n4487), .A2(n7128), .ZN(n5447) );
  NAND2_X1 U6937 ( .A1(n5448), .A2(n5447), .ZN(n7125) );
  NAND2_X1 U6938 ( .A1(n9136), .A2(n5816), .ZN(n5450) );
  OR2_X1 U6939 ( .A1(n5767), .A2(n7128), .ZN(n5449) );
  NAND2_X1 U6940 ( .A1(n5450), .A2(n5449), .ZN(n5451) );
  XNOR2_X1 U6941 ( .A(n5451), .B(n7043), .ZN(n7124) );
  OAI21_X1 U6942 ( .B1(n7127), .B2(n7125), .A(n7124), .ZN(n5453) );
  NAND2_X1 U6943 ( .A1(n7127), .A2(n7125), .ZN(n5452) );
  NAND2_X1 U6944 ( .A1(n5453), .A2(n5452), .ZN(n7315) );
  NAND2_X1 U6945 ( .A1(n5325), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5461) );
  INV_X1 U6946 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5454) );
  OR2_X1 U6947 ( .A1(n8832), .A2(n5454), .ZN(n5460) );
  NAND2_X1 U6948 ( .A1(n5456), .A2(n5455), .ZN(n5457) );
  NAND2_X1 U6949 ( .A1(n5483), .A2(n5457), .ZN(n7324) );
  OR2_X1 U6950 ( .A1(n5856), .A2(n7324), .ZN(n5459) );
  INV_X1 U6951 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7082) );
  OR2_X1 U6952 ( .A1(n6526), .A2(n7082), .ZN(n5458) );
  NAND4_X1 U6953 ( .A1(n5461), .A2(n5460), .A3(n5459), .A4(n5458), .ZN(n9135)
         );
  NAND2_X1 U6954 ( .A1(n9135), .A2(n5816), .ZN(n5470) );
  AND2_X1 U6955 ( .A1(n5463), .A2(n5462), .ZN(n5480) );
  OR2_X1 U6956 ( .A1(n5480), .A2(n5464), .ZN(n5465) );
  XNOR2_X1 U6957 ( .A(n5465), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6835) );
  INV_X1 U6958 ( .A(n6835), .ZN(n6534) );
  NAND2_X1 U6959 ( .A1(n6533), .A2(n8866), .ZN(n5468) );
  OR2_X1 U6960 ( .A1(n4485), .A2(n9680), .ZN(n5467) );
  OAI211_X1 U6961 ( .C1(n4482), .C2(n6534), .A(n5468), .B(n5467), .ZN(n7322)
         );
  NAND2_X1 U6962 ( .A1(n7322), .A2(n5817), .ZN(n5469) );
  NAND2_X1 U6963 ( .A1(n5470), .A2(n5469), .ZN(n5471) );
  XNOR2_X1 U6964 ( .A(n5471), .B(n5749), .ZN(n5473) );
  AOI22_X1 U6965 ( .A1(n9135), .A2(n5278), .B1(n5491), .B2(n7322), .ZN(n5472)
         );
  NAND2_X1 U6966 ( .A1(n5473), .A2(n5472), .ZN(n5475) );
  OR2_X1 U6967 ( .A1(n5473), .A2(n5472), .ZN(n5474) );
  NAND2_X1 U6968 ( .A1(n5475), .A2(n5474), .ZN(n7314) );
  NAND2_X1 U6969 ( .A1(n6552), .A2(n8866), .ZN(n5482) );
  INV_X1 U6970 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U6971 ( .A1(n5480), .A2(n5479), .ZN(n5522) );
  NAND2_X1 U6972 ( .A1(n5522), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5501) );
  XNOR2_X1 U6973 ( .A(n5501), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6873) );
  AOI22_X1 U6974 ( .A1(n5673), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6545), .B2(
        n6873), .ZN(n5481) );
  NAND2_X1 U6975 ( .A1(n5325), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U6976 ( .A1(n5483), .A2(n6840), .ZN(n5484) );
  NAND2_X1 U6977 ( .A1(n5508), .A2(n5484), .ZN(n7495) );
  OR2_X1 U6978 ( .A1(n5856), .A2(n7495), .ZN(n5487) );
  INV_X1 U6979 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7178) );
  OR2_X1 U6980 ( .A1(n6526), .A2(n7178), .ZN(n5486) );
  INV_X1 U6981 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6831) );
  OR2_X1 U6982 ( .A1(n8832), .A2(n6831), .ZN(n5485) );
  NAND4_X1 U6983 ( .A1(n5488), .A2(n5487), .A3(n5486), .A4(n5485), .ZN(n9134)
         );
  NAND2_X1 U6984 ( .A1(n9134), .A2(n5816), .ZN(n5489) );
  OAI21_X1 U6985 ( .B1(n10002), .B2(n5767), .A(n5489), .ZN(n5490) );
  XNOR2_X1 U6986 ( .A(n5490), .B(n7043), .ZN(n5494) );
  OR2_X1 U6987 ( .A1(n10002), .A2(n4487), .ZN(n5493) );
  NAND2_X1 U6988 ( .A1(n9134), .A2(n5278), .ZN(n5492) );
  NAND2_X1 U6989 ( .A1(n5493), .A2(n5492), .ZN(n5495) );
  NAND2_X1 U6990 ( .A1(n5494), .A2(n5495), .ZN(n7497) );
  INV_X1 U6991 ( .A(n5494), .ZN(n5497) );
  INV_X1 U6992 ( .A(n5495), .ZN(n5496) );
  NAND2_X1 U6993 ( .A1(n5497), .A2(n5496), .ZN(n7496) );
  INV_X1 U6994 ( .A(n7465), .ZN(n5516) );
  XNOR2_X1 U6995 ( .A(n5499), .B(n5498), .ZN(n6555) );
  NAND2_X1 U6996 ( .A1(n6555), .A2(n8866), .ZN(n5505) );
  INV_X1 U6997 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U6998 ( .A1(n5501), .A2(n5500), .ZN(n5502) );
  NAND2_X1 U6999 ( .A1(n5502), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5503) );
  XNOR2_X1 U7000 ( .A(n5503), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7063) );
  AOI22_X1 U7001 ( .A1(n5673), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6545), .B2(
        n7063), .ZN(n5504) );
  NAND2_X1 U7002 ( .A1(n5325), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5513) );
  INV_X1 U7003 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5506) );
  OR2_X1 U7004 ( .A1(n8832), .A2(n5506), .ZN(n5512) );
  AND2_X1 U7005 ( .A1(n5508), .A2(n5507), .ZN(n5509) );
  OR2_X1 U7006 ( .A1(n5509), .A2(n5527), .ZN(n7471) );
  OR2_X1 U7007 ( .A1(n5856), .A2(n7471), .ZN(n5511) );
  INV_X1 U7008 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7293) );
  OR2_X1 U7009 ( .A1(n6526), .A2(n7293), .ZN(n5510) );
  OAI22_X1 U7010 ( .A1(n7558), .A2(n5767), .B1(n7639), .B2(n4487), .ZN(n5514)
         );
  XNOR2_X1 U7011 ( .A(n5514), .B(n7043), .ZN(n5518) );
  OAI22_X1 U7012 ( .A1(n7558), .A2(n4487), .B1(n7639), .B2(n5812), .ZN(n5517)
         );
  XNOR2_X1 U7013 ( .A(n5518), .B(n5517), .ZN(n7464) );
  NAND2_X1 U7014 ( .A1(n5516), .A2(n5515), .ZN(n7466) );
  NAND2_X1 U7015 ( .A1(n5518), .A2(n5517), .ZN(n5519) );
  AND2_X2 U7016 ( .A1(n7466), .A2(n5519), .ZN(n7635) );
  XNOR2_X1 U7017 ( .A(n5521), .B(n5520), .ZN(n6603) );
  NAND2_X1 U7018 ( .A1(n6603), .A2(n8866), .ZN(n5525) );
  NAND2_X1 U7019 ( .A1(n5544), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5523) );
  XNOR2_X1 U7020 ( .A(n5523), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7068) );
  AOI22_X1 U7021 ( .A1(n5673), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6545), .B2(
        n7068), .ZN(n5524) );
  NAND2_X1 U7022 ( .A1(n10020), .A2(n5817), .ZN(n5535) );
  NAND2_X1 U7023 ( .A1(n5325), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5533) );
  INV_X1 U7024 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n5526) );
  OR2_X1 U7025 ( .A1(n6526), .A2(n5526), .ZN(n5532) );
  OR2_X1 U7026 ( .A1(n5527), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5528) );
  NAND2_X1 U7027 ( .A1(n5549), .A2(n5528), .ZN(n10018) );
  OR2_X1 U7028 ( .A1(n5856), .A2(n10018), .ZN(n5531) );
  INV_X1 U7029 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5529) );
  OR2_X1 U7030 ( .A1(n8832), .A2(n5529), .ZN(n5530) );
  OR2_X1 U7031 ( .A1(n7555), .A2(n4487), .ZN(n5534) );
  NAND2_X1 U7032 ( .A1(n5535), .A2(n5534), .ZN(n5536) );
  XNOR2_X1 U7033 ( .A(n5536), .B(n7043), .ZN(n5538) );
  NOR2_X1 U7034 ( .A1(n7555), .A2(n5812), .ZN(n5537) );
  AOI21_X1 U7035 ( .B1(n10020), .B2(n5816), .A(n5537), .ZN(n5539) );
  XNOR2_X1 U7036 ( .A(n5538), .B(n5539), .ZN(n7636) );
  INV_X1 U7037 ( .A(n5538), .ZN(n5540) );
  NAND2_X1 U7038 ( .A1(n5540), .A2(n5539), .ZN(n5541) );
  XNOR2_X1 U7039 ( .A(n5543), .B(n5542), .ZN(n6639) );
  NAND2_X1 U7040 ( .A1(n6639), .A2(n8866), .ZN(n5547) );
  NOR2_X1 U7041 ( .A1(n5544), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5563) );
  OR2_X1 U7042 ( .A1(n5563), .A2(n5464), .ZN(n5545) );
  XNOR2_X1 U7043 ( .A(n5545), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7407) );
  AOI22_X1 U7044 ( .A1(n5673), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6545), .B2(
        n7407), .ZN(n5546) );
  NAND2_X1 U7045 ( .A1(n9516), .A2(n5817), .ZN(n5556) );
  NAND2_X1 U7046 ( .A1(n5325), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5554) );
  INV_X1 U7047 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7403) );
  OR2_X1 U7048 ( .A1(n6526), .A2(n7403), .ZN(n5553) );
  NAND2_X1 U7049 ( .A1(n5549), .A2(n5548), .ZN(n5550) );
  NAND2_X1 U7050 ( .A1(n5571), .A2(n5550), .ZN(n7650) );
  OR2_X1 U7051 ( .A1(n5856), .A2(n7650), .ZN(n5552) );
  INV_X1 U7052 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7399) );
  OR2_X1 U7053 ( .A1(n8832), .A2(n7399), .ZN(n5551) );
  NAND4_X1 U7054 ( .A1(n5554), .A2(n5553), .A3(n5552), .A4(n5551), .ZN(n10013)
         );
  NAND2_X1 U7055 ( .A1(n10013), .A2(n5816), .ZN(n5555) );
  NAND2_X1 U7056 ( .A1(n5556), .A2(n5555), .ZN(n5557) );
  XNOR2_X1 U7057 ( .A(n5557), .B(n5749), .ZN(n7645) );
  AND2_X1 U7058 ( .A1(n10013), .A2(n5278), .ZN(n5558) );
  AOI21_X1 U7059 ( .B1(n9516), .B2(n5816), .A(n5558), .ZN(n7644) );
  AND2_X1 U7060 ( .A1(n7645), .A2(n7644), .ZN(n5559) );
  XNOR2_X1 U7061 ( .A(n5561), .B(n5560), .ZN(n6680) );
  NAND2_X1 U7062 ( .A1(n6680), .A2(n8866), .ZN(n5569) );
  AND2_X1 U7063 ( .A1(n5563), .A2(n5562), .ZN(n5602) );
  OR2_X1 U7064 ( .A1(n5602), .A2(n5464), .ZN(n5566) );
  INV_X1 U7065 ( .A(n5566), .ZN(n5564) );
  NAND2_X1 U7066 ( .A1(n5564), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5567) );
  NAND2_X1 U7067 ( .A1(n5566), .A2(n5565), .ZN(n5584) );
  AND2_X1 U7068 ( .A1(n5567), .A2(n5584), .ZN(n7400) );
  AOI22_X1 U7069 ( .A1(n5673), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6545), .B2(
        n7400), .ZN(n5568) );
  NAND2_X1 U7070 ( .A1(n8897), .A2(n5817), .ZN(n5578) );
  NAND2_X1 U7071 ( .A1(n5325), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5576) );
  INV_X1 U7072 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n5570) );
  OR2_X1 U7073 ( .A1(n8832), .A2(n5570), .ZN(n5575) );
  AND2_X1 U7074 ( .A1(n5571), .A2(n7409), .ZN(n5572) );
  OR2_X1 U7075 ( .A1(n5572), .A2(n5589), .ZN(n7697) );
  OR2_X1 U7076 ( .A1(n5856), .A2(n7697), .ZN(n5574) );
  INV_X1 U7077 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7562) );
  OR2_X1 U7078 ( .A1(n6526), .A2(n7562), .ZN(n5573) );
  NAND4_X1 U7079 ( .A1(n5576), .A2(n5575), .A3(n5574), .A4(n5573), .ZN(n9132)
         );
  NAND2_X1 U7080 ( .A1(n9132), .A2(n5816), .ZN(n5577) );
  NAND2_X1 U7081 ( .A1(n5578), .A2(n5577), .ZN(n5579) );
  XNOR2_X1 U7082 ( .A(n5579), .B(n7043), .ZN(n7690) );
  NAND2_X1 U7083 ( .A1(n8897), .A2(n5816), .ZN(n5581) );
  NAND2_X1 U7084 ( .A1(n9132), .A2(n5278), .ZN(n5580) );
  NAND2_X1 U7085 ( .A1(n5581), .A2(n5580), .ZN(n5597) );
  AND2_X1 U7086 ( .A1(n7690), .A2(n5597), .ZN(n5623) );
  XNOR2_X1 U7087 ( .A(n5583), .B(n5582), .ZN(n6814) );
  NAND2_X1 U7088 ( .A1(n6814), .A2(n8866), .ZN(n5587) );
  NAND2_X1 U7089 ( .A1(n5584), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5585) );
  XNOR2_X1 U7090 ( .A(n5585), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10117) );
  AOI22_X1 U7091 ( .A1(n5673), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6545), .B2(
        n10117), .ZN(n5586) );
  NAND2_X1 U7092 ( .A1(n7804), .A2(n5817), .ZN(n5595) );
  NAND2_X1 U7093 ( .A1(n5325), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5593) );
  INV_X1 U7094 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7751) );
  OR2_X1 U7095 ( .A1(n6526), .A2(n7751), .ZN(n5592) );
  INV_X1 U7096 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n5588) );
  OR2_X1 U7097 ( .A1(n8832), .A2(n5588), .ZN(n5591) );
  OAI21_X1 U7098 ( .B1(n5589), .B2(P1_REG3_REG_15__SCAN_IN), .A(n5607), .ZN(
        n7802) );
  OR2_X1 U7099 ( .A1(n5856), .A2(n7802), .ZN(n5590) );
  NAND4_X1 U7100 ( .A1(n5593), .A2(n5592), .A3(n5591), .A4(n5590), .ZN(n9131)
         );
  NAND2_X1 U7101 ( .A1(n9131), .A2(n5816), .ZN(n5594) );
  NAND2_X1 U7102 ( .A1(n5595), .A2(n5594), .ZN(n5596) );
  XNOR2_X1 U7103 ( .A(n5596), .B(n7043), .ZN(n5622) );
  INV_X1 U7104 ( .A(n7690), .ZN(n5598) );
  INV_X1 U7105 ( .A(n5597), .ZN(n7689) );
  NAND2_X1 U7106 ( .A1(n5598), .A2(n7689), .ZN(n5621) );
  XNOR2_X1 U7107 ( .A(n5600), .B(n5599), .ZN(n6882) );
  NAND2_X1 U7108 ( .A1(n6882), .A2(n8866), .ZN(n5605) );
  NOR2_X1 U7109 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5601) );
  NAND2_X1 U7110 ( .A1(n5602), .A2(n5601), .ZN(n5634) );
  NAND2_X1 U7111 ( .A1(n5634), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5603) );
  XNOR2_X1 U7112 ( .A(n5603), .B(P1_IR_REG_16__SCAN_IN), .ZN(n10128) );
  AOI22_X1 U7113 ( .A1(n5673), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6545), .B2(
        n10128), .ZN(n5604) );
  NAND2_X1 U7114 ( .A1(n9507), .A2(n5817), .ZN(n5615) );
  NAND2_X1 U7115 ( .A1(n5853), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5613) );
  INV_X1 U7116 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n5606) );
  OR2_X1 U7117 ( .A1(n5855), .A2(n5606), .ZN(n5612) );
  AND2_X1 U7118 ( .A1(n5607), .A2(n7813), .ZN(n5608) );
  OR2_X1 U7119 ( .A1(n5608), .A2(n5638), .ZN(n7712) );
  OR2_X1 U7120 ( .A1(n5856), .A2(n7712), .ZN(n5611) );
  INV_X1 U7121 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n5609) );
  OR2_X1 U7122 ( .A1(n6526), .A2(n5609), .ZN(n5610) );
  OR2_X1 U7123 ( .A1(n7747), .A2(n4487), .ZN(n5614) );
  NAND2_X1 U7124 ( .A1(n5615), .A2(n5614), .ZN(n5616) );
  XNOR2_X1 U7125 ( .A(n5616), .B(n5749), .ZN(n5619) );
  NOR2_X1 U7126 ( .A1(n7747), .A2(n5812), .ZN(n5617) );
  AOI21_X1 U7127 ( .B1(n9507), .B2(n5816), .A(n5617), .ZN(n5618) );
  NAND2_X1 U7128 ( .A1(n5619), .A2(n5618), .ZN(n5631) );
  OR2_X1 U7129 ( .A1(n5619), .A2(n5618), .ZN(n5620) );
  AND2_X1 U7130 ( .A1(n5631), .A2(n5620), .ZN(n7808) );
  AND2_X1 U7131 ( .A1(n7809), .A2(n7808), .ZN(n5630) );
  NAND2_X1 U7132 ( .A1(n7692), .A2(n5621), .ZN(n5627) );
  INV_X1 U7133 ( .A(n5622), .ZN(n5625) );
  INV_X1 U7134 ( .A(n5623), .ZN(n5624) );
  AND2_X1 U7135 ( .A1(n5625), .A2(n5624), .ZN(n5626) );
  NAND2_X1 U7136 ( .A1(n5627), .A2(n5626), .ZN(n7797) );
  NAND2_X1 U7137 ( .A1(n7804), .A2(n5816), .ZN(n5629) );
  NAND2_X1 U7138 ( .A1(n9131), .A2(n5278), .ZN(n5628) );
  NAND2_X1 U7139 ( .A1(n5629), .A2(n5628), .ZN(n7799) );
  NAND2_X1 U7140 ( .A1(n7797), .A2(n7799), .ZN(n7810) );
  NAND2_X1 U7141 ( .A1(n5630), .A2(n7810), .ZN(n7807) );
  NAND2_X1 U7142 ( .A1(n7807), .A2(n5631), .ZN(n8746) );
  NAND2_X1 U7143 ( .A1(n6885), .A2(n8866), .ZN(n5637) );
  OR2_X1 U7144 ( .A1(n5634), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U7145 ( .A1(n5635), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5670) );
  XNOR2_X1 U7146 ( .A(n5670), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9177) );
  AOI22_X1 U7147 ( .A1(n5673), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6545), .B2(
        n9177), .ZN(n5636) );
  NAND2_X1 U7148 ( .A1(n9500), .A2(n5817), .ZN(n5646) );
  NAND2_X1 U7149 ( .A1(n5325), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5644) );
  INV_X1 U7150 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9185) );
  OR2_X1 U7151 ( .A1(n8832), .A2(n9185), .ZN(n5643) );
  OR2_X1 U7152 ( .A1(n5638), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5639) );
  NAND2_X1 U7153 ( .A1(n5677), .A2(n5639), .ZN(n9415) );
  OR2_X1 U7154 ( .A1(n5856), .A2(n9415), .ZN(n5642) );
  INV_X1 U7155 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n5640) );
  OR2_X1 U7156 ( .A1(n6526), .A2(n5640), .ZN(n5641) );
  NAND4_X1 U7157 ( .A1(n5644), .A2(n5643), .A3(n5642), .A4(n5641), .ZN(n9130)
         );
  NAND2_X1 U7158 ( .A1(n9130), .A2(n5816), .ZN(n5645) );
  NAND2_X1 U7159 ( .A1(n5646), .A2(n5645), .ZN(n5647) );
  XNOR2_X1 U7160 ( .A(n5647), .B(n7043), .ZN(n5649) );
  AND2_X1 U7161 ( .A1(n9130), .A2(n5278), .ZN(n5648) );
  AOI21_X1 U7162 ( .B1(n9500), .B2(n5816), .A(n5648), .ZN(n5650) );
  XNOR2_X1 U7163 ( .A(n5649), .B(n5650), .ZN(n8747) );
  INV_X1 U7164 ( .A(n5649), .ZN(n5651) );
  NAND2_X1 U7165 ( .A1(n5651), .A2(n5650), .ZN(n5652) );
  XNOR2_X1 U7166 ( .A(n5654), .B(n5653), .ZN(n7054) );
  NAND2_X1 U7167 ( .A1(n7054), .A2(n8866), .ZN(n5656) );
  INV_X1 U7168 ( .A(n9332), .ZN(n10206) );
  AOI22_X1 U7169 ( .A1(n5673), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10206), 
        .B2(n6545), .ZN(n5655) );
  NAND2_X1 U7170 ( .A1(n9491), .A2(n5817), .ZN(n5664) );
  AND2_X1 U7171 ( .A1(n5679), .A2(n5657), .ZN(n5658) );
  OR2_X1 U7172 ( .A1(n5658), .A2(n5699), .ZN(n9401) );
  OR2_X1 U7173 ( .A1(n5856), .A2(n9401), .ZN(n5662) );
  NAND2_X1 U7174 ( .A1(n5325), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5661) );
  INV_X1 U7175 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9187) );
  OR2_X1 U7176 ( .A1(n8832), .A2(n9187), .ZN(n5660) );
  INV_X1 U7177 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9402) );
  OR2_X1 U7178 ( .A1(n6526), .A2(n9402), .ZN(n5659) );
  NAND4_X1 U7179 ( .A1(n5662), .A2(n5661), .A3(n5660), .A4(n5659), .ZN(n9203)
         );
  NAND2_X1 U7180 ( .A1(n9203), .A2(n5816), .ZN(n5663) );
  NAND2_X1 U7181 ( .A1(n5664), .A2(n5663), .ZN(n5665) );
  XNOR2_X1 U7182 ( .A(n5665), .B(n7043), .ZN(n5689) );
  NAND2_X1 U7183 ( .A1(n9491), .A2(n5816), .ZN(n5667) );
  NAND2_X1 U7184 ( .A1(n9203), .A2(n5278), .ZN(n5666) );
  NAND2_X1 U7185 ( .A1(n5667), .A2(n5666), .ZN(n5690) );
  NAND2_X1 U7186 ( .A1(n5689), .A2(n5690), .ZN(n8723) );
  XNOR2_X1 U7187 ( .A(n5669), .B(n5668), .ZN(n6975) );
  NAND2_X1 U7188 ( .A1(n6975), .A2(n8866), .ZN(n5675) );
  INV_X1 U7189 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9907) );
  NAND2_X1 U7190 ( .A1(n5670), .A2(n9907), .ZN(n5671) );
  NAND2_X1 U7191 ( .A1(n5671), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5672) );
  XNOR2_X1 U7192 ( .A(n5672), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9176) );
  AOI22_X1 U7193 ( .A1(n6545), .A2(n9176), .B1(n5673), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U7194 ( .A1(n8796), .A2(n5817), .ZN(n5685) );
  NAND2_X1 U7195 ( .A1(n5325), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5683) );
  INV_X1 U7196 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9186) );
  OR2_X1 U7197 ( .A1(n8832), .A2(n9186), .ZN(n5682) );
  NAND2_X1 U7198 ( .A1(n5677), .A2(n5676), .ZN(n5678) );
  NAND2_X1 U7199 ( .A1(n5679), .A2(n5678), .ZN(n8803) );
  OR2_X1 U7200 ( .A1(n5856), .A2(n8803), .ZN(n5681) );
  INV_X1 U7201 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9174) );
  OR2_X1 U7202 ( .A1(n6526), .A2(n9174), .ZN(n5680) );
  OR2_X1 U7203 ( .A1(n9411), .A2(n4487), .ZN(n5684) );
  NAND2_X1 U7204 ( .A1(n5685), .A2(n5684), .ZN(n5686) );
  XNOR2_X1 U7205 ( .A(n5686), .B(n5749), .ZN(n8720) );
  NOR2_X1 U7206 ( .A1(n9411), .A2(n5812), .ZN(n5687) );
  AOI21_X1 U7207 ( .B1(n8796), .B2(n5816), .A(n5687), .ZN(n8719) );
  NAND3_X1 U7208 ( .A1(n8723), .A2(n8719), .A3(n8720), .ZN(n5693) );
  INV_X1 U7209 ( .A(n5689), .ZN(n5692) );
  INV_X1 U7210 ( .A(n5690), .ZN(n5691) );
  NAND2_X1 U7211 ( .A1(n5692), .A2(n5691), .ZN(n8722) );
  AND2_X1 U7212 ( .A1(n5693), .A2(n8722), .ZN(n5694) );
  XNOR2_X1 U7213 ( .A(n5696), .B(n5695), .ZN(n7259) );
  NAND2_X1 U7214 ( .A1(n7259), .A2(n8866), .ZN(n5698) );
  OR2_X1 U7215 ( .A1(n4484), .A2(n7280), .ZN(n5697) );
  NAND2_X1 U7216 ( .A1(n9486), .A2(n5817), .ZN(n5706) );
  NOR2_X1 U7217 ( .A1(n5699), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5700) );
  OR2_X1 U7218 ( .A1(n5718), .A2(n5700), .ZN(n9388) );
  OR2_X1 U7219 ( .A1(n9388), .A2(n5856), .ZN(n5704) );
  NAND2_X1 U7220 ( .A1(n5325), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U7221 ( .A1(n5853), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5702) );
  INV_X1 U7222 ( .A(n6526), .ZN(n8828) );
  NAND2_X1 U7223 ( .A1(n8828), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5701) );
  NAND4_X1 U7224 ( .A1(n5704), .A2(n5703), .A3(n5702), .A4(n5701), .ZN(n9206)
         );
  NAND2_X1 U7225 ( .A1(n9206), .A2(n5816), .ZN(n5705) );
  NAND2_X1 U7226 ( .A1(n5706), .A2(n5705), .ZN(n5707) );
  XNOR2_X1 U7227 ( .A(n5707), .B(n7043), .ZN(n5710) );
  NAND2_X1 U7228 ( .A1(n9486), .A2(n5816), .ZN(n5709) );
  NAND2_X1 U7229 ( .A1(n9206), .A2(n5278), .ZN(n5708) );
  NAND2_X1 U7230 ( .A1(n5709), .A2(n5708), .ZN(n5711) );
  NAND2_X1 U7231 ( .A1(n5710), .A2(n5711), .ZN(n8765) );
  NAND2_X1 U7232 ( .A1(n8764), .A2(n8765), .ZN(n8763) );
  INV_X1 U7233 ( .A(n5710), .ZN(n5713) );
  INV_X1 U7234 ( .A(n5711), .ZN(n5712) );
  NAND2_X1 U7235 ( .A1(n5713), .A2(n5712), .ZN(n8767) );
  XNOR2_X1 U7236 ( .A(n5715), .B(n5714), .ZN(n7281) );
  NAND2_X1 U7237 ( .A1(n7281), .A2(n8866), .ZN(n5717) );
  INV_X1 U7238 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n9702) );
  OR2_X1 U7239 ( .A1(n4485), .A2(n9702), .ZN(n5716) );
  NAND2_X1 U7240 ( .A1(n9481), .A2(n5817), .ZN(n5726) );
  NOR2_X1 U7241 ( .A1(n5718), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5719) );
  OR2_X1 U7242 ( .A1(n5737), .A2(n5719), .ZN(n9373) );
  NAND2_X1 U7243 ( .A1(n8828), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5720) );
  OAI21_X1 U7244 ( .B1(n9373), .B2(n5856), .A(n5720), .ZN(n5724) );
  INV_X1 U7245 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5722) );
  NAND2_X1 U7246 ( .A1(n5325), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5721) );
  OAI21_X1 U7247 ( .B1(n5722), .B2(n8832), .A(n5721), .ZN(n5723) );
  NAND2_X1 U7248 ( .A1(n9361), .A2(n5816), .ZN(n5725) );
  NAND2_X1 U7249 ( .A1(n5726), .A2(n5725), .ZN(n5727) );
  XNOR2_X1 U7250 ( .A(n5727), .B(n7043), .ZN(n5729) );
  AND2_X1 U7251 ( .A1(n9361), .A2(n5278), .ZN(n5728) );
  AOI21_X1 U7252 ( .B1(n9481), .B2(n5816), .A(n5728), .ZN(n5730) );
  XNOR2_X1 U7253 ( .A(n5729), .B(n5730), .ZN(n8731) );
  INV_X1 U7254 ( .A(n5729), .ZN(n5731) );
  AND2_X1 U7255 ( .A1(n5731), .A2(n5730), .ZN(n5732) );
  AOI21_X1 U7256 ( .B1(n8732), .B2(n8731), .A(n5732), .ZN(n5751) );
  XNOR2_X1 U7257 ( .A(n5734), .B(n5733), .ZN(n7372) );
  NAND2_X1 U7258 ( .A1(n7372), .A2(n8866), .ZN(n5736) );
  OR2_X1 U7259 ( .A1(n4484), .A2(n7373), .ZN(n5735) );
  OR2_X1 U7260 ( .A1(n9358), .A2(n4487), .ZN(n5748) );
  OR2_X1 U7261 ( .A1(n5737), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5739) );
  AND2_X1 U7262 ( .A1(n5739), .A2(n5738), .ZN(n9356) );
  NAND2_X1 U7263 ( .A1(n9356), .A2(n5740), .ZN(n5746) );
  INV_X1 U7264 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5743) );
  NAND2_X1 U7265 ( .A1(n8828), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5742) );
  NAND2_X1 U7266 ( .A1(n5325), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5741) );
  OAI211_X1 U7267 ( .C1(n8832), .C2(n5743), .A(n5742), .B(n5741), .ZN(n5744)
         );
  INV_X1 U7268 ( .A(n5744), .ZN(n5745) );
  OR2_X1 U7269 ( .A1(n9371), .A2(n5812), .ZN(n5747) );
  NAND2_X1 U7270 ( .A1(n5748), .A2(n5747), .ZN(n5752) );
  NAND2_X1 U7271 ( .A1(n5751), .A2(n5752), .ZN(n8779) );
  OAI22_X1 U7272 ( .A1(n9358), .A2(n5767), .B1(n9371), .B2(n4487), .ZN(n5750)
         );
  XNOR2_X1 U7273 ( .A(n5750), .B(n5749), .ZN(n8777) );
  NAND2_X1 U7274 ( .A1(n8779), .A2(n8777), .ZN(n8776) );
  INV_X1 U7275 ( .A(n5751), .ZN(n5754) );
  INV_X1 U7276 ( .A(n5752), .ZN(n5753) );
  NAND2_X1 U7277 ( .A1(n5754), .A2(n5753), .ZN(n8778) );
  NAND2_X1 U7278 ( .A1(n7435), .A2(n8866), .ZN(n5758) );
  OR2_X1 U7279 ( .A1(n4485), .A2(n7434), .ZN(n5757) );
  NAND2_X1 U7280 ( .A1(n5853), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5766) );
  INV_X1 U7281 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n5759) );
  OR2_X1 U7282 ( .A1(n5855), .A2(n5759), .ZN(n5765) );
  OAI21_X1 U7283 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n5761), .A(n5760), .ZN(
        n9342) );
  OR2_X1 U7284 ( .A1(n5856), .A2(n9342), .ZN(n5764) );
  INV_X1 U7285 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n5762) );
  OR2_X1 U7286 ( .A1(n6526), .A2(n5762), .ZN(n5763) );
  NAND4_X1 U7287 ( .A1(n5766), .A2(n5765), .A3(n5764), .A4(n5763), .ZN(n9362)
         );
  OAI22_X1 U7288 ( .A1(n9345), .A2(n5767), .B1(n8836), .B2(n4487), .ZN(n5768)
         );
  XOR2_X1 U7289 ( .A(n7043), .B(n5768), .Z(n5769) );
  OAI22_X1 U7290 ( .A1(n9345), .A2(n4487), .B1(n8836), .B2(n5812), .ZN(n8712)
         );
  XOR2_X1 U7291 ( .A(n5771), .B(n5770), .Z(n8755) );
  XNOR2_X1 U7292 ( .A(n5775), .B(n5774), .ZN(n7629) );
  NAND2_X1 U7293 ( .A1(n7629), .A2(n8866), .ZN(n5777) );
  OR2_X1 U7294 ( .A1(n4485), .A2(n9859), .ZN(n5776) );
  INV_X1 U7295 ( .A(n9305), .ZN(n9306) );
  NAND2_X1 U7296 ( .A1(n5325), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5786) );
  INV_X1 U7297 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9308) );
  OR2_X1 U7298 ( .A1(n6526), .A2(n9308), .ZN(n5785) );
  INV_X1 U7299 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5778) );
  NAND2_X1 U7300 ( .A1(n5779), .A2(n5778), .ZN(n5780) );
  NAND2_X1 U7301 ( .A1(n5781), .A2(n5780), .ZN(n9307) );
  OR2_X1 U7302 ( .A1(n5856), .A2(n9307), .ZN(n5784) );
  INV_X1 U7303 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n5782) );
  OR2_X1 U7304 ( .A1(n8832), .A2(n5782), .ZN(n5783) );
  OAI22_X1 U7305 ( .A1(n9306), .A2(n4487), .B1(n9218), .B2(n5812), .ZN(n5791)
         );
  NAND2_X1 U7306 ( .A1(n9305), .A2(n5817), .ZN(n5788) );
  OR2_X1 U7307 ( .A1(n9218), .A2(n4487), .ZN(n5787) );
  NAND2_X1 U7308 ( .A1(n5788), .A2(n5787), .ZN(n5789) );
  XNOR2_X1 U7309 ( .A(n5789), .B(n7043), .ZN(n5790) );
  XOR2_X1 U7310 ( .A(n5791), .B(n5790), .Z(n8739) );
  INV_X1 U7311 ( .A(n5790), .ZN(n5793) );
  INV_X1 U7312 ( .A(n5791), .ZN(n5792) );
  XNOR2_X1 U7313 ( .A(n5794), .B(n5795), .ZN(n8814) );
  NAND2_X1 U7314 ( .A1(n5797), .A2(n5796), .ZN(n5799) );
  MUX2_X1 U7315 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7875), .Z(n6277) );
  INV_X1 U7316 ( .A(SI_28_), .ZN(n9681) );
  XNOR2_X1 U7317 ( .A(n6277), .B(n9681), .ZN(n6275) );
  NAND2_X1 U7318 ( .A1(n8149), .A2(n8866), .ZN(n5801) );
  INV_X1 U7319 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9878) );
  OR2_X1 U7320 ( .A1(n4484), .A2(n9878), .ZN(n5800) );
  NAND2_X1 U7321 ( .A1(n9444), .A2(n5816), .ZN(n5814) );
  NAND2_X1 U7322 ( .A1(n5853), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5811) );
  INV_X1 U7323 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n5802) );
  OR2_X1 U7324 ( .A1(n5855), .A2(n5802), .ZN(n5810) );
  INV_X1 U7325 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5803) );
  OAI21_X1 U7326 ( .B1(n5804), .B2(n8705), .A(n5803), .ZN(n5807) );
  INV_X1 U7327 ( .A(n5804), .ZN(n5806) );
  AND2_X1 U7328 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5805) );
  NAND2_X1 U7329 ( .A1(n5806), .A2(n5805), .ZN(n9252) );
  NAND2_X1 U7330 ( .A1(n5807), .A2(n9252), .ZN(n9262) );
  OR2_X1 U7331 ( .A1(n5856), .A2(n9262), .ZN(n5809) );
  INV_X1 U7332 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9263) );
  OR2_X1 U7333 ( .A1(n6526), .A2(n9263), .ZN(n5808) );
  OR2_X1 U7334 ( .A1(n5812), .A2(n9275), .ZN(n5813) );
  NAND2_X1 U7335 ( .A1(n5814), .A2(n5813), .ZN(n5815) );
  XNOR2_X1 U7336 ( .A(n5815), .B(n7043), .ZN(n5819) );
  INV_X1 U7337 ( .A(n9275), .ZN(n9248) );
  AOI22_X1 U7338 ( .A1(n9444), .A2(n5817), .B1(n5816), .B2(n9248), .ZN(n5818)
         );
  XNOR2_X1 U7339 ( .A(n5819), .B(n5818), .ZN(n5873) );
  INV_X1 U7340 ( .A(n5873), .ZN(n5844) );
  INV_X1 U7341 ( .A(n5820), .ZN(n7553) );
  INV_X1 U7342 ( .A(n7764), .ZN(n5823) );
  INV_X1 U7343 ( .A(n5821), .ZN(n7632) );
  NAND3_X1 U7344 ( .A1(n7632), .A2(P1_B_REG_SCAN_IN), .A3(n7553), .ZN(n5822)
         );
  OAI211_X1 U7345 ( .C1(P1_B_REG_SCAN_IN), .C2(n7553), .A(n5823), .B(n5822), 
        .ZN(n6608) );
  OR2_X1 U7346 ( .A1(n6608), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5824) );
  NAND2_X1 U7347 ( .A1(n7764), .A2(n7632), .ZN(n6519) );
  NAND2_X1 U7348 ( .A1(n5824), .A2(n6519), .ZN(n6939) );
  NOR4_X1 U7349 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5828) );
  NOR4_X1 U7350 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5827) );
  NOR4_X1 U7351 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5826) );
  NOR4_X1 U7352 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5825) );
  AND4_X1 U7353 ( .A1(n5828), .A2(n5827), .A3(n5826), .A4(n5825), .ZN(n5834)
         );
  NOR2_X1 U7354 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n5832) );
  NOR4_X1 U7355 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5831) );
  NOR4_X1 U7356 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5830) );
  NOR4_X1 U7357 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5829) );
  AND4_X1 U7358 ( .A1(n5832), .A2(n5831), .A3(n5830), .A4(n5829), .ZN(n5833)
         );
  NAND2_X1 U7359 ( .A1(n5834), .A2(n5833), .ZN(n6605) );
  INV_X1 U7360 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9688) );
  NOR2_X1 U7361 ( .A1(n6605), .A2(n9688), .ZN(n5835) );
  OR2_X1 U7362 ( .A1(n6608), .A2(n5835), .ZN(n5836) );
  NAND2_X1 U7363 ( .A1(n7764), .A2(n7553), .ZN(n9551) );
  NAND2_X1 U7364 ( .A1(n5836), .A2(n9551), .ZN(n6618) );
  NOR2_X1 U7365 ( .A1(n6939), .A2(n6618), .ZN(n5847) );
  INV_X1 U7366 ( .A(n5837), .ZN(n5838) );
  NAND2_X1 U7367 ( .A1(n5838), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5840) );
  XNOR2_X1 U7368 ( .A(n5840), .B(n5839), .ZN(n7432) );
  AND2_X1 U7369 ( .A1(n7432), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5841) );
  AND2_X1 U7370 ( .A1(n5847), .A2(n9122), .ZN(n5849) );
  INV_X1 U7371 ( .A(n5849), .ZN(n5843) );
  NAND2_X1 U7372 ( .A1(n8938), .A2(n9076), .ZN(n6614) );
  NAND2_X1 U7373 ( .A1(n9125), .A2(n6927), .ZN(n9067) );
  NAND2_X1 U7374 ( .A1(n10304), .A2(n9067), .ZN(n5842) );
  NAND2_X1 U7375 ( .A1(n5844), .A2(n8812), .ZN(n5878) );
  NAND2_X1 U7376 ( .A1(n8702), .A2(n5845), .ZN(n5872) );
  AND2_X1 U7377 ( .A1(n5873), .A2(n5065), .ZN(n5846) );
  NAND2_X1 U7378 ( .A1(n5879), .A2(n5846), .ZN(n5877) );
  NOR2_X1 U7379 ( .A1(n6614), .A2(n9437), .ZN(n10201) );
  INV_X1 U7380 ( .A(n5847), .ZN(n5864) );
  NAND3_X1 U7381 ( .A1(n10201), .A2(n9122), .A3(n5864), .ZN(n5867) );
  OR2_X1 U7382 ( .A1(n9067), .A2(n9116), .ZN(n5862) );
  NAND2_X1 U7383 ( .A1(n9122), .A2(n5862), .ZN(n6619) );
  INV_X1 U7384 ( .A(n6619), .ZN(n5848) );
  AND2_X1 U7385 ( .A1(n5867), .A2(n5848), .ZN(n8795) );
  OR2_X1 U7386 ( .A1(n6936), .A2(n6922), .ZN(n7044) );
  INV_X1 U7387 ( .A(n7044), .ZN(n9121) );
  AND2_X1 U7388 ( .A1(n5849), .A2(n9121), .ZN(n5851) );
  INV_X1 U7389 ( .A(n5850), .ZN(n10049) );
  NAND2_X1 U7390 ( .A1(n5851), .A2(n10049), .ZN(n8819) );
  INV_X1 U7391 ( .A(n5851), .ZN(n5852) );
  OR2_X1 U7392 ( .A1(n5852), .A2(n10049), .ZN(n8805) );
  INV_X2 U7393 ( .A(n8805), .ZN(n8817) );
  NAND2_X1 U7394 ( .A1(n5853), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5861) );
  INV_X1 U7395 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5854) );
  OR2_X1 U7396 ( .A1(n5855), .A2(n5854), .ZN(n5860) );
  OR2_X1 U7397 ( .A1(n5856), .A2(n9252), .ZN(n5859) );
  INV_X1 U7398 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n5857) );
  OR2_X1 U7399 ( .A1(n6526), .A2(n5857), .ZN(n5858) );
  INV_X1 U7400 ( .A(n9258), .ZN(n9129) );
  AOI22_X1 U7401 ( .A1(n8817), .A2(n9129), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n5871) );
  AND3_X1 U7402 ( .A1(n5863), .A2(n7432), .A3(n5862), .ZN(n5865) );
  NAND2_X1 U7403 ( .A1(n5864), .A2(n10304), .ZN(n6629) );
  NAND2_X1 U7404 ( .A1(n5865), .A2(n6629), .ZN(n5866) );
  NAND2_X1 U7405 ( .A1(n5866), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5868) );
  INV_X1 U7406 ( .A(n8804), .ZN(n8821) );
  INV_X1 U7407 ( .A(n9262), .ZN(n5869) );
  NAND2_X1 U7408 ( .A1(n8821), .A2(n5869), .ZN(n5870) );
  OAI211_X1 U7409 ( .C1(n9259), .C2(n8819), .A(n5871), .B(n5870), .ZN(n5875)
         );
  NOR3_X1 U7410 ( .A1(n5873), .A2(n8773), .A3(n5872), .ZN(n5874) );
  AOI211_X1 U7411 ( .C1(n8791), .C2(n9444), .A(n5875), .B(n5874), .ZN(n5876)
         );
  OAI211_X1 U7412 ( .C1(n5879), .C2(n5878), .A(n5877), .B(n5876), .ZN(P1_U3218) );
  NOR2_X2 U7413 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5943) );
  NOR2_X1 U7414 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5883) );
  NAND3_X1 U7415 ( .A1(n4523), .A2(n5995), .A3(n5885), .ZN(n5928) );
  NOR2_X1 U7416 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5889) );
  NOR2_X1 U7417 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5888) );
  NOR2_X1 U7418 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5887) );
  NOR2_X1 U7419 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5886) );
  INV_X1 U7420 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5890) );
  INV_X1 U7421 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5891) );
  INV_X1 U7422 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5893) );
  NAND2_X2 U7423 ( .A1(n5896), .A2(n5946), .ZN(n6043) );
  NAND2_X1 U7424 ( .A1(n7549), .A2(n7885), .ZN(n5898) );
  NAND2_X4 U7425 ( .A1(n5946), .A2(n7875), .ZN(n7886) );
  INV_X1 U7426 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7550) );
  OR2_X1 U7427 ( .A1(n7886), .A2(n7550), .ZN(n5897) );
  NAND3_X1 U7428 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n6009) );
  INV_X1 U7429 ( .A(n6009), .ZN(n5899) );
  INV_X1 U7430 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n6090) );
  INV_X1 U7431 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9929) );
  INV_X1 U7432 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9926) );
  INV_X1 U7433 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9871) );
  INV_X1 U7434 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9900) );
  INV_X1 U7435 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n7904) );
  NAND2_X1 U7436 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(P2_REG3_REG_24__SCAN_IN), 
        .ZN(n5909) );
  INV_X1 U7437 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9903) );
  INV_X1 U7438 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5910) );
  OAI21_X1 U7439 ( .B1(n6222), .B2(n9903), .A(n5910), .ZN(n5911) );
  AND2_X1 U7440 ( .A1(n6233), .A2(n5911), .ZN(n8430) );
  INV_X1 U7441 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5913) );
  INV_X1 U7442 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5914) );
  INV_X1 U7443 ( .A(n5921), .ZN(n5920) );
  INV_X1 U7444 ( .A(n4488), .ZN(n6262) );
  NAND2_X4 U7445 ( .A1(n5920), .A2(n7912), .ZN(n5962) );
  INV_X1 U7446 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n5926) );
  NAND2_X1 U7447 ( .A1(n5950), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5925) );
  NAND2_X1 U7448 ( .A1(n5923), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5924) );
  OAI211_X1 U7449 ( .C1(n5962), .C2(n5926), .A(n5925), .B(n5924), .ZN(n5927)
         );
  AOI21_X1 U7450 ( .B1(n8430), .B2(n6262), .A(n5927), .ZN(n8210) );
  NAND2_X1 U7451 ( .A1(n7054), .A2(n7885), .ZN(n5930) );
  INV_X2 U7452 ( .A(n7886), .ZN(n5996) );
  BUF_X1 U7453 ( .A(n5928), .Z(n6158) );
  AOI22_X1 U7454 ( .A1(n5996), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n10367), 
        .B2(n6538), .ZN(n5929) );
  INV_X1 U7455 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U7456 ( .A1(n6186), .A2(n5931), .ZN(n5932) );
  NAND2_X1 U7457 ( .A1(n6194), .A2(n5932), .ZN(n8523) );
  OR2_X1 U7458 ( .A1(n8523), .A2(n4488), .ZN(n5937) );
  INV_X1 U7459 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8616) );
  NAND2_X1 U7460 ( .A1(n6353), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5934) );
  NAND2_X1 U7461 ( .A1(n5950), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5933) );
  OAI211_X1 U7462 ( .C1(n8616), .C2(n6016), .A(n5934), .B(n5933), .ZN(n5935)
         );
  INV_X1 U7463 ( .A(n5935), .ZN(n5936) );
  INV_X1 U7464 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6662) );
  INV_X1 U7465 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9841) );
  OR2_X1 U7466 ( .A1(n5974), .A2(n9841), .ZN(n5941) );
  NAND2_X1 U7467 ( .A1(n5950), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5940) );
  INV_X1 U7468 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n5938) );
  INV_X1 U7469 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6515) );
  OR2_X1 U7470 ( .A1(n7886), .A2(n6515), .ZN(n5949) );
  OR2_X1 U7471 ( .A1(n6043), .A2(n6514), .ZN(n5948) );
  NAND2_X1 U7472 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5942) );
  MUX2_X1 U7473 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5942), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5945) );
  INV_X1 U7474 ( .A(n5943), .ZN(n5944) );
  OR2_X1 U7475 ( .A1(n5946), .A2(n9981), .ZN(n5947) );
  OR2_X2 U7476 ( .A1(n8261), .A2(n7903), .ZN(n7938) );
  INV_X1 U7477 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5951) );
  OR2_X1 U7478 ( .A1(n5973), .A2(n5951), .ZN(n5957) );
  INV_X1 U7479 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5952) );
  INV_X1 U7480 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5953) );
  OR2_X1 U7481 ( .A1(n5962), .A2(n5953), .ZN(n5955) );
  INV_X1 U7482 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9752) );
  OR2_X1 U7483 ( .A1(n5974), .A2(n9752), .ZN(n5954) );
  INV_X1 U7484 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10335) );
  INV_X1 U7485 ( .A(SI_0_), .ZN(n5958) );
  OR2_X1 U7486 ( .A1(n7875), .A2(n5958), .ZN(n5960) );
  INV_X1 U7487 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5959) );
  XNOR2_X1 U7488 ( .A(n5960), .B(n5959), .ZN(n8687) );
  MUX2_X1 U7489 ( .A(n10335), .B(n8687), .S(n5946), .Z(n10430) );
  INV_X1 U7490 ( .A(n10430), .ZN(n7119) );
  NAND2_X1 U7491 ( .A1(n8262), .A2(n7119), .ZN(n7097) );
  NAND2_X1 U7492 ( .A1(n7087), .A2(n7097), .ZN(n7096) );
  INV_X1 U7493 ( .A(n7903), .ZN(n7098) );
  OR2_X1 U7494 ( .A1(n8261), .A2(n7098), .ZN(n5961) );
  NAND2_X1 U7495 ( .A1(n7096), .A2(n5961), .ZN(n6740) );
  NAND2_X1 U7496 ( .A1(n5950), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5966) );
  INV_X1 U7497 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9860) );
  OR2_X1 U7498 ( .A1(n5974), .A2(n9860), .ZN(n5965) );
  INV_X1 U7499 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6661) );
  OR2_X1 U7500 ( .A1(n4483), .A2(n6661), .ZN(n5964) );
  INV_X1 U7501 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7101) );
  OR2_X1 U7502 ( .A1(n7886), .A2(n6518), .ZN(n5970) );
  OR2_X1 U7503 ( .A1(n6043), .A2(n6517), .ZN(n5969) );
  OR2_X1 U7504 ( .A1(n5943), .A2(n5917), .ZN(n5967) );
  XNOR2_X1 U7505 ( .A(n5967), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9993) );
  INV_X1 U7506 ( .A(n9993), .ZN(n6516) );
  AND3_X2 U7507 ( .A1(n5970), .A2(n5969), .A3(n5968), .ZN(n6755) );
  OR2_X2 U7508 ( .A1(n5971), .A2(n6755), .ZN(n7937) );
  NAND2_X1 U7509 ( .A1(n5971), .A2(n6755), .ZN(n7940) );
  NAND2_X1 U7510 ( .A1(n6740), .A2(n8099), .ZN(n6739) );
  INV_X1 U7511 ( .A(n6755), .ZN(n7106) );
  OR2_X1 U7512 ( .A1(n5971), .A2(n7106), .ZN(n5972) );
  NAND2_X1 U7513 ( .A1(n6739), .A2(n5972), .ZN(n6854) );
  INV_X2 U7514 ( .A(n5973), .ZN(n6559) );
  NAND2_X1 U7515 ( .A1(n6559), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5979) );
  OR2_X1 U7516 ( .A1(n4488), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5978) );
  INV_X1 U7517 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6660) );
  OR2_X1 U7518 ( .A1(n4483), .A2(n6660), .ZN(n5977) );
  INV_X1 U7519 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5975) );
  OR2_X1 U7520 ( .A1(n5962), .A2(n5975), .ZN(n5976) );
  OR2_X1 U7521 ( .A1(n6043), .A2(n6506), .ZN(n5983) );
  OR2_X1 U7522 ( .A1(n7886), .A2(n4610), .ZN(n5982) );
  NAND2_X1 U7523 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4522), .ZN(n5980) );
  XNOR2_X1 U7524 ( .A(n5980), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6720) );
  INV_X1 U7525 ( .A(n6720), .ZN(n6500) );
  OR2_X1 U7526 ( .A1(n5946), .A2(n6500), .ZN(n5981) );
  NAND2_X1 U7527 ( .A1(n8260), .A2(n6865), .ZN(n7959) );
  NAND2_X1 U7528 ( .A1(n6854), .A2(n7953), .ZN(n6853) );
  OR2_X1 U7529 ( .A1(n8260), .A2(n5984), .ZN(n5986) );
  NAND2_X1 U7530 ( .A1(n6853), .A2(n5986), .ZN(n6818) );
  NAND2_X1 U7531 ( .A1(n6559), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5994) );
  INV_X1 U7532 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6914) );
  NAND2_X1 U7533 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5987) );
  NAND2_X1 U7534 ( .A1(n6914), .A2(n5987), .ZN(n5988) );
  NAND2_X1 U7535 ( .A1(n6009), .A2(n5988), .ZN(n10362) );
  OR2_X1 U7536 ( .A1(n4488), .A2(n10362), .ZN(n5993) );
  INV_X1 U7537 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5989) );
  INV_X1 U7538 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5990) );
  OR2_X1 U7539 ( .A1(n5962), .A2(n5990), .ZN(n5991) );
  OR2_X1 U7540 ( .A1(n6502), .A2(n6043), .ZN(n5998) );
  NAND2_X1 U7541 ( .A1(n5995), .A2(n6021), .ZN(n6047) );
  NAND2_X1 U7542 ( .A1(n6047), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6001) );
  XNOR2_X1 U7543 ( .A(n6001), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6732) );
  AOI22_X1 U7544 ( .A1(n5996), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6538), .B2(
        n6732), .ZN(n5997) );
  AND2_X2 U7545 ( .A1(n5998), .A2(n5997), .ZN(n10437) );
  OR2_X1 U7546 ( .A1(n8258), .A2(n10437), .ZN(n7935) );
  NAND2_X1 U7547 ( .A1(n7935), .A2(n7960), .ZN(n6332) );
  INV_X1 U7548 ( .A(n6026), .ZN(n5999) );
  OR2_X1 U7549 ( .A1(n6332), .A2(n5999), .ZN(n10344) );
  OR2_X1 U7550 ( .A1(n6508), .A2(n6043), .ZN(n6007) );
  INV_X1 U7551 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U7552 ( .A1(n6001), .A2(n6000), .ZN(n6002) );
  NAND2_X1 U7553 ( .A1(n6002), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6004) );
  INV_X1 U7554 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U7555 ( .A1(n6004), .A2(n6003), .ZN(n6032) );
  OR2_X1 U7556 ( .A1(n6004), .A2(n6003), .ZN(n6005) );
  INV_X1 U7557 ( .A(n10347), .ZN(n10444) );
  NAND2_X1 U7558 ( .A1(n6353), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6014) );
  INV_X1 U7559 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n6008) );
  OR2_X1 U7560 ( .A1(n5973), .A2(n6008), .ZN(n6013) );
  INV_X1 U7561 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9848) );
  NAND2_X1 U7562 ( .A1(n6009), .A2(n9848), .ZN(n6010) );
  NAND2_X1 U7563 ( .A1(n6037), .A2(n6010), .ZN(n8228) );
  OR2_X1 U7564 ( .A1(n4488), .A2(n8228), .ZN(n6012) );
  INV_X1 U7565 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6659) );
  OR2_X1 U7566 ( .A1(n4483), .A2(n6659), .ZN(n6011) );
  NAND2_X1 U7567 ( .A1(n6015), .A2(n4509), .ZN(n6027) );
  NAND2_X1 U7568 ( .A1(n6353), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6020) );
  NAND2_X1 U7569 ( .A1(n6559), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6019) );
  XNOR2_X1 U7570 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7110) );
  INV_X1 U7571 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6665) );
  OR2_X1 U7572 ( .A1(n4483), .A2(n6665), .ZN(n6017) );
  NAND4_X1 U7573 ( .A1(n6020), .A2(n6019), .A3(n6018), .A4(n6017), .ZN(n8259)
         );
  OR2_X1 U7574 ( .A1(n6498), .A2(n6043), .ZN(n6025) );
  OR2_X1 U7575 ( .A1(n7886), .A2(n6499), .ZN(n6024) );
  OR2_X1 U7576 ( .A1(n5995), .A2(n5917), .ZN(n6022) );
  XNOR2_X1 U7577 ( .A(n6022), .B(n6021), .ZN(n6666) );
  OR2_X1 U7578 ( .A1(n5946), .A2(n6666), .ZN(n6023) );
  OR2_X1 U7579 ( .A1(n8259), .A2(n6824), .ZN(n7930) );
  NAND2_X1 U7580 ( .A1(n8259), .A2(n6824), .ZN(n7958) );
  NAND2_X1 U7581 ( .A1(n7930), .A2(n7958), .ZN(n8101) );
  NAND3_X1 U7582 ( .A1(n6818), .A2(n6027), .A3(n8101), .ZN(n6029) );
  INV_X1 U7583 ( .A(n6824), .ZN(n7115) );
  OR2_X1 U7584 ( .A1(n8259), .A2(n7115), .ZN(n10355) );
  AND2_X1 U7585 ( .A1(n10355), .A2(n6026), .ZN(n10342) );
  NAND2_X1 U7586 ( .A1(n6027), .A2(n5063), .ZN(n6028) );
  NAND2_X1 U7587 ( .A1(n6029), .A2(n6028), .ZN(n6031) );
  OR2_X1 U7588 ( .A1(n10444), .A2(n7966), .ZN(n6030) );
  NAND2_X1 U7589 ( .A1(n6031), .A2(n6030), .ZN(n6953) );
  OR2_X1 U7590 ( .A1(n6512), .A2(n6043), .ZN(n6035) );
  NAND2_X1 U7591 ( .A1(n6032), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6033) );
  XNOR2_X1 U7592 ( .A(n6033), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6763) );
  AOI22_X1 U7593 ( .A1(n5996), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6538), .B2(
        n6763), .ZN(n6034) );
  NAND2_X1 U7594 ( .A1(n6035), .A2(n6034), .ZN(n7252) );
  NAND2_X1 U7595 ( .A1(n6559), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6042) );
  INV_X1 U7596 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7249) );
  OR2_X1 U7597 ( .A1(n5962), .A2(n7249), .ZN(n6041) );
  INV_X1 U7598 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6036) );
  NAND2_X1 U7599 ( .A1(n6037), .A2(n6036), .ZN(n6038) );
  NAND2_X1 U7600 ( .A1(n6052), .A2(n6038), .ZN(n7248) );
  OR2_X1 U7601 ( .A1(n4488), .A2(n7248), .ZN(n6040) );
  INV_X1 U7602 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6671) );
  OR2_X1 U7603 ( .A1(n6016), .A2(n6671), .ZN(n6039) );
  OR2_X1 U7604 ( .A1(n7252), .A2(n8225), .ZN(n7968) );
  NAND2_X1 U7605 ( .A1(n7252), .A2(n8225), .ZN(n7969) );
  NAND2_X1 U7606 ( .A1(n7968), .A2(n7969), .ZN(n8107) );
  INV_X1 U7607 ( .A(n8107), .ZN(n6954) );
  INV_X1 U7608 ( .A(n8225), .ZN(n8256) );
  INV_X1 U7609 ( .A(n7135), .ZN(n6058) );
  OR2_X1 U7610 ( .A1(n6523), .A2(n6043), .ZN(n6050) );
  NAND2_X1 U7611 ( .A1(n6044), .A2(n6045), .ZN(n6046) );
  NAND2_X1 U7612 ( .A1(n6060), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6048) );
  XNOR2_X1 U7613 ( .A(n6048), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6980) );
  AOI22_X1 U7614 ( .A1(n5996), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6538), .B2(
        n6980), .ZN(n6049) );
  NAND2_X1 U7615 ( .A1(n6050), .A2(n6049), .ZN(n7975) );
  NAND2_X1 U7616 ( .A1(n6353), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6057) );
  INV_X1 U7617 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6051) );
  OR2_X1 U7618 ( .A1(n5973), .A2(n6051), .ZN(n6056) );
  INV_X1 U7619 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9842) );
  NAND2_X1 U7620 ( .A1(n6052), .A2(n9842), .ZN(n6053) );
  NAND2_X1 U7621 ( .A1(n6064), .A2(n6053), .ZN(n7144) );
  OR2_X1 U7622 ( .A1(n4488), .A2(n7144), .ZN(n6055) );
  INV_X1 U7623 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6990) );
  OR2_X1 U7624 ( .A1(n4483), .A2(n6990), .ZN(n6054) );
  NAND4_X1 U7625 ( .A1(n6057), .A2(n6056), .A3(n6055), .A4(n6054), .ZN(n8255)
         );
  NAND2_X1 U7626 ( .A1(n6058), .A2(n4486), .ZN(n7137) );
  NAND2_X1 U7627 ( .A1(n7975), .A2(n8255), .ZN(n6059) );
  NAND2_X1 U7628 ( .A1(n6533), .A2(n7885), .ZN(n6062) );
  NOR2_X1 U7629 ( .A1(n6060), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n6103) );
  OR2_X1 U7630 ( .A1(n6103), .A2(n5917), .ZN(n6071) );
  XNOR2_X1 U7631 ( .A(n6071), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8272) );
  AOI22_X1 U7632 ( .A1(n5996), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6538), .B2(
        n8272), .ZN(n6061) );
  NAND2_X1 U7633 ( .A1(n6062), .A2(n6061), .ZN(n7356) );
  NAND2_X1 U7634 ( .A1(n6559), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6069) );
  INV_X1 U7635 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7350) );
  OR2_X1 U7636 ( .A1(n5962), .A2(n7350), .ZN(n6068) );
  INV_X1 U7637 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U7638 ( .A1(n6064), .A2(n6063), .ZN(n6065) );
  NAND2_X1 U7639 ( .A1(n6075), .A2(n6065), .ZN(n7857) );
  OR2_X1 U7640 ( .A1(n4488), .A2(n7857), .ZN(n6067) );
  INV_X1 U7641 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6986) );
  OR2_X1 U7642 ( .A1(n6016), .A2(n6986), .ZN(n6066) );
  OR2_X1 U7643 ( .A1(n7356), .A2(n7263), .ZN(n7988) );
  AND2_X1 U7644 ( .A1(n7356), .A2(n7263), .ZN(n7979) );
  INV_X1 U7645 ( .A(n7979), .ZN(n7981) );
  INV_X1 U7646 ( .A(n7263), .ZN(n8254) );
  OR2_X1 U7647 ( .A1(n7356), .A2(n8254), .ZN(n6070) );
  INV_X1 U7648 ( .A(n7269), .ZN(n6082) );
  NAND2_X1 U7649 ( .A1(n6552), .A2(n7885), .ZN(n6074) );
  INV_X1 U7650 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U7651 ( .A1(n6071), .A2(n6101), .ZN(n6072) );
  NAND2_X1 U7652 ( .A1(n6072), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6084) );
  XNOR2_X1 U7653 ( .A(n6084), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7188) );
  AOI22_X1 U7654 ( .A1(n5996), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6538), .B2(
        n7188), .ZN(n6073) );
  INV_X1 U7655 ( .A(n7274), .ZN(n10454) );
  NAND2_X1 U7656 ( .A1(n6559), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6080) );
  INV_X1 U7657 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7272) );
  OR2_X1 U7658 ( .A1(n5962), .A2(n7272), .ZN(n6079) );
  NAND2_X1 U7659 ( .A1(n6075), .A2(n9692), .ZN(n6076) );
  NAND2_X1 U7660 ( .A1(n6091), .A2(n6076), .ZN(n7271) );
  OR2_X1 U7661 ( .A1(n4488), .A2(n7271), .ZN(n6078) );
  INV_X1 U7662 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6992) );
  OR2_X1 U7663 ( .A1(n6016), .A2(n6992), .ZN(n6077) );
  INV_X1 U7664 ( .A(n7346), .ZN(n8253) );
  NAND2_X1 U7665 ( .A1(n7274), .A2(n7346), .ZN(n7986) );
  NAND2_X1 U7666 ( .A1(n6082), .A2(n6081), .ZN(n7267) );
  NAND2_X1 U7667 ( .A1(n7274), .A2(n8253), .ZN(n6083) );
  NAND2_X1 U7668 ( .A1(n7267), .A2(n6083), .ZN(n7374) );
  NAND2_X1 U7669 ( .A1(n6555), .A2(n7885), .ZN(n6088) );
  INV_X1 U7670 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6100) );
  NAND2_X1 U7671 ( .A1(n6084), .A2(n6100), .ZN(n6085) );
  NAND2_X1 U7672 ( .A1(n6085), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6086) );
  XNOR2_X1 U7673 ( .A(n6086), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7307) );
  AOI22_X1 U7674 ( .A1(n5996), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6538), .B2(
        n7307), .ZN(n6087) );
  NAND2_X1 U7675 ( .A1(n6088), .A2(n6087), .ZN(n7382) );
  NAND2_X1 U7676 ( .A1(n6559), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6096) );
  INV_X1 U7677 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6089) );
  OR2_X1 U7678 ( .A1(n5962), .A2(n6089), .ZN(n6095) );
  NAND2_X1 U7679 ( .A1(n6091), .A2(n6090), .ZN(n6092) );
  NAND2_X1 U7680 ( .A1(n6109), .A2(n6092), .ZN(n7438) );
  OR2_X1 U7681 ( .A1(n4488), .A2(n7438), .ZN(n6094) );
  INV_X1 U7682 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7187) );
  OR2_X1 U7683 ( .A1(n6016), .A2(n7187), .ZN(n6093) );
  OR2_X1 U7684 ( .A1(n7382), .A2(n7364), .ZN(n7994) );
  NAND2_X1 U7685 ( .A1(n7382), .A2(n7364), .ZN(n8001) );
  NAND2_X1 U7686 ( .A1(n7994), .A2(n8001), .ZN(n8112) );
  NAND2_X1 U7687 ( .A1(n7374), .A2(n8112), .ZN(n6098) );
  INV_X1 U7688 ( .A(n7364), .ZN(n8252) );
  NAND2_X1 U7689 ( .A1(n7382), .A2(n8252), .ZN(n6097) );
  NAND2_X1 U7690 ( .A1(n6098), .A2(n6097), .ZN(n7360) );
  NAND2_X1 U7691 ( .A1(n6603), .A2(n7885), .ZN(n6106) );
  INV_X1 U7692 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6099) );
  AND3_X1 U7693 ( .A1(n6101), .A2(n6100), .A3(n6099), .ZN(n6102) );
  AND2_X1 U7694 ( .A1(n6103), .A2(n6102), .ZN(n6118) );
  OR2_X1 U7695 ( .A1(n6118), .A2(n5917), .ZN(n6104) );
  XNOR2_X1 U7696 ( .A(n6104), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7450) );
  AOI22_X1 U7697 ( .A1(n5996), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6538), .B2(
        n7450), .ZN(n6105) );
  NAND2_X1 U7698 ( .A1(n6353), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6115) );
  INV_X1 U7699 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n6107) );
  OR2_X1 U7700 ( .A1(n5973), .A2(n6107), .ZN(n6114) );
  INV_X1 U7701 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U7702 ( .A1(n6109), .A2(n6108), .ZN(n6110) );
  NAND2_X1 U7703 ( .A1(n6122), .A2(n6110), .ZN(n7365) );
  OR2_X1 U7704 ( .A1(n4488), .A2(n7365), .ZN(n6113) );
  INV_X1 U7705 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6111) );
  OR2_X1 U7706 ( .A1(n6016), .A2(n6111), .ZN(n6112) );
  NAND2_X1 U7707 ( .A1(n8003), .A2(n8004), .ZN(n7998) );
  NAND2_X1 U7708 ( .A1(n7993), .A2(n7998), .ZN(n8114) );
  INV_X1 U7709 ( .A(n8114), .ZN(n7359) );
  NAND2_X1 U7710 ( .A1(n6639), .A2(n7885), .ZN(n6120) );
  NAND2_X1 U7711 ( .A1(n6118), .A2(n6117), .ZN(n6162) );
  NAND2_X1 U7712 ( .A1(n6162), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6129) );
  XNOR2_X1 U7713 ( .A(n6129), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7575) );
  AOI22_X1 U7714 ( .A1(n5996), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6538), .B2(
        n7575), .ZN(n6119) );
  NAND2_X1 U7715 ( .A1(n6559), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6127) );
  INV_X1 U7716 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7426) );
  OR2_X1 U7717 ( .A1(n5962), .A2(n7426), .ZN(n6126) );
  INV_X1 U7718 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6121) );
  NAND2_X1 U7719 ( .A1(n6122), .A2(n6121), .ZN(n6123) );
  NAND2_X1 U7720 ( .A1(n6137), .A2(n6123), .ZN(n7425) );
  OR2_X1 U7721 ( .A1(n4488), .A2(n7425), .ZN(n6125) );
  INV_X1 U7722 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7601) );
  OR2_X1 U7723 ( .A1(n6016), .A2(n7601), .ZN(n6124) );
  OR2_X1 U7724 ( .A1(n7424), .A2(n7543), .ZN(n8009) );
  NAND2_X1 U7725 ( .A1(n7424), .A2(n7543), .ZN(n7539) );
  NAND2_X1 U7726 ( .A1(n8009), .A2(n7539), .ZN(n8115) );
  INV_X1 U7727 ( .A(n8115), .ZN(n7419) );
  INV_X1 U7728 ( .A(n7543), .ZN(n8251) );
  NAND2_X1 U7729 ( .A1(n7424), .A2(n8251), .ZN(n6128) );
  NAND2_X1 U7730 ( .A1(n6680), .A2(n7885), .ZN(n6135) );
  INV_X1 U7731 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U7732 ( .A1(n6129), .A2(n6160), .ZN(n6130) );
  NAND2_X1 U7733 ( .A1(n6130), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6132) );
  NAND2_X1 U7734 ( .A1(n6132), .A2(n6131), .ZN(n6145) );
  OR2_X1 U7735 ( .A1(n6132), .A2(n6131), .ZN(n6133) );
  AOI22_X1 U7736 ( .A1(n5996), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6538), .B2(
        n8278), .ZN(n6134) );
  NAND2_X1 U7737 ( .A1(n6559), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6142) );
  INV_X1 U7738 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6136) );
  OR2_X1 U7739 ( .A1(n5962), .A2(n6136), .ZN(n6141) );
  NAND2_X1 U7740 ( .A1(n6137), .A2(n9929), .ZN(n6138) );
  NAND2_X1 U7741 ( .A1(n6150), .A2(n6138), .ZN(n7479) );
  OR2_X1 U7742 ( .A1(n4488), .A2(n7479), .ZN(n6140) );
  INV_X1 U7743 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8281) );
  OR2_X1 U7744 ( .A1(n6016), .A2(n8281), .ZN(n6139) );
  NAND2_X1 U7745 ( .A1(n8643), .A2(n7591), .ZN(n8010) );
  INV_X1 U7746 ( .A(n7591), .ZN(n8250) );
  OR2_X1 U7747 ( .A1(n8643), .A2(n8250), .ZN(n6143) );
  NAND2_X1 U7748 ( .A1(n6144), .A2(n6143), .ZN(n7526) );
  NAND2_X1 U7749 ( .A1(n6814), .A2(n7885), .ZN(n6148) );
  NAND2_X1 U7750 ( .A1(n6145), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6146) );
  XNOR2_X1 U7751 ( .A(n6146), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8291) );
  AOI22_X1 U7752 ( .A1(n8291), .A2(n6538), .B1(n5996), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7753 ( .A1(n6559), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6156) );
  INV_X1 U7754 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7527) );
  OR2_X1 U7755 ( .A1(n5962), .A2(n7527), .ZN(n6155) );
  INV_X1 U7756 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7757 ( .A1(n6150), .A2(n6149), .ZN(n6151) );
  NAND2_X1 U7758 ( .A1(n6167), .A2(n6151), .ZN(n7590) );
  OR2_X1 U7759 ( .A1(n4488), .A2(n7590), .ZN(n6154) );
  INV_X1 U7760 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n6152) );
  OR2_X1 U7761 ( .A1(n6016), .A2(n6152), .ZN(n6153) );
  NAND2_X1 U7762 ( .A1(n8638), .A2(n7672), .ZN(n8018) );
  NAND2_X1 U7763 ( .A1(n7526), .A2(n8017), .ZN(n7525) );
  INV_X1 U7764 ( .A(n7672), .ZN(n8249) );
  OR2_X1 U7765 ( .A1(n8638), .A2(n8249), .ZN(n6157) );
  NAND2_X1 U7766 ( .A1(n7525), .A2(n6157), .ZN(n7668) );
  NAND2_X1 U7767 ( .A1(n6882), .A2(n7885), .ZN(n6166) );
  INV_X1 U7768 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6159) );
  NAND3_X1 U7769 ( .A1(n6160), .A2(n6131), .A3(n6159), .ZN(n6161) );
  OAI21_X1 U7770 ( .B1(n6162), .B2(n6161), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6163) );
  MUX2_X1 U7771 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6163), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n6164) );
  AND2_X1 U7772 ( .A1(n6158), .A2(n6164), .ZN(n8313) );
  AOI22_X1 U7773 ( .A1(n5996), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6538), .B2(
        n8313), .ZN(n6165) );
  NAND2_X1 U7774 ( .A1(n6167), .A2(n9926), .ZN(n6168) );
  NAND2_X1 U7775 ( .A1(n6175), .A2(n6168), .ZN(n7677) );
  INV_X1 U7776 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n6169) );
  OAI22_X1 U7777 ( .A1(n7677), .A2(n4488), .B1(n6016), .B2(n6169), .ZN(n6172)
         );
  INV_X1 U7778 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7678) );
  NAND2_X1 U7779 ( .A1(n6559), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6170) );
  OAI21_X1 U7780 ( .B1(n7678), .B2(n5962), .A(n6170), .ZN(n6171) );
  NAND2_X1 U7781 ( .A1(n7683), .A2(n7729), .ZN(n8025) );
  NAND2_X1 U7782 ( .A1(n8024), .A2(n8025), .ZN(n8022) );
  INV_X1 U7783 ( .A(n8022), .ZN(n8118) );
  NAND2_X1 U7784 ( .A1(n6158), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6173) );
  XNOR2_X1 U7785 ( .A(n6173), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8324) );
  AOI22_X1 U7786 ( .A1(n5996), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6538), .B2(
        n8324), .ZN(n6174) );
  INV_X1 U7787 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9949) );
  NAND2_X1 U7788 ( .A1(n6175), .A2(n9949), .ZN(n6176) );
  NAND2_X1 U7789 ( .A1(n6184), .A2(n6176), .ZN(n7738) );
  OR2_X1 U7790 ( .A1(n7738), .A2(n4488), .ZN(n6179) );
  AOI22_X1 U7791 ( .A1(n6353), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n6559), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n6178) );
  NAND2_X1 U7792 ( .A1(n5923), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U7793 ( .A1(n7737), .A2(n7828), .ZN(n8029) );
  INV_X1 U7794 ( .A(n7828), .ZN(n8542) );
  NAND2_X1 U7795 ( .A1(n6975), .A2(n7885), .ZN(n6183) );
  NAND2_X1 U7796 ( .A1(n4566), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6181) );
  XNOR2_X1 U7797 ( .A(n6181), .B(n4939), .ZN(n8344) );
  INV_X1 U7798 ( .A(n8344), .ZN(n8329) );
  AOI22_X1 U7799 ( .A1(n5996), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6538), .B2(
        n8329), .ZN(n6182) );
  INV_X1 U7800 ( .A(n8618), .ZN(n8538) );
  NAND2_X1 U7801 ( .A1(n6184), .A2(n9871), .ZN(n6185) );
  AND2_X1 U7802 ( .A1(n6186), .A2(n6185), .ZN(n8535) );
  NAND2_X1 U7803 ( .A1(n8535), .A2(n6262), .ZN(n6189) );
  AOI22_X1 U7804 ( .A1(n6353), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n6559), .B2(
        P2_REG0_REG_18__SCAN_IN), .ZN(n6188) );
  INV_X1 U7805 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8343) );
  OR2_X1 U7806 ( .A1(n6016), .A2(n8343), .ZN(n6187) );
  NAND2_X1 U7807 ( .A1(n8530), .A2(n5058), .ZN(n6191) );
  INV_X1 U7808 ( .A(n8514), .ZN(n8247) );
  NAND2_X1 U7809 ( .A1(n6191), .A2(n6190), .ZN(n8506) );
  INV_X1 U7810 ( .A(n8498), .ZN(n8545) );
  NAND2_X1 U7811 ( .A1(n7259), .A2(n7885), .ZN(n6193) );
  OR2_X1 U7812 ( .A1(n7886), .A2(n7260), .ZN(n6192) );
  NAND2_X1 U7813 ( .A1(n6194), .A2(n9900), .ZN(n6195) );
  AND2_X1 U7814 ( .A1(n6203), .A2(n6195), .ZN(n8493) );
  INV_X1 U7815 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U7816 ( .A1(n6559), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6197) );
  NAND2_X1 U7817 ( .A1(n5923), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6196) );
  OAI211_X1 U7818 ( .C1(n5962), .C2(n6198), .A(n6197), .B(n6196), .ZN(n6199)
         );
  AOI21_X1 U7819 ( .B1(n8493), .B2(n6262), .A(n6199), .ZN(n8516) );
  NAND2_X1 U7820 ( .A1(n8608), .A2(n8516), .ZN(n8046) );
  NAND2_X1 U7821 ( .A1(n8048), .A2(n8046), .ZN(n8496) );
  INV_X1 U7822 ( .A(n8496), .ZN(n8490) );
  INV_X1 U7823 ( .A(n8608), .ZN(n8495) );
  NAND2_X1 U7824 ( .A1(n7281), .A2(n7885), .ZN(n6201) );
  INV_X1 U7825 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7282) );
  OR2_X1 U7826 ( .A1(n7886), .A2(n7282), .ZN(n6200) );
  INV_X1 U7827 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6202) );
  NAND2_X1 U7828 ( .A1(n6203), .A2(n6202), .ZN(n6204) );
  NAND2_X1 U7829 ( .A1(n6213), .A2(n6204), .ZN(n8479) );
  OR2_X1 U7830 ( .A1(n8479), .A2(n4488), .ZN(n6210) );
  INV_X1 U7831 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U7832 ( .A1(n6559), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U7833 ( .A1(n5923), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6205) );
  OAI211_X1 U7834 ( .C1(n6207), .C2(n5962), .A(n6206), .B(n6205), .ZN(n6208)
         );
  INV_X1 U7835 ( .A(n6208), .ZN(n6209) );
  NAND2_X1 U7836 ( .A1(n7372), .A2(n7885), .ZN(n6212) );
  OR2_X1 U7837 ( .A1(n7886), .A2(n7915), .ZN(n6211) );
  NAND2_X1 U7838 ( .A1(n6213), .A2(n7904), .ZN(n6214) );
  NAND2_X1 U7839 ( .A1(n6222), .A2(n6214), .ZN(n8469) );
  OR2_X1 U7840 ( .A1(n8469), .A2(n4488), .ZN(n6219) );
  INV_X1 U7841 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8470) );
  NAND2_X1 U7842 ( .A1(n5923), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U7843 ( .A1(n6559), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6215) );
  OAI211_X1 U7844 ( .C1(n5962), .C2(n8470), .A(n6216), .B(n6215), .ZN(n6217)
         );
  INV_X1 U7845 ( .A(n6217), .ZN(n6218) );
  NAND2_X1 U7846 ( .A1(n8467), .A2(n8179), .ZN(n8054) );
  NAND2_X1 U7847 ( .A1(n8444), .A2(n8054), .ZN(n8463) );
  INV_X1 U7848 ( .A(n8467), .ZN(n8667) );
  AOI22_X1 U7849 ( .A1(n8464), .A2(n8463), .B1(n8179), .B2(n8667), .ZN(n8450)
         );
  NAND2_X1 U7850 ( .A1(n7435), .A2(n7885), .ZN(n6221) );
  OR2_X1 U7851 ( .A1(n7886), .A2(n7437), .ZN(n6220) );
  XNOR2_X1 U7852 ( .A(n6222), .B(P2_REG3_REG_23__SCAN_IN), .ZN(n8453) );
  NAND2_X1 U7853 ( .A1(n8453), .A2(n6262), .ZN(n6228) );
  INV_X1 U7854 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U7855 ( .A1(n5950), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U7856 ( .A1(n5923), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6223) );
  OAI211_X1 U7857 ( .C1(n5962), .C2(n6225), .A(n6224), .B(n6223), .ZN(n6226)
         );
  INV_X1 U7858 ( .A(n6226), .ZN(n6227) );
  NAND2_X1 U7859 ( .A1(n6228), .A2(n6227), .ZN(n8436) );
  XNOR2_X1 U7860 ( .A(n8593), .B(n8436), .ZN(n8446) );
  INV_X1 U7861 ( .A(n8446), .ZN(n8449) );
  INV_X1 U7862 ( .A(n8593), .ZN(n8455) );
  INV_X1 U7863 ( .A(n8436), .ZN(n6346) );
  NAND2_X1 U7864 ( .A1(n8593), .A2(n8436), .ZN(n6229) );
  NAND2_X1 U7865 ( .A1(n8451), .A2(n6229), .ZN(n8426) );
  NAND2_X1 U7866 ( .A1(n8587), .A2(n8210), .ZN(n8059) );
  NAND2_X1 U7867 ( .A1(n7629), .A2(n7885), .ZN(n6231) );
  OR2_X1 U7868 ( .A1(n7886), .A2(n7631), .ZN(n6230) );
  INV_X1 U7869 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9690) );
  NAND2_X1 U7870 ( .A1(n6233), .A2(n9690), .ZN(n6234) );
  NAND2_X1 U7871 ( .A1(n6247), .A2(n6234), .ZN(n8413) );
  OR2_X1 U7872 ( .A1(n8413), .A2(n4488), .ZN(n6240) );
  INV_X1 U7873 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U7874 ( .A1(n5923), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7875 ( .A1(n5950), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6235) );
  OAI211_X1 U7876 ( .C1(n5962), .C2(n6237), .A(n6236), .B(n6235), .ZN(n6238)
         );
  INV_X1 U7877 ( .A(n6238), .ZN(n6239) );
  NAND2_X1 U7878 ( .A1(n8583), .A2(n6241), .ZN(n8067) );
  NAND2_X1 U7879 ( .A1(n7686), .A2(n7885), .ZN(n6244) );
  OR2_X1 U7880 ( .A1(n7886), .A2(n7687), .ZN(n6243) );
  INV_X1 U7881 ( .A(n6247), .ZN(n6245) );
  NAND2_X1 U7882 ( .A1(n6245), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6256) );
  INV_X1 U7883 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6246) );
  NAND2_X1 U7884 ( .A1(n6247), .A2(n6246), .ZN(n6248) );
  NAND2_X1 U7885 ( .A1(n6256), .A2(n6248), .ZN(n8398) );
  OR2_X1 U7886 ( .A1(n8398), .A2(n4488), .ZN(n6253) );
  INV_X1 U7887 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8399) );
  NAND2_X1 U7888 ( .A1(n5923), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6250) );
  NAND2_X1 U7889 ( .A1(n5950), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6249) );
  OAI211_X1 U7890 ( .C1(n5962), .C2(n8399), .A(n6250), .B(n6249), .ZN(n6251)
         );
  INV_X1 U7891 ( .A(n6251), .ZN(n6252) );
  NAND2_X1 U7892 ( .A1(n8397), .A2(n8204), .ZN(n8069) );
  NAND2_X1 U7893 ( .A1(n7761), .A2(n7885), .ZN(n6255) );
  OR2_X1 U7894 ( .A1(n7886), .A2(n7762), .ZN(n6254) );
  INV_X1 U7895 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8168) );
  NAND2_X1 U7896 ( .A1(n6256), .A2(n8168), .ZN(n6257) );
  INV_X1 U7897 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n6260) );
  NAND2_X1 U7898 ( .A1(n6559), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6259) );
  NAND2_X1 U7899 ( .A1(n5923), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6258) );
  OAI211_X1 U7900 ( .C1(n6260), .C2(n5962), .A(n6259), .B(n6258), .ZN(n6261)
         );
  NAND2_X1 U7901 ( .A1(n8572), .A2(n8371), .ZN(n8072) );
  INV_X1 U7902 ( .A(n8371), .ZN(n8244) );
  NAND2_X1 U7903 ( .A1(n8149), .A2(n7885), .ZN(n6264) );
  INV_X1 U7904 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7769) );
  OR2_X1 U7905 ( .A1(n7886), .A2(n7769), .ZN(n6263) );
  INV_X1 U7906 ( .A(n6267), .ZN(n6265) );
  NAND2_X1 U7907 ( .A1(n6265), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6361) );
  INV_X1 U7908 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6266) );
  NAND2_X1 U7909 ( .A1(n6267), .A2(n6266), .ZN(n6268) );
  NAND2_X1 U7910 ( .A1(n6361), .A2(n6268), .ZN(n8197) );
  INV_X1 U7911 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n6271) );
  NAND2_X1 U7912 ( .A1(n5923), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U7913 ( .A1(n5950), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6269) );
  OAI211_X1 U7914 ( .C1(n5962), .C2(n6271), .A(n6270), .B(n6269), .ZN(n6272)
         );
  INV_X1 U7915 ( .A(n6272), .ZN(n6273) );
  AOI21_X1 U7916 ( .B1(n8362), .B2(n8369), .A(n5059), .ZN(n6289) );
  INV_X1 U7917 ( .A(n6277), .ZN(n6278) );
  INV_X1 U7918 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7911) );
  INV_X1 U7919 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9718) );
  MUX2_X1 U7920 ( .A(n7911), .B(n9718), .S(n7875), .Z(n7871) );
  XNOR2_X1 U7921 ( .A(n7871), .B(SI_29_), .ZN(n6279) );
  NAND2_X1 U7922 ( .A1(n8833), .A2(n7885), .ZN(n6281) );
  OR2_X1 U7923 ( .A1(n7886), .A2(n7911), .ZN(n6280) );
  OR2_X1 U7924 ( .A1(n6361), .A2(n4488), .ZN(n6287) );
  INV_X1 U7925 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n6284) );
  NAND2_X1 U7926 ( .A1(n5950), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6283) );
  NAND2_X1 U7927 ( .A1(n5923), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6282) );
  OAI211_X1 U7928 ( .C1(n6284), .C2(n5962), .A(n6283), .B(n6282), .ZN(n6285)
         );
  INV_X1 U7929 ( .A(n6285), .ZN(n6286) );
  INV_X1 U7930 ( .A(n8125), .ZN(n6288) );
  XNOR2_X1 U7931 ( .A(n6289), .B(n6288), .ZN(n8566) );
  NOR4_X1 U7932 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6298) );
  INV_X1 U7933 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n10422) );
  INV_X1 U7934 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10421) );
  INV_X1 U7935 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n10420) );
  INV_X1 U7936 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n10419) );
  NAND4_X1 U7937 ( .A1(n10422), .A2(n10421), .A3(n10420), .A4(n10419), .ZN(
        n6295) );
  NOR4_X1 U7938 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6293) );
  NOR4_X1 U7939 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6292) );
  NOR4_X1 U7940 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6291) );
  NOR4_X1 U7941 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6290) );
  NAND4_X1 U7942 ( .A1(n6293), .A2(n6292), .A3(n6291), .A4(n6290), .ZN(n6294)
         );
  NOR4_X1 U7943 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n6295), .A4(n6294), .ZN(n6297) );
  NOR4_X1 U7944 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n6296) );
  NAND3_X1 U7945 ( .A1(n6298), .A2(n6297), .A3(n6296), .ZN(n6313) );
  NAND2_X1 U7946 ( .A1(n6299), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6300) );
  MUX2_X1 U7947 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6300), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6301) );
  NAND2_X1 U7948 ( .A1(n6301), .A2(n5894), .ZN(n7688) );
  NAND2_X1 U7949 ( .A1(n6302), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6304) );
  MUX2_X1 U7950 ( .A(n6304), .B(P2_IR_REG_31__SCAN_IN), .S(n6303), .Z(n6305)
         );
  NAND2_X1 U7951 ( .A1(n6305), .A2(n6299), .ZN(n7630) );
  INV_X1 U7952 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6306) );
  INV_X1 U7953 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U7954 ( .A1(n6320), .A2(n6319), .ZN(n6308) );
  NAND2_X1 U7955 ( .A1(n6308), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6315) );
  INV_X1 U7956 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6314) );
  NAND2_X1 U7957 ( .A1(n6315), .A2(n6314), .ZN(n6317) );
  NAND2_X1 U7958 ( .A1(n6317), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6310) );
  INV_X1 U7959 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6309) );
  XNOR2_X1 U7960 ( .A(n7551), .B(P2_B_REG_SCAN_IN), .ZN(n6311) );
  AND2_X1 U7961 ( .A1(n6313), .A2(n10391), .ZN(n6435) );
  OR2_X1 U7962 ( .A1(n6315), .A2(n6314), .ZN(n6316) );
  NAND2_X1 U7963 ( .A1(n6317), .A2(n6316), .ZN(n6537) );
  AND2_X1 U7964 ( .A1(n6537), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6318) );
  INV_X1 U7965 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6321) );
  OR2_X1 U7966 ( .A1(n6349), .A2(n8131), .ZN(n6649) );
  NAND2_X1 U7967 ( .A1(n4552), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6322) );
  MUX2_X1 U7968 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6322), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n6323) );
  NOR2_X1 U7969 ( .A1(n8103), .A2(n10367), .ZN(n6451) );
  NOR2_X1 U7970 ( .A1(n6649), .A2(n6451), .ZN(n6446) );
  OR2_X1 U7971 ( .A1(n10390), .A2(n6446), .ZN(n6324) );
  NOR2_X1 U7972 ( .A1(n6435), .A2(n6324), .ZN(n6736) );
  NAND2_X1 U7973 ( .A1(n7551), .A2(n7688), .ZN(n10423) );
  INV_X1 U7974 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6325) );
  NAND2_X1 U7975 ( .A1(n10391), .A2(n6325), .ZN(n6326) );
  NAND2_X1 U7976 ( .A1(n6736), .A2(n6750), .ZN(n6328) );
  INV_X1 U7977 ( .A(n10391), .ZN(n6327) );
  NAND2_X1 U7978 ( .A1(n7630), .A2(n7688), .ZN(n10426) );
  OAI21_X1 U7979 ( .B1(P2_D_REG_1__SCAN_IN), .B2(n6327), .A(n10426), .ZN(n6735) );
  OR2_X1 U7980 ( .A1(n6328), .A2(n6735), .ZN(n6360) );
  INV_X1 U7981 ( .A(n8103), .ZN(n8129) );
  NAND2_X1 U7982 ( .A1(n7944), .A2(n8129), .ZN(n8140) );
  XNOR2_X1 U7983 ( .A(n6349), .B(n8140), .ZN(n6329) );
  OR2_X1 U7984 ( .A1(n6329), .A2(n10367), .ZN(n7676) );
  OR2_X1 U7985 ( .A1(n8140), .A2(n8350), .ZN(n7138) );
  NAND2_X1 U7986 ( .A1(n7676), .A2(n7138), .ZN(n10375) );
  NAND2_X1 U7987 ( .A1(n10376), .A2(n10375), .ZN(n8553) );
  OR2_X1 U7988 ( .A1(n8566), .A2(n8553), .ZN(n6370) );
  INV_X1 U7989 ( .A(n8262), .ZN(n6330) );
  NAND2_X1 U7990 ( .A1(n6330), .A2(n7119), .ZN(n6809) );
  NAND2_X1 U7991 ( .A1(n6809), .A2(n7938), .ZN(n7942) );
  NAND2_X1 U7992 ( .A1(n7942), .A2(n7945), .ZN(n6742) );
  OAI21_X1 U7993 ( .B1(n6742), .B2(n8099), .A(n7937), .ZN(n6857) );
  NAND2_X1 U7994 ( .A1(n6857), .A2(n8104), .ZN(n6331) );
  NAND2_X1 U7995 ( .A1(n6331), .A2(n7931), .ZN(n6819) );
  OAI21_X1 U7996 ( .B1(n6819), .B2(n8101), .A(n7958), .ZN(n10371) );
  NAND2_X1 U7997 ( .A1(n10371), .A2(n10370), .ZN(n10368) );
  NAND2_X1 U7998 ( .A1(n10368), .A2(n7960), .ZN(n10338) );
  XNOR2_X1 U7999 ( .A(n7966), .B(n10347), .ZN(n10345) );
  NAND2_X1 U8000 ( .A1(n7966), .A2(n10347), .ZN(n7934) );
  OAI21_X1 U8001 ( .B1(n10338), .B2(n10345), .A(n7934), .ZN(n6955) );
  INV_X1 U8002 ( .A(n8255), .ZN(n7858) );
  AOI21_X1 U8003 ( .B1(n7345), .B2(n7988), .A(n7979), .ZN(n7261) );
  NAND2_X1 U8004 ( .A1(n7261), .A2(n7986), .ZN(n7375) );
  NOR2_X1 U8005 ( .A1(n8112), .A2(n7984), .ZN(n6333) );
  NAND2_X1 U8006 ( .A1(n7375), .A2(n6333), .ZN(n7361) );
  INV_X1 U8007 ( .A(n8001), .ZN(n6334) );
  NOR2_X1 U8008 ( .A1(n8114), .A2(n6334), .ZN(n6335) );
  NAND2_X1 U8009 ( .A1(n7361), .A2(n6335), .ZN(n6336) );
  INV_X1 U8010 ( .A(n7539), .ZN(n8015) );
  NAND2_X1 U8011 ( .A1(n6338), .A2(n8024), .ZN(n7728) );
  NAND2_X1 U8012 ( .A1(n8618), .A2(n8514), .ZN(n8041) );
  OR2_X1 U8013 ( .A1(n8521), .A2(n8498), .ZN(n8042) );
  NAND2_X1 U8014 ( .A1(n8521), .A2(n8498), .ZN(n8045) );
  NAND2_X1 U8015 ( .A1(n8042), .A2(n8045), .ZN(n8508) );
  INV_X1 U8016 ( .A(n8508), .ZN(n6339) );
  AND2_X1 U8017 ( .A1(n8507), .A2(n6339), .ZN(n6340) );
  XNOR2_X1 U8018 ( .A(n8603), .B(n8499), .ZN(n8483) );
  INV_X1 U8019 ( .A(n8483), .ZN(n6342) );
  NAND2_X1 U8020 ( .A1(n8603), .A2(n8499), .ZN(n8050) );
  NAND2_X1 U8021 ( .A1(n6343), .A2(n8050), .ZN(n8459) );
  AND2_X1 U8022 ( .A1(n8444), .A2(n8446), .ZN(n6345) );
  NAND2_X1 U8023 ( .A1(n8593), .A2(n6346), .ZN(n8060) );
  NAND2_X1 U8024 ( .A1(n8435), .A2(n8434), .ZN(n8433) );
  NAND2_X1 U8025 ( .A1(n8433), .A2(n8062), .ZN(n8417) );
  INV_X1 U8026 ( .A(n8402), .ZN(n6347) );
  NOR2_X1 U8027 ( .A1(n8394), .A2(n6347), .ZN(n6348) );
  INV_X1 U8028 ( .A(n8069), .ZN(n8387) );
  INV_X1 U8029 ( .A(n6349), .ZN(n8141) );
  NAND2_X1 U8030 ( .A1(n7944), .A2(n8103), .ZN(n7925) );
  NAND2_X1 U8031 ( .A1(n8128), .A2(n7925), .ZN(n10369) );
  INV_X1 U8032 ( .A(n6350), .ZN(n8138) );
  INV_X1 U8033 ( .A(P2_B_REG_SCAN_IN), .ZN(n9869) );
  NOR2_X1 U8034 ( .A1(n6351), .A2(n9869), .ZN(n6352) );
  NOR2_X1 U8035 ( .A1(n8515), .A2(n6352), .ZN(n7891) );
  NAND2_X1 U8036 ( .A1(n6353), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U8037 ( .A1(n6559), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6355) );
  NAND2_X1 U8038 ( .A1(n5923), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6354) );
  AND3_X1 U8039 ( .A1(n6356), .A2(n6355), .A3(n6354), .ZN(n7920) );
  INV_X1 U8040 ( .A(n7920), .ZN(n8241) );
  NAND2_X1 U8041 ( .A1(n7891), .A2(n8241), .ZN(n6357) );
  NOR2_X1 U8042 ( .A1(n8565), .A2(n8548), .ZN(n6368) );
  INV_X1 U8043 ( .A(n8572), .ZN(n8384) );
  NAND2_X1 U8044 ( .A1(n7903), .A2(n10430), .ZN(n7093) );
  NAND2_X1 U8045 ( .A1(n6855), .A2(n6824), .ZN(n10358) );
  OR2_X2 U8046 ( .A1(n10358), .A2(n10363), .ZN(n10359) );
  NOR2_X4 U8047 ( .A1(n10359), .A2(n10347), .ZN(n10349) );
  INV_X1 U8048 ( .A(n7252), .ZN(n6963) );
  INV_X1 U8049 ( .A(n7975), .ZN(n10448) );
  INV_X1 U8050 ( .A(n7382), .ZN(n7441) );
  INV_X1 U8051 ( .A(n8003), .ZN(n10461) );
  NAND2_X1 U8052 ( .A1(n7380), .A2(n10461), .ZN(n7423) );
  INV_X1 U8053 ( .A(n7683), .ZN(n8629) );
  AND2_X2 U8054 ( .A1(n7735), .A2(n6180), .ZN(n8531) );
  OR2_X2 U8055 ( .A1(n8477), .A2(n8467), .ZN(n8465) );
  NAND2_X1 U8056 ( .A1(n8432), .A2(n8452), .ZN(n8427) );
  NOR2_X2 U8057 ( .A1(n8562), .A2(n8363), .ZN(n8357) );
  AOI21_X1 U8058 ( .B1(n8562), .B2(n8363), .A(n8357), .ZN(n8563) );
  NOR2_X1 U8059 ( .A1(n6360), .A2(n10367), .ZN(n10383) );
  INV_X1 U8060 ( .A(n8562), .ZN(n6364) );
  NOR2_X1 U8061 ( .A1(n10431), .A2(n8129), .ZN(n10364) );
  INV_X1 U8062 ( .A(n6361), .ZN(n6362) );
  INV_X1 U8063 ( .A(n8468), .ZN(n10379) );
  AOI22_X1 U8064 ( .A1(n6362), .A2(n10379), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n8548), .ZN(n6363) );
  OAI21_X1 U8065 ( .B1(n6364), .B2(n8537), .A(n6363), .ZN(n6365) );
  AOI21_X1 U8066 ( .B1(n8563), .B2(n8551), .A(n6365), .ZN(n6366) );
  INV_X1 U8067 ( .A(n6366), .ZN(n6367) );
  NAND2_X1 U8068 ( .A1(n6370), .A2(n6369), .ZN(P2_U3267) );
  NAND2_X1 U8069 ( .A1(n6371), .A2(n7432), .ZN(n6489) );
  OR2_X2 U8070 ( .A1(n6489), .A2(P1_U3084), .ZN(n9138) );
  NAND2_X1 U8071 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6537), .ZN(n10425) );
  INV_X2 U8072 ( .A(n8245), .ZN(P2_U3966) );
  INV_X1 U8073 ( .A(n7432), .ZN(n6372) );
  OR2_X1 U8074 ( .A1(n9067), .A2(n6372), .ZN(n6373) );
  NAND2_X1 U8075 ( .A1(n6489), .A2(n6373), .ZN(n6547) );
  OR2_X1 U8076 ( .A1(n6547), .A2(n6545), .ZN(n6374) );
  NAND2_X1 U8077 ( .A1(n6374), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8078 ( .A(n8097), .ZN(n6375) );
  XNOR2_X1 U8079 ( .A(n7424), .B(n7853), .ZN(n6377) );
  OR2_X2 U8080 ( .A1(n10462), .A2(n10367), .ZN(n7926) );
  INV_X2 U8081 ( .A(n7926), .ZN(n8186) );
  NOR2_X1 U8082 ( .A1(n7543), .A2(n8186), .ZN(n6378) );
  NAND2_X1 U8083 ( .A1(n6377), .A2(n6378), .ZN(n7483) );
  INV_X1 U8084 ( .A(n6377), .ZN(n7476) );
  INV_X1 U8085 ( .A(n6378), .ZN(n6379) );
  NAND2_X1 U8086 ( .A1(n7476), .A2(n6379), .ZN(n6380) );
  NAND2_X1 U8087 ( .A1(n7483), .A2(n6380), .ZN(n6441) );
  NAND2_X1 U8088 ( .A1(n8261), .A2(n7926), .ZN(n6381) );
  NAND2_X1 U8089 ( .A1(n6382), .A2(n6381), .ZN(n6385) );
  NAND2_X1 U8090 ( .A1(n8262), .A2(n7926), .ZN(n6384) );
  MUX2_X1 U8091 ( .A(n4490), .B(n6384), .S(n7119), .Z(n6772) );
  NAND2_X1 U8092 ( .A1(n6771), .A2(n6385), .ZN(n6789) );
  XNOR2_X1 U8093 ( .A(n4490), .B(n6755), .ZN(n6387) );
  NAND2_X1 U8094 ( .A1(n5971), .A2(n7926), .ZN(n6386) );
  XNOR2_X1 U8095 ( .A(n6387), .B(n6386), .ZN(n6788) );
  AND2_X1 U8096 ( .A1(n8260), .A2(n7926), .ZN(n6389) );
  XNOR2_X1 U8097 ( .A(n4490), .B(n6865), .ZN(n6391) );
  XNOR2_X1 U8098 ( .A(n6389), .B(n6391), .ZN(n6794) );
  INV_X1 U8099 ( .A(n6389), .ZN(n6390) );
  OR2_X1 U8100 ( .A1(n6391), .A2(n6390), .ZN(n6392) );
  XNOR2_X1 U8101 ( .A(n7115), .B(n4490), .ZN(n6802) );
  NAND2_X1 U8102 ( .A1(n8259), .A2(n7926), .ZN(n6801) );
  NAND2_X1 U8103 ( .A1(n6393), .A2(n6801), .ZN(n6395) );
  OR2_X1 U8104 ( .A1(n6804), .A2(n6802), .ZN(n6394) );
  NAND2_X1 U8105 ( .A1(n6395), .A2(n6394), .ZN(n6888) );
  INV_X1 U8106 ( .A(n6888), .ZN(n6406) );
  XNOR2_X1 U8107 ( .A(n10437), .B(n4490), .ZN(n8223) );
  NAND2_X1 U8108 ( .A1(n8258), .A2(n7926), .ZN(n6396) );
  OR2_X1 U8109 ( .A1(n8223), .A2(n6396), .ZN(n6405) );
  NAND2_X1 U8110 ( .A1(n8223), .A2(n6396), .ZN(n6397) );
  NAND2_X1 U8111 ( .A1(n6405), .A2(n6397), .ZN(n6911) );
  XNOR2_X1 U8112 ( .A(n10347), .B(n4490), .ZN(n6404) );
  INV_X1 U8113 ( .A(n6404), .ZN(n6398) );
  OR2_X1 U8114 ( .A1(n7966), .A2(n8186), .ZN(n6403) );
  OR2_X1 U8115 ( .A1(n6911), .A2(n4519), .ZN(n6889) );
  XNOR2_X1 U8116 ( .A(n7252), .B(n4490), .ZN(n6399) );
  NOR2_X1 U8117 ( .A1(n8225), .A2(n8186), .ZN(n6400) );
  NAND2_X1 U8118 ( .A1(n6399), .A2(n6400), .ZN(n6407) );
  INV_X1 U8119 ( .A(n6399), .ZN(n6905) );
  INV_X1 U8120 ( .A(n6400), .ZN(n6401) );
  NAND2_X1 U8121 ( .A1(n6905), .A2(n6401), .ZN(n6402) );
  NAND2_X1 U8122 ( .A1(n6407), .A2(n6402), .ZN(n6894) );
  XNOR2_X1 U8123 ( .A(n6404), .B(n6403), .ZN(n8234) );
  AND2_X1 U8124 ( .A1(n8234), .A2(n6405), .ZN(n8231) );
  OR2_X1 U8125 ( .A1(n4519), .A2(n8231), .ZN(n6890) );
  NAND2_X1 U8126 ( .A1(n6892), .A2(n6407), .ZN(n6412) );
  XNOR2_X1 U8127 ( .A(n7975), .B(n4490), .ZN(n7862) );
  AND2_X1 U8128 ( .A1(n8255), .A2(n7926), .ZN(n6408) );
  NAND2_X1 U8129 ( .A1(n7862), .A2(n6408), .ZN(n6413) );
  INV_X1 U8130 ( .A(n7862), .ZN(n6410) );
  INV_X1 U8131 ( .A(n6408), .ZN(n6409) );
  NAND2_X1 U8132 ( .A1(n6410), .A2(n6409), .ZN(n6411) );
  AND2_X1 U8133 ( .A1(n6413), .A2(n6411), .ZN(n6903) );
  XNOR2_X1 U8134 ( .A(n7356), .B(n7720), .ZN(n6417) );
  NOR2_X1 U8135 ( .A1(n7263), .A2(n8186), .ZN(n6415) );
  XNOR2_X1 U8136 ( .A(n6417), .B(n6415), .ZN(n7865) );
  INV_X1 U8137 ( .A(n6415), .ZN(n6416) );
  NAND2_X1 U8138 ( .A1(n6417), .A2(n6416), .ZN(n6418) );
  XNOR2_X1 U8139 ( .A(n7274), .B(n4489), .ZN(n6419) );
  NOR2_X1 U8140 ( .A1(n7346), .A2(n8186), .ZN(n6420) );
  NAND2_X1 U8141 ( .A1(n6419), .A2(n6420), .ZN(n6423) );
  INV_X1 U8142 ( .A(n6419), .ZN(n7154) );
  INV_X1 U8143 ( .A(n6420), .ZN(n6421) );
  NAND2_X1 U8144 ( .A1(n7154), .A2(n6421), .ZN(n6422) );
  AND2_X1 U8145 ( .A1(n6423), .A2(n6422), .ZN(n7049) );
  XNOR2_X1 U8146 ( .A(n7382), .B(n7853), .ZN(n6424) );
  NOR2_X1 U8147 ( .A1(n7364), .A2(n8186), .ZN(n6425) );
  NAND2_X1 U8148 ( .A1(n6424), .A2(n6425), .ZN(n6429) );
  INV_X1 U8149 ( .A(n6424), .ZN(n7328) );
  INV_X1 U8150 ( .A(n6425), .ZN(n6426) );
  NAND2_X1 U8151 ( .A1(n7328), .A2(n6426), .ZN(n6427) );
  AND2_X1 U8152 ( .A1(n6429), .A2(n6427), .ZN(n7152) );
  XNOR2_X1 U8153 ( .A(n8003), .B(n7720), .ZN(n6433) );
  NOR2_X1 U8154 ( .A1(n8004), .A2(n8186), .ZN(n6431) );
  XNOR2_X1 U8155 ( .A(n6433), .B(n6431), .ZN(n7340) );
  AND2_X1 U8156 ( .A1(n7340), .A2(n6429), .ZN(n6430) );
  INV_X1 U8157 ( .A(n6431), .ZN(n6432) );
  NAND2_X1 U8158 ( .A1(n6433), .A2(n6432), .ZN(n6434) );
  INV_X1 U8159 ( .A(n6435), .ZN(n6436) );
  NAND2_X1 U8160 ( .A1(n6436), .A2(n6737), .ZN(n6437) );
  NOR2_X1 U8161 ( .A1(n6735), .A2(n6437), .ZN(n6443) );
  INV_X1 U8162 ( .A(n10390), .ZN(n6438) );
  OR2_X1 U8163 ( .A1(n10431), .A2(n6451), .ZN(n10460) );
  AND2_X1 U8164 ( .A1(n10460), .A2(n6649), .ZN(n6439) );
  INV_X1 U8165 ( .A(n7485), .ZN(n7478) );
  AOI211_X1 U8166 ( .C1(n6441), .C2(n6440), .A(n8211), .B(n7478), .ZN(n6457)
         );
  NAND2_X1 U8167 ( .A1(n6450), .A2(n10364), .ZN(n6442) );
  INV_X1 U8168 ( .A(n7424), .ZN(n7606) );
  NOR2_X1 U8169 ( .A1(n8220), .A2(n7606), .ZN(n6456) );
  INV_X1 U8170 ( .A(n6443), .ZN(n6444) );
  NAND2_X1 U8171 ( .A1(n6444), .A2(n6734), .ZN(n6449) );
  INV_X1 U8172 ( .A(n6537), .ZN(n6445) );
  NOR2_X1 U8173 ( .A1(n6446), .A2(n6445), .ZN(n6447) );
  AND2_X1 U8174 ( .A1(n6650), .A2(n6447), .ZN(n6448) );
  NAND2_X1 U8175 ( .A1(n6449), .A2(n6448), .ZN(n6770) );
  OAI22_X1 U8176 ( .A1(n8206), .A2(n7425), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6121), .ZN(n6455) );
  INV_X1 U8177 ( .A(n6450), .ZN(n6453) );
  INV_X1 U8178 ( .A(n6451), .ZN(n6452) );
  OAI22_X1 U8179 ( .A1(n8004), .A2(n7859), .B1(n7827), .B2(n7591), .ZN(n6454)
         );
  OR4_X1 U8180 ( .A1(n6457), .A2(n6456), .A3(n6455), .A4(n6454), .ZN(P2_U3236)
         );
  AND2_X1 U8181 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7318) );
  NAND2_X1 U8182 ( .A1(n6835), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6458) );
  OAI21_X1 U8183 ( .B1(n6835), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6458), .ZN(
        n6470) );
  NOR2_X1 U8184 ( .A1(n10080), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6459) );
  AOI21_X1 U8185 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n10080), .A(n6459), .ZN(
        n10083) );
  NOR2_X1 U8186 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6573), .ZN(n6460) );
  AOI21_X1 U8187 ( .B1(n6573), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6460), .ZN(
        n6571) );
  OR2_X1 U8188 ( .A1(n6588), .A2(n6461), .ZN(n6467) );
  NOR2_X1 U8189 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9156), .ZN(n6462) );
  AOI21_X1 U8190 ( .B1(n9156), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6462), .ZN(
        n9153) );
  INV_X1 U8191 ( .A(n6505), .ZN(n9143) );
  AND2_X1 U8192 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n10048) );
  NAND2_X1 U8193 ( .A1(n6599), .A2(n10048), .ZN(n6598) );
  INV_X1 U8194 ( .A(n6602), .ZN(n6474) );
  NAND2_X1 U8195 ( .A1(n6474), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6463) );
  NAND2_X1 U8196 ( .A1(n6598), .A2(n6463), .ZN(n10042) );
  NAND2_X1 U8197 ( .A1(n10053), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6464) );
  OAI21_X1 U8198 ( .B1(n10053), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6464), .ZN(
        n10044) );
  INV_X1 U8199 ( .A(n10044), .ZN(n6465) );
  AOI21_X1 U8200 ( .B1(n10053), .B2(P1_REG2_REG_2__SCAN_IN), .A(n10043), .ZN(
        n9141) );
  XNOR2_X1 U8201 ( .A(n6505), .B(n7215), .ZN(n9140) );
  NOR2_X1 U8202 ( .A1(n9141), .A2(n9140), .ZN(n9139) );
  MUX2_X1 U8203 ( .A(n5345), .B(P1_REG2_REG_4__SCAN_IN), .S(n10069), .Z(n10065) );
  NAND2_X1 U8204 ( .A1(n9153), .A2(n9154), .ZN(n9152) );
  OAI21_X1 U8205 ( .B1(n9156), .B2(P1_REG2_REG_5__SCAN_IN), .A(n9152), .ZN(
        n6582) );
  MUX2_X1 U8206 ( .A(n6461), .B(P1_REG2_REG_6__SCAN_IN), .S(n6588), .Z(n6584)
         );
  INV_X1 U8207 ( .A(n6584), .ZN(n6466) );
  NAND2_X1 U8208 ( .A1(n6571), .A2(n6570), .ZN(n6569) );
  OAI21_X1 U8209 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6573), .A(n6569), .ZN(
        n10084) );
  NAND2_X1 U8210 ( .A1(n10083), .A2(n10084), .ZN(n10082) );
  OAI21_X1 U8211 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n10080), .A(n10082), .ZN(
        n6469) );
  NOR2_X1 U8212 ( .A1(n6469), .A2(n6470), .ZN(n6834) );
  NOR2_X1 U8213 ( .A1(n6547), .A2(P1_U3084), .ZN(n6487) );
  INV_X1 U8214 ( .A(n6468), .ZN(n9193) );
  NAND2_X1 U8215 ( .A1(n6487), .A2(n9193), .ZN(n9189) );
  OR2_X1 U8216 ( .A1(n9189), .A2(n5850), .ZN(n10159) );
  AOI211_X1 U8217 ( .C1(n6470), .C2(n6469), .A(n6834), .B(n10159), .ZN(n6493)
         );
  NAND2_X1 U8218 ( .A1(n10080), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6483) );
  MUX2_X1 U8219 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6471), .S(n10080), .Z(n10088) );
  NOR2_X1 U8220 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6573), .ZN(n6482) );
  NAND2_X1 U8221 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n9156), .ZN(n6479) );
  MUX2_X1 U8222 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6472), .S(n9156), .Z(n9159)
         );
  OR2_X1 U8223 ( .A1(n10069), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6478) );
  AOI22_X1 U8224 ( .A1(n10069), .A2(n5344), .B1(P1_REG1_REG_4__SCAN_IN), .B2(
        n6497), .ZN(n10071) );
  MUX2_X1 U8225 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6590), .S(n6602), .Z(n6473)
         );
  NAND2_X1 U8226 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n6589) );
  NOR2_X1 U8227 ( .A1(n6473), .A2(n6589), .ZN(n6591) );
  AOI21_X1 U8228 ( .B1(n6474), .B2(P1_REG1_REG_1__SCAN_IN), .A(n6591), .ZN(
        n10055) );
  MUX2_X1 U8229 ( .A(n10054), .B(P1_REG1_REG_2__SCAN_IN), .S(n10053), .Z(n6475) );
  NAND2_X1 U8230 ( .A1(n10053), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9145) );
  MUX2_X1 U8231 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6476), .S(n6505), .Z(n9144)
         );
  NOR2_X1 U8232 ( .A1(n10071), .A2(n10072), .ZN(n10070) );
  INV_X1 U8233 ( .A(n10070), .ZN(n6477) );
  MUX2_X1 U8234 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6480), .S(n6588), .Z(n6578)
         );
  MUX2_X1 U8235 ( .A(n6481), .B(P1_REG1_REG_7__SCAN_IN), .S(n6573), .Z(n6566)
         );
  NOR2_X1 U8236 ( .A1(n6565), .A2(n6566), .ZN(n6564) );
  AOI22_X1 U8237 ( .A1(n6835), .A2(n5454), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6534), .ZN(n6484) );
  AOI21_X1 U8238 ( .B1(n6485), .B2(n6484), .A(n6829), .ZN(n6488) );
  NOR2_X1 U8239 ( .A1(n5850), .A2(n9193), .ZN(n6486) );
  NAND2_X1 U8240 ( .A1(n6487), .A2(n6486), .ZN(n10169) );
  NOR2_X1 U8241 ( .A1(n6488), .A2(n10169), .ZN(n6492) );
  INV_X1 U8242 ( .A(n6489), .ZN(n6490) );
  NOR2_X1 U8243 ( .A1(P1_U3083), .A2(n6490), .ZN(n10079) );
  INV_X1 U8244 ( .A(n10079), .ZN(n10172) );
  INV_X1 U8245 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10507) );
  OR2_X1 U8246 ( .A1(n9189), .A2(n10049), .ZN(n10163) );
  OAI22_X1 U8247 ( .A1(n10172), .A2(n10507), .B1(n6534), .B2(n10163), .ZN(
        n6491) );
  OR4_X1 U8248 ( .A1(n7318), .A2(n6493), .A3(n6492), .A4(n6491), .ZN(P1_U3250)
         );
  XNOR2_X1 U8249 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  OR2_X1 U8250 ( .A1(n7875), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8686) );
  AND2_X1 U8251 ( .A1(n7875), .A2(P2_U3152), .ZN(n8684) );
  AOI22_X1 U8252 ( .A1(n6732), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n8684), .ZN(n6494) );
  OAI21_X1 U8253 ( .B1(n6502), .B2(n8686), .A(n6494), .ZN(P2_U3353) );
  AND2_X1 U8254 ( .A1(n7875), .A2(P1_U3084), .ZN(n7431) );
  INV_X2 U8255 ( .A(n7431), .ZN(n9560) );
  OR2_X1 U8256 ( .A1(n7875), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9562) );
  OAI222_X1 U8257 ( .A1(P1_U3084), .A2(n10059), .B1(n9560), .B2(n6517), .C1(
        n6495), .C2(n9562), .ZN(P1_U3351) );
  OAI222_X1 U8258 ( .A1(P1_U3084), .A2(n6497), .B1(n9560), .B2(n6498), .C1(
        n6496), .C2(n9562), .ZN(P1_U3349) );
  INV_X2 U8259 ( .A(n8684), .ZN(n8148) );
  OAI222_X1 U8260 ( .A1(n8148), .A2(n6499), .B1(n8686), .B2(n6498), .C1(
        P2_U3152), .C2(n6666), .ZN(P2_U3354) );
  OAI222_X1 U8261 ( .A1(n8148), .A2(n4610), .B1(n8686), .B2(n6506), .C1(
        P2_U3152), .C2(n6500), .ZN(P2_U3355) );
  OAI222_X1 U8262 ( .A1(P1_U3084), .A2(n6503), .B1(n9560), .B2(n6502), .C1(
        n6501), .C2(n9562), .ZN(P1_U3348) );
  INV_X1 U8263 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6504) );
  INV_X1 U8264 ( .A(n6694), .ZN(n6670) );
  OAI222_X1 U8265 ( .A1(n8148), .A2(n6504), .B1(n8686), .B2(n6508), .C1(
        P2_U3152), .C2(n6670), .ZN(P2_U3352) );
  INV_X1 U8266 ( .A(n9562), .ZN(n6886) );
  INV_X1 U8267 ( .A(n6886), .ZN(n9553) );
  OAI222_X1 U8268 ( .A1(n9553), .A2(n6507), .B1(n9560), .B2(n6506), .C1(
        P1_U3084), .C2(n6505), .ZN(P1_U3350) );
  OAI222_X1 U8269 ( .A1(n9553), .A2(n9755), .B1(n9560), .B2(n6508), .C1(
        P1_U3084), .C2(n6588), .ZN(P1_U3347) );
  OAI222_X1 U8270 ( .A1(n9553), .A2(n6509), .B1(n9560), .B2(n6514), .C1(
        P1_U3084), .C2(n6602), .ZN(P1_U3352) );
  OAI222_X1 U8271 ( .A1(n9553), .A2(n6511), .B1(n9560), .B2(n6512), .C1(
        P1_U3084), .C2(n6510), .ZN(P1_U3346) );
  INV_X1 U8272 ( .A(n8686), .ZN(n7766) );
  INV_X1 U8273 ( .A(n7766), .ZN(n7914) );
  INV_X1 U8274 ( .A(n6763), .ZN(n6677) );
  OAI222_X1 U8275 ( .A1(n8148), .A2(n6513), .B1(n7914), .B2(n6512), .C1(
        P2_U3152), .C2(n6677), .ZN(P2_U3351) );
  OAI222_X1 U8276 ( .A1(n8148), .A2(n6515), .B1(n7914), .B2(n6514), .C1(
        P2_U3152), .C2(n9981), .ZN(P2_U3357) );
  OAI222_X1 U8277 ( .A1(n8148), .A2(n6518), .B1(n7914), .B2(n6517), .C1(
        P2_U3152), .C2(n6516), .ZN(P2_U3356) );
  NAND2_X1 U8278 ( .A1(n9122), .A2(n6608), .ZN(n10247) );
  INV_X1 U8279 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9854) );
  INV_X1 U8280 ( .A(n6519), .ZN(n6520) );
  AOI22_X1 U8281 ( .A1(n10247), .A2(n9854), .B1(n6520), .B2(n9122), .ZN(
        P1_U3441) );
  OAI222_X1 U8282 ( .A1(n9553), .A2(n6522), .B1(n9560), .B2(n6523), .C1(
        P1_U3084), .C2(n6521), .ZN(P1_U3345) );
  INV_X1 U8283 ( .A(n6980), .ZN(n6989) );
  OAI222_X1 U8284 ( .A1(n8148), .A2(n6524), .B1(n7914), .B2(n6523), .C1(
        P2_U3152), .C2(n6989), .ZN(P2_U3350) );
  INV_X1 U8285 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6531) );
  INV_X1 U8286 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U8287 ( .A1(n5325), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6528) );
  INV_X1 U8288 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6525) );
  OR2_X1 U8289 ( .A1(n6526), .A2(n6525), .ZN(n6527) );
  OAI211_X1 U8290 ( .C1(n8832), .C2(n6529), .A(n6528), .B(n6527), .ZN(n9194)
         );
  NAND2_X1 U8291 ( .A1(P1_U4006), .A2(n9194), .ZN(n6530) );
  OAI21_X1 U8292 ( .B1(P1_U4006), .B2(n6531), .A(n6530), .ZN(P1_U3586) );
  NAND2_X1 U8293 ( .A1(P1_U4006), .A2(n6932), .ZN(n6532) );
  OAI21_X1 U8294 ( .B1(P1_U4006), .B2(n5959), .A(n6532), .ZN(P1_U3555) );
  INV_X1 U8295 ( .A(n6533), .ZN(n6535) );
  OAI222_X1 U8296 ( .A1(n9553), .A2(n9680), .B1(n9560), .B2(n6535), .C1(n6534), 
        .C2(P1_U3084), .ZN(P1_U3344) );
  INV_X1 U8297 ( .A(n8272), .ZN(n6991) );
  OAI222_X1 U8298 ( .A1(n8148), .A2(n6536), .B1(n7914), .B2(n6535), .C1(n6991), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  NOR2_X1 U8299 ( .A1(n6537), .A2(P2_U3152), .ZN(n8143) );
  INV_X1 U8300 ( .A(n8143), .ZN(n8145) );
  NAND2_X1 U8301 ( .A1(n10390), .A2(n8145), .ZN(n6539) );
  NAND2_X1 U8302 ( .A1(n6539), .A2(n6538), .ZN(n6541) );
  OR2_X1 U8303 ( .A1(n10390), .A2(n6649), .ZN(n6540) );
  NAND2_X1 U8304 ( .A1(n6541), .A2(n6540), .ZN(n10333) );
  NOR2_X1 U8305 ( .A1(P2_U3966), .A2(n10333), .ZN(P2_U3151) );
  INV_X1 U8306 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6551) );
  AOI21_X1 U8307 ( .B1(n9193), .B2(n6542), .A(n5850), .ZN(n10052) );
  INV_X1 U8308 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6624) );
  AND2_X1 U8309 ( .A1(n6468), .A2(n6624), .ZN(n6543) );
  OAI21_X1 U8310 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n6543), .A(n10052), .ZN(
        n6544) );
  OAI21_X1 U8311 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n10052), .A(n6544), .ZN(
        n6546) );
  NOR4_X1 U8312 ( .A1(n6547), .A2(n6546), .A3(n6545), .A4(P1_U3084), .ZN(n6549) );
  INV_X1 U8313 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9908) );
  NOR3_X1 U8314 ( .A1(n10169), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n9908), .ZN(
        n6548) );
  AOI211_X1 U8315 ( .C1(P1_REG3_REG_0__SCAN_IN), .C2(P1_U3084), .A(n6549), .B(
        n6548), .ZN(n6550) );
  OAI21_X1 U8316 ( .B1(n10172), .B2(n6551), .A(n6550), .ZN(P1_U3241) );
  INV_X1 U8317 ( .A(n6552), .ZN(n6553) );
  OAI222_X1 U8318 ( .A1(n9553), .A2(n9750), .B1(n9560), .B2(n6553), .C1(n4720), 
        .C2(P1_U3084), .ZN(P1_U3343) );
  INV_X1 U8319 ( .A(n7188), .ZN(n6997) );
  OAI222_X1 U8320 ( .A1(n8148), .A2(n6554), .B1(n7914), .B2(n6553), .C1(n6997), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U8321 ( .A(n6555), .ZN(n6556) );
  INV_X1 U8322 ( .A(n7063), .ZN(n7058) );
  OAI222_X1 U8323 ( .A1(n9553), .A2(n9934), .B1(n9560), .B2(n6556), .C1(n7058), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  INV_X1 U8324 ( .A(n7307), .ZN(n7183) );
  OAI222_X1 U8325 ( .A1(n8148), .A2(n6557), .B1(n7914), .B2(n6556), .C1(n7183), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  NAND2_X1 U8326 ( .A1(n8245), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6558) );
  OAI21_X1 U8327 ( .B1(n8516), .B2(n8245), .A(n6558), .ZN(P2_U3572) );
  INV_X1 U8328 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6563) );
  INV_X1 U8329 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n7890) );
  NAND2_X1 U8330 ( .A1(n5923), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6561) );
  NAND2_X1 U8331 ( .A1(n6559), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6560) );
  OAI211_X1 U8332 ( .C1(n5962), .C2(n7890), .A(n6561), .B(n6560), .ZN(n7919)
         );
  NAND2_X1 U8333 ( .A1(P2_U3966), .A2(n7919), .ZN(n6562) );
  OAI21_X1 U8334 ( .B1(P2_U3966), .B2(n6563), .A(n6562), .ZN(P2_U3583) );
  AND2_X1 U8335 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8694) );
  AOI21_X1 U8336 ( .B1(n6566), .B2(n6565), .A(n6564), .ZN(n6567) );
  NOR2_X1 U8337 ( .A1(n10169), .A2(n6567), .ZN(n6568) );
  AOI211_X1 U8338 ( .C1(n10079), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n8694), .B(
        n6568), .ZN(n6575) );
  INV_X1 U8339 ( .A(n10159), .ZN(n10086) );
  OAI21_X1 U8340 ( .B1(n6571), .B2(n6570), .A(n6569), .ZN(n6572) );
  AOI22_X1 U8341 ( .A1(n6573), .A2(n10129), .B1(n10086), .B2(n6572), .ZN(n6574) );
  NAND2_X1 U8342 ( .A1(n6575), .A2(n6574), .ZN(P1_U3248) );
  INV_X1 U8343 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6576) );
  NOR2_X1 U8344 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6576), .ZN(n7007) );
  AOI21_X1 U8345 ( .B1(n6579), .B2(n6578), .A(n6577), .ZN(n6580) );
  NOR2_X1 U8346 ( .A1(n10169), .A2(n6580), .ZN(n6581) );
  AOI211_X1 U8347 ( .C1(n10079), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n7007), .B(
        n6581), .ZN(n6587) );
  INV_X1 U8348 ( .A(n6582), .ZN(n6585) );
  OAI211_X1 U8349 ( .C1(n6585), .C2(n6584), .A(n10086), .B(n6583), .ZN(n6586)
         );
  OAI211_X1 U8350 ( .C1(n10163), .C2(n6588), .A(n6587), .B(n6586), .ZN(
        P1_U3247) );
  INV_X1 U8351 ( .A(n6589), .ZN(n6594) );
  MUX2_X1 U8352 ( .A(n6590), .B(P1_REG1_REG_1__SCAN_IN), .S(n6602), .Z(n6593)
         );
  INV_X1 U8353 ( .A(n10169), .ZN(n10147) );
  INV_X1 U8354 ( .A(n6591), .ZN(n6592) );
  OAI211_X1 U8355 ( .C1(n6594), .C2(n6593), .A(n10147), .B(n6592), .ZN(n6595)
         );
  OAI21_X1 U8356 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6596), .A(n6595), .ZN(n6597) );
  AOI21_X1 U8357 ( .B1(n10079), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n6597), .ZN(
        n6601) );
  OAI211_X1 U8358 ( .C1(n6599), .C2(n10048), .A(n10086), .B(n6598), .ZN(n6600)
         );
  OAI211_X1 U8359 ( .C1(n10163), .C2(n6602), .A(n6601), .B(n6600), .ZN(
        P1_U3242) );
  INV_X1 U8360 ( .A(n6603), .ZN(n6625) );
  AOI22_X1 U8361 ( .A1(n7450), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n8684), .ZN(n6604) );
  OAI21_X1 U8362 ( .B1(n6625), .B2(n8686), .A(n6604), .ZN(P2_U3346) );
  INV_X1 U8363 ( .A(n6605), .ZN(n6606) );
  NOR2_X1 U8364 ( .A1(n6608), .A2(n6606), .ZN(n6607) );
  NOR2_X1 U8365 ( .A1(n6619), .A2(n6607), .ZN(n6610) );
  OAI21_X1 U8366 ( .B1(n6608), .B2(P1_D_REG_0__SCAN_IN), .A(n9551), .ZN(n6609)
         );
  AND2_X1 U8367 ( .A1(n6610), .A2(n6609), .ZN(n6941) );
  INV_X1 U8368 ( .A(n9437), .ZN(n6926) );
  AND2_X2 U8369 ( .A1(n6941), .A2(n6620), .ZN(n10315) );
  INV_X1 U8370 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6617) );
  INV_X1 U8371 ( .A(n6946), .ZN(n6615) );
  AND2_X1 U8372 ( .A1(n6932), .A2(n6615), .ZN(n9077) );
  NOR2_X1 U8373 ( .A1(n7014), .A2(n9077), .ZN(n8841) );
  NAND2_X1 U8374 ( .A1(n7044), .A2(n6614), .ZN(n6612) );
  INV_X1 U8375 ( .A(n6920), .ZN(n6611) );
  OR2_X1 U8376 ( .A1(n9067), .A2(n10049), .ZN(n10183) );
  OAI22_X1 U8377 ( .A1(n8841), .A2(n6612), .B1(n6611), .B2(n10183), .ZN(n6949)
         );
  INV_X1 U8378 ( .A(n6949), .ZN(n6613) );
  OAI21_X1 U8379 ( .B1(n6615), .B2(n6614), .A(n6613), .ZN(n6622) );
  NAND2_X1 U8380 ( .A1(n6622), .A2(n10315), .ZN(n6616) );
  OAI21_X1 U8381 ( .B1(n10315), .B2(n6617), .A(n6616), .ZN(P1_U3454) );
  NOR2_X1 U8382 ( .A1(n6619), .A2(n6618), .ZN(n6621) );
  AND2_X2 U8383 ( .A1(n6621), .A2(n6620), .ZN(n10326) );
  NAND2_X1 U8384 ( .A1(n6622), .A2(n10326), .ZN(n6623) );
  OAI21_X1 U8385 ( .B1(n10326), .B2(n6624), .A(n6623), .ZN(P1_U3523) );
  INV_X1 U8386 ( .A(n7068), .ZN(n7398) );
  OAI222_X1 U8387 ( .A1(n9553), .A2(n9728), .B1(n9560), .B2(n6625), .C1(
        P1_U3084), .C2(n7398), .ZN(P1_U3341) );
  OAI21_X1 U8388 ( .B1(n6628), .B2(n6627), .A(n6626), .ZN(n10046) );
  AOI22_X1 U8389 ( .A1(n8817), .A2(n6920), .B1(n10046), .B2(n8812), .ZN(n6631)
         );
  NAND2_X1 U8390 ( .A1(n8795), .A2(n6629), .ZN(n8790) );
  AOI22_X1 U8391 ( .A1(n8791), .A2(n6946), .B1(n8790), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n6630) );
  NAND2_X1 U8392 ( .A1(n6631), .A2(n6630), .ZN(P1_U3230) );
  NAND2_X1 U8393 ( .A1(n6632), .A2(n6633), .ZN(n6635) );
  XNOR2_X1 U8394 ( .A(n6635), .B(n6634), .ZN(n6638) );
  INV_X1 U8395 ( .A(n8819), .ZN(n8808) );
  AOI22_X1 U8396 ( .A1(n8808), .A2(n6932), .B1(n8817), .B2(n7020), .ZN(n6637)
         );
  AOI22_X1 U8397 ( .A1(n8791), .A2(n7030), .B1(n8790), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n6636) );
  OAI211_X1 U8398 ( .C1(n6638), .C2(n8773), .A(n6637), .B(n6636), .ZN(P1_U3220) );
  INV_X1 U8399 ( .A(n7407), .ZN(n10104) );
  INV_X1 U8400 ( .A(n6639), .ZN(n6640) );
  OAI222_X1 U8401 ( .A1(P1_U3084), .A2(n10104), .B1(n9560), .B2(n6640), .C1(
        n9738), .C2(n9562), .ZN(P1_U3340) );
  INV_X1 U8402 ( .A(n7575), .ZN(n7571) );
  OAI222_X1 U8403 ( .A1(n8148), .A2(n6641), .B1(n7914), .B2(n6640), .C1(n7571), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8404 ( .A(n6666), .ZN(n6707) );
  INV_X1 U8405 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6642) );
  MUX2_X1 U8406 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6642), .S(n6666), .Z(n6703)
         );
  INV_X1 U8407 ( .A(n9981), .ZN(n6643) );
  AOI22_X1 U8408 ( .A1(n6643), .A2(n5938), .B1(P2_REG2_REG_1__SCAN_IN), .B2(
        n9981), .ZN(n9977) );
  NOR3_X1 U8409 ( .A1(n10335), .A2(n5953), .A3(n9977), .ZN(n9975) );
  AOI21_X1 U8410 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n6643), .A(n9975), .ZN(
        n9991) );
  NAND2_X1 U8411 ( .A1(n9993), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6644) );
  OAI21_X1 U8412 ( .B1(n9993), .B2(P2_REG2_REG_2__SCAN_IN), .A(n6644), .ZN(
        n9990) );
  NOR2_X1 U8413 ( .A1(n9991), .A2(n9990), .ZN(n9989) );
  NAND2_X1 U8414 ( .A1(n6720), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6645) );
  OAI21_X1 U8415 ( .B1(n6720), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6645), .ZN(
        n6716) );
  AOI21_X1 U8416 ( .B1(n6707), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6702), .ZN(
        n6729) );
  NAND2_X1 U8417 ( .A1(n6732), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6646) );
  OAI21_X1 U8418 ( .B1(n6732), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6646), .ZN(
        n6728) );
  INV_X1 U8419 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6647) );
  AOI22_X1 U8420 ( .A1(n6694), .A2(n6647), .B1(P2_REG2_REG_6__SCAN_IN), .B2(
        n6670), .ZN(n6690) );
  NAND2_X1 U8421 ( .A1(n6763), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6648) );
  OAI21_X1 U8422 ( .B1(n6763), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6648), .ZN(
        n6655) );
  NOR2_X1 U8423 ( .A1(n6656), .A2(n6655), .ZN(n6762) );
  INV_X1 U8424 ( .A(n6649), .ZN(n6652) );
  OR2_X1 U8425 ( .A1(n6350), .A2(P2_U3152), .ZN(n7767) );
  OR2_X1 U8426 ( .A1(n6650), .A2(n7767), .ZN(n6651) );
  OAI211_X1 U8427 ( .C1(n10390), .C2(n6652), .A(n8145), .B(n6651), .ZN(n6653)
         );
  AND2_X1 U8428 ( .A1(n6653), .A2(n5946), .ZN(n6672) );
  NOR2_X1 U8429 ( .A1(n6350), .A2(n6351), .ZN(n6654) );
  NAND2_X1 U8430 ( .A1(n6657), .A2(n6654), .ZN(n9988) );
  AOI211_X1 U8431 ( .C1(n6656), .C2(n6655), .A(n6762), .B(n9988), .ZN(n6679)
         );
  NAND2_X1 U8432 ( .A1(n6657), .A2(n6350), .ZN(n10327) );
  NOR2_X1 U8433 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6036), .ZN(n6658) );
  AOI21_X1 U8434 ( .B1(n10333), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6658), .ZN(
        n6676) );
  MUX2_X1 U8435 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6659), .S(n6694), .Z(n6684)
         );
  NAND2_X1 U8436 ( .A1(n6732), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6669) );
  NAND2_X1 U8437 ( .A1(n6720), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6664) );
  MUX2_X1 U8438 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6660), .S(n6720), .Z(n6710)
         );
  NAND2_X1 U8439 ( .A1(n9993), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6663) );
  MUX2_X1 U8440 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6661), .S(n9993), .Z(n9996)
         );
  MUX2_X1 U8441 ( .A(n6662), .B(P2_REG1_REG_1__SCAN_IN), .S(n9981), .Z(n9984)
         );
  NAND3_X1 U8442 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n9984), .ZN(n9983) );
  OAI21_X1 U8443 ( .B1(n9981), .B2(n6662), .A(n9983), .ZN(n9997) );
  NAND2_X1 U8444 ( .A1(n9996), .A2(n9997), .ZN(n9995) );
  NAND2_X1 U8445 ( .A1(n6663), .A2(n9995), .ZN(n6711) );
  NAND2_X1 U8446 ( .A1(n6710), .A2(n6711), .ZN(n6709) );
  NAND2_X1 U8447 ( .A1(n6664), .A2(n6709), .ZN(n6698) );
  MUX2_X1 U8448 ( .A(n6665), .B(P2_REG1_REG_4__SCAN_IN), .S(n6666), .Z(n6697)
         );
  NAND2_X1 U8449 ( .A1(n6698), .A2(n6697), .ZN(n6696) );
  OAI21_X1 U8450 ( .B1(n6665), .B2(n6666), .A(n6696), .ZN(n6722) );
  MUX2_X1 U8451 ( .A(n5989), .B(P2_REG1_REG_5__SCAN_IN), .S(n6732), .Z(n6723)
         );
  INV_X1 U8452 ( .A(n6723), .ZN(n6667) );
  NAND2_X1 U8453 ( .A1(n6722), .A2(n6667), .ZN(n6668) );
  NAND2_X1 U8454 ( .A1(n6669), .A2(n6668), .ZN(n6685) );
  NAND2_X1 U8455 ( .A1(n6684), .A2(n6685), .ZN(n6683) );
  OAI21_X1 U8456 ( .B1(n6670), .B2(n6659), .A(n6683), .ZN(n6674) );
  MUX2_X1 U8457 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6671), .S(n6763), .Z(n6673)
         );
  NAND2_X1 U8458 ( .A1(n6672), .A2(n6351), .ZN(n10328) );
  INV_X1 U8459 ( .A(n10328), .ZN(n10330) );
  NAND2_X1 U8460 ( .A1(n6673), .A2(n6674), .ZN(n6756) );
  OAI211_X1 U8461 ( .C1(n6674), .C2(n6673), .A(n10330), .B(n6756), .ZN(n6675)
         );
  OAI211_X1 U8462 ( .C1(n10327), .C2(n6677), .A(n6676), .B(n6675), .ZN(n6678)
         );
  OR2_X1 U8463 ( .A1(n6679), .A2(n6678), .ZN(P2_U3252) );
  INV_X1 U8464 ( .A(n6680), .ZN(n6681) );
  INV_X1 U8465 ( .A(n7400), .ZN(n9179) );
  OAI222_X1 U8466 ( .A1(n9553), .A2(n9703), .B1(n9560), .B2(n6681), .C1(n9179), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U8467 ( .A(n8278), .ZN(n8282) );
  OAI222_X1 U8468 ( .A1(n8148), .A2(n6682), .B1(n7914), .B2(n6681), .C1(n8282), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8469 ( .A(n10327), .ZN(n9994) );
  OAI21_X1 U8470 ( .B1(n6685), .B2(n6684), .A(n6683), .ZN(n6688) );
  NOR2_X1 U8471 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9848), .ZN(n6686) );
  AOI21_X1 U8472 ( .B1(n10333), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n6686), .ZN(
        n6687) );
  OAI21_X1 U8473 ( .B1(n10328), .B2(n6688), .A(n6687), .ZN(n6693) );
  AOI211_X1 U8474 ( .C1(n6691), .C2(n6690), .A(n6689), .B(n9988), .ZN(n6692)
         );
  AOI211_X1 U8475 ( .C1(n9994), .C2(n6694), .A(n6693), .B(n6692), .ZN(n6695)
         );
  INV_X1 U8476 ( .A(n6695), .ZN(P2_U3251) );
  OAI21_X1 U8477 ( .B1(n6698), .B2(n6697), .A(n6696), .ZN(n6701) );
  INV_X1 U8478 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9902) );
  NOR2_X1 U8479 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9902), .ZN(n6699) );
  AOI21_X1 U8480 ( .B1(n10333), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6699), .ZN(
        n6700) );
  OAI21_X1 U8481 ( .B1(n10328), .B2(n6701), .A(n6700), .ZN(n6706) );
  AOI211_X1 U8482 ( .C1(n6704), .C2(n6703), .A(n6702), .B(n9988), .ZN(n6705)
         );
  AOI211_X1 U8483 ( .C1(n9994), .C2(n6707), .A(n6706), .B(n6705), .ZN(n6708)
         );
  INV_X1 U8484 ( .A(n6708), .ZN(P2_U3249) );
  OAI21_X1 U8485 ( .B1(n6711), .B2(n6710), .A(n6709), .ZN(n6714) );
  INV_X1 U8486 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10378) );
  NOR2_X1 U8487 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10378), .ZN(n6712) );
  AOI21_X1 U8488 ( .B1(n10333), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n6712), .ZN(
        n6713) );
  OAI21_X1 U8489 ( .B1(n10328), .B2(n6714), .A(n6713), .ZN(n6719) );
  AOI211_X1 U8490 ( .C1(n6717), .C2(n6716), .A(n6715), .B(n9988), .ZN(n6718)
         );
  AOI211_X1 U8491 ( .C1(n9994), .C2(n6720), .A(n6719), .B(n6718), .ZN(n6721)
         );
  INV_X1 U8492 ( .A(n6721), .ZN(P2_U3248) );
  XOR2_X1 U8493 ( .A(n6723), .B(n6722), .Z(n6726) );
  NOR2_X1 U8494 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6914), .ZN(n6724) );
  AOI21_X1 U8495 ( .B1(n10333), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6724), .ZN(
        n6725) );
  OAI21_X1 U8496 ( .B1(n10328), .B2(n6726), .A(n6725), .ZN(n6731) );
  AOI211_X1 U8497 ( .C1(n6729), .C2(n6728), .A(n6727), .B(n9988), .ZN(n6730)
         );
  AOI211_X1 U8498 ( .C1(n9994), .C2(n6732), .A(n6731), .B(n6730), .ZN(n6733)
         );
  INV_X1 U8499 ( .A(n6733), .ZN(P2_U3250) );
  AND2_X2 U8500 ( .A1(n6751), .A2(n6737), .ZN(n10477) );
  NAND2_X1 U8501 ( .A1(n10477), .A2(n8644), .ZN(n8628) );
  NOR2_X1 U8502 ( .A1(n8103), .A2(n8350), .ZN(n6738) );
  NAND2_X1 U8503 ( .A1(n6349), .A2(n6738), .ZN(n8633) );
  OAI21_X1 U8504 ( .B1(n6740), .B2(n8099), .A(n6739), .ZN(n7107) );
  NAND2_X1 U8505 ( .A1(n7093), .A2(n7106), .ZN(n6741) );
  NAND3_X1 U8506 ( .A1(n6856), .A2(n10360), .A3(n6741), .ZN(n7102) );
  INV_X1 U8507 ( .A(n7102), .ZN(n6748) );
  XNOR2_X1 U8508 ( .A(n6742), .B(n8099), .ZN(n6743) );
  NAND2_X1 U8509 ( .A1(n6743), .A2(n10369), .ZN(n6747) );
  NAND2_X1 U8510 ( .A1(n8260), .A2(n8544), .ZN(n6745) );
  NAND2_X1 U8511 ( .A1(n8261), .A2(n8543), .ZN(n6744) );
  NAND2_X1 U8512 ( .A1(n6745), .A2(n6744), .ZN(n6790) );
  INV_X1 U8513 ( .A(n6790), .ZN(n6746) );
  NAND2_X1 U8514 ( .A1(n6747), .A2(n6746), .ZN(n7105) );
  AOI211_X1 U8515 ( .C1(n10466), .C2(n7107), .A(n6748), .B(n7105), .ZN(n6752)
         );
  MUX2_X1 U8516 ( .A(n6661), .B(n6752), .S(n10477), .Z(n6749) );
  OAI21_X1 U8517 ( .B1(n6755), .B2(n8628), .A(n6749), .ZN(P2_U3522) );
  AND2_X2 U8518 ( .A1(n6751), .A2(n6750), .ZN(n10469) );
  NAND2_X1 U8519 ( .A1(n10469), .A2(n8644), .ZN(n8678) );
  INV_X1 U8520 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6753) );
  MUX2_X1 U8521 ( .A(n6753), .B(n6752), .S(n10469), .Z(n6754) );
  OAI21_X1 U8522 ( .B1(n6755), .B2(n8678), .A(n6754), .ZN(P2_U3457) );
  NOR2_X1 U8523 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9842), .ZN(n6761) );
  NAND2_X1 U8524 ( .A1(n6763), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6757) );
  AND2_X1 U8525 ( .A1(n6757), .A2(n6756), .ZN(n6759) );
  MUX2_X1 U8526 ( .A(n6990), .B(P2_REG1_REG_8__SCAN_IN), .S(n6980), .Z(n6758)
         );
  NOR2_X1 U8527 ( .A1(n6759), .A2(n6758), .ZN(n6987) );
  AOI211_X1 U8528 ( .C1(n6759), .C2(n6758), .A(n10328), .B(n6987), .ZN(n6760)
         );
  AOI211_X1 U8529 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n10333), .A(n6761), .B(
        n6760), .ZN(n6769) );
  XNOR2_X1 U8530 ( .A(n6980), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n6765) );
  INV_X1 U8531 ( .A(n6765), .ZN(n6767) );
  INV_X1 U8532 ( .A(n6764), .ZN(n6766) );
  OAI211_X1 U8533 ( .C1(n6767), .C2(n6766), .A(n10331), .B(n6979), .ZN(n6768)
         );
  OAI211_X1 U8534 ( .C1(n10327), .C2(n6989), .A(n6769), .B(n6768), .ZN(
        P2_U3253) );
  NOR2_X1 U8535 ( .A1(n6770), .A2(P2_U3152), .ZN(n6787) );
  INV_X1 U8536 ( .A(n8211), .ZN(n8235) );
  NAND2_X1 U8537 ( .A1(n5971), .A2(n8544), .ZN(n6774) );
  NAND2_X1 U8538 ( .A1(n8262), .A2(n8543), .ZN(n6773) );
  NAND2_X1 U8539 ( .A1(n6774), .A2(n6773), .ZN(n7090) );
  AOI22_X1 U8540 ( .A1(n8235), .A2(n6775), .B1(n8227), .B2(n7090), .ZN(n6777)
         );
  NAND2_X1 U8541 ( .A1(n8230), .A2(n7098), .ZN(n6776) );
  OAI211_X1 U8542 ( .C1(n6787), .C2(n9841), .A(n6777), .B(n6776), .ZN(P2_U3224) );
  OAI21_X1 U8543 ( .B1(n6780), .B2(n6779), .A(n6778), .ZN(n6785) );
  NAND2_X1 U8544 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9150) );
  INV_X1 U8545 ( .A(n9150), .ZN(n6781) );
  AOI21_X1 U8546 ( .B1(n8808), .B2(n7020), .A(n6781), .ZN(n6783) );
  AOI22_X1 U8547 ( .A1(n8817), .A2(n9137), .B1(n8791), .B2(n7220), .ZN(n6782)
         );
  OAI211_X1 U8548 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n8804), .A(n6783), .B(
        n6782), .ZN(n6784) );
  AOI21_X1 U8549 ( .B1(n6785), .B2(n8812), .A(n6784), .ZN(n6786) );
  INV_X1 U8550 ( .A(n6786), .ZN(P1_U3216) );
  INV_X1 U8551 ( .A(n6787), .ZN(n6811) );
  AOI22_X1 U8552 ( .A1(n6811), .A2(P2_REG3_REG_2__SCAN_IN), .B1(n7106), .B2(
        n8230), .ZN(n6793) );
  XOR2_X1 U8553 ( .A(n6789), .B(n6788), .Z(n6791) );
  AOI22_X1 U8554 ( .A1(n8235), .A2(n6791), .B1(n8227), .B2(n6790), .ZN(n6792)
         );
  NAND2_X1 U8555 ( .A1(n6793), .A2(n6792), .ZN(P2_U3239) );
  XNOR2_X1 U8556 ( .A(n6795), .B(n6794), .ZN(n6800) );
  AOI22_X1 U8557 ( .A1(n5984), .A2(n8230), .B1(n8229), .B2(n10378), .ZN(n6799)
         );
  INV_X1 U8558 ( .A(n8259), .ZN(n6797) );
  INV_X1 U8559 ( .A(n5971), .ZN(n6796) );
  OAI22_X1 U8560 ( .A1(n6797), .A2(n8515), .B1(n6796), .B2(n8513), .ZN(n6860)
         );
  AOI22_X1 U8561 ( .A1(n8227), .A2(n6860), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        P2_U3152), .ZN(n6798) );
  OAI211_X1 U8562 ( .C1(n8211), .C2(n6800), .A(n6799), .B(n6798), .ZN(P2_U3220) );
  XNOR2_X1 U8563 ( .A(n6802), .B(n6801), .ZN(n6803) );
  XNOR2_X1 U8564 ( .A(n6804), .B(n6803), .ZN(n6808) );
  INV_X1 U8565 ( .A(n7110), .ZN(n6805) );
  AOI22_X1 U8566 ( .A1(n7115), .A2(n8230), .B1(n8229), .B2(n6805), .ZN(n6807)
         );
  INV_X1 U8567 ( .A(n8258), .ZN(n8226) );
  OAI22_X1 U8568 ( .A1(n5985), .A2(n8513), .B1(n8226), .B2(n8515), .ZN(n6820)
         );
  AOI22_X1 U8569 ( .A1(n8227), .A2(n6820), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n6806) );
  OAI211_X1 U8570 ( .C1(n8211), .C2(n6808), .A(n6807), .B(n6806), .ZN(P2_U3232) );
  NAND2_X1 U8571 ( .A1(n8262), .A2(n10430), .ZN(n7943) );
  AOI22_X1 U8572 ( .A1(n8216), .A2(n8261), .B1(n7119), .B2(n8230), .ZN(n6813)
         );
  OAI21_X1 U8573 ( .B1(n10430), .B2(n7926), .A(n6809), .ZN(n6810) );
  AOI22_X1 U8574 ( .A1(n6811), .A2(P2_REG3_REG_0__SCAN_IN), .B1(n8235), .B2(
        n6810), .ZN(n6812) );
  OAI211_X1 U8575 ( .C1(n8224), .C2(n7943), .A(n6813), .B(n6812), .ZN(P2_U3234) );
  INV_X1 U8576 ( .A(n6814), .ZN(n6816) );
  INV_X1 U8577 ( .A(n8291), .ZN(n8297) );
  OAI222_X1 U8578 ( .A1(n8148), .A2(n6815), .B1(n7914), .B2(n6816), .C1(
        P2_U3152), .C2(n8297), .ZN(P2_U3343) );
  INV_X1 U8579 ( .A(n10117), .ZN(n9180) );
  OAI222_X1 U8580 ( .A1(n9553), .A2(n9899), .B1(n9560), .B2(n6816), .C1(
        P1_U3084), .C2(n9180), .ZN(P1_U3338) );
  NAND2_X1 U8581 ( .A1(n8245), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6817) );
  OAI21_X1 U8582 ( .B1(n8204), .B2(n8245), .A(n6817), .ZN(P2_U3578) );
  NAND2_X1 U8583 ( .A1(n6818), .A2(n8101), .ZN(n10356) );
  OAI21_X1 U8584 ( .B1(n6818), .B2(n8101), .A(n10356), .ZN(n7116) );
  OAI211_X1 U8585 ( .C1(n6855), .C2(n6824), .A(n10358), .B(n10360), .ZN(n7111)
         );
  INV_X1 U8586 ( .A(n7111), .ZN(n6822) );
  INV_X1 U8587 ( .A(n10369), .ZN(n8510) );
  AOI211_X1 U8588 ( .C1(n8101), .C2(n6819), .A(n8510), .B(n4569), .ZN(n6821)
         );
  OR2_X1 U8589 ( .A1(n6821), .A2(n6820), .ZN(n7114) );
  AOI211_X1 U8590 ( .C1(n10466), .C2(n7116), .A(n6822), .B(n7114), .ZN(n6828)
         );
  INV_X1 U8591 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6823) );
  OAI22_X1 U8592 ( .A1(n8678), .A2(n6824), .B1(n10469), .B2(n6823), .ZN(n6825)
         );
  INV_X1 U8593 ( .A(n6825), .ZN(n6826) );
  OAI21_X1 U8594 ( .B1(n6828), .B2(n10468), .A(n6826), .ZN(P2_U3463) );
  INV_X1 U8595 ( .A(n8628), .ZN(n8556) );
  AOI22_X1 U8596 ( .A1(n8556), .A2(n7115), .B1(n10475), .B2(
        P2_REG1_REG_4__SCAN_IN), .ZN(n6827) );
  OAI21_X1 U8597 ( .B1(n6828), .B2(n10475), .A(n6827), .ZN(P2_U3524) );
  NOR2_X1 U8598 ( .A1(n6835), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6830) );
  NOR2_X1 U8599 ( .A1(n6830), .A2(n6829), .ZN(n6833) );
  MUX2_X1 U8600 ( .A(n6831), .B(P1_REG1_REG_10__SCAN_IN), .S(n6873), .Z(n6832)
         );
  NOR2_X1 U8601 ( .A1(n6833), .A2(n6832), .ZN(n6869) );
  AOI21_X1 U8602 ( .B1(n6833), .B2(n6832), .A(n6869), .ZN(n6843) );
  NAND2_X1 U8603 ( .A1(n6873), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6836) );
  OAI21_X1 U8604 ( .B1(n6873), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6836), .ZN(
        n6837) );
  AOI211_X1 U8605 ( .C1(n6838), .C2(n6837), .A(n6872), .B(n10159), .ZN(n6839)
         );
  AOI21_X1 U8606 ( .B1(n10129), .B2(n6873), .A(n6839), .ZN(n6842) );
  NOR2_X1 U8607 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6840), .ZN(n7491) );
  AOI21_X1 U8608 ( .B1(n10079), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n7491), .ZN(
        n6841) );
  OAI211_X1 U8609 ( .C1(n6843), .C2(n10169), .A(n6842), .B(n6841), .ZN(
        P1_U3251) );
  INV_X1 U8610 ( .A(n6844), .ZN(n6848) );
  OAI21_X1 U8611 ( .B1(n6848), .B2(n6846), .A(n6845), .ZN(n6847) );
  OAI211_X1 U8612 ( .C1(n6849), .C2(n6848), .A(n8812), .B(n6847), .ZN(n6852)
         );
  AND2_X1 U8613 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10075) );
  INV_X1 U8614 ( .A(n10224), .ZN(n10181) );
  OAI22_X1 U8615 ( .A1(n8805), .A2(n10181), .B1(n8824), .B2(n10270), .ZN(n6850) );
  AOI211_X1 U8616 ( .C1(n8808), .C2(n10225), .A(n10075), .B(n6850), .ZN(n6851)
         );
  OAI211_X1 U8617 ( .C1(n8804), .C2(n10238), .A(n6852), .B(n6851), .ZN(
        P1_U3228) );
  INV_X1 U8618 ( .A(n8633), .ZN(n10453) );
  OAI21_X1 U8619 ( .B1(n6854), .B2(n7953), .A(n6853), .ZN(n10385) );
  AOI211_X1 U8620 ( .C1(n5984), .C2(n6856), .A(n10462), .B(n6855), .ZN(n10382)
         );
  INV_X1 U8621 ( .A(n7676), .ZN(n6861) );
  XNOR2_X1 U8622 ( .A(n6857), .B(n7953), .ZN(n6858) );
  NOR2_X1 U8623 ( .A1(n6858), .A2(n8510), .ZN(n6859) );
  AOI211_X1 U8624 ( .C1(n6861), .C2(n10385), .A(n6860), .B(n6859), .ZN(n10388)
         );
  INV_X1 U8625 ( .A(n10388), .ZN(n6862) );
  AOI211_X1 U8626 ( .C1(n10453), .C2(n10385), .A(n10382), .B(n6862), .ZN(n6868) );
  AOI22_X1 U8627 ( .A1(n8556), .A2(n5984), .B1(n10475), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n6863) );
  OAI21_X1 U8628 ( .B1(n6868), .B2(n10475), .A(n6863), .ZN(P2_U3523) );
  INV_X1 U8629 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6864) );
  OAI22_X1 U8630 ( .A1(n8678), .A2(n6865), .B1(n10469), .B2(n6864), .ZN(n6866)
         );
  INV_X1 U8631 ( .A(n6866), .ZN(n6867) );
  OAI21_X1 U8632 ( .B1(n6868), .B2(n10468), .A(n6867), .ZN(P2_U3460) );
  AOI21_X1 U8633 ( .B1(n4720), .B2(n6831), .A(n6869), .ZN(n6871) );
  AOI22_X1 U8634 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n7058), .B1(n7063), .B2(
        n5506), .ZN(n6870) );
  NOR2_X1 U8635 ( .A1(n6871), .A2(n6870), .ZN(n7057) );
  AOI21_X1 U8636 ( .B1(n6871), .B2(n6870), .A(n7057), .ZN(n6881) );
  AOI22_X1 U8637 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n7063), .B1(n7058), .B2(
        n7293), .ZN(n6875) );
  OAI21_X1 U8638 ( .B1(n6875), .B2(n6874), .A(n7062), .ZN(n6879) );
  INV_X1 U8639 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6877) );
  NAND2_X1 U8640 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7468) );
  NAND2_X1 U8641 ( .A1(n10129), .A2(n7063), .ZN(n6876) );
  OAI211_X1 U8642 ( .C1(n10172), .C2(n6877), .A(n7468), .B(n6876), .ZN(n6878)
         );
  AOI21_X1 U8643 ( .B1(n6879), .B2(n10086), .A(n6878), .ZN(n6880) );
  OAI21_X1 U8644 ( .B1(n6881), .B2(n10169), .A(n6880), .ZN(P1_U3252) );
  INV_X1 U8645 ( .A(n6882), .ZN(n6884) );
  INV_X1 U8646 ( .A(n8313), .ZN(n8304) );
  OAI222_X1 U8647 ( .A1(n8148), .A2(n6883), .B1(n7914), .B2(n6884), .C1(n8304), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  INV_X1 U8648 ( .A(n10128), .ZN(n9184) );
  OAI222_X1 U8649 ( .A1(n9553), .A2(n9726), .B1(n9560), .B2(n6884), .C1(n9184), 
        .C2(P1_U3084), .ZN(P1_U3337) );
  INV_X1 U8650 ( .A(n6885), .ZN(n6944) );
  AOI22_X1 U8651 ( .A1(n9177), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n6886), .ZN(n6887) );
  OAI21_X1 U8652 ( .B1(n6944), .B2(n9560), .A(n6887), .ZN(P1_U3336) );
  OR2_X1 U8653 ( .A1(n6888), .A2(n6889), .ZN(n6891) );
  AND2_X1 U8654 ( .A1(n6891), .A2(n6890), .ZN(n6895) );
  INV_X1 U8655 ( .A(n6892), .ZN(n6893) );
  AOI211_X1 U8656 ( .C1(n6895), .C2(n6894), .A(n8211), .B(n6893), .ZN(n6900)
         );
  AOI22_X1 U8657 ( .A1(n8216), .A2(n8255), .B1(n7252), .B2(n8230), .ZN(n6898)
         );
  INV_X1 U8658 ( .A(n7248), .ZN(n6896) );
  AOI22_X1 U8659 ( .A1(n8229), .A2(n6896), .B1(P2_REG3_REG_7__SCAN_IN), .B2(
        P2_U3152), .ZN(n6897) );
  OAI211_X1 U8660 ( .C1(n7859), .C2(n7966), .A(n6898), .B(n6897), .ZN(n6899)
         );
  OR2_X1 U8661 ( .A1(n6900), .A2(n6899), .ZN(P2_U3215) );
  OAI22_X1 U8662 ( .A1(n8206), .A2(n7144), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9842), .ZN(n6902) );
  OAI22_X1 U8663 ( .A1(n7827), .A2(n7263), .B1(n10448), .B2(n8220), .ZN(n6901)
         );
  AOI211_X1 U8664 ( .C1(n8217), .C2(n8256), .A(n6902), .B(n6901), .ZN(n6909)
         );
  INV_X1 U8665 ( .A(n6903), .ZN(n6904) );
  AOI21_X1 U8666 ( .B1(n6892), .B2(n6904), .A(n8211), .ZN(n6907) );
  NOR3_X1 U8667 ( .A1(n8224), .A2(n6905), .A3(n8225), .ZN(n6906) );
  OAI21_X1 U8668 ( .B1(n6907), .B2(n6906), .A(n7864), .ZN(n6908) );
  NAND2_X1 U8669 ( .A1(n6909), .A2(n6908), .ZN(P2_U3223) );
  OR2_X1 U8670 ( .A1(n6888), .A2(n6911), .ZN(n8233) );
  INV_X1 U8671 ( .A(n8233), .ZN(n6910) );
  AOI211_X1 U8672 ( .C1(n6911), .C2(n6888), .A(n8211), .B(n6910), .ZN(n6917)
         );
  INV_X1 U8673 ( .A(n8227), .ZN(n8169) );
  OR2_X1 U8674 ( .A1(n7966), .A2(n8515), .ZN(n6913) );
  NAND2_X1 U8675 ( .A1(n8259), .A2(n8543), .ZN(n6912) );
  AND2_X1 U8676 ( .A1(n6913), .A2(n6912), .ZN(n10372) );
  OAI22_X1 U8677 ( .A1(n8169), .A2(n10372), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6914), .ZN(n6916) );
  OAI22_X1 U8678 ( .A1(n10437), .A2(n8220), .B1(n8206), .B2(n10362), .ZN(n6915) );
  OR3_X1 U8679 ( .A1(n6917), .A2(n6916), .A3(n6915), .ZN(P2_U3229) );
  INV_X1 U8680 ( .A(n6918), .ZN(n6919) );
  INV_X1 U8681 ( .A(n10237), .ZN(n10203) );
  NAND2_X1 U8682 ( .A1(n7013), .A2(n6921), .ZN(n7032) );
  OAI21_X1 U8683 ( .B1(n8843), .B2(n6921), .A(n7032), .ZN(n10248) );
  OR2_X1 U8684 ( .A1(n6922), .A2(n7080), .ZN(n6925) );
  OR2_X1 U8685 ( .A1(n6923), .A2(n9076), .ZN(n6924) );
  NAND2_X1 U8686 ( .A1(n6925), .A2(n6924), .ZN(n10184) );
  INV_X1 U8687 ( .A(n10184), .ZN(n10235) );
  XNOR2_X1 U8688 ( .A(n7015), .B(n7014), .ZN(n6930) );
  NAND2_X1 U8689 ( .A1(n9125), .A2(n10206), .ZN(n6929) );
  NAND2_X1 U8690 ( .A1(n6927), .A2(n6926), .ZN(n6928) );
  INV_X1 U8691 ( .A(n10228), .ZN(n9424) );
  NAND2_X1 U8692 ( .A1(n6930), .A2(n9424), .ZN(n6934) );
  INV_X1 U8693 ( .A(n9067), .ZN(n6931) );
  AOI22_X1 U8694 ( .A1(n10226), .A2(n6932), .B1(n7020), .B2(n10223), .ZN(n6933) );
  OAI211_X1 U8695 ( .C1(n10248), .C2(n10235), .A(n6934), .B(n6933), .ZN(n10252) );
  INV_X1 U8696 ( .A(n7205), .ZN(n6935) );
  AOI211_X1 U8697 ( .C1(n6946), .C2(n7030), .A(n10306), .B(n6935), .ZN(n10249)
         );
  NOR2_X1 U8698 ( .A1(n10248), .A2(n6936), .ZN(n6937) );
  MUX2_X1 U8699 ( .A(n10249), .B(n6937), .S(n10206), .Z(n6938) );
  AOI211_X1 U8700 ( .C1(n10203), .C2(P1_REG3_REG_1__SCAN_IN), .A(n10252), .B(
        n6938), .ZN(n6943) );
  INV_X1 U8701 ( .A(n6939), .ZN(n6940) );
  NAND2_X1 U8702 ( .A1(n6941), .A2(n6940), .ZN(n7027) );
  INV_X2 U8703 ( .A(n10215), .ZN(n9403) );
  AOI22_X1 U8704 ( .A1(n10187), .A2(n7030), .B1(n10215), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n6942) );
  OAI21_X1 U8705 ( .B1(n6943), .B2(n10215), .A(n6942), .ZN(P1_U3290) );
  INV_X1 U8706 ( .A(n8324), .ZN(n8328) );
  OAI222_X1 U8707 ( .A1(n8148), .A2(n6945), .B1(n7914), .B2(n6944), .C1(n8328), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  OAI21_X1 U8708 ( .B1(n10221), .B2(n10187), .A(n6946), .ZN(n6951) );
  NOR2_X1 U8709 ( .A1(n10237), .A2(n6947), .ZN(n6948) );
  OAI21_X1 U8710 ( .B1(n6949), .B2(n6948), .A(n9403), .ZN(n6950) );
  OAI211_X1 U8711 ( .C1(n6542), .C2(n9403), .A(n6951), .B(n6950), .ZN(P1_U3291) );
  NOR2_X1 U8712 ( .A1(n10349), .A2(n6963), .ZN(n6952) );
  OR2_X1 U8713 ( .A1(n7146), .A2(n6952), .ZN(n7247) );
  XNOR2_X1 U8714 ( .A(n6953), .B(n6954), .ZN(n7257) );
  NAND2_X1 U8715 ( .A1(n7257), .A2(n10466), .ZN(n6959) );
  AOI21_X1 U8716 ( .B1(n6955), .B2(n8107), .A(n8510), .ZN(n6958) );
  OR2_X1 U8717 ( .A1(n6955), .A2(n8107), .ZN(n6957) );
  OAI22_X1 U8718 ( .A1(n7858), .A2(n8515), .B1(n7966), .B2(n8513), .ZN(n6956)
         );
  AOI21_X1 U8719 ( .B1(n6958), .B2(n6957), .A(n6956), .ZN(n7255) );
  OAI211_X1 U8720 ( .C1(n10462), .C2(n7247), .A(n6959), .B(n7255), .ZN(n6965)
         );
  INV_X1 U8721 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6960) );
  OAI22_X1 U8722 ( .A1(n8678), .A2(n6963), .B1(n10469), .B2(n6960), .ZN(n6961)
         );
  AOI21_X1 U8723 ( .B1(n6965), .B2(n10469), .A(n6961), .ZN(n6962) );
  INV_X1 U8724 ( .A(n6962), .ZN(P2_U3472) );
  OAI22_X1 U8725 ( .A1(n8628), .A2(n6963), .B1(n10477), .B2(n6671), .ZN(n6964)
         );
  AOI21_X1 U8726 ( .B1(n6965), .B2(n10477), .A(n6964), .ZN(n6966) );
  INV_X1 U8727 ( .A(n6966), .ZN(P2_U3527) );
  INV_X1 U8728 ( .A(n10202), .ZN(n6974) );
  XNOR2_X1 U8729 ( .A(n7001), .B(n6967), .ZN(n6968) );
  NAND2_X1 U8730 ( .A1(n6968), .A2(n6969), .ZN(n7000) );
  OAI21_X1 U8731 ( .B1(n6969), .B2(n6968), .A(n7000), .ZN(n6970) );
  NAND2_X1 U8732 ( .A1(n6970), .A2(n8812), .ZN(n6973) );
  AND2_X1 U8733 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9157) );
  INV_X1 U8734 ( .A(n9137), .ZN(n10210) );
  OAI22_X1 U8735 ( .A1(n8824), .A2(n10278), .B1(n8819), .B2(n10210), .ZN(n6971) );
  AOI211_X1 U8736 ( .C1(n8817), .C2(n10204), .A(n9157), .B(n6971), .ZN(n6972)
         );
  OAI211_X1 U8737 ( .C1(n8804), .C2(n6974), .A(n6973), .B(n6972), .ZN(P1_U3225) );
  INV_X1 U8738 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6976) );
  INV_X1 U8739 ( .A(n6975), .ZN(n6977) );
  INV_X1 U8740 ( .A(n9176), .ZN(n10162) );
  OAI222_X1 U8741 ( .A1(n9562), .A2(n6976), .B1(n9560), .B2(n6977), .C1(
        P1_U3084), .C2(n10162), .ZN(P1_U3335) );
  INV_X1 U8742 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6978) );
  OAI222_X1 U8743 ( .A1(n8148), .A2(n6978), .B1(n8686), .B2(n6977), .C1(
        P2_U3152), .C2(n8344), .ZN(P2_U3340) );
  NAND2_X1 U8744 ( .A1(n8272), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6981) );
  OAI21_X1 U8745 ( .B1(n8272), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6981), .ZN(
        n8264) );
  AOI21_X1 U8746 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n8272), .A(n8263), .ZN(
        n6984) );
  NAND2_X1 U8747 ( .A1(n7188), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6982) );
  OAI21_X1 U8748 ( .B1(n7188), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6982), .ZN(
        n6983) );
  AOI211_X1 U8749 ( .C1(n6984), .C2(n6983), .A(n7184), .B(n9988), .ZN(n6999)
         );
  NOR2_X1 U8750 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9692), .ZN(n6985) );
  AOI21_X1 U8751 ( .B1(n10333), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n6985), .ZN(
        n6996) );
  MUX2_X1 U8752 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n6986), .S(n8272), .Z(n8270)
         );
  INV_X1 U8753 ( .A(n6987), .ZN(n6988) );
  OAI21_X1 U8754 ( .B1(n6990), .B2(n6989), .A(n6988), .ZN(n8271) );
  NAND2_X1 U8755 ( .A1(n8270), .A2(n8271), .ZN(n8269) );
  OAI21_X1 U8756 ( .B1(n6991), .B2(n6986), .A(n8269), .ZN(n6994) );
  MUX2_X1 U8757 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n6992), .S(n7188), .Z(n6993)
         );
  NAND2_X1 U8758 ( .A1(n6993), .A2(n6994), .ZN(n7189) );
  OAI211_X1 U8759 ( .C1(n6994), .C2(n6993), .A(n10330), .B(n7189), .ZN(n6995)
         );
  OAI211_X1 U8760 ( .C1(n10327), .C2(n6997), .A(n6996), .B(n6995), .ZN(n6998)
         );
  OR2_X1 U8761 ( .A1(n6999), .A2(n6998), .ZN(P2_U3255) );
  OAI21_X1 U8762 ( .B1(n7002), .B2(n7001), .A(n7000), .ZN(n7006) );
  XNOR2_X1 U8763 ( .A(n7004), .B(n7003), .ZN(n7005) );
  XNOR2_X1 U8764 ( .A(n7006), .B(n7005), .ZN(n7012) );
  NOR2_X1 U8765 ( .A1(n10189), .A2(n10304), .ZN(n10283) );
  AOI21_X1 U8766 ( .B1(n8795), .B2(n10283), .A(n7007), .ZN(n7008) );
  OAI21_X1 U8767 ( .B1(n8819), .B2(n10181), .A(n7008), .ZN(n7010) );
  NOR2_X1 U8768 ( .A1(n8804), .A2(n10185), .ZN(n7009) );
  AOI211_X1 U8769 ( .C1(n8817), .C2(n10174), .A(n7010), .B(n7009), .ZN(n7011)
         );
  OAI21_X1 U8770 ( .B1(n7012), .B2(n8773), .A(n7011), .ZN(P1_U3237) );
  INV_X1 U8771 ( .A(n7013), .ZN(n7015) );
  NAND2_X1 U8772 ( .A1(n7015), .A2(n7014), .ZN(n7017) );
  NAND2_X1 U8773 ( .A1(n7020), .A2(n10257), .ZN(n9080) );
  NAND2_X1 U8774 ( .A1(n7021), .A2(n9082), .ZN(n7221) );
  NAND2_X1 U8775 ( .A1(n10225), .A2(n10264), .ZN(n8902) );
  NAND2_X1 U8776 ( .A1(n9083), .A2(n8902), .ZN(n7035) );
  INV_X1 U8777 ( .A(n7035), .ZN(n8839) );
  OR2_X1 U8778 ( .A1(n9137), .A2(n10270), .ZN(n8907) );
  INV_X1 U8779 ( .A(n8907), .ZN(n9090) );
  NAND2_X1 U8780 ( .A1(n9137), .A2(n10270), .ZN(n10227) );
  OR2_X1 U8781 ( .A1(n10204), .A2(n10189), .ZN(n7042) );
  OR2_X1 U8782 ( .A1(n10224), .A2(n10278), .ZN(n10176) );
  NAND2_X1 U8783 ( .A1(n7042), .A2(n10176), .ZN(n9089) );
  AND2_X1 U8784 ( .A1(n10224), .A2(n10278), .ZN(n8904) );
  NAND2_X1 U8785 ( .A1(n8904), .A2(n7042), .ZN(n7022) );
  NAND2_X1 U8786 ( .A1(n10204), .A2(n10189), .ZN(n8908) );
  OR2_X1 U8787 ( .A1(n10174), .A2(n10292), .ZN(n8936) );
  NAND2_X1 U8788 ( .A1(n10174), .A2(n10292), .ZN(n8935) );
  NAND2_X1 U8789 ( .A1(n8936), .A2(n8935), .ZN(n7072) );
  OAI21_X1 U8790 ( .B1(n7024), .B2(n7023), .A(n7075), .ZN(n7025) );
  AOI222_X1 U8791 ( .A1(n9424), .A2(n7025), .B1(n9136), .B2(n10223), .C1(
        n10204), .C2(n10226), .ZN(n10291) );
  INV_X1 U8792 ( .A(n10292), .ZN(n8695) );
  OAI22_X1 U8793 ( .A1(n9403), .A2(n7026), .B1(n8696), .B2(n10237), .ZN(n7029)
         );
  NAND2_X1 U8794 ( .A1(n7216), .A2(n10264), .ZN(n10217) );
  OAI211_X1 U8795 ( .C1(n10191), .C2(n10292), .A(n10198), .B(n7239), .ZN(
        n10290) );
  NOR2_X1 U8796 ( .A1(n7027), .A2(n10206), .ZN(n10024) );
  INV_X1 U8797 ( .A(n10024), .ZN(n7565) );
  NOR2_X1 U8798 ( .A1(n10290), .A2(n7565), .ZN(n7028) );
  AOI211_X1 U8799 ( .C1(n10187), .C2(n8695), .A(n7029), .B(n7028), .ZN(n7046)
         );
  NAND2_X1 U8800 ( .A1(n6920), .A2(n7030), .ZN(n7031) );
  OR2_X1 U8801 ( .A1(n7020), .A2(n7018), .ZN(n7034) );
  NAND2_X1 U8802 ( .A1(n7214), .A2(n7035), .ZN(n7037) );
  OR2_X1 U8803 ( .A1(n10225), .A2(n7220), .ZN(n7036) );
  NAND2_X1 U8804 ( .A1(n7037), .A2(n7036), .ZN(n10216) );
  NAND2_X1 U8805 ( .A1(n8907), .A2(n10227), .ZN(n10229) );
  NAND2_X1 U8806 ( .A1(n10216), .A2(n10229), .ZN(n7040) );
  OR2_X1 U8807 ( .A1(n9137), .A2(n7038), .ZN(n7039) );
  NAND2_X1 U8808 ( .A1(n7040), .A2(n7039), .ZN(n10196) );
  XNOR2_X1 U8809 ( .A(n10224), .B(n10200), .ZN(n10208) );
  INV_X1 U8810 ( .A(n10208), .ZN(n7041) );
  NAND2_X1 U8811 ( .A1(n7042), .A2(n8908), .ZN(n10178) );
  INV_X1 U8812 ( .A(n10189), .ZN(n10188) );
  XNOR2_X1 U8813 ( .A(n7073), .B(n7072), .ZN(n10294) );
  AND2_X1 U8814 ( .A1(n7044), .A2(n7043), .ZN(n10213) );
  NAND2_X1 U8815 ( .A1(n9403), .A2(n10213), .ZN(n9428) );
  INV_X1 U8816 ( .A(n9428), .ZN(n7790) );
  NAND2_X1 U8817 ( .A1(n10294), .A2(n7790), .ZN(n7045) );
  OAI211_X1 U8818 ( .C1(n10291), .C2(n10215), .A(n7046), .B(n7045), .ZN(
        P1_U3284) );
  OAI211_X1 U8819 ( .C1(n7049), .C2(n7048), .A(n7047), .B(n8235), .ZN(n7053)
         );
  OAI22_X1 U8820 ( .A1(n8206), .A2(n7271), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9692), .ZN(n7051) );
  OAI22_X1 U8821 ( .A1(n7364), .A2(n7827), .B1(n7859), .B2(n7263), .ZN(n7050)
         );
  AOI211_X1 U8822 ( .C1(n7274), .C2(n8230), .A(n7051), .B(n7050), .ZN(n7052)
         );
  NAND2_X1 U8823 ( .A1(n7053), .A2(n7052), .ZN(P2_U3219) );
  INV_X1 U8824 ( .A(n7054), .ZN(n7056) );
  OAI222_X1 U8825 ( .A1(n8148), .A2(n7055), .B1(n8686), .B2(n7056), .C1(
        P2_U3152), .C2(n8350), .ZN(P2_U3339) );
  OAI222_X1 U8826 ( .A1(n9562), .A2(n9748), .B1(n9560), .B2(n7056), .C1(n9332), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  AOI21_X1 U8827 ( .B1(n5506), .B2(n7058), .A(n7057), .ZN(n7060) );
  AOI22_X1 U8828 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n7398), .B1(n7068), .B2(
        n5529), .ZN(n7059) );
  NOR2_X1 U8829 ( .A1(n7060), .A2(n7059), .ZN(n7397) );
  AOI21_X1 U8830 ( .B1(n7060), .B2(n7059), .A(n7397), .ZN(n7070) );
  INV_X1 U8831 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7061) );
  NAND2_X1 U8832 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7638) );
  OAI21_X1 U8833 ( .B1(n10172), .B2(n7061), .A(n7638), .ZN(n7067) );
  OAI21_X1 U8834 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7063), .A(n7062), .ZN(
        n7065) );
  NAND2_X1 U8835 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7068), .ZN(n7406) );
  OAI21_X1 U8836 ( .B1(n7068), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7406), .ZN(
        n7064) );
  NOR2_X1 U8837 ( .A1(n7064), .A2(n7065), .ZN(n7404) );
  AOI211_X1 U8838 ( .C1(n7065), .C2(n7064), .A(n7404), .B(n10159), .ZN(n7066)
         );
  AOI211_X1 U8839 ( .C1(n10129), .C2(n7068), .A(n7067), .B(n7066), .ZN(n7069)
         );
  OAI21_X1 U8840 ( .B1(n7070), .B2(n10169), .A(n7069), .ZN(P1_U3253) );
  NOR2_X1 U8841 ( .A1(n10174), .A2(n8695), .ZN(n7071) );
  OR2_X1 U8842 ( .A1(n9136), .A2(n7128), .ZN(n8940) );
  NAND2_X1 U8843 ( .A1(n9136), .A2(n7128), .ZN(n7231) );
  NAND2_X1 U8844 ( .A1(n8940), .A2(n7231), .ZN(n8845) );
  NAND2_X1 U8845 ( .A1(n7228), .A2(n8845), .ZN(n7230) );
  INV_X1 U8846 ( .A(n7128), .ZN(n7244) );
  NAND2_X1 U8847 ( .A1(n9136), .A2(n7244), .ZN(n7074) );
  NAND2_X1 U8848 ( .A1(n7230), .A2(n7074), .ZN(n7163) );
  INV_X1 U8849 ( .A(n7322), .ZN(n10305) );
  OR2_X1 U8850 ( .A1(n9135), .A2(n10305), .ZN(n8949) );
  NAND2_X1 U8851 ( .A1(n9135), .A2(n10305), .ZN(n8943) );
  AND2_X1 U8852 ( .A1(n8949), .A2(n8943), .ZN(n8846) );
  XNOR2_X1 U8853 ( .A(n7163), .B(n8846), .ZN(n10310) );
  NAND2_X1 U8854 ( .A1(n7168), .A2(n7231), .ZN(n7076) );
  XNOR2_X1 U8855 ( .A(n7076), .B(n8846), .ZN(n7078) );
  AOI22_X1 U8856 ( .A1(n10226), .A2(n9136), .B1(n9134), .B2(n10223), .ZN(n7077) );
  OAI21_X1 U8857 ( .B1(n7078), .B2(n10228), .A(n7077), .ZN(n7079) );
  AOI21_X1 U8858 ( .B1(n10310), .B2(n10184), .A(n7079), .ZN(n10312) );
  NAND3_X1 U8859 ( .A1(n9403), .A2(n7080), .A3(n10206), .ZN(n7759) );
  INV_X1 U8860 ( .A(n7759), .ZN(n10222) );
  NAND2_X1 U8861 ( .A1(n7241), .A2(n7322), .ZN(n7081) );
  NAND2_X1 U8862 ( .A1(n7176), .A2(n7081), .ZN(n10307) );
  INV_X1 U8863 ( .A(n10221), .ZN(n7754) );
  OAI22_X1 U8864 ( .A1(n9403), .A2(n7082), .B1(n7324), .B2(n10237), .ZN(n7083)
         );
  AOI21_X1 U8865 ( .B1(n10187), .B2(n7322), .A(n7083), .ZN(n7084) );
  OAI21_X1 U8866 ( .B1(n10307), .B2(n7754), .A(n7084), .ZN(n7085) );
  AOI21_X1 U8867 ( .B1(n10310), .B2(n10222), .A(n7085), .ZN(n7086) );
  OAI21_X1 U8868 ( .B1(n10312), .B2(n10215), .A(n7086), .ZN(P1_U3282) );
  INV_X1 U8869 ( .A(n7087), .ZN(n8105) );
  INV_X1 U8870 ( .A(n6809), .ZN(n7088) );
  XNOR2_X1 U8871 ( .A(n8105), .B(n7088), .ZN(n7089) );
  NAND2_X1 U8872 ( .A1(n7089), .A2(n10369), .ZN(n7092) );
  INV_X1 U8873 ( .A(n7090), .ZN(n7091) );
  NAND2_X1 U8874 ( .A1(n7092), .A2(n7091), .ZN(n7896) );
  NOR2_X1 U8875 ( .A1(n10376), .A2(n5938), .ZN(n7095) );
  INV_X1 U8876 ( .A(n10383), .ZN(n8361) );
  OAI211_X1 U8877 ( .C1(n7903), .C2(n10430), .A(n10360), .B(n7093), .ZN(n7895)
         );
  OAI22_X1 U8878 ( .A1(n8361), .A2(n7895), .B1(n9841), .B2(n8468), .ZN(n7094)
         );
  AOI211_X1 U8879 ( .C1(n10376), .C2(n7896), .A(n7095), .B(n7094), .ZN(n7100)
         );
  OAI21_X1 U8880 ( .B1(n7087), .B2(n7097), .A(n7096), .ZN(n7898) );
  AOI22_X1 U8881 ( .A1(n10352), .A2(n7898), .B1(n10381), .B2(n7098), .ZN(n7099) );
  NAND2_X1 U8882 ( .A1(n7100), .A2(n7099), .ZN(P2_U3295) );
  NOR2_X1 U8883 ( .A1(n10376), .A2(n7101), .ZN(n7104) );
  OAI22_X1 U8884 ( .A1(n8361), .A2(n7102), .B1(n9860), .B2(n8468), .ZN(n7103)
         );
  AOI211_X1 U8885 ( .C1(n10376), .C2(n7105), .A(n7104), .B(n7103), .ZN(n7109)
         );
  AOI22_X1 U8886 ( .A1(n10352), .A2(n7107), .B1(n10381), .B2(n7106), .ZN(n7108) );
  NAND2_X1 U8887 ( .A1(n7109), .A2(n7108), .ZN(P2_U3294) );
  NOR2_X1 U8888 ( .A1(n10376), .A2(n6642), .ZN(n7113) );
  OAI22_X1 U8889 ( .A1(n8361), .A2(n7111), .B1(n7110), .B2(n8468), .ZN(n7112)
         );
  AOI211_X1 U8890 ( .C1(n10376), .C2(n7114), .A(n7113), .B(n7112), .ZN(n7118)
         );
  AOI22_X1 U8891 ( .A1(n10352), .A2(n7116), .B1(n10381), .B2(n7115), .ZN(n7117) );
  NAND2_X1 U8892 ( .A1(n7118), .A2(n7117), .ZN(P2_U3292) );
  NAND2_X1 U8893 ( .A1(n6809), .A2(n7943), .ZN(n8100) );
  INV_X1 U8894 ( .A(n8100), .ZN(n10433) );
  OAI21_X1 U8895 ( .B1(n8551), .B2(n10381), .A(n7119), .ZN(n7123) );
  AOI22_X1 U8896 ( .A1(n8100), .A2(n10369), .B1(n8544), .B2(n8261), .ZN(n10429) );
  OAI21_X1 U8897 ( .B1(n9752), .B2(n8468), .A(n10429), .ZN(n7121) );
  NOR2_X1 U8898 ( .A1(n10376), .A2(n5953), .ZN(n7120) );
  AOI21_X1 U8899 ( .B1(n10376), .B2(n7121), .A(n7120), .ZN(n7122) );
  OAI211_X1 U8900 ( .C1(n10433), .C2(n8553), .A(n7123), .B(n7122), .ZN(
        P2_U3296) );
  XOR2_X1 U8901 ( .A(n7125), .B(n7124), .Z(n7126) );
  XNOR2_X1 U8902 ( .A(n7127), .B(n7126), .ZN(n7134) );
  OR2_X1 U8903 ( .A1(n7128), .A2(n10304), .ZN(n10298) );
  INV_X1 U8904 ( .A(n10298), .ZN(n7129) );
  AOI22_X1 U8905 ( .A1(n8817), .A2(n9135), .B1(n7129), .B2(n8795), .ZN(n7133)
         );
  INV_X1 U8906 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7130) );
  NOR2_X1 U8907 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7130), .ZN(n10081) );
  NOR2_X1 U8908 ( .A1(n8804), .A2(n7237), .ZN(n7131) );
  AOI211_X1 U8909 ( .C1(n8808), .C2(n10174), .A(n10081), .B(n7131), .ZN(n7132)
         );
  OAI211_X1 U8910 ( .C1(n7134), .C2(n8773), .A(n7133), .B(n7132), .ZN(P1_U3219) );
  NAND2_X1 U8911 ( .A1(n7135), .A2(n8108), .ZN(n7136) );
  NAND2_X1 U8912 ( .A1(n7137), .A2(n7136), .ZN(n10447) );
  OR2_X1 U8913 ( .A1(n10389), .A2(n7138), .ZN(n10380) );
  OAI21_X1 U8914 ( .B1(n7140), .B2(n8108), .A(n7139), .ZN(n7142) );
  OAI22_X1 U8915 ( .A1(n8225), .A2(n8513), .B1(n7263), .B2(n8515), .ZN(n7141)
         );
  AOI21_X1 U8916 ( .B1(n7142), .B2(n10369), .A(n7141), .ZN(n7143) );
  OAI21_X1 U8917 ( .B1(n10447), .B2(n7676), .A(n7143), .ZN(n10450) );
  NAND2_X1 U8918 ( .A1(n10450), .A2(n10376), .ZN(n7151) );
  INV_X1 U8919 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7145) );
  OAI22_X1 U8920 ( .A1(n10376), .A2(n7145), .B1(n7144), .B2(n8468), .ZN(n7149)
         );
  INV_X1 U8921 ( .A(n8551), .ZN(n7894) );
  OR2_X1 U8922 ( .A1(n7146), .A2(n10448), .ZN(n7147) );
  NAND2_X1 U8923 ( .A1(n7351), .A2(n7147), .ZN(n10449) );
  NOR2_X1 U8924 ( .A1(n7894), .A2(n10449), .ZN(n7148) );
  AOI211_X1 U8925 ( .C1(n10381), .C2(n7975), .A(n7149), .B(n7148), .ZN(n7150)
         );
  OAI211_X1 U8926 ( .C1(n10447), .C2(n10380), .A(n7151), .B(n7150), .ZN(
        P2_U3288) );
  INV_X1 U8927 ( .A(n7152), .ZN(n7153) );
  AOI21_X1 U8928 ( .B1(n7047), .B2(n7153), .A(n8211), .ZN(n7157) );
  NOR3_X1 U8929 ( .A1(n8224), .A2(n7154), .A3(n7346), .ZN(n7156) );
  OAI21_X1 U8930 ( .B1(n7157), .B2(n7156), .A(n7155), .ZN(n7161) );
  OAI22_X1 U8931 ( .A1(n8206), .A2(n7438), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6090), .ZN(n7159) );
  OAI22_X1 U8932 ( .A1(n7346), .A2(n7859), .B1(n7827), .B2(n8004), .ZN(n7158)
         );
  AOI211_X1 U8933 ( .C1(n7382), .C2(n8230), .A(n7159), .B(n7158), .ZN(n7160)
         );
  NAND2_X1 U8934 ( .A1(n7161), .A2(n7160), .ZN(P2_U3238) );
  OR2_X1 U8935 ( .A1(n9135), .A2(n7322), .ZN(n7162) );
  NAND2_X1 U8936 ( .A1(n9135), .A2(n7322), .ZN(n7164) );
  NAND2_X1 U8937 ( .A1(n10002), .A2(n9134), .ZN(n8953) );
  NAND2_X1 U8938 ( .A1(n7166), .A2(n8848), .ZN(n7167) );
  NAND2_X1 U8939 ( .A1(n7285), .A2(n7167), .ZN(n10004) );
  AND2_X1 U8940 ( .A1(n7231), .A2(n8943), .ZN(n8884) );
  NAND2_X1 U8941 ( .A1(n7169), .A2(n8949), .ZN(n7170) );
  INV_X1 U8942 ( .A(n8953), .ZN(n8889) );
  AOI21_X1 U8943 ( .B1(n7170), .B2(n7165), .A(n10228), .ZN(n7171) );
  OAI21_X1 U8944 ( .B1(n7287), .B2(n8889), .A(n7171), .ZN(n7173) );
  INV_X1 U8945 ( .A(n7639), .ZN(n10014) );
  AOI22_X1 U8946 ( .A1(n10014), .A2(n10223), .B1(n10226), .B2(n9135), .ZN(
        n7172) );
  NAND2_X1 U8947 ( .A1(n7173), .A2(n7172), .ZN(n7174) );
  AOI21_X1 U8948 ( .B1(n10004), .B2(n10184), .A(n7174), .ZN(n10006) );
  NAND2_X1 U8949 ( .A1(n7176), .A2(n7503), .ZN(n7175) );
  NAND2_X1 U8950 ( .A1(n7175), .A2(n10198), .ZN(n7177) );
  OR2_X1 U8951 ( .A1(n7177), .A2(n7291), .ZN(n10001) );
  OAI22_X1 U8952 ( .A1(n9403), .A2(n7178), .B1(n7495), .B2(n10237), .ZN(n7179)
         );
  AOI21_X1 U8953 ( .B1(n10187), .B2(n7503), .A(n7179), .ZN(n7180) );
  OAI21_X1 U8954 ( .B1(n10001), .B2(n7565), .A(n7180), .ZN(n7181) );
  AOI21_X1 U8955 ( .B1(n10004), .B2(n10222), .A(n7181), .ZN(n7182) );
  OAI21_X1 U8956 ( .B1(n10006), .B2(n10215), .A(n7182), .ZN(P1_U3281) );
  AOI22_X1 U8957 ( .A1(n7307), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n6089), .B2(
        n7183), .ZN(n7186) );
  OAI21_X1 U8958 ( .B1(n7186), .B2(n7185), .A(n7306), .ZN(n7198) );
  MUX2_X1 U8959 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n7187), .S(n7307), .Z(n7192)
         );
  NAND2_X1 U8960 ( .A1(n7188), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7190) );
  NAND2_X1 U8961 ( .A1(n7190), .A2(n7189), .ZN(n7191) );
  NAND2_X1 U8962 ( .A1(n7192), .A2(n7191), .ZN(n7298) );
  OAI21_X1 U8963 ( .B1(n7192), .B2(n7191), .A(n7298), .ZN(n7196) );
  NAND2_X1 U8964 ( .A1(n9994), .A2(n7307), .ZN(n7195) );
  NOR2_X1 U8965 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6090), .ZN(n7193) );
  AOI21_X1 U8966 ( .B1(n10333), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7193), .ZN(
        n7194) );
  OAI211_X1 U8967 ( .C1(n10328), .C2(n7196), .A(n7195), .B(n7194), .ZN(n7197)
         );
  AOI21_X1 U8968 ( .B1(n10331), .B2(n7198), .A(n7197), .ZN(n7199) );
  INV_X1 U8969 ( .A(n7199), .ZN(P2_U3256) );
  INV_X1 U8970 ( .A(n7200), .ZN(n7201) );
  AOI21_X1 U8971 ( .B1(n8838), .B2(n7202), .A(n7201), .ZN(n10256) );
  OAI22_X1 U8972 ( .A1(n9403), .A2(n7204), .B1(n7203), .B2(n10237), .ZN(n7208)
         );
  AND2_X1 U8973 ( .A1(n7018), .A2(n7205), .ZN(n7206) );
  OR2_X1 U8974 ( .A1(n7206), .A2(n7216), .ZN(n10258) );
  NOR2_X1 U8975 ( .A1(n7754), .A2(n10258), .ZN(n7207) );
  AOI211_X1 U8976 ( .C1(n10187), .C2(n7018), .A(n7208), .B(n7207), .ZN(n7213)
         );
  AOI22_X1 U8977 ( .A1(n10226), .A2(n6920), .B1(n10225), .B2(n10223), .ZN(
        n7211) );
  NAND2_X1 U8978 ( .A1(n7209), .A2(n9424), .ZN(n7210) );
  OAI211_X1 U8979 ( .C1(n10256), .C2(n10235), .A(n7211), .B(n7210), .ZN(n10259) );
  NAND2_X1 U8980 ( .A1(n10259), .A2(n9403), .ZN(n7212) );
  OAI211_X1 U8981 ( .C1(n10256), .C2(n7759), .A(n7213), .B(n7212), .ZN(
        P1_U3289) );
  XNOR2_X1 U8982 ( .A(n7214), .B(n8839), .ZN(n10263) );
  OAI22_X1 U8983 ( .A1(n9403), .A2(n7215), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10237), .ZN(n7219) );
  OR2_X1 U8984 ( .A1(n7216), .A2(n10264), .ZN(n7217) );
  NAND2_X1 U8985 ( .A1(n10217), .A2(n7217), .ZN(n10265) );
  NOR2_X1 U8986 ( .A1(n7754), .A2(n10265), .ZN(n7218) );
  AOI211_X1 U8987 ( .C1(n10187), .C2(n7220), .A(n7219), .B(n7218), .ZN(n7227)
         );
  AOI22_X1 U8988 ( .A1(n10226), .A2(n7020), .B1(n9137), .B2(n10223), .ZN(n7225) );
  OAI21_X1 U8989 ( .B1(n8839), .B2(n7221), .A(n7222), .ZN(n7223) );
  NAND2_X1 U8990 ( .A1(n7223), .A2(n9424), .ZN(n7224) );
  OAI211_X1 U8991 ( .C1(n10263), .C2(n10235), .A(n7225), .B(n7224), .ZN(n10266) );
  NAND2_X1 U8992 ( .A1(n10266), .A2(n9403), .ZN(n7226) );
  OAI211_X1 U8993 ( .C1(n10263), .C2(n7759), .A(n7227), .B(n7226), .ZN(
        P1_U3288) );
  OR2_X1 U8994 ( .A1(n7228), .A2(n8845), .ZN(n7229) );
  NAND2_X1 U8995 ( .A1(n7230), .A2(n7229), .ZN(n10297) );
  AOI22_X1 U8996 ( .A1(n10223), .A2(n9135), .B1(n10174), .B2(n10226), .ZN(
        n7236) );
  INV_X1 U8997 ( .A(n7231), .ZN(n8942) );
  INV_X1 U8998 ( .A(n7232), .ZN(n7233) );
  AOI21_X1 U8999 ( .B1(n7233), .B2(n8845), .A(n10228), .ZN(n7234) );
  OAI21_X1 U9000 ( .B1(n8942), .B2(n7168), .A(n7234), .ZN(n7235) );
  OAI211_X1 U9001 ( .C1(n10297), .C2(n10235), .A(n7236), .B(n7235), .ZN(n10300) );
  NAND2_X1 U9002 ( .A1(n10300), .A2(n9403), .ZN(n7246) );
  OAI22_X1 U9003 ( .A1(n9403), .A2(n7238), .B1(n7237), .B2(n10237), .ZN(n7243)
         );
  NAND2_X1 U9004 ( .A1(n7239), .A2(n7244), .ZN(n7240) );
  NAND2_X1 U9005 ( .A1(n7241), .A2(n7240), .ZN(n10299) );
  NOR2_X1 U9006 ( .A1(n10299), .A2(n7754), .ZN(n7242) );
  AOI211_X1 U9007 ( .C1(n10187), .C2(n7244), .A(n7243), .B(n7242), .ZN(n7245)
         );
  OAI211_X1 U9008 ( .C1(n10297), .C2(n7759), .A(n7246), .B(n7245), .ZN(
        P1_U3283) );
  INV_X1 U9009 ( .A(n7247), .ZN(n7251) );
  OAI22_X1 U9010 ( .A1(n10376), .A2(n7249), .B1(n7248), .B2(n8468), .ZN(n7250)
         );
  AOI21_X1 U9011 ( .B1(n8551), .B2(n7251), .A(n7250), .ZN(n7254) );
  NAND2_X1 U9012 ( .A1(n10381), .A2(n7252), .ZN(n7253) );
  OAI211_X1 U9013 ( .C1(n7255), .C2(n10389), .A(n7254), .B(n7253), .ZN(n7256)
         );
  AOI21_X1 U9014 ( .B1(n10352), .B2(n7257), .A(n7256), .ZN(n7258) );
  INV_X1 U9015 ( .A(n7258), .ZN(P2_U3289) );
  INV_X1 U9016 ( .A(n7259), .ZN(n7279) );
  OAI222_X1 U9017 ( .A1(n8148), .A2(n7260), .B1(n8686), .B2(n7279), .C1(n8129), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  XNOR2_X1 U9018 ( .A(n7261), .B(n6081), .ZN(n7262) );
  NAND2_X1 U9019 ( .A1(n7262), .A2(n10369), .ZN(n7266) );
  OAI22_X1 U9020 ( .A1(n7364), .A2(n8515), .B1(n7263), .B2(n8513), .ZN(n7264)
         );
  INV_X1 U9021 ( .A(n7264), .ZN(n7265) );
  NAND2_X1 U9022 ( .A1(n7266), .A2(n7265), .ZN(n10457) );
  INV_X1 U9023 ( .A(n10457), .ZN(n7278) );
  INV_X1 U9024 ( .A(n7267), .ZN(n7268) );
  AOI21_X1 U9025 ( .B1(n8111), .B2(n7269), .A(n7268), .ZN(n10458) );
  AND2_X1 U9026 ( .A1(n7352), .A2(n7274), .ZN(n7270) );
  OR2_X1 U9027 ( .A1(n7270), .A2(n7379), .ZN(n10455) );
  OAI22_X1 U9028 ( .A1(n10376), .A2(n7272), .B1(n7271), .B2(n8468), .ZN(n7273)
         );
  AOI21_X1 U9029 ( .B1(n10381), .B2(n7274), .A(n7273), .ZN(n7275) );
  OAI21_X1 U9030 ( .B1(n7894), .B2(n10455), .A(n7275), .ZN(n7276) );
  AOI21_X1 U9031 ( .B1(n10458), .B2(n10352), .A(n7276), .ZN(n7277) );
  OAI21_X1 U9032 ( .B1(n8548), .B2(n7278), .A(n7277), .ZN(P2_U3286) );
  OAI222_X1 U9033 ( .A1(n9562), .A2(n7280), .B1(P1_U3084), .B2(n9437), .C1(
        n9560), .C2(n7279), .ZN(P1_U3333) );
  INV_X1 U9034 ( .A(n7281), .ZN(n7283) );
  OAI222_X1 U9035 ( .A1(n8148), .A2(n7282), .B1(n8686), .B2(n7283), .C1(n8131), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  OAI222_X1 U9036 ( .A1(n9562), .A2(n9702), .B1(P1_U3084), .B2(n9076), .C1(
        n9560), .C2(n7283), .ZN(P1_U3332) );
  OR2_X1 U9037 ( .A1(n9134), .A2(n7503), .ZN(n7284) );
  NAND2_X1 U9038 ( .A1(n7285), .A2(n7284), .ZN(n7559) );
  XNOR2_X1 U9039 ( .A(n7558), .B(n7639), .ZN(n8971) );
  INV_X1 U9040 ( .A(n8971), .ZN(n7286) );
  XNOR2_X1 U9041 ( .A(n7559), .B(n7286), .ZN(n9522) );
  XNOR2_X1 U9042 ( .A(n7554), .B(n8971), .ZN(n7289) );
  INV_X1 U9043 ( .A(n7555), .ZN(n9133) );
  AOI22_X1 U9044 ( .A1(n9133), .A2(n10223), .B1(n10226), .B2(n9134), .ZN(n7288) );
  OAI21_X1 U9045 ( .B1(n7289), .B2(n10228), .A(n7288), .ZN(n7290) );
  AOI21_X1 U9046 ( .B1(n9522), .B2(n10184), .A(n7290), .ZN(n9527) );
  INV_X1 U9047 ( .A(n7291), .ZN(n7292) );
  NAND2_X1 U9048 ( .A1(n7291), .A2(n7558), .ZN(n7563) );
  INV_X1 U9049 ( .A(n7563), .ZN(n10022) );
  AOI21_X1 U9050 ( .B1(n9523), .B2(n7292), .A(n10022), .ZN(n9525) );
  NOR2_X1 U9051 ( .A1(n10239), .A2(n7558), .ZN(n7295) );
  OAI22_X1 U9052 ( .A1(n9403), .A2(n7293), .B1(n7471), .B2(n10237), .ZN(n7294)
         );
  AOI211_X1 U9053 ( .C1(n9525), .C2(n10221), .A(n7295), .B(n7294), .ZN(n7297)
         );
  NAND2_X1 U9054 ( .A1(n9522), .A2(n10222), .ZN(n7296) );
  OAI211_X1 U9055 ( .C1(n9527), .C2(n10215), .A(n7297), .B(n7296), .ZN(
        P1_U3280) );
  INV_X1 U9056 ( .A(n7450), .ZN(n7453) );
  INV_X1 U9057 ( .A(n7298), .ZN(n7299) );
  AOI21_X1 U9058 ( .B1(n7307), .B2(P2_REG1_REG_11__SCAN_IN), .A(n7299), .ZN(
        n7301) );
  MUX2_X1 U9059 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6111), .S(n7450), .Z(n7300)
         );
  NAND2_X1 U9060 ( .A1(n7301), .A2(n7300), .ZN(n7455) );
  OAI21_X1 U9061 ( .B1(n7301), .B2(n7300), .A(n7455), .ZN(n7305) );
  NAND2_X1 U9062 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7333) );
  INV_X1 U9063 ( .A(n7333), .ZN(n7304) );
  INV_X1 U9064 ( .A(n10333), .ZN(n7581) );
  INV_X1 U9065 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7302) );
  NOR2_X1 U9066 ( .A1(n7581), .A2(n7302), .ZN(n7303) );
  AOI211_X1 U9067 ( .C1(n10330), .C2(n7305), .A(n7304), .B(n7303), .ZN(n7313)
         );
  XNOR2_X1 U9068 ( .A(n7450), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n7309) );
  INV_X1 U9069 ( .A(n7309), .ZN(n7311) );
  INV_X1 U9070 ( .A(n7308), .ZN(n7310) );
  OAI211_X1 U9071 ( .C1(n7311), .C2(n7310), .A(n10331), .B(n7449), .ZN(n7312)
         );
  OAI211_X1 U9072 ( .C1(n10327), .C2(n7453), .A(n7313), .B(n7312), .ZN(
        P2_U3257) );
  NAND2_X1 U9073 ( .A1(n7315), .A2(n7314), .ZN(n7316) );
  AOI21_X1 U9074 ( .B1(n7317), .B2(n7316), .A(n8773), .ZN(n7327) );
  INV_X1 U9075 ( .A(n9136), .ZN(n7321) );
  NAND2_X1 U9076 ( .A1(n8817), .A2(n9134), .ZN(n7320) );
  INV_X1 U9077 ( .A(n7318), .ZN(n7319) );
  OAI211_X1 U9078 ( .C1(n7321), .C2(n8819), .A(n7320), .B(n7319), .ZN(n7326)
         );
  NAND2_X1 U9079 ( .A1(n8791), .A2(n7322), .ZN(n7323) );
  OAI21_X1 U9080 ( .B1(n8804), .B2(n7324), .A(n7323), .ZN(n7325) );
  OR3_X1 U9081 ( .A1(n7327), .A2(n7326), .A3(n7325), .ZN(P1_U3229) );
  INV_X1 U9082 ( .A(n7155), .ZN(n7330) );
  NOR3_X1 U9083 ( .A1(n8224), .A2(n7328), .A3(n7364), .ZN(n7329) );
  AOI21_X1 U9084 ( .B1(n7330), .B2(n8235), .A(n7329), .ZN(n7341) );
  NAND2_X1 U9085 ( .A1(n8217), .A2(n8252), .ZN(n7335) );
  NAND2_X1 U9086 ( .A1(n8216), .A2(n8251), .ZN(n7334) );
  INV_X1 U9087 ( .A(n7365), .ZN(n7331) );
  NAND2_X1 U9088 ( .A1(n8229), .A2(n7331), .ZN(n7332) );
  NAND4_X1 U9089 ( .A1(n7335), .A2(n7334), .A3(n7333), .A4(n7332), .ZN(n7338)
         );
  NOR2_X1 U9090 ( .A1(n7336), .A2(n8211), .ZN(n7337) );
  AOI211_X1 U9091 ( .C1(n8003), .C2(n8230), .A(n7338), .B(n7337), .ZN(n7339)
         );
  OAI21_X1 U9092 ( .B1(n7341), .B2(n7340), .A(n7339), .ZN(P2_U3226) );
  INV_X1 U9093 ( .A(n7342), .ZN(n7343) );
  AOI21_X1 U9094 ( .B1(n8110), .B2(n7344), .A(n7343), .ZN(n7390) );
  XNOR2_X1 U9095 ( .A(n7345), .B(n8110), .ZN(n7349) );
  OAI22_X1 U9096 ( .A1(n7858), .A2(n8513), .B1(n7346), .B2(n8515), .ZN(n7348)
         );
  NOR2_X1 U9097 ( .A1(n7390), .A2(n7676), .ZN(n7347) );
  AOI211_X1 U9098 ( .C1(n7349), .C2(n10369), .A(n7348), .B(n7347), .ZN(n7389)
         );
  OR2_X1 U9099 ( .A1(n7389), .A2(n10389), .ZN(n7358) );
  OAI22_X1 U9100 ( .A1(n10376), .A2(n7350), .B1(n7857), .B2(n8468), .ZN(n7355)
         );
  INV_X1 U9101 ( .A(n7351), .ZN(n7353) );
  OAI211_X1 U9102 ( .C1(n7353), .C2(n4765), .A(n10360), .B(n7352), .ZN(n7388)
         );
  NOR2_X1 U9103 ( .A1(n8361), .A2(n7388), .ZN(n7354) );
  AOI211_X1 U9104 ( .C1(n10381), .C2(n7356), .A(n7355), .B(n7354), .ZN(n7357)
         );
  OAI211_X1 U9105 ( .C1(n7390), .C2(n10380), .A(n7358), .B(n7357), .ZN(
        P2_U3287) );
  XNOR2_X1 U9106 ( .A(n7360), .B(n7359), .ZN(n10467) );
  INV_X1 U9107 ( .A(n10467), .ZN(n7371) );
  NAND2_X1 U9108 ( .A1(n7361), .A2(n8001), .ZN(n7362) );
  XNOR2_X1 U9109 ( .A(n7362), .B(n8114), .ZN(n7363) );
  OAI222_X1 U9110 ( .A1(n8515), .A2(n7543), .B1(n8513), .B2(n7364), .C1(n7363), 
        .C2(n8510), .ZN(n10464) );
  OAI21_X1 U9111 ( .B1(n7380), .B2(n10461), .A(n7423), .ZN(n10463) );
  INV_X1 U9112 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7366) );
  OAI22_X1 U9113 ( .A1(n10376), .A2(n7366), .B1(n7365), .B2(n8468), .ZN(n7367)
         );
  AOI21_X1 U9114 ( .B1(n10381), .B2(n8003), .A(n7367), .ZN(n7368) );
  OAI21_X1 U9115 ( .B1(n10463), .B2(n7894), .A(n7368), .ZN(n7369) );
  AOI21_X1 U9116 ( .B1(n10464), .B2(n10376), .A(n7369), .ZN(n7370) );
  OAI21_X1 U9117 ( .B1(n8553), .B2(n7371), .A(n7370), .ZN(P2_U3284) );
  INV_X1 U9118 ( .A(n7372), .ZN(n7913) );
  OAI222_X1 U9119 ( .A1(n9562), .A2(n7373), .B1(n9560), .B2(n7913), .C1(n8938), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  XNOR2_X1 U9120 ( .A(n7374), .B(n8112), .ZN(n7447) );
  INV_X1 U9121 ( .A(n7375), .ZN(n7376) );
  OAI21_X1 U9122 ( .B1(n7376), .B2(n7984), .A(n8112), .ZN(n7377) );
  NAND2_X1 U9123 ( .A1(n7377), .A2(n7361), .ZN(n7378) );
  AOI222_X1 U9124 ( .A1(n10369), .A2(n7378), .B1(n4870), .B2(n8544), .C1(n8253), .C2(n8543), .ZN(n7442) );
  INV_X1 U9125 ( .A(n7379), .ZN(n7381) );
  AOI21_X1 U9126 ( .B1(n7382), .B2(n7381), .A(n7380), .ZN(n7445) );
  AOI22_X1 U9127 ( .A1(n7445), .A2(n10360), .B1(n8644), .B2(n7382), .ZN(n7383)
         );
  OAI211_X1 U9128 ( .C1(n10432), .C2(n7447), .A(n7442), .B(n7383), .ZN(n7385)
         );
  NAND2_X1 U9129 ( .A1(n7385), .A2(n10477), .ZN(n7384) );
  OAI21_X1 U9130 ( .B1(n10477), .B2(n7187), .A(n7384), .ZN(P2_U3531) );
  INV_X1 U9131 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7387) );
  NAND2_X1 U9132 ( .A1(n7385), .A2(n10469), .ZN(n7386) );
  OAI21_X1 U9133 ( .B1(n10469), .B2(n7387), .A(n7386), .ZN(P2_U3484) );
  OAI211_X1 U9134 ( .C1(n7390), .C2(n8633), .A(n7389), .B(n7388), .ZN(n7395)
         );
  OAI22_X1 U9135 ( .A1(n8628), .A2(n4765), .B1(n10477), .B2(n6986), .ZN(n7391)
         );
  AOI21_X1 U9136 ( .B1(n7395), .B2(n10477), .A(n7391), .ZN(n7392) );
  INV_X1 U9137 ( .A(n7392), .ZN(P2_U3529) );
  INV_X1 U9138 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7393) );
  OAI22_X1 U9139 ( .A1(n8678), .A2(n4765), .B1(n10469), .B2(n7393), .ZN(n7394)
         );
  AOI21_X1 U9140 ( .B1(n7395), .B2(n10469), .A(n7394), .ZN(n7396) );
  INV_X1 U9141 ( .A(n7396), .ZN(P2_U3478) );
  AOI21_X1 U9142 ( .B1(n5529), .B2(n7398), .A(n7397), .ZN(n10108) );
  MUX2_X1 U9143 ( .A(n7399), .B(P1_REG1_REG_13__SCAN_IN), .S(n7407), .Z(n10107) );
  NOR2_X1 U9144 ( .A1(n10108), .A2(n10107), .ZN(n10106) );
  AOI21_X1 U9145 ( .B1(n7399), .B2(n10104), .A(n10106), .ZN(n7402) );
  AOI22_X1 U9146 ( .A1(n7400), .A2(n5570), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n9179), .ZN(n7401) );
  NOR2_X1 U9147 ( .A1(n7402), .A2(n7401), .ZN(n9178) );
  AOI21_X1 U9148 ( .B1(n7402), .B2(n7401), .A(n9178), .ZN(n7415) );
  XNOR2_X1 U9149 ( .A(n7407), .B(n7403), .ZN(n10094) );
  INV_X1 U9150 ( .A(n7404), .ZN(n7405) );
  NAND2_X1 U9151 ( .A1(n7406), .A2(n7405), .ZN(n10095) );
  NAND2_X1 U9152 ( .A1(n7408), .A2(n7562), .ZN(n9167) );
  OAI21_X1 U9153 ( .B1(n7408), .B2(n7562), .A(n9167), .ZN(n7413) );
  NAND2_X1 U9154 ( .A1(n10079), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n7411) );
  NOR2_X1 U9155 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7409), .ZN(n7695) );
  INV_X1 U9156 ( .A(n7695), .ZN(n7410) );
  OAI211_X1 U9157 ( .C1(n10163), .C2(n9179), .A(n7411), .B(n7410), .ZN(n7412)
         );
  AOI21_X1 U9158 ( .B1(n7413), .B2(n10086), .A(n7412), .ZN(n7414) );
  OAI21_X1 U9159 ( .B1(n7415), .B2(n10169), .A(n7414), .ZN(P1_U3255) );
  NAND2_X1 U9160 ( .A1(n7416), .A2(n7419), .ZN(n7417) );
  NAND2_X1 U9161 ( .A1(n7418), .A2(n7417), .ZN(n7597) );
  OAI21_X1 U9162 ( .B1(n4506), .B2(n7419), .A(n7540), .ZN(n7421) );
  OAI22_X1 U9163 ( .A1(n8004), .A2(n8513), .B1(n7591), .B2(n8515), .ZN(n7420)
         );
  AOI21_X1 U9164 ( .B1(n7421), .B2(n10369), .A(n7420), .ZN(n7422) );
  OAI21_X1 U9165 ( .B1(n7597), .B2(n7676), .A(n7422), .ZN(n7598) );
  NAND2_X1 U9166 ( .A1(n7598), .A2(n10376), .ZN(n7430) );
  AOI211_X1 U9167 ( .C1(n7424), .C2(n7423), .A(n10462), .B(n4764), .ZN(n7599)
         );
  NOR2_X1 U9168 ( .A1(n7606), .A2(n8537), .ZN(n7428) );
  OAI22_X1 U9169 ( .A1(n10376), .A2(n7426), .B1(n7425), .B2(n8468), .ZN(n7427)
         );
  AOI211_X1 U9170 ( .C1(n7599), .C2(n10383), .A(n7428), .B(n7427), .ZN(n7429)
         );
  OAI211_X1 U9171 ( .C1(n7597), .C2(n10380), .A(n7430), .B(n7429), .ZN(
        P2_U3283) );
  NAND2_X1 U9172 ( .A1(n7435), .A2(n7431), .ZN(n7433) );
  NOR2_X1 U9173 ( .A1(n7432), .A2(P1_U3084), .ZN(n9117) );
  INV_X1 U9174 ( .A(n9117), .ZN(n9124) );
  OAI211_X1 U9175 ( .C1(n7434), .C2(n9553), .A(n7433), .B(n9124), .ZN(P1_U3330) );
  NAND2_X1 U9176 ( .A1(n7435), .A2(n7766), .ZN(n7436) );
  OAI211_X1 U9177 ( .C1(n7437), .C2(n8148), .A(n7436), .B(n8145), .ZN(P2_U3335) );
  INV_X1 U9178 ( .A(n7438), .ZN(n7439) );
  AOI22_X1 U9179 ( .A1(n10389), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7439), .B2(
        n10379), .ZN(n7440) );
  OAI21_X1 U9180 ( .B1(n7441), .B2(n8537), .A(n7440), .ZN(n7444) );
  NOR2_X1 U9181 ( .A1(n7442), .A2(n8548), .ZN(n7443) );
  AOI211_X1 U9182 ( .C1(n7445), .C2(n8551), .A(n7444), .B(n7443), .ZN(n7446)
         );
  OAI21_X1 U9183 ( .B1(n8553), .B2(n7447), .A(n7446), .ZN(P2_U3285) );
  NOR2_X1 U9184 ( .A1(n7575), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7448) );
  AOI21_X1 U9185 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n7575), .A(n7448), .ZN(
        n7452) );
  OAI21_X1 U9186 ( .B1(n7452), .B2(n7451), .A(n7574), .ZN(n7462) );
  NAND2_X1 U9187 ( .A1(n7453), .A2(n6111), .ZN(n7454) );
  AOI22_X1 U9188 ( .A1(n7575), .A2(n7601), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7571), .ZN(n7456) );
  NOR2_X1 U9189 ( .A1(n7457), .A2(n7456), .ZN(n7570) );
  AOI21_X1 U9190 ( .B1(n7457), .B2(n7456), .A(n7570), .ZN(n7460) );
  NAND2_X1 U9191 ( .A1(n9994), .A2(n7575), .ZN(n7459) );
  AOI22_X1 U9192 ( .A1(n10333), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3152), .ZN(n7458) );
  OAI211_X1 U9193 ( .C1(n7460), .C2(n10328), .A(n7459), .B(n7458), .ZN(n7461)
         );
  AOI21_X1 U9194 ( .B1(n10331), .B2(n7462), .A(n7461), .ZN(n7463) );
  INV_X1 U9195 ( .A(n7463), .ZN(P2_U3258) );
  AOI21_X1 U9196 ( .B1(n7465), .B2(n7464), .A(n8773), .ZN(n7467) );
  NAND2_X1 U9197 ( .A1(n7467), .A2(n7466), .ZN(n7475) );
  INV_X1 U9198 ( .A(n9134), .ZN(n7470) );
  NAND2_X1 U9199 ( .A1(n8817), .A2(n9133), .ZN(n7469) );
  OAI211_X1 U9200 ( .C1(n7470), .C2(n8819), .A(n7469), .B(n7468), .ZN(n7473)
         );
  NOR2_X1 U9201 ( .A1(n8804), .A2(n7471), .ZN(n7472) );
  NOR2_X1 U9202 ( .A1(n7473), .A2(n7472), .ZN(n7474) );
  OAI211_X1 U9203 ( .C1(n7558), .C2(n8824), .A(n7475), .B(n7474), .ZN(P1_U3234) );
  NOR3_X1 U9204 ( .A1(n7476), .A2(n7543), .A3(n8224), .ZN(n7477) );
  AOI21_X1 U9205 ( .B1(n7478), .B2(n8235), .A(n7477), .ZN(n7490) );
  XNOR2_X1 U9206 ( .A(n8643), .B(n7720), .ZN(n7507) );
  NOR2_X1 U9207 ( .A1(n7591), .A2(n8186), .ZN(n7505) );
  XNOR2_X1 U9208 ( .A(n7507), .B(n7505), .ZN(n7489) );
  NAND2_X1 U9209 ( .A1(n8217), .A2(n8251), .ZN(n7482) );
  NAND2_X1 U9210 ( .A1(n8216), .A2(n8249), .ZN(n7481) );
  NAND2_X1 U9211 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7579) );
  INV_X1 U9212 ( .A(n7479), .ZN(n7536) );
  NAND2_X1 U9213 ( .A1(n8229), .A2(n7536), .ZN(n7480) );
  NAND4_X1 U9214 ( .A1(n7482), .A2(n7481), .A3(n7579), .A4(n7480), .ZN(n7487)
         );
  AND2_X1 U9215 ( .A1(n7489), .A2(n7483), .ZN(n7484) );
  NOR2_X1 U9216 ( .A1(n7509), .A2(n8211), .ZN(n7486) );
  AOI211_X1 U9217 ( .C1(n8643), .C2(n8230), .A(n7487), .B(n7486), .ZN(n7488)
         );
  OAI21_X1 U9218 ( .B1(n7490), .B2(n7489), .A(n7488), .ZN(P2_U3217) );
  AOI21_X1 U9219 ( .B1(n8817), .B2(n10014), .A(n7491), .ZN(n7494) );
  INV_X1 U9220 ( .A(n9135), .ZN(n7492) );
  OR2_X1 U9221 ( .A1(n8819), .A2(n7492), .ZN(n7493) );
  OAI211_X1 U9222 ( .C1(n8804), .C2(n7495), .A(n7494), .B(n7493), .ZN(n7502)
         );
  NAND2_X1 U9223 ( .A1(n7497), .A2(n7496), .ZN(n7498) );
  XNOR2_X1 U9224 ( .A(n7499), .B(n7498), .ZN(n7500) );
  NOR2_X1 U9225 ( .A1(n7500), .A2(n8773), .ZN(n7501) );
  AOI211_X1 U9226 ( .C1(n8791), .C2(n7503), .A(n7502), .B(n7501), .ZN(n7504)
         );
  INV_X1 U9227 ( .A(n7504), .ZN(P1_U3215) );
  INV_X1 U9228 ( .A(n7505), .ZN(n7506) );
  NAND2_X1 U9229 ( .A1(n7507), .A2(n7506), .ZN(n7508) );
  XNOR2_X1 U9230 ( .A(n7683), .B(n7853), .ZN(n7622) );
  AND2_X1 U9231 ( .A1(n8248), .A2(n7926), .ZN(n7511) );
  NOR2_X1 U9232 ( .A1(n7672), .A2(n8186), .ZN(n7510) );
  XNOR2_X1 U9233 ( .A(n8638), .B(n7853), .ZN(n7587) );
  AOI22_X1 U9234 ( .A1(n7622), .A2(n7511), .B1(n7510), .B2(n7587), .ZN(n7515)
         );
  INV_X1 U9235 ( .A(n7587), .ZN(n7618) );
  INV_X1 U9236 ( .A(n7510), .ZN(n7619) );
  INV_X1 U9237 ( .A(n7511), .ZN(n7621) );
  AOI21_X1 U9238 ( .B1(n7618), .B2(n7619), .A(n7621), .ZN(n7513) );
  NAND2_X1 U9239 ( .A1(n7619), .A2(n7621), .ZN(n7512) );
  OAI22_X1 U9240 ( .A1(n7622), .A2(n7513), .B1(n7587), .B2(n7512), .ZN(n7514)
         );
  NAND2_X1 U9241 ( .A1(n8542), .A2(n7926), .ZN(n7516) );
  NOR2_X1 U9242 ( .A1(n7823), .A2(n7516), .ZN(n7659) );
  AOI21_X1 U9243 ( .B1(n7823), .B2(n7516), .A(n7659), .ZN(n7517) );
  OAI211_X1 U9244 ( .C1(n7518), .C2(n7517), .A(n7822), .B(n8235), .ZN(n7522)
         );
  OAI22_X1 U9245 ( .A1(n8206), .A2(n7738), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9949), .ZN(n7520) );
  OAI22_X1 U9246 ( .A1(n8514), .A2(n7827), .B1(n7859), .B2(n7729), .ZN(n7519)
         );
  AOI211_X1 U9247 ( .C1(n7737), .C2(n8230), .A(n7520), .B(n7519), .ZN(n7521)
         );
  NAND2_X1 U9248 ( .A1(n7522), .A2(n7521), .ZN(P2_U3230) );
  XNOR2_X1 U9249 ( .A(n7523), .B(n8017), .ZN(n7524) );
  AOI222_X1 U9250 ( .A1(n10369), .A2(n7524), .B1(n8250), .B2(n8543), .C1(n8248), .C2(n8544), .ZN(n8641) );
  OAI21_X1 U9251 ( .B1(n7526), .B2(n8017), .A(n7525), .ZN(n8637) );
  NAND2_X1 U9252 ( .A1(n8637), .A2(n10352), .ZN(n7531) );
  AOI21_X1 U9253 ( .B1(n8638), .B2(n7533), .A(n7679), .ZN(n8639) );
  INV_X1 U9254 ( .A(n8638), .ZN(n7596) );
  NOR2_X1 U9255 ( .A1(n7596), .A2(n8537), .ZN(n7529) );
  OAI22_X1 U9256 ( .A1(n10376), .A2(n7527), .B1(n7590), .B2(n8468), .ZN(n7528)
         );
  AOI211_X1 U9257 ( .C1(n8639), .C2(n8551), .A(n7529), .B(n7528), .ZN(n7530)
         );
  OAI211_X1 U9258 ( .C1(n8641), .C2(n10389), .A(n7531), .B(n7530), .ZN(
        P2_U3281) );
  XNOR2_X1 U9259 ( .A(n7532), .B(n8014), .ZN(n8648) );
  INV_X1 U9260 ( .A(n7533), .ZN(n7534) );
  AOI21_X1 U9261 ( .B1(n8643), .B2(n7535), .A(n7534), .ZN(n8645) );
  AOI22_X1 U9262 ( .A1(n10389), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7536), .B2(
        n10379), .ZN(n7537) );
  OAI21_X1 U9263 ( .B1(n4763), .B2(n8537), .A(n7537), .ZN(n7547) );
  INV_X1 U9264 ( .A(n7538), .ZN(n7542) );
  AOI21_X1 U9265 ( .B1(n7540), .B2(n7539), .A(n4812), .ZN(n7541) );
  NOR3_X1 U9266 ( .A1(n7542), .A2(n7541), .A3(n8510), .ZN(n7545) );
  OAI22_X1 U9267 ( .A1(n7672), .A2(n8515), .B1(n7543), .B2(n8513), .ZN(n7544)
         );
  NOR2_X1 U9268 ( .A1(n7545), .A2(n7544), .ZN(n8647) );
  NOR2_X1 U9269 ( .A1(n8647), .A2(n8548), .ZN(n7546) );
  AOI211_X1 U9270 ( .C1(n8645), .C2(n8551), .A(n7547), .B(n7546), .ZN(n7548)
         );
  OAI21_X1 U9271 ( .B1(n8553), .B2(n8648), .A(n7548), .ZN(P2_U3282) );
  INV_X1 U9272 ( .A(n7549), .ZN(n7552) );
  OAI222_X1 U9273 ( .A1(P2_U3152), .A2(n7551), .B1(n8686), .B2(n7552), .C1(
        n7550), .C2(n8148), .ZN(P2_U3334) );
  OAI222_X1 U9274 ( .A1(P1_U3084), .A2(n7553), .B1(n9560), .B2(n7552), .C1(
        n9928), .C2(n9562), .ZN(P1_U3329) );
  XNOR2_X1 U9275 ( .A(n8897), .B(n8976), .ZN(n8853) );
  NAND2_X1 U9276 ( .A1(n9523), .A2(n7639), .ZN(n8960) );
  NOR2_X1 U9277 ( .A1(n9523), .A2(n7639), .ZN(n8890) );
  NAND2_X1 U9278 ( .A1(n10011), .A2(n8962), .ZN(n7556) );
  NAND2_X1 U9279 ( .A1(n10020), .A2(n7555), .ZN(n8961) );
  NAND2_X1 U9280 ( .A1(n7556), .A2(n8961), .ZN(n7613) );
  INV_X1 U9281 ( .A(n10013), .ZN(n7693) );
  OR2_X1 U9282 ( .A1(n9516), .A2(n7693), .ZN(n8894) );
  NAND2_X1 U9283 ( .A1(n9516), .A2(n7693), .ZN(n8965) );
  NAND2_X1 U9284 ( .A1(n7613), .A2(n8850), .ZN(n7612) );
  XOR2_X1 U9285 ( .A(n8853), .B(n7706), .Z(n7557) );
  AOI222_X1 U9286 ( .A1(n9424), .A2(n7557), .B1(n9131), .B2(n10223), .C1(
        n10013), .C2(n10226), .ZN(n10028) );
  NAND2_X1 U9287 ( .A1(n7558), .A2(n7639), .ZN(n7560) );
  NOR2_X1 U9288 ( .A1(n9516), .A2(n10013), .ZN(n7561) );
  INV_X1 U9289 ( .A(n9516), .ZN(n7611) );
  XOR2_X1 U9290 ( .A(n8853), .B(n7701), .Z(n10031) );
  NAND2_X1 U9291 ( .A1(n10031), .A2(n7790), .ZN(n7569) );
  OAI22_X1 U9292 ( .A1(n9403), .A2(n7562), .B1(n7697), .B2(n10237), .ZN(n7567)
         );
  INV_X1 U9293 ( .A(n7753), .ZN(n7564) );
  OAI211_X1 U9294 ( .C1(n10029), .C2(n7608), .A(n7564), .B(n10198), .ZN(n10027) );
  NOR2_X1 U9295 ( .A1(n10027), .A2(n7565), .ZN(n7566) );
  AOI211_X1 U9296 ( .C1(n10187), .C2(n8897), .A(n7567), .B(n7566), .ZN(n7568)
         );
  OAI211_X1 U9297 ( .C1(n10215), .C2(n10028), .A(n7569), .B(n7568), .ZN(
        P1_U3277) );
  AOI21_X1 U9298 ( .B1(n7571), .B2(n7601), .A(n7570), .ZN(n7573) );
  AOI22_X1 U9299 ( .A1(n8278), .A2(n8281), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n8282), .ZN(n7572) );
  NOR2_X1 U9300 ( .A1(n7573), .A2(n7572), .ZN(n8280) );
  AOI21_X1 U9301 ( .B1(n7573), .B2(n7572), .A(n8280), .ZN(n7585) );
  AOI22_X1 U9302 ( .A1(n8278), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n6136), .B2(
        n8282), .ZN(n7577) );
  NAND2_X1 U9303 ( .A1(n7577), .A2(n7576), .ZN(n8277) );
  OAI21_X1 U9304 ( .B1(n7577), .B2(n7576), .A(n8277), .ZN(n7578) );
  NAND2_X1 U9305 ( .A1(n7578), .A2(n10331), .ZN(n7584) );
  INV_X1 U9306 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7580) );
  OAI21_X1 U9307 ( .B1(n7581), .B2(n7580), .A(n7579), .ZN(n7582) );
  AOI21_X1 U9308 ( .B1(n9994), .B2(n8278), .A(n7582), .ZN(n7583) );
  OAI211_X1 U9309 ( .C1(n7585), .C2(n10328), .A(n7584), .B(n7583), .ZN(
        P2_U3259) );
  INV_X1 U9310 ( .A(n8224), .ZN(n8175) );
  NAND2_X1 U9311 ( .A1(n8175), .A2(n8249), .ZN(n7589) );
  NAND2_X1 U9312 ( .A1(n8235), .A2(n7619), .ZN(n7588) );
  XNOR2_X1 U9313 ( .A(n7586), .B(n7587), .ZN(n7620) );
  MUX2_X1 U9314 ( .A(n7589), .B(n7588), .S(n7620), .Z(n7595) );
  NOR2_X1 U9315 ( .A1(n8206), .A2(n7590), .ZN(n7593) );
  OAI22_X1 U9316 ( .A1(n7729), .A2(n7827), .B1(n7859), .B2(n7591), .ZN(n7592)
         );
  AOI211_X1 U9317 ( .C1(P2_REG3_REG_15__SCAN_IN), .C2(P2_U3152), .A(n7593), 
        .B(n7592), .ZN(n7594) );
  OAI211_X1 U9318 ( .C1(n7596), .C2(n8220), .A(n7595), .B(n7594), .ZN(P2_U3243) );
  INV_X1 U9319 ( .A(n7597), .ZN(n7600) );
  AOI211_X1 U9320 ( .C1(n7600), .C2(n10453), .A(n7599), .B(n7598), .ZN(n7603)
         );
  MUX2_X1 U9321 ( .A(n7601), .B(n7603), .S(n10477), .Z(n7602) );
  OAI21_X1 U9322 ( .B1(n7606), .B2(n8628), .A(n7602), .ZN(P2_U3533) );
  INV_X1 U9323 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7604) );
  MUX2_X1 U9324 ( .A(n7604), .B(n7603), .S(n10469), .Z(n7605) );
  OAI21_X1 U9325 ( .B1(n7606), .B2(n8678), .A(n7605), .ZN(P2_U3490) );
  XNOR2_X1 U9326 ( .A(n7607), .B(n8850), .ZN(n9521) );
  AOI21_X1 U9327 ( .B1(n9516), .B2(n10021), .A(n7608), .ZN(n9517) );
  INV_X1 U9328 ( .A(n7650), .ZN(n7609) );
  AOI22_X1 U9329 ( .A1(n10215), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7609), .B2(
        n10203), .ZN(n7610) );
  OAI21_X1 U9330 ( .B1(n10239), .B2(n7611), .A(n7610), .ZN(n7616) );
  OAI21_X1 U9331 ( .B1(n8850), .B2(n7613), .A(n7612), .ZN(n7614) );
  AOI222_X1 U9332 ( .A1(n9424), .A2(n7614), .B1(n9132), .B2(n10223), .C1(n9133), .C2(n10226), .ZN(n9519) );
  NOR2_X1 U9333 ( .A1(n9519), .A2(n10215), .ZN(n7615) );
  AOI211_X1 U9334 ( .C1(n9517), .C2(n10221), .A(n7616), .B(n7615), .ZN(n7617)
         );
  OAI21_X1 U9335 ( .B1(n9428), .B2(n9521), .A(n7617), .ZN(P1_U3278) );
  AOI22_X1 U9336 ( .A1(n7620), .A2(n7619), .B1(n7618), .B2(n7586), .ZN(n7624)
         );
  XNOR2_X1 U9337 ( .A(n7622), .B(n7621), .ZN(n7623) );
  XNOR2_X1 U9338 ( .A(n7624), .B(n7623), .ZN(n7628) );
  AOI22_X1 U9339 ( .A1(n8217), .A2(n8249), .B1(n8216), .B2(n8542), .ZN(n7625)
         );
  NAND2_X1 U9340 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8303) );
  OAI211_X1 U9341 ( .C1(n7677), .C2(n8206), .A(n7625), .B(n8303), .ZN(n7626)
         );
  AOI21_X1 U9342 ( .B1(n7683), .B2(n8230), .A(n7626), .ZN(n7627) );
  OAI21_X1 U9343 ( .B1(n7628), .B2(n8211), .A(n7627), .ZN(P2_U3228) );
  INV_X1 U9344 ( .A(n7629), .ZN(n7633) );
  OAI222_X1 U9345 ( .A1(n8148), .A2(n7631), .B1(n8686), .B2(n7633), .C1(
        P2_U3152), .C2(n7630), .ZN(P2_U3333) );
  OAI222_X1 U9346 ( .A1(n9562), .A2(n9859), .B1(n9560), .B2(n7633), .C1(
        P1_U3084), .C2(n7632), .ZN(P1_U3328) );
  INV_X1 U9347 ( .A(n10020), .ZN(n10033) );
  OAI21_X1 U9348 ( .B1(n7636), .B2(n7635), .A(n7634), .ZN(n7637) );
  NAND2_X1 U9349 ( .A1(n7637), .A2(n8812), .ZN(n7643) );
  OAI21_X1 U9350 ( .B1(n8819), .B2(n7639), .A(n7638), .ZN(n7641) );
  NOR2_X1 U9351 ( .A1(n8804), .A2(n10018), .ZN(n7640) );
  AOI211_X1 U9352 ( .C1(n8817), .C2(n10013), .A(n7641), .B(n7640), .ZN(n7642)
         );
  OAI211_X1 U9353 ( .C1(n10033), .C2(n8824), .A(n7643), .B(n7642), .ZN(
        P1_U3222) );
  XNOR2_X1 U9354 ( .A(n7645), .B(n7644), .ZN(n7646) );
  XNOR2_X1 U9355 ( .A(n7647), .B(n7646), .ZN(n7653) );
  AND2_X1 U9356 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10101) );
  AOI21_X1 U9357 ( .B1(n8808), .B2(n9133), .A(n10101), .ZN(n7649) );
  NAND2_X1 U9358 ( .A1(n8817), .A2(n9132), .ZN(n7648) );
  OAI211_X1 U9359 ( .C1(n8804), .C2(n7650), .A(n7649), .B(n7648), .ZN(n7651)
         );
  AOI21_X1 U9360 ( .B1(n8791), .B2(n9516), .A(n7651), .ZN(n7652) );
  OAI21_X1 U9361 ( .B1(n7653), .B2(n8773), .A(n7652), .ZN(P1_U3232) );
  XNOR2_X1 U9362 ( .A(n8521), .B(n7720), .ZN(n7654) );
  NAND2_X1 U9363 ( .A1(n8545), .A2(n7926), .ZN(n7656) );
  INV_X1 U9364 ( .A(n7654), .ZN(n7658) );
  NOR2_X1 U9365 ( .A1(n8224), .A2(n8498), .ZN(n7655) );
  AOI22_X1 U9366 ( .A1(n7717), .A2(n8235), .B1(n7658), .B2(n7655), .ZN(n7663)
         );
  INV_X1 U9367 ( .A(n7656), .ZN(n7657) );
  NAND2_X1 U9368 ( .A1(n7658), .A2(n7657), .ZN(n7718) );
  NAND3_X1 U9369 ( .A1(n4605), .A2(n8235), .A3(n7718), .ZN(n7662) );
  XNOR2_X1 U9370 ( .A(n8618), .B(n7853), .ZN(n7661) );
  NOR2_X1 U9371 ( .A1(n8514), .A2(n8186), .ZN(n7660) );
  XNOR2_X1 U9372 ( .A(n7661), .B(n7660), .ZN(n7821) );
  MUX2_X1 U9373 ( .A(n7663), .B(n7662), .S(n7719), .Z(n7667) );
  NOR2_X1 U9374 ( .A1(n8206), .A2(n8523), .ZN(n7665) );
  OAI22_X1 U9375 ( .A1(n8514), .A2(n7859), .B1(n7827), .B2(n8516), .ZN(n7664)
         );
  AOI211_X1 U9376 ( .C1(P2_REG3_REG_19__SCAN_IN), .C2(P2_U3152), .A(n7665), 
        .B(n7664), .ZN(n7666) );
  OAI211_X1 U9377 ( .C1(n8673), .C2(n8220), .A(n7667), .B(n7666), .ZN(P2_U3221) );
  AND2_X1 U9378 ( .A1(n7668), .A2(n8118), .ZN(n7670) );
  OR2_X1 U9379 ( .A1(n7670), .A2(n7669), .ZN(n8634) );
  XNOR2_X1 U9380 ( .A(n7671), .B(n8022), .ZN(n7674) );
  OAI22_X1 U9381 ( .A1(n7828), .A2(n8515), .B1(n7672), .B2(n8513), .ZN(n7673)
         );
  AOI21_X1 U9382 ( .B1(n7674), .B2(n10369), .A(n7673), .ZN(n7675) );
  OAI21_X1 U9383 ( .B1(n8634), .B2(n7676), .A(n7675), .ZN(n8636) );
  NAND2_X1 U9384 ( .A1(n8636), .A2(n10376), .ZN(n7685) );
  OAI22_X1 U9385 ( .A1(n10376), .A2(n7678), .B1(n7677), .B2(n8468), .ZN(n7682)
         );
  NOR2_X1 U9386 ( .A1(n7679), .A2(n8629), .ZN(n7680) );
  OR2_X1 U9387 ( .A1(n7735), .A2(n7680), .ZN(n8630) );
  NOR2_X1 U9388 ( .A1(n8630), .A2(n7894), .ZN(n7681) );
  AOI211_X1 U9389 ( .C1(n10381), .C2(n7683), .A(n7682), .B(n7681), .ZN(n7684)
         );
  OAI211_X1 U9390 ( .C1(n8634), .C2(n10380), .A(n7685), .B(n7684), .ZN(
        P2_U3280) );
  INV_X1 U9391 ( .A(n7686), .ZN(n7763) );
  OAI222_X1 U9392 ( .A1(P2_U3152), .A2(n7688), .B1(n8686), .B2(n7763), .C1(
        n7687), .C2(n8148), .ZN(P2_U3332) );
  XNOR2_X1 U9393 ( .A(n7690), .B(n7689), .ZN(n7691) );
  XNOR2_X1 U9394 ( .A(n7692), .B(n7691), .ZN(n7700) );
  NOR2_X1 U9395 ( .A1(n8819), .A2(n7693), .ZN(n7694) );
  AOI211_X1 U9396 ( .C1(n8817), .C2(n9131), .A(n7695), .B(n7694), .ZN(n7696)
         );
  OAI21_X1 U9397 ( .B1(n8804), .B2(n7697), .A(n7696), .ZN(n7698) );
  AOI21_X1 U9398 ( .B1(n8791), .B2(n8897), .A(n7698), .ZN(n7699) );
  OAI21_X1 U9399 ( .B1(n7700), .B2(n8773), .A(n7699), .ZN(P1_U3213) );
  AOI21_X1 U9400 ( .B1(n9132), .B2(n8897), .A(n7701), .ZN(n7703) );
  NAND2_X1 U9401 ( .A1(n7745), .A2(n7704), .ZN(n7705) );
  INV_X1 U9402 ( .A(n9131), .ZN(n7815) );
  NAND2_X1 U9403 ( .A1(n9507), .A2(n7747), .ZN(n8993) );
  NAND2_X1 U9404 ( .A1(n8992), .A2(n8993), .ZN(n8988) );
  XNOR2_X1 U9405 ( .A(n7787), .B(n8988), .ZN(n9509) );
  INV_X1 U9406 ( .A(n9130), .ZN(n7788) );
  INV_X1 U9407 ( .A(n10226), .ZN(n10209) );
  OR2_X1 U9408 ( .A1(n8897), .A2(n8976), .ZN(n8969) );
  AND2_X1 U9409 ( .A1(n9510), .A2(n9131), .ZN(n8986) );
  NAND2_X1 U9410 ( .A1(n7804), .A2(n7815), .ZN(n8898) );
  INV_X1 U9411 ( .A(n8988), .ZN(n8855) );
  XNOR2_X1 U9412 ( .A(n7780), .B(n8855), .ZN(n7710) );
  OAI222_X1 U9413 ( .A1(n10183), .A2(n7788), .B1(n10209), .B2(n7815), .C1(
        n7710), .C2(n10228), .ZN(n9505) );
  INV_X1 U9414 ( .A(n9507), .ZN(n7820) );
  INV_X1 U9415 ( .A(n9414), .ZN(n7711) );
  AOI211_X1 U9416 ( .C1(n9507), .C2(n7752), .A(n10306), .B(n7711), .ZN(n9506)
         );
  NAND2_X1 U9417 ( .A1(n9506), .A2(n10024), .ZN(n7714) );
  INV_X1 U9418 ( .A(n7712), .ZN(n7817) );
  AOI22_X1 U9419 ( .A1(n10215), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n7817), .B2(
        n10203), .ZN(n7713) );
  OAI211_X1 U9420 ( .C1(n7820), .C2(n10239), .A(n7714), .B(n7713), .ZN(n7715)
         );
  AOI21_X1 U9421 ( .B1(n9505), .B2(n9403), .A(n7715), .ZN(n7716) );
  OAI21_X1 U9422 ( .B1(n9509), .B2(n9428), .A(n7716), .ZN(P1_U3275) );
  XNOR2_X1 U9423 ( .A(n8608), .B(n7720), .ZN(n7770) );
  NOR2_X1 U9424 ( .A1(n8516), .A2(n8186), .ZN(n7772) );
  XNOR2_X1 U9425 ( .A(n7770), .B(n7772), .ZN(n7773) );
  XNOR2_X1 U9426 ( .A(n7774), .B(n7773), .ZN(n7725) );
  INV_X1 U9427 ( .A(n8493), .ZN(n7721) );
  OAI22_X1 U9428 ( .A1(n8206), .A2(n7721), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9900), .ZN(n7723) );
  OAI22_X1 U9429 ( .A1(n8498), .A2(n7859), .B1(n7827), .B2(n8499), .ZN(n7722)
         );
  AOI211_X1 U9430 ( .C1(n8608), .C2(n8230), .A(n7723), .B(n7722), .ZN(n7724)
         );
  OAI21_X1 U9431 ( .B1(n7725), .B2(n8211), .A(n7724), .ZN(P2_U3235) );
  OAI211_X1 U9432 ( .C1(n7728), .C2(n7727), .A(n7726), .B(n10369), .ZN(n7732)
         );
  OAI22_X1 U9433 ( .A1(n8514), .A2(n8515), .B1(n7729), .B2(n8513), .ZN(n7730)
         );
  INV_X1 U9434 ( .A(n7730), .ZN(n7731) );
  NAND2_X1 U9435 ( .A1(n7732), .A2(n7731), .ZN(n8623) );
  INV_X1 U9436 ( .A(n8623), .ZN(n7744) );
  OAI21_X1 U9437 ( .B1(n7734), .B2(n8120), .A(n7733), .ZN(n8625) );
  NAND2_X1 U9438 ( .A1(n8625), .A2(n10352), .ZN(n7743) );
  INV_X1 U9439 ( .A(n7735), .ZN(n7736) );
  AOI211_X1 U9440 ( .C1(n7737), .C2(n7736), .A(n10462), .B(n8531), .ZN(n8624)
         );
  NOR2_X1 U9441 ( .A1(n10389), .A2(n10367), .ZN(n8522) );
  NOR2_X1 U9442 ( .A1(n6180), .A2(n8537), .ZN(n7741) );
  INV_X1 U9443 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n7739) );
  OAI22_X1 U9444 ( .A1(n10376), .A2(n7739), .B1(n7738), .B2(n8468), .ZN(n7740)
         );
  AOI211_X1 U9445 ( .C1(n8624), .C2(n8522), .A(n7741), .B(n7740), .ZN(n7742)
         );
  OAI211_X1 U9446 ( .C1(n10389), .C2(n7744), .A(n7743), .B(n7742), .ZN(
        P2_U3279) );
  XOR2_X1 U9447 ( .A(n7745), .B(n8985), .Z(n9514) );
  INV_X1 U9448 ( .A(n9514), .ZN(n7760) );
  XOR2_X1 U9449 ( .A(n7746), .B(n8985), .Z(n7750) );
  NAND2_X1 U9450 ( .A1(n9514), .A2(n10184), .ZN(n7749) );
  INV_X1 U9451 ( .A(n7747), .ZN(n9421) );
  AOI22_X1 U9452 ( .A1(n9421), .A2(n10223), .B1(n10226), .B2(n9132), .ZN(n7748) );
  OAI211_X1 U9453 ( .C1(n10228), .C2(n7750), .A(n7749), .B(n7748), .ZN(n9512)
         );
  NAND2_X1 U9454 ( .A1(n9512), .A2(n9403), .ZN(n7758) );
  OAI22_X1 U9455 ( .A1(n9403), .A2(n7751), .B1(n7802), .B2(n10237), .ZN(n7756)
         );
  OAI21_X1 U9456 ( .B1(n9510), .B2(n7753), .A(n7752), .ZN(n9511) );
  NOR2_X1 U9457 ( .A1(n9511), .A2(n7754), .ZN(n7755) );
  AOI211_X1 U9458 ( .C1(n10187), .C2(n7804), .A(n7756), .B(n7755), .ZN(n7757)
         );
  OAI211_X1 U9459 ( .C1(n7760), .C2(n7759), .A(n7758), .B(n7757), .ZN(P1_U3276) );
  INV_X1 U9460 ( .A(n7761), .ZN(n7765) );
  OAI222_X1 U9461 ( .A1(n8148), .A2(n7762), .B1(n8686), .B2(n7765), .C1(n6351), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  OAI222_X1 U9462 ( .A1(P1_U3084), .A2(n7764), .B1(n9560), .B2(n7763), .C1(
        n9940), .C2(n9562), .ZN(P1_U3327) );
  OAI222_X1 U9463 ( .A1(n9562), .A2(n9946), .B1(P1_U3084), .B2(n6468), .C1(
        n9560), .C2(n7765), .ZN(P1_U3326) );
  NAND2_X1 U9464 ( .A1(n8149), .A2(n7766), .ZN(n7768) );
  OAI211_X1 U9465 ( .C1(n8148), .C2(n7769), .A(n7768), .B(n7767), .ZN(P2_U3330) );
  INV_X1 U9466 ( .A(n7770), .ZN(n7771) );
  XNOR2_X1 U9467 ( .A(n8482), .B(n7853), .ZN(n7840) );
  NAND2_X1 U9468 ( .A1(n8246), .A2(n7926), .ZN(n7839) );
  XNOR2_X1 U9469 ( .A(n7840), .B(n7839), .ZN(n7841) );
  XNOR2_X1 U9470 ( .A(n7842), .B(n7841), .ZN(n7778) );
  OAI22_X1 U9471 ( .A1(n8179), .A2(n8515), .B1(n8516), .B2(n8513), .ZN(n8485)
         );
  AOI22_X1 U9472 ( .A1(n8227), .A2(n8485), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n7775) );
  OAI21_X1 U9473 ( .B1(n8479), .B2(n8206), .A(n7775), .ZN(n7776) );
  AOI21_X1 U9474 ( .B1(n8603), .B2(n8230), .A(n7776), .ZN(n7777) );
  OAI21_X1 U9475 ( .B1(n7778), .B2(n8211), .A(n7777), .ZN(P2_U3225) );
  INV_X1 U9476 ( .A(n8992), .ZN(n7779) );
  NAND2_X1 U9477 ( .A1(n9500), .A2(n7788), .ZN(n8883) );
  INV_X1 U9478 ( .A(n8883), .ZN(n7781) );
  OR2_X1 U9479 ( .A1(n9500), .A2(n7788), .ZN(n8874) );
  OAI21_X1 U9480 ( .B1(n9420), .B2(n7781), .A(n8874), .ZN(n7782) );
  OR2_X1 U9481 ( .A1(n8796), .A2(n9411), .ZN(n9009) );
  NAND2_X1 U9482 ( .A1(n8796), .A2(n9411), .ZN(n9226) );
  NAND2_X1 U9483 ( .A1(n9009), .A2(n9226), .ZN(n8856) );
  XNOR2_X1 U9484 ( .A(n7782), .B(n8856), .ZN(n7783) );
  NAND2_X1 U9485 ( .A1(n7783), .A2(n9424), .ZN(n7785) );
  AOI22_X1 U9486 ( .A1(n10223), .A2(n9203), .B1(n9130), .B2(n10226), .ZN(n7784) );
  INV_X1 U9487 ( .A(n9500), .ZN(n9418) );
  OR2_X1 U9488 ( .A1(n7789), .A2(n8856), .ZN(n9495) );
  NAND3_X1 U9489 ( .A1(n9495), .A2(n9494), .A3(n7790), .ZN(n7796) );
  OAI22_X1 U9490 ( .A1(n9403), .A2(n9174), .B1(n8803), .B2(n10237), .ZN(n7794)
         );
  INV_X1 U9491 ( .A(n8796), .ZN(n9201) );
  OAI21_X1 U9492 ( .B1(n4559), .B2(n9201), .A(n10198), .ZN(n7791) );
  OR2_X1 U9493 ( .A1(n7791), .A2(n9396), .ZN(n9496) );
  INV_X1 U9494 ( .A(n9406), .ZN(n7792) );
  NOR2_X1 U9495 ( .A1(n9496), .A2(n7792), .ZN(n7793) );
  AOI211_X1 U9496 ( .C1(n10187), .C2(n8796), .A(n7794), .B(n7793), .ZN(n7795)
         );
  OAI211_X1 U9497 ( .C1(n10215), .C2(n9498), .A(n7796), .B(n7795), .ZN(
        P1_U3273) );
  NAND2_X1 U9498 ( .A1(n7809), .A2(n7797), .ZN(n7798) );
  XOR2_X1 U9499 ( .A(n7799), .B(n7798), .Z(n7806) );
  AND2_X1 U9500 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10116) );
  NOR2_X1 U9501 ( .A1(n8819), .A2(n8976), .ZN(n7800) );
  AOI211_X1 U9502 ( .C1(n8817), .C2(n9421), .A(n10116), .B(n7800), .ZN(n7801)
         );
  OAI21_X1 U9503 ( .B1(n7802), .B2(n8804), .A(n7801), .ZN(n7803) );
  AOI21_X1 U9504 ( .B1(n8791), .B2(n7804), .A(n7803), .ZN(n7805) );
  OAI21_X1 U9505 ( .B1(n7806), .B2(n8773), .A(n7805), .ZN(P1_U3239) );
  INV_X1 U9506 ( .A(n7807), .ZN(n7812) );
  AOI21_X1 U9507 ( .B1(n7810), .B2(n7809), .A(n7808), .ZN(n7811) );
  OAI21_X1 U9508 ( .B1(n7812), .B2(n7811), .A(n8812), .ZN(n7819) );
  NOR2_X1 U9509 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7813), .ZN(n10127) );
  AOI21_X1 U9510 ( .B1(n8817), .B2(n9130), .A(n10127), .ZN(n7814) );
  OAI21_X1 U9511 ( .B1(n7815), .B2(n8819), .A(n7814), .ZN(n7816) );
  AOI21_X1 U9512 ( .B1(n7817), .B2(n8821), .A(n7816), .ZN(n7818) );
  OAI211_X1 U9513 ( .C1(n7820), .C2(n8824), .A(n7819), .B(n7818), .ZN(P1_U3224) );
  AOI21_X1 U9514 ( .B1(n7822), .B2(n7821), .A(n8211), .ZN(n7825) );
  NOR3_X1 U9515 ( .A1(n7823), .A2(n7828), .A3(n8224), .ZN(n7824) );
  NOR2_X1 U9516 ( .A1(n7825), .A2(n7824), .ZN(n7833) );
  INV_X1 U9517 ( .A(n8535), .ZN(n7826) );
  OAI22_X1 U9518 ( .A1(n8206), .A2(n7826), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9871), .ZN(n7830) );
  OAI22_X1 U9519 ( .A1(n7828), .A2(n7859), .B1(n7827), .B2(n8498), .ZN(n7829)
         );
  AOI211_X1 U9520 ( .C1(n8618), .C2(n8230), .A(n7830), .B(n7829), .ZN(n7831)
         );
  OAI21_X1 U9521 ( .B1(n7833), .B2(n7832), .A(n7831), .ZN(P2_U3240) );
  OR2_X1 U9522 ( .A1(n8371), .A2(n8515), .ZN(n7835) );
  NAND2_X1 U9523 ( .A1(n8437), .A2(n8543), .ZN(n7834) );
  AND2_X1 U9524 ( .A1(n7835), .A2(n7834), .ZN(n8406) );
  INV_X1 U9525 ( .A(n8406), .ZN(n7836) );
  AOI22_X1 U9526 ( .A1(n7836), .A2(n8227), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n7837) );
  OAI21_X1 U9527 ( .B1(n8398), .B2(n8206), .A(n7837), .ZN(n7856) );
  XNOR2_X1 U9528 ( .A(n8397), .B(n7853), .ZN(n8160) );
  NOR2_X1 U9529 ( .A1(n8204), .A2(n8186), .ZN(n7838) );
  NAND2_X1 U9530 ( .A1(n8160), .A2(n7838), .ZN(n8162) );
  OAI21_X1 U9531 ( .B1(n8160), .B2(n7838), .A(n8162), .ZN(n7855) );
  XNOR2_X1 U9532 ( .A(n8467), .B(n7853), .ZN(n7846) );
  INV_X1 U9533 ( .A(n7846), .ZN(n7843) );
  XNOR2_X1 U9534 ( .A(n7847), .B(n7843), .ZN(n7907) );
  NAND2_X1 U9535 ( .A1(n7844), .A2(n7926), .ZN(n7845) );
  NAND2_X1 U9536 ( .A1(n7907), .A2(n7845), .ZN(n7910) );
  OR2_X1 U9537 ( .A1(n7847), .A2(n7846), .ZN(n7848) );
  NAND2_X1 U9538 ( .A1(n8436), .A2(n7926), .ZN(n8174) );
  XNOR2_X1 U9539 ( .A(n8587), .B(n7853), .ZN(n7852) );
  NOR2_X1 U9540 ( .A1(n8210), .A2(n8186), .ZN(n8212) );
  XOR2_X1 U9541 ( .A(n7853), .B(n8583), .Z(n8201) );
  NAND2_X1 U9542 ( .A1(n8437), .A2(n7926), .ZN(n8200) );
  NAND2_X1 U9543 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n8267) );
  OAI21_X1 U9544 ( .B1(n8206), .B2(n7857), .A(n8267), .ZN(n7861) );
  OAI22_X1 U9545 ( .A1(n7859), .A2(n7858), .B1(n4765), .B2(n8220), .ZN(n7860)
         );
  AOI211_X1 U9546 ( .C1(n8216), .C2(n8253), .A(n7861), .B(n7860), .ZN(n7869)
         );
  NAND3_X1 U9547 ( .A1(n8175), .A2(n7862), .A3(n8255), .ZN(n7863) );
  OAI21_X1 U9548 ( .B1(n7864), .B2(n8211), .A(n7863), .ZN(n7867) );
  INV_X1 U9549 ( .A(n7865), .ZN(n7866) );
  NAND2_X1 U9550 ( .A1(n7867), .A2(n7866), .ZN(n7868) );
  OAI211_X1 U9551 ( .C1(n8211), .C2(n7870), .A(n7869), .B(n7868), .ZN(P2_U3233) );
  INV_X1 U9552 ( .A(SI_29_), .ZN(n9677) );
  AND2_X1 U9553 ( .A1(n7871), .A2(n9677), .ZN(n7873) );
  INV_X1 U9554 ( .A(n7871), .ZN(n7872) );
  MUX2_X1 U9555 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n7875), .Z(n7876) );
  NAND2_X1 U9556 ( .A1(n7877), .A2(n7876), .ZN(n7878) );
  MUX2_X1 U9557 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7875), .Z(n7879) );
  XNOR2_X1 U9558 ( .A(n7879), .B(SI_31_), .ZN(n7880) );
  NAND2_X1 U9559 ( .A1(n8682), .A2(n7885), .ZN(n7883) );
  OR2_X1 U9560 ( .A1(n7886), .A2(n6531), .ZN(n7882) );
  NAND2_X1 U9561 ( .A1(n8825), .A2(n7885), .ZN(n7888) );
  INV_X1 U9562 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8147) );
  OR2_X1 U9563 ( .A1(n7886), .A2(n8147), .ZN(n7887) );
  NOR2_X1 U9564 ( .A1(n10376), .A2(n7890), .ZN(n7892) );
  NAND2_X1 U9565 ( .A1(n7919), .A2(n7891), .ZN(n8558) );
  NOR2_X1 U9566 ( .A1(n10389), .A2(n8558), .ZN(n8359) );
  AOI211_X1 U9567 ( .C1(n7922), .C2(n10381), .A(n7892), .B(n8359), .ZN(n7893)
         );
  OAI21_X1 U9568 ( .B1(n8554), .B2(n7894), .A(n7893), .ZN(P2_U3265) );
  INV_X1 U9569 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7899) );
  INV_X1 U9570 ( .A(n7895), .ZN(n7897) );
  AOI211_X1 U9571 ( .C1(n10466), .C2(n7898), .A(n7897), .B(n7896), .ZN(n7901)
         );
  MUX2_X1 U9572 ( .A(n7899), .B(n7901), .S(n10469), .Z(n7900) );
  OAI21_X1 U9573 ( .B1(n7903), .B2(n8678), .A(n7900), .ZN(P2_U3454) );
  MUX2_X1 U9574 ( .A(n6662), .B(n7901), .S(n10477), .Z(n7902) );
  OAI21_X1 U9575 ( .B1(n7903), .B2(n8628), .A(n7902), .ZN(P2_U3521) );
  NOR2_X1 U9576 ( .A1(n8206), .A2(n8469), .ZN(n7906) );
  AOI22_X1 U9577 ( .A1(n8436), .A2(n8544), .B1(n8543), .B2(n8246), .ZN(n8461)
         );
  OAI22_X1 U9578 ( .A1(n8169), .A2(n8461), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7904), .ZN(n7905) );
  AOI211_X1 U9579 ( .C1(n8467), .C2(n8230), .A(n7906), .B(n7905), .ZN(n7909)
         );
  OR3_X1 U9580 ( .A1(n7907), .A2(n8179), .A3(n8224), .ZN(n7908) );
  OAI211_X1 U9581 ( .C1(n7910), .C2(n8211), .A(n7909), .B(n7908), .ZN(P2_U3237) );
  INV_X1 U9582 ( .A(n8833), .ZN(n9559) );
  OAI222_X1 U9583 ( .A1(n7912), .A2(P2_U3152), .B1(n7914), .B2(n9559), .C1(
        n7911), .C2(n8148), .ZN(P2_U3329) );
  OAI222_X1 U9584 ( .A1(n8148), .A2(n7915), .B1(n7914), .B2(n7913), .C1(
        P2_U3152), .C2(n6349), .ZN(P2_U3336) );
  INV_X1 U9585 ( .A(n7916), .ZN(n7918) );
  NOR2_X1 U9586 ( .A1(n8355), .A2(n7920), .ZN(n8088) );
  OAI22_X1 U9587 ( .A1(n7916), .A2(n8088), .B1(n8131), .B2(n7919), .ZN(n7917)
         );
  OAI21_X1 U9588 ( .B1(n7918), .B2(n8355), .A(n7917), .ZN(n7923) );
  INV_X1 U9589 ( .A(n7919), .ZN(n7921) );
  NAND2_X1 U9590 ( .A1(n8355), .A2(n7920), .ZN(n8080) );
  AOI21_X1 U9591 ( .B1(n7923), .B2(n8127), .A(n8090), .ZN(n7924) );
  XNOR2_X1 U9592 ( .A(n7924), .B(n8350), .ZN(n8136) );
  INV_X1 U9593 ( .A(n7927), .ZN(n8013) );
  NAND2_X1 U9594 ( .A1(n7930), .A2(n7935), .ZN(n7929) );
  NAND2_X1 U9595 ( .A1(n7958), .A2(n7960), .ZN(n7928) );
  MUX2_X1 U9596 ( .A(n7929), .B(n7928), .S(n8093), .Z(n7957) );
  INV_X1 U9597 ( .A(n7930), .ZN(n7933) );
  INV_X1 U9598 ( .A(n7931), .ZN(n7932) );
  NOR2_X1 U9599 ( .A1(n7933), .A2(n7932), .ZN(n7936) );
  OAI211_X1 U9600 ( .C1(n7957), .C2(n7936), .A(n7935), .B(n7934), .ZN(n7956)
         );
  INV_X1 U9601 ( .A(n7937), .ZN(n7949) );
  INV_X1 U9602 ( .A(n7938), .ZN(n7939) );
  AOI211_X1 U9603 ( .C1(n7945), .C2(n7943), .A(n7949), .B(n7939), .ZN(n7941)
         );
  INV_X1 U9604 ( .A(n7940), .ZN(n7946) );
  NOR2_X1 U9605 ( .A1(n7941), .A2(n7946), .ZN(n7952) );
  INV_X1 U9606 ( .A(n7945), .ZN(n7947) );
  NOR3_X1 U9607 ( .A1(n7948), .A2(n7947), .A3(n7946), .ZN(n7950) );
  NOR2_X1 U9608 ( .A1(n7950), .A2(n7949), .ZN(n7951) );
  MUX2_X1 U9609 ( .A(n7952), .B(n7951), .S(n8093), .Z(n7954) );
  NOR3_X1 U9610 ( .A1(n7954), .A2(n7957), .A3(n7953), .ZN(n7955) );
  AOI21_X1 U9611 ( .B1(n8093), .B2(n7956), .A(n7955), .ZN(n7965) );
  NOR2_X1 U9612 ( .A1(n7966), .A2(n10347), .ZN(n7964) );
  AOI21_X1 U9613 ( .B1(n7959), .B2(n7958), .A(n7957), .ZN(n7962) );
  INV_X1 U9614 ( .A(n7960), .ZN(n7961) );
  NOR3_X1 U9615 ( .A1(n7962), .A2(n7961), .A3(n7964), .ZN(n7963) );
  OAI22_X1 U9616 ( .A1(n7965), .A2(n7964), .B1(n7963), .B2(n8093), .ZN(n7974)
         );
  INV_X1 U9617 ( .A(n7966), .ZN(n8257) );
  NOR2_X1 U9618 ( .A1(n8257), .A2(n8093), .ZN(n7967) );
  AOI21_X1 U9619 ( .B1(n7967), .B2(n10347), .A(n8107), .ZN(n7973) );
  INV_X1 U9620 ( .A(n7968), .ZN(n7971) );
  INV_X1 U9621 ( .A(n7969), .ZN(n7970) );
  MUX2_X1 U9622 ( .A(n7971), .B(n7970), .S(n8093), .Z(n7972) );
  AOI211_X1 U9623 ( .C1(n7974), .C2(n7973), .A(n4486), .B(n7972), .ZN(n7980)
         );
  NOR2_X1 U9624 ( .A1(n10448), .A2(n8093), .ZN(n7977) );
  INV_X1 U9625 ( .A(n8093), .ZN(n8089) );
  NOR2_X1 U9626 ( .A1(n7975), .A2(n8089), .ZN(n7976) );
  MUX2_X1 U9627 ( .A(n7977), .B(n7976), .S(n8255), .Z(n7978) );
  NOR3_X1 U9628 ( .A1(n7980), .A2(n7979), .A3(n7978), .ZN(n7985) );
  INV_X1 U9629 ( .A(n7988), .ZN(n7983) );
  AOI21_X1 U9630 ( .B1(n7986), .B2(n7981), .A(n8089), .ZN(n7982) );
  NAND2_X1 U9631 ( .A1(n8001), .A2(n7986), .ZN(n7991) );
  INV_X1 U9632 ( .A(n7986), .ZN(n7989) );
  OAI211_X1 U9633 ( .C1(n7989), .C2(n7988), .A(n7994), .B(n7987), .ZN(n7990)
         );
  INV_X1 U9634 ( .A(n8002), .ZN(n7997) );
  INV_X1 U9635 ( .A(n7993), .ZN(n7996) );
  INV_X1 U9636 ( .A(n7994), .ZN(n7995) );
  INV_X1 U9637 ( .A(n7998), .ZN(n7999) );
  NOR2_X1 U9638 ( .A1(n8000), .A2(n7999), .ZN(n8007) );
  OAI21_X1 U9639 ( .B1(n4525), .B2(n4870), .A(n8005), .ZN(n8006) );
  MUX2_X1 U9640 ( .A(n8007), .B(n8006), .S(n8093), .Z(n8008) );
  NOR2_X1 U9641 ( .A1(n8008), .A2(n8115), .ZN(n8016) );
  NAND2_X1 U9642 ( .A1(n4812), .A2(n8009), .ZN(n8011) );
  OAI21_X1 U9643 ( .B1(n8016), .B2(n8011), .A(n8010), .ZN(n8012) );
  INV_X1 U9644 ( .A(n8018), .ZN(n8021) );
  INV_X1 U9645 ( .A(n8019), .ZN(n8020) );
  MUX2_X1 U9646 ( .A(n8021), .B(n8020), .S(n8093), .Z(n8023) );
  INV_X1 U9647 ( .A(n8024), .ZN(n8027) );
  INV_X1 U9648 ( .A(n8025), .ZN(n8026) );
  MUX2_X1 U9649 ( .A(n8027), .B(n8026), .S(n8093), .Z(n8028) );
  NAND2_X1 U9650 ( .A1(n8041), .A2(n8029), .ZN(n8032) );
  INV_X1 U9651 ( .A(n8030), .ZN(n8031) );
  MUX2_X1 U9652 ( .A(n8032), .B(n8031), .S(n8093), .Z(n8033) );
  NOR2_X1 U9653 ( .A1(n8034), .A2(n8033), .ZN(n8044) );
  INV_X1 U9654 ( .A(n8507), .ZN(n8035) );
  OAI21_X1 U9655 ( .B1(n8044), .B2(n8035), .A(n8045), .ZN(n8036) );
  NAND3_X1 U9656 ( .A1(n8036), .A2(n8048), .A3(n8042), .ZN(n8037) );
  NAND3_X1 U9657 ( .A1(n8037), .A2(n8046), .A3(n8050), .ZN(n8040) );
  INV_X1 U9658 ( .A(n8444), .ZN(n8055) );
  NOR2_X1 U9659 ( .A1(n8603), .A2(n8499), .ZN(n8049) );
  NOR2_X1 U9660 ( .A1(n8055), .A2(n8049), .ZN(n8039) );
  INV_X1 U9661 ( .A(n8054), .ZN(n8038) );
  INV_X1 U9662 ( .A(n8041), .ZN(n8043) );
  OAI211_X1 U9663 ( .C1(n8044), .C2(n8043), .A(n8042), .B(n8507), .ZN(n8047)
         );
  NAND3_X1 U9664 ( .A1(n8047), .A2(n8046), .A3(n8045), .ZN(n8053) );
  NOR2_X1 U9665 ( .A1(n8049), .A2(n4945), .ZN(n8052) );
  INV_X1 U9666 ( .A(n8050), .ZN(n8051) );
  AOI21_X1 U9667 ( .B1(n8053), .B2(n8052), .A(n8051), .ZN(n8056) );
  OAI21_X1 U9668 ( .B1(n8056), .B2(n8055), .A(n8054), .ZN(n8057) );
  OAI21_X1 U9669 ( .B1(n8089), .B2(n8060), .A(n8059), .ZN(n8061) );
  INV_X1 U9670 ( .A(n8062), .ZN(n8064) );
  AOI21_X1 U9671 ( .B1(n8455), .B2(n8436), .A(n8064), .ZN(n8063) );
  NAND3_X1 U9672 ( .A1(n8587), .A2(n8210), .A3(n8089), .ZN(n8065) );
  OAI211_X1 U9673 ( .C1(n8402), .C2(n8093), .A(n8066), .B(n8071), .ZN(n8070)
         );
  NAND2_X1 U9674 ( .A1(n8069), .A2(n8067), .ZN(n8068) );
  AOI22_X1 U9675 ( .A1(n8070), .A2(n8069), .B1(n8093), .B2(n8068), .ZN(n8076)
         );
  OAI21_X1 U9676 ( .B1(n8089), .B2(n8071), .A(n4636), .ZN(n8075) );
  MUX2_X1 U9677 ( .A(n8073), .B(n8072), .S(n8093), .Z(n8074) );
  OAI211_X1 U9678 ( .C1(n8076), .C2(n8075), .A(n4964), .B(n8074), .ZN(n8079)
         );
  NAND3_X1 U9679 ( .A1(n8367), .A2(n8243), .A3(n8093), .ZN(n8078) );
  NAND3_X1 U9680 ( .A1(n8567), .A2(n8187), .A3(n8089), .ZN(n8077) );
  NAND4_X1 U9681 ( .A1(n8079), .A2(n8125), .A3(n8078), .A4(n8077), .ZN(n8087)
         );
  INV_X1 U9682 ( .A(n8080), .ZN(n8084) );
  MUX2_X1 U9683 ( .A(n4962), .B(n8082), .S(n8093), .Z(n8083) );
  NOR3_X1 U9684 ( .A1(n8088), .A2(n8084), .A3(n8083), .ZN(n8086) );
  AOI22_X1 U9685 ( .A1(n8087), .A2(n8086), .B1(n8089), .B2(n8085), .ZN(n8091)
         );
  OAI22_X1 U9686 ( .A1(n8091), .A2(n8090), .B1(n8126), .B2(n8089), .ZN(n8096)
         );
  INV_X1 U9687 ( .A(n8092), .ZN(n8094) );
  NAND2_X1 U9688 ( .A1(n8094), .A2(n8093), .ZN(n8095) );
  INV_X1 U9689 ( .A(n8434), .ZN(n8123) );
  NOR3_X1 U9690 ( .A1(n8101), .A2(n8100), .A3(n8099), .ZN(n8102) );
  NAND4_X1 U9691 ( .A1(n8105), .A2(n8104), .A3(n8103), .A4(n8102), .ZN(n8106)
         );
  NOR4_X1 U9692 ( .A1(n10345), .A2(n8107), .A3(n8106), .A4(n6332), .ZN(n8109)
         );
  NAND4_X1 U9693 ( .A1(n8111), .A2(n8110), .A3(n8109), .A4(n8108), .ZN(n8113)
         );
  NOR4_X1 U9694 ( .A1(n8115), .A2(n8114), .A3(n8113), .A4(n8112), .ZN(n8116)
         );
  NAND4_X1 U9695 ( .A1(n8118), .A2(n8117), .A3(n4812), .A4(n8116), .ZN(n8119)
         );
  NOR4_X1 U9696 ( .A1(n8508), .A2(n4944), .A3(n8120), .A4(n8119), .ZN(n8121)
         );
  NAND4_X1 U9697 ( .A1(n6344), .A2(n8490), .A3(n8121), .A4(n6342), .ZN(n8122)
         );
  NOR4_X1 U9698 ( .A1(n4798), .A2(n8123), .A3(n8449), .A4(n8122), .ZN(n8124)
         );
  XNOR2_X1 U9699 ( .A(n5066), .B(n8350), .ZN(n8132) );
  INV_X1 U9700 ( .A(n8128), .ZN(n8130) );
  AOI22_X1 U9701 ( .A1(n8132), .A2(n8131), .B1(n8130), .B2(n8129), .ZN(n8134)
         );
  INV_X1 U9702 ( .A(n6351), .ZN(n8137) );
  NAND3_X1 U9703 ( .A1(n8138), .A2(n8137), .A3(n8350), .ZN(n8139) );
  NOR3_X1 U9704 ( .A1(n10390), .A2(n8140), .A3(n8139), .ZN(n8142) );
  MUX2_X1 U9705 ( .A(n8143), .B(n8142), .S(n8141), .Z(n8144) );
  OAI22_X1 U9706 ( .A1(n8146), .A2(n8145), .B1(n8144), .B2(n9869), .ZN(
        P2_U3244) );
  INV_X1 U9707 ( .A(n8825), .ZN(n8152) );
  OAI222_X1 U9708 ( .A1(n8148), .A2(n8147), .B1(n8686), .B2(n8152), .C1(n5921), 
        .C2(P2_U3152), .ZN(P2_U3328) );
  INV_X1 U9709 ( .A(n8149), .ZN(n8150) );
  OAI222_X1 U9710 ( .A1(n9562), .A2(n9878), .B1(P1_U3084), .B2(n5850), .C1(
        n9560), .C2(n8150), .ZN(P1_U3325) );
  INV_X1 U9711 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9737) );
  OAI222_X1 U9712 ( .A1(n9553), .A2(n9737), .B1(n9560), .B2(n8152), .C1(n8151), 
        .C2(P1_U3084), .ZN(P1_U3323) );
  XNOR2_X1 U9713 ( .A(n8572), .B(n7853), .ZN(n8153) );
  NOR2_X1 U9714 ( .A1(n8371), .A2(n8186), .ZN(n8154) );
  NAND2_X1 U9715 ( .A1(n8153), .A2(n8154), .ZN(n8184) );
  INV_X1 U9716 ( .A(n8153), .ZN(n8156) );
  INV_X1 U9717 ( .A(n8154), .ZN(n8155) );
  NAND2_X1 U9718 ( .A1(n8156), .A2(n8155), .ZN(n8157) );
  INV_X1 U9719 ( .A(n8163), .ZN(n8158) );
  AOI21_X1 U9720 ( .B1(n8159), .B2(n8158), .A(n8211), .ZN(n8167) );
  INV_X1 U9721 ( .A(n8160), .ZN(n8161) );
  NOR3_X1 U9722 ( .A1(n8161), .A2(n8204), .A3(n8224), .ZN(n8166) );
  INV_X1 U9723 ( .A(n8162), .ZN(n8164) );
  OAI21_X1 U9724 ( .B1(n8167), .B2(n8166), .A(n8185), .ZN(n8173) );
  OAI22_X1 U9725 ( .A1(n8187), .A2(n8515), .B1(n8204), .B2(n8513), .ZN(n8388)
         );
  INV_X1 U9726 ( .A(n8388), .ZN(n8170) );
  OAI22_X1 U9727 ( .A1(n8170), .A2(n8169), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8168), .ZN(n8171) );
  AOI21_X1 U9728 ( .B1(n8382), .B2(n8229), .A(n8171), .ZN(n8172) );
  OAI211_X1 U9729 ( .C1(n8384), .C2(n8220), .A(n8173), .B(n8172), .ZN(P2_U3216) );
  NAND2_X1 U9730 ( .A1(n8235), .A2(n8174), .ZN(n8178) );
  NAND2_X1 U9731 ( .A1(n8175), .A2(n8436), .ZN(n8177) );
  MUX2_X1 U9732 ( .A(n8178), .B(n8177), .S(n8176), .Z(n8183) );
  AOI22_X1 U9733 ( .A1(n8229), .A2(n8453), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8182) );
  AOI22_X1 U9734 ( .A1(n8216), .A2(n4801), .B1(n8217), .B2(n7844), .ZN(n8181)
         );
  NAND2_X1 U9735 ( .A1(n8593), .A2(n8230), .ZN(n8180) );
  NAND4_X1 U9736 ( .A1(n8183), .A2(n8182), .A3(n8181), .A4(n8180), .ZN(
        P2_U3218) );
  NOR2_X1 U9737 ( .A1(n8187), .A2(n8186), .ZN(n8188) );
  XNOR2_X1 U9738 ( .A(n8188), .B(n7853), .ZN(n8190) );
  INV_X1 U9739 ( .A(n8190), .ZN(n8191) );
  NOR3_X1 U9740 ( .A1(n8367), .A2(n8230), .A3(n8191), .ZN(n8189) );
  AOI21_X1 U9741 ( .B1(n8367), .B2(n8191), .A(n8189), .ZN(n8196) );
  OAI21_X1 U9742 ( .B1(n8367), .B2(n8220), .A(n8211), .ZN(n8195) );
  NOR3_X1 U9743 ( .A1(n8367), .A2(n8190), .A3(n8230), .ZN(n8193) );
  NOR2_X1 U9744 ( .A1(n8567), .A2(n8191), .ZN(n8192) );
  INV_X1 U9745 ( .A(n8197), .ZN(n8365) );
  AOI22_X1 U9746 ( .A1(n8365), .A2(n8229), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n8199) );
  INV_X1 U9747 ( .A(n8372), .ZN(n8242) );
  AOI22_X1 U9748 ( .A1(n8216), .A2(n8242), .B1(n8244), .B2(n8217), .ZN(n8198)
         );
  XNOR2_X1 U9749 ( .A(n8201), .B(n8200), .ZN(n8202) );
  XNOR2_X1 U9750 ( .A(n8203), .B(n8202), .ZN(n8209) );
  OAI22_X1 U9751 ( .A1(n8204), .A2(n8515), .B1(n8210), .B2(n8513), .ZN(n8419)
         );
  AOI22_X1 U9752 ( .A1(n8419), .A2(n8227), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8205) );
  OAI21_X1 U9753 ( .B1(n8413), .B2(n8206), .A(n8205), .ZN(n8207) );
  AOI21_X1 U9754 ( .B1(n8583), .B2(n8230), .A(n8207), .ZN(n8208) );
  OAI21_X1 U9755 ( .B1(n8209), .B2(n8211), .A(n8208), .ZN(P2_U3227) );
  NOR2_X1 U9756 ( .A1(n8224), .A2(n8210), .ZN(n8215) );
  NOR2_X1 U9757 ( .A1(n8212), .A2(n8211), .ZN(n8214) );
  MUX2_X1 U9758 ( .A(n8215), .B(n8214), .S(n8213), .Z(n8222) );
  AOI22_X1 U9759 ( .A1(n8229), .A2(n8430), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n8219) );
  AOI22_X1 U9760 ( .A1(n8217), .A2(n8436), .B1(n8216), .B2(n8437), .ZN(n8218)
         );
  OAI211_X1 U9761 ( .C1(n8432), .C2(n8220), .A(n8219), .B(n8218), .ZN(n8221)
         );
  OR2_X1 U9762 ( .A1(n8222), .A2(n8221), .ZN(P2_U3231) );
  OR4_X1 U9763 ( .A1(n8224), .A2(n8223), .A3(n8226), .A4(n8234), .ZN(n8240) );
  OAI22_X1 U9764 ( .A1(n8226), .A2(n8513), .B1(n8225), .B2(n8515), .ZN(n10339)
         );
  AOI22_X1 U9765 ( .A1(n8227), .A2(n10339), .B1(P2_REG3_REG_6__SCAN_IN), .B2(
        P2_U3152), .ZN(n8239) );
  INV_X1 U9766 ( .A(n8228), .ZN(n10341) );
  AOI22_X1 U9767 ( .A1(n10347), .A2(n8230), .B1(n8229), .B2(n10341), .ZN(n8238) );
  NAND2_X1 U9768 ( .A1(n8233), .A2(n8231), .ZN(n8232) );
  OAI21_X1 U9769 ( .B1(n8234), .B2(n8233), .A(n8232), .ZN(n8236) );
  NAND2_X1 U9770 ( .A1(n8236), .A2(n8235), .ZN(n8237) );
  NAND4_X1 U9771 ( .A1(n8240), .A2(n8239), .A3(n8238), .A4(n8237), .ZN(
        P2_U3241) );
  MUX2_X1 U9772 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8241), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9773 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8242), .S(P2_U3966), .Z(
        P2_U3581) );
  MUX2_X1 U9774 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8243), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U9775 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8244), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U9776 ( .A(n8437), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8245), .Z(
        P2_U3577) );
  MUX2_X1 U9777 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n4801), .S(P2_U3966), .Z(
        P2_U3576) );
  MUX2_X1 U9778 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8436), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U9779 ( .A(n7844), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8245), .Z(
        P2_U3574) );
  MUX2_X1 U9780 ( .A(n8246), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8245), .Z(
        P2_U3573) );
  MUX2_X1 U9781 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8545), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9782 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8247), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9783 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8542), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9784 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8248), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9785 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8249), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9786 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8250), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9787 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8251), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9788 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n4870), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U9789 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8252), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U9790 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8253), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U9791 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8254), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U9792 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8255), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U9793 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8256), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U9794 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8257), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U9795 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8258), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U9796 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8259), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U9797 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8260), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U9798 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n5971), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U9799 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8261), .S(P2_U3966), .Z(
        P2_U3553) );
  MUX2_X1 U9800 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8262), .S(P2_U3966), .Z(
        P2_U3552) );
  AOI211_X1 U9801 ( .C1(n8265), .C2(n8264), .A(n8263), .B(n9988), .ZN(n8266)
         );
  INV_X1 U9802 ( .A(n8266), .ZN(n8276) );
  INV_X1 U9803 ( .A(n8267), .ZN(n8268) );
  AOI21_X1 U9804 ( .B1(n10333), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8268), .ZN(
        n8275) );
  OAI211_X1 U9805 ( .C1(n8271), .C2(n8270), .A(n10330), .B(n8269), .ZN(n8274)
         );
  NAND2_X1 U9806 ( .A1(n9994), .A2(n8272), .ZN(n8273) );
  NAND4_X1 U9807 ( .A1(n8276), .A2(n8275), .A3(n8274), .A4(n8273), .ZN(
        P2_U3254) );
  OAI21_X1 U9808 ( .B1(n8278), .B2(P2_REG2_REG_14__SCAN_IN), .A(n8277), .ZN(
        n8296) );
  XNOR2_X1 U9809 ( .A(n8291), .B(n8296), .ZN(n8279) );
  NAND2_X1 U9810 ( .A1(n8279), .A2(n7527), .ZN(n8298) );
  OAI21_X1 U9811 ( .B1(n8279), .B2(n7527), .A(n8298), .ZN(n8288) );
  AOI21_X1 U9812 ( .B1(n8282), .B2(n8281), .A(n8280), .ZN(n8290) );
  XNOR2_X1 U9813 ( .A(n8290), .B(n8297), .ZN(n8283) );
  NAND2_X1 U9814 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8283), .ZN(n8292) );
  OAI211_X1 U9815 ( .C1(n8283), .C2(P2_REG1_REG_15__SCAN_IN), .A(n10330), .B(
        n8292), .ZN(n8286) );
  AND2_X1 U9816 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8284) );
  AOI21_X1 U9817 ( .B1(n10333), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8284), .ZN(
        n8285) );
  OAI211_X1 U9818 ( .C1(n10327), .C2(n8297), .A(n8286), .B(n8285), .ZN(n8287)
         );
  AOI21_X1 U9819 ( .B1(n8288), .B2(n10331), .A(n8287), .ZN(n8289) );
  INV_X1 U9820 ( .A(n8289), .ZN(P2_U3260) );
  NAND2_X1 U9821 ( .A1(n8291), .A2(n8290), .ZN(n8293) );
  NAND2_X1 U9822 ( .A1(n8293), .A2(n8292), .ZN(n8295) );
  XNOR2_X1 U9823 ( .A(n8313), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8294) );
  NOR2_X1 U9824 ( .A1(n8295), .A2(n8294), .ZN(n8316) );
  AOI21_X1 U9825 ( .B1(n8295), .B2(n8294), .A(n8316), .ZN(n8309) );
  NAND2_X1 U9826 ( .A1(n8297), .A2(n8296), .ZN(n8299) );
  XNOR2_X1 U9827 ( .A(n8313), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n8300) );
  AOI211_X1 U9828 ( .C1(n8301), .C2(n8300), .A(n9988), .B(n8310), .ZN(n8302)
         );
  INV_X1 U9829 ( .A(n8302), .ZN(n8308) );
  INV_X1 U9830 ( .A(n8303), .ZN(n8306) );
  NOR2_X1 U9831 ( .A1(n10327), .A2(n8304), .ZN(n8305) );
  AOI211_X1 U9832 ( .C1(P2_ADDR_REG_16__SCAN_IN), .C2(n10333), .A(n8306), .B(
        n8305), .ZN(n8307) );
  OAI211_X1 U9833 ( .C1(n8309), .C2(n10328), .A(n8308), .B(n8307), .ZN(
        P2_U3261) );
  NAND2_X1 U9834 ( .A1(n8324), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8311) );
  OAI21_X1 U9835 ( .B1(n8324), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8311), .ZN(
        n8312) );
  AOI211_X1 U9836 ( .C1(n4562), .C2(n8312), .A(n8323), .B(n9988), .ZN(n8322)
         );
  NOR2_X1 U9837 ( .A1(n8313), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8315) );
  XNOR2_X1 U9838 ( .A(n8324), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8314) );
  OAI21_X1 U9839 ( .B1(n8316), .B2(n8315), .A(n8314), .ZN(n8317) );
  OR3_X1 U9840 ( .A1(n8316), .A2(n8315), .A3(n8314), .ZN(n8327) );
  NAND3_X1 U9841 ( .A1(n8317), .A2(n10330), .A3(n8327), .ZN(n8320) );
  NOR2_X1 U9842 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9949), .ZN(n8318) );
  AOI21_X1 U9843 ( .B1(n10333), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8318), .ZN(
        n8319) );
  OAI211_X1 U9844 ( .C1(n10327), .C2(n8328), .A(n8320), .B(n8319), .ZN(n8321)
         );
  OR2_X1 U9845 ( .A1(n8322), .A2(n8321), .ZN(P2_U3262) );
  XNOR2_X1 U9846 ( .A(n8338), .B(n8344), .ZN(n8326) );
  INV_X1 U9847 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8325) );
  NOR2_X1 U9848 ( .A1(n8325), .A2(n8326), .ZN(n8339) );
  AOI211_X1 U9849 ( .C1(n8326), .C2(n8325), .A(n8339), .B(n9988), .ZN(n8337)
         );
  INV_X1 U9850 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8626) );
  OAI21_X1 U9851 ( .B1(n8626), .B2(n8328), .A(n8327), .ZN(n8331) );
  XNOR2_X1 U9852 ( .A(n8329), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8330) );
  NOR2_X1 U9853 ( .A1(n8331), .A2(n8330), .ZN(n8342) );
  AOI21_X1 U9854 ( .B1(n8331), .B2(n8330), .A(n8342), .ZN(n8332) );
  NOR2_X1 U9855 ( .A1(n8332), .A2(n10328), .ZN(n8336) );
  NOR2_X1 U9856 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9871), .ZN(n8333) );
  AOI21_X1 U9857 ( .B1(n10333), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8333), .ZN(
        n8334) );
  OAI21_X1 U9858 ( .B1(n10327), .B2(n8344), .A(n8334), .ZN(n8335) );
  OR3_X1 U9859 ( .A1(n8337), .A2(n8336), .A3(n8335), .ZN(P2_U3263) );
  NOR2_X1 U9860 ( .A1(n8338), .A2(n8344), .ZN(n8340) );
  NOR2_X1 U9861 ( .A1(n8340), .A2(n8339), .ZN(n8341) );
  XNOR2_X1 U9862 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8341), .ZN(n8349) );
  INV_X1 U9863 ( .A(n8349), .ZN(n8347) );
  AOI21_X1 U9864 ( .B1(n8344), .B2(n8343), .A(n8342), .ZN(n8345) );
  XNOR2_X1 U9865 ( .A(n8616), .B(n8345), .ZN(n8348) );
  OAI21_X1 U9866 ( .B1(n8348), .B2(n10328), .A(n10327), .ZN(n8346) );
  AOI21_X1 U9867 ( .B1(n8347), .B2(n10331), .A(n8346), .ZN(n8352) );
  AOI22_X1 U9868 ( .A1(n8349), .A2(n10331), .B1(n10330), .B2(n8348), .ZN(n8351) );
  MUX2_X1 U9869 ( .A(n8352), .B(n8351), .S(n8350), .Z(n8354) );
  NAND2_X1 U9870 ( .A1(n10333), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8353) );
  OAI211_X1 U9871 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n5931), .A(n8354), .B(n8353), .ZN(P2_U3264) );
  OAI211_X1 U9872 ( .C1(n7889), .C2(n8357), .A(n10360), .B(n8356), .ZN(n8559)
         );
  NOR2_X1 U9873 ( .A1(n7889), .A2(n8537), .ZN(n8358) );
  AOI211_X1 U9874 ( .C1(n10389), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8359), .B(
        n8358), .ZN(n8360) );
  OAI21_X1 U9875 ( .B1(n8361), .B2(n8559), .A(n8360), .ZN(P2_U3266) );
  XNOR2_X1 U9876 ( .A(n8362), .B(n4964), .ZN(n8571) );
  INV_X1 U9877 ( .A(n8363), .ZN(n8364) );
  AOI21_X1 U9878 ( .B1(n8567), .B2(n8379), .A(n8364), .ZN(n8568) );
  AOI22_X1 U9879 ( .A1(n8365), .A2(n10379), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n8548), .ZN(n8366) );
  OAI21_X1 U9880 ( .B1(n8367), .B2(n8537), .A(n8366), .ZN(n8376) );
  AOI211_X1 U9881 ( .C1(n8370), .C2(n8369), .A(n8510), .B(n8368), .ZN(n8374)
         );
  OAI22_X1 U9882 ( .A1(n8372), .A2(n8515), .B1(n8371), .B2(n8513), .ZN(n8373)
         );
  NOR2_X1 U9883 ( .A1(n8374), .A2(n8373), .ZN(n8570) );
  NOR2_X1 U9884 ( .A1(n8570), .A2(n8548), .ZN(n8375) );
  AOI211_X1 U9885 ( .C1(n8551), .C2(n8568), .A(n8376), .B(n8375), .ZN(n8377)
         );
  OAI21_X1 U9886 ( .B1(n8571), .B2(n8553), .A(n8377), .ZN(P2_U3268) );
  XNOR2_X1 U9887 ( .A(n8378), .B(n8386), .ZN(n8576) );
  INV_X1 U9888 ( .A(n8396), .ZN(n8381) );
  INV_X1 U9889 ( .A(n8379), .ZN(n8380) );
  AOI21_X1 U9890 ( .B1(n8572), .B2(n8381), .A(n8380), .ZN(n8573) );
  AOI22_X1 U9891 ( .A1(P2_REG2_REG_27__SCAN_IN), .A2(n10389), .B1(n8382), .B2(
        n10379), .ZN(n8383) );
  OAI21_X1 U9892 ( .B1(n8384), .B2(n8537), .A(n8383), .ZN(n8392) );
  NOR2_X1 U9893 ( .A1(n8385), .A2(n8510), .ZN(n8390) );
  OAI21_X1 U9894 ( .B1(n8404), .B2(n8387), .A(n8386), .ZN(n8389) );
  AOI21_X1 U9895 ( .B1(n8390), .B2(n8389), .A(n8388), .ZN(n8575) );
  NOR2_X1 U9896 ( .A1(n8575), .A2(n8548), .ZN(n8391) );
  AOI211_X1 U9897 ( .C1(n8551), .C2(n8573), .A(n8392), .B(n8391), .ZN(n8393)
         );
  OAI21_X1 U9898 ( .B1(n8576), .B2(n8553), .A(n8393), .ZN(P2_U3269) );
  XNOR2_X1 U9899 ( .A(n8395), .B(n8394), .ZN(n8579) );
  INV_X1 U9900 ( .A(n8579), .ZN(n8410) );
  AOI211_X1 U9901 ( .C1(n8397), .C2(n8412), .A(n10462), .B(n8396), .ZN(n8578)
         );
  NOR2_X1 U9902 ( .A1(n8660), .A2(n8537), .ZN(n8401) );
  OAI22_X1 U9903 ( .A1(n10376), .A2(n8399), .B1(n8398), .B2(n8468), .ZN(n8400)
         );
  AOI211_X1 U9904 ( .C1(n8578), .C2(n8522), .A(n8401), .B(n8400), .ZN(n8409)
         );
  AOI21_X1 U9905 ( .B1(n8420), .B2(n8402), .A(n4791), .ZN(n8403) );
  NAND2_X1 U9906 ( .A1(n8405), .A2(n10369), .ZN(n8407) );
  NAND2_X1 U9907 ( .A1(n8407), .A2(n8406), .ZN(n8577) );
  NAND2_X1 U9908 ( .A1(n8577), .A2(n10376), .ZN(n8408) );
  OAI211_X1 U9909 ( .C1(n8410), .C2(n8553), .A(n8409), .B(n8408), .ZN(P2_U3270) );
  XNOR2_X1 U9910 ( .A(n8411), .B(n4798), .ZN(n8586) );
  AOI211_X1 U9911 ( .C1(n8583), .C2(n8427), .A(n10462), .B(n6359), .ZN(n8582)
         );
  INV_X1 U9912 ( .A(n8583), .ZN(n8416) );
  INV_X1 U9913 ( .A(n8413), .ZN(n8414) );
  AOI22_X1 U9914 ( .A1(n8548), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8414), .B2(
        n10379), .ZN(n8415) );
  OAI21_X1 U9915 ( .B1(n8416), .B2(n8537), .A(n8415), .ZN(n8423) );
  INV_X1 U9916 ( .A(n8417), .ZN(n8418) );
  AOI21_X1 U9917 ( .B1(n8418), .B2(n4798), .A(n8510), .ZN(n8421) );
  AOI21_X1 U9918 ( .B1(n8421), .B2(n8420), .A(n8419), .ZN(n8585) );
  NOR2_X1 U9919 ( .A1(n8585), .A2(n8548), .ZN(n8422) );
  AOI211_X1 U9920 ( .C1(n8522), .C2(n8582), .A(n8423), .B(n8422), .ZN(n8424)
         );
  OAI21_X1 U9921 ( .B1(n8586), .B2(n8553), .A(n8424), .ZN(P2_U3271) );
  AOI21_X1 U9922 ( .B1(n8434), .B2(n8426), .A(n8425), .ZN(n8591) );
  INV_X1 U9923 ( .A(n8452), .ZN(n8429) );
  INV_X1 U9924 ( .A(n8427), .ZN(n8428) );
  AOI21_X1 U9925 ( .B1(n8587), .B2(n8429), .A(n8428), .ZN(n8588) );
  AOI22_X1 U9926 ( .A1(n10389), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8430), .B2(
        n10379), .ZN(n8431) );
  OAI21_X1 U9927 ( .B1(n8432), .B2(n8537), .A(n8431), .ZN(n8441) );
  OAI211_X1 U9928 ( .C1(n8435), .C2(n8434), .A(n8433), .B(n10369), .ZN(n8439)
         );
  AOI22_X1 U9929 ( .A1(n8437), .A2(n8544), .B1(n8543), .B2(n8436), .ZN(n8438)
         );
  NOR2_X1 U9930 ( .A1(n8590), .A2(n10389), .ZN(n8440) );
  AOI211_X1 U9931 ( .C1(n8588), .C2(n8551), .A(n8441), .B(n8440), .ZN(n8442)
         );
  OAI21_X1 U9932 ( .B1(n8591), .B2(n8553), .A(n8442), .ZN(P2_U3272) );
  AND2_X1 U9933 ( .A1(n8443), .A2(n8444), .ZN(n8447) );
  OAI21_X1 U9934 ( .B1(n8447), .B2(n8446), .A(n8445), .ZN(n8448) );
  AOI222_X1 U9935 ( .A1(n10369), .A2(n8448), .B1(n7844), .B2(n8543), .C1(n4801), .C2(n8544), .ZN(n8596) );
  OR2_X1 U9936 ( .A1(n8450), .A2(n8449), .ZN(n8592) );
  NAND3_X1 U9937 ( .A1(n8592), .A2(n8451), .A3(n10352), .ZN(n8458) );
  AOI21_X1 U9938 ( .B1(n8593), .B2(n8465), .A(n8452), .ZN(n8594) );
  AOI22_X1 U9939 ( .A1(n10389), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8453), .B2(
        n10379), .ZN(n8454) );
  OAI21_X1 U9940 ( .B1(n8455), .B2(n8537), .A(n8454), .ZN(n8456) );
  AOI21_X1 U9941 ( .B1(n8594), .B2(n8551), .A(n8456), .ZN(n8457) );
  OAI211_X1 U9942 ( .C1(n10389), .C2(n8596), .A(n8458), .B(n8457), .ZN(
        P2_U3273) );
  NAND2_X1 U9943 ( .A1(n8459), .A2(n8463), .ZN(n8460) );
  NAND3_X1 U9944 ( .A1(n8443), .A2(n10369), .A3(n8460), .ZN(n8462) );
  NAND2_X1 U9945 ( .A1(n8462), .A2(n8461), .ZN(n8598) );
  INV_X1 U9946 ( .A(n8598), .ZN(n8475) );
  XNOR2_X1 U9947 ( .A(n8464), .B(n8463), .ZN(n8600) );
  NAND2_X1 U9948 ( .A1(n8600), .A2(n10352), .ZN(n8474) );
  INV_X1 U9949 ( .A(n8465), .ZN(n8466) );
  AOI211_X1 U9950 ( .C1(n8467), .C2(n8477), .A(n10462), .B(n8466), .ZN(n8599)
         );
  NOR2_X1 U9951 ( .A1(n8667), .A2(n8537), .ZN(n8472) );
  OAI22_X1 U9952 ( .A1(n10376), .A2(n8470), .B1(n8469), .B2(n8468), .ZN(n8471)
         );
  AOI211_X1 U9953 ( .C1(n8599), .C2(n10383), .A(n8472), .B(n8471), .ZN(n8473)
         );
  OAI211_X1 U9954 ( .C1(n8548), .C2(n8475), .A(n8474), .B(n8473), .ZN(P2_U3274) );
  XNOR2_X1 U9955 ( .A(n8476), .B(n8483), .ZN(n8607) );
  INV_X1 U9956 ( .A(n8477), .ZN(n8478) );
  AOI21_X1 U9957 ( .B1(n8603), .B2(n4774), .A(n8478), .ZN(n8604) );
  INV_X1 U9958 ( .A(n8479), .ZN(n8480) );
  AOI22_X1 U9959 ( .A1(n10389), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8480), .B2(
        n10379), .ZN(n8481) );
  OAI21_X1 U9960 ( .B1(n8482), .B2(n8537), .A(n8481), .ZN(n8488) );
  XNOR2_X1 U9961 ( .A(n8484), .B(n8483), .ZN(n8486) );
  AOI21_X1 U9962 ( .B1(n8486), .B2(n10369), .A(n8485), .ZN(n8606) );
  NOR2_X1 U9963 ( .A1(n8606), .A2(n10389), .ZN(n8487) );
  AOI211_X1 U9964 ( .C1(n8604), .C2(n8551), .A(n8488), .B(n8487), .ZN(n8489)
         );
  OAI21_X1 U9965 ( .B1(n8607), .B2(n8553), .A(n8489), .ZN(P2_U3275) );
  XNOR2_X1 U9966 ( .A(n8491), .B(n8490), .ZN(n8612) );
  AOI21_X1 U9967 ( .B1(n8608), .B2(n8519), .A(n8492), .ZN(n8609) );
  AOI22_X1 U9968 ( .A1(n8548), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8493), .B2(
        n10379), .ZN(n8494) );
  OAI21_X1 U9969 ( .B1(n8495), .B2(n8537), .A(n8494), .ZN(n8504) );
  AOI21_X1 U9970 ( .B1(n8497), .B2(n8496), .A(n8510), .ZN(n8502) );
  OAI22_X1 U9971 ( .A1(n8499), .A2(n8515), .B1(n8498), .B2(n8513), .ZN(n8500)
         );
  AOI21_X1 U9972 ( .B1(n8502), .B2(n8501), .A(n8500), .ZN(n8611) );
  NOR2_X1 U9973 ( .A1(n8611), .A2(n10389), .ZN(n8503) );
  AOI211_X1 U9974 ( .C1(n8609), .C2(n8551), .A(n8504), .B(n8503), .ZN(n8505)
         );
  OAI21_X1 U9975 ( .B1(n8612), .B2(n8553), .A(n8505), .ZN(P2_U3276) );
  XNOR2_X1 U9976 ( .A(n8506), .B(n8508), .ZN(n8615) );
  INV_X1 U9977 ( .A(n8615), .ZN(n8529) );
  NAND2_X1 U9978 ( .A1(n8539), .A2(n8507), .ZN(n8509) );
  NAND2_X1 U9979 ( .A1(n8509), .A2(n8508), .ZN(n8511) );
  AOI21_X1 U9980 ( .B1(n8512), .B2(n8511), .A(n8510), .ZN(n8518) );
  OAI22_X1 U9981 ( .A1(n8516), .A2(n8515), .B1(n8514), .B2(n8513), .ZN(n8517)
         );
  OR2_X1 U9982 ( .A1(n8518), .A2(n8517), .ZN(n8613) );
  INV_X1 U9983 ( .A(n8519), .ZN(n8520) );
  AOI211_X1 U9984 ( .C1(n8521), .C2(n8532), .A(n10462), .B(n8520), .ZN(n8614)
         );
  NAND2_X1 U9985 ( .A1(n8614), .A2(n8522), .ZN(n8526) );
  INV_X1 U9986 ( .A(n8523), .ZN(n8524) );
  AOI22_X1 U9987 ( .A1(n8548), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8524), .B2(
        n10379), .ZN(n8525) );
  OAI211_X1 U9988 ( .C1(n8673), .C2(n8537), .A(n8526), .B(n8525), .ZN(n8527)
         );
  AOI21_X1 U9989 ( .B1(n8613), .B2(n10376), .A(n8527), .ZN(n8528) );
  OAI21_X1 U9990 ( .B1(n8529), .B2(n8553), .A(n8528), .ZN(P2_U3277) );
  XNOR2_X1 U9991 ( .A(n8530), .B(n8540), .ZN(n8622) );
  INV_X1 U9992 ( .A(n8531), .ZN(n8534) );
  INV_X1 U9993 ( .A(n8532), .ZN(n8533) );
  AOI21_X1 U9994 ( .B1(n8618), .B2(n8534), .A(n8533), .ZN(n8619) );
  AOI22_X1 U9995 ( .A1(n10389), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8535), .B2(
        n10379), .ZN(n8536) );
  OAI21_X1 U9996 ( .B1(n8538), .B2(n8537), .A(n8536), .ZN(n8550) );
  OAI211_X1 U9997 ( .C1(n8541), .C2(n8540), .A(n8539), .B(n10369), .ZN(n8547)
         );
  AOI22_X1 U9998 ( .A1(n8545), .A2(n8544), .B1(n8543), .B2(n8542), .ZN(n8546)
         );
  NOR2_X1 U9999 ( .A1(n8621), .A2(n8548), .ZN(n8549) );
  AOI211_X1 U10000 ( .C1(n8619), .C2(n8551), .A(n8550), .B(n8549), .ZN(n8552)
         );
  OAI21_X1 U10001 ( .B1(n8622), .B2(n8553), .A(n8552), .ZN(P2_U3278) );
  MUX2_X1 U10002 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8649), .S(n10477), .Z(
        n8555) );
  AOI21_X1 U10003 ( .B1(n8556), .B2(n7922), .A(n8555), .ZN(n8557) );
  INV_X1 U10004 ( .A(n8557), .ZN(P2_U3551) );
  AND2_X1 U10005 ( .A1(n8559), .A2(n8558), .ZN(n8652) );
  INV_X1 U10006 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8560) );
  MUX2_X1 U10007 ( .A(n8652), .B(n8560), .S(n10475), .Z(n8561) );
  OAI21_X1 U10008 ( .B1(n7889), .B2(n8628), .A(n8561), .ZN(P2_U3550) );
  AOI22_X1 U10009 ( .A1(n8563), .A2(n10360), .B1(n8644), .B2(n8562), .ZN(n8564) );
  MUX2_X1 U10010 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8654), .S(n10477), .Z(
        P2_U3549) );
  AOI22_X1 U10011 ( .A1(n8568), .A2(n10360), .B1(n8644), .B2(n8567), .ZN(n8569) );
  OAI211_X1 U10012 ( .C1(n8571), .C2(n10432), .A(n8570), .B(n8569), .ZN(n8655)
         );
  MUX2_X1 U10013 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8655), .S(n10477), .Z(
        P2_U3548) );
  AOI22_X1 U10014 ( .A1(n8573), .A2(n10360), .B1(n8644), .B2(n8572), .ZN(n8574) );
  OAI211_X1 U10015 ( .C1(n8576), .C2(n10432), .A(n8575), .B(n8574), .ZN(n8656)
         );
  MUX2_X1 U10016 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8656), .S(n10477), .Z(
        P2_U3547) );
  INV_X1 U10017 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8580) );
  AOI211_X1 U10018 ( .C1(n8579), .C2(n10466), .A(n8578), .B(n8577), .ZN(n8657)
         );
  MUX2_X1 U10019 ( .A(n8580), .B(n8657), .S(n10477), .Z(n8581) );
  OAI21_X1 U10020 ( .B1(n8660), .B2(n8628), .A(n8581), .ZN(P2_U3546) );
  AOI21_X1 U10021 ( .B1(n8644), .B2(n8583), .A(n8582), .ZN(n8584) );
  OAI211_X1 U10022 ( .C1(n8586), .C2(n10432), .A(n8585), .B(n8584), .ZN(n8661)
         );
  MUX2_X1 U10023 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8661), .S(n10477), .Z(
        P2_U3545) );
  AOI22_X1 U10024 ( .A1(n8588), .A2(n10360), .B1(n8644), .B2(n8587), .ZN(n8589) );
  OAI211_X1 U10025 ( .C1(n8591), .C2(n10432), .A(n8590), .B(n8589), .ZN(n8662)
         );
  MUX2_X1 U10026 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8662), .S(n10477), .Z(
        P2_U3544) );
  NAND3_X1 U10027 ( .A1(n8592), .A2(n8451), .A3(n10466), .ZN(n8597) );
  AOI22_X1 U10028 ( .A1(n8594), .A2(n10360), .B1(n8644), .B2(n8593), .ZN(n8595) );
  NAND3_X1 U10029 ( .A1(n8597), .A2(n8596), .A3(n8595), .ZN(n8663) );
  MUX2_X1 U10030 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8663), .S(n10477), .Z(
        P2_U3543) );
  INV_X1 U10031 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8601) );
  AOI211_X1 U10032 ( .C1(n8600), .C2(n10466), .A(n8599), .B(n8598), .ZN(n8664)
         );
  MUX2_X1 U10033 ( .A(n8601), .B(n8664), .S(n10477), .Z(n8602) );
  OAI21_X1 U10034 ( .B1(n8667), .B2(n8628), .A(n8602), .ZN(P2_U3542) );
  AOI22_X1 U10035 ( .A1(n8604), .A2(n10360), .B1(n8644), .B2(n8603), .ZN(n8605) );
  OAI211_X1 U10036 ( .C1(n8607), .C2(n10432), .A(n8606), .B(n8605), .ZN(n8668)
         );
  MUX2_X1 U10037 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8668), .S(n10477), .Z(
        P2_U3541) );
  AOI22_X1 U10038 ( .A1(n8609), .A2(n10360), .B1(n8644), .B2(n8608), .ZN(n8610) );
  OAI211_X1 U10039 ( .C1(n8612), .C2(n10432), .A(n8611), .B(n8610), .ZN(n8669)
         );
  MUX2_X1 U10040 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8669), .S(n10477), .Z(
        P2_U3540) );
  AOI211_X1 U10041 ( .C1(n8615), .C2(n10466), .A(n8614), .B(n8613), .ZN(n8670)
         );
  MUX2_X1 U10042 ( .A(n8616), .B(n8670), .S(n10477), .Z(n8617) );
  OAI21_X1 U10043 ( .B1(n8673), .B2(n8628), .A(n8617), .ZN(P2_U3539) );
  AOI22_X1 U10044 ( .A1(n8619), .A2(n10360), .B1(n8644), .B2(n8618), .ZN(n8620) );
  OAI211_X1 U10045 ( .C1(n8622), .C2(n10432), .A(n8621), .B(n8620), .ZN(n8674)
         );
  MUX2_X1 U10046 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8674), .S(n10477), .Z(
        P2_U3538) );
  AOI211_X1 U10047 ( .C1(n8625), .C2(n10466), .A(n8624), .B(n8623), .ZN(n8675)
         );
  MUX2_X1 U10048 ( .A(n8626), .B(n8675), .S(n10477), .Z(n8627) );
  OAI21_X1 U10049 ( .B1(n6180), .B2(n8628), .A(n8627), .ZN(P2_U3537) );
  OAI22_X1 U10050 ( .A1(n8630), .A2(n10462), .B1(n8629), .B2(n10460), .ZN(
        n8631) );
  INV_X1 U10051 ( .A(n8631), .ZN(n8632) );
  OAI21_X1 U10052 ( .B1(n8634), .B2(n8633), .A(n8632), .ZN(n8635) );
  OR2_X1 U10053 ( .A1(n8636), .A2(n8635), .ZN(n8679) );
  MUX2_X1 U10054 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8679), .S(n10477), .Z(
        P2_U3536) );
  INV_X1 U10055 ( .A(n8637), .ZN(n8642) );
  AOI22_X1 U10056 ( .A1(n8639), .A2(n10360), .B1(n8644), .B2(n8638), .ZN(n8640) );
  OAI211_X1 U10057 ( .C1(n8642), .C2(n10432), .A(n8641), .B(n8640), .ZN(n8680)
         );
  MUX2_X1 U10058 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8680), .S(n10477), .Z(
        P2_U3535) );
  AOI22_X1 U10059 ( .A1(n8645), .A2(n10360), .B1(n8644), .B2(n8643), .ZN(n8646) );
  OAI211_X1 U10060 ( .C1(n8648), .C2(n10432), .A(n8647), .B(n8646), .ZN(n8681)
         );
  MUX2_X1 U10061 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8681), .S(n10477), .Z(
        P2_U3534) );
  INV_X1 U10062 ( .A(n8678), .ZN(n8650) );
  INV_X1 U10063 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8651) );
  MUX2_X1 U10064 ( .A(n8652), .B(n8651), .S(n10468), .Z(n8653) );
  OAI21_X1 U10065 ( .B1(n7889), .B2(n8678), .A(n8653), .ZN(P2_U3518) );
  MUX2_X1 U10066 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8654), .S(n10469), .Z(
        P2_U3517) );
  MUX2_X1 U10067 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8655), .S(n10469), .Z(
        P2_U3516) );
  MUX2_X1 U10068 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8656), .S(n10469), .Z(
        P2_U3515) );
  INV_X1 U10069 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8658) );
  MUX2_X1 U10070 ( .A(n8658), .B(n8657), .S(n10469), .Z(n8659) );
  OAI21_X1 U10071 ( .B1(n8660), .B2(n8678), .A(n8659), .ZN(P2_U3514) );
  MUX2_X1 U10072 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8661), .S(n10469), .Z(
        P2_U3513) );
  MUX2_X1 U10073 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8662), .S(n10469), .Z(
        P2_U3512) );
  MUX2_X1 U10074 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8663), .S(n10469), .Z(
        P2_U3511) );
  INV_X1 U10075 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8665) );
  MUX2_X1 U10076 ( .A(n8665), .B(n8664), .S(n10469), .Z(n8666) );
  OAI21_X1 U10077 ( .B1(n8667), .B2(n8678), .A(n8666), .ZN(P2_U3510) );
  MUX2_X1 U10078 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8668), .S(n10469), .Z(
        P2_U3509) );
  MUX2_X1 U10079 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8669), .S(n10469), .Z(
        P2_U3508) );
  INV_X1 U10080 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8671) );
  MUX2_X1 U10081 ( .A(n8671), .B(n8670), .S(n10469), .Z(n8672) );
  OAI21_X1 U10082 ( .B1(n8673), .B2(n8678), .A(n8672), .ZN(P2_U3507) );
  MUX2_X1 U10083 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8674), .S(n10469), .Z(
        P2_U3505) );
  INV_X1 U10084 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8676) );
  MUX2_X1 U10085 ( .A(n8676), .B(n8675), .S(n10469), .Z(n8677) );
  OAI21_X1 U10086 ( .B1(n6180), .B2(n8678), .A(n8677), .ZN(P2_U3502) );
  MUX2_X1 U10087 ( .A(n8679), .B(P2_REG0_REG_16__SCAN_IN), .S(n10468), .Z(
        P2_U3499) );
  MUX2_X1 U10088 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8680), .S(n10469), .Z(
        P2_U3496) );
  MUX2_X1 U10089 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8681), .S(n10469), .Z(
        P2_U3493) );
  INV_X1 U10090 ( .A(n8682), .ZN(n9558) );
  NOR4_X1 U10091 ( .A1(n5916), .A2(P2_IR_REG_30__SCAN_IN), .A3(n5917), .A4(
        P2_U3152), .ZN(n8683) );
  AOI21_X1 U10092 ( .B1(n8684), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8683), .ZN(
        n8685) );
  OAI21_X1 U10093 ( .B1(n9558), .B2(n8686), .A(n8685), .ZN(P2_U3327) );
  INV_X1 U10094 ( .A(n8687), .ZN(n8688) );
  MUX2_X1 U10095 ( .A(n8688), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10096 ( .A(n8690), .B(n8689), .ZN(n8691) );
  XNOR2_X1 U10097 ( .A(n8692), .B(n8691), .ZN(n8693) );
  NAND2_X1 U10098 ( .A1(n8693), .A2(n8812), .ZN(n8700) );
  AOI21_X1 U10099 ( .B1(n8817), .B2(n9136), .A(n8694), .ZN(n8699) );
  AOI22_X1 U10100 ( .A1(n8808), .A2(n10204), .B1(n8791), .B2(n8695), .ZN(n8698) );
  OR2_X1 U10101 ( .A1(n8804), .A2(n8696), .ZN(n8697) );
  NAND4_X1 U10102 ( .A1(n8700), .A2(n8699), .A3(n8698), .A4(n8697), .ZN(
        P1_U3211) );
  XNOR2_X1 U10103 ( .A(n8702), .B(n8701), .ZN(n8703) );
  XNOR2_X1 U10104 ( .A(n8704), .B(n8703), .ZN(n8710) );
  OAI22_X1 U10105 ( .A1(n8819), .A2(n9317), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8705), .ZN(n8706) );
  AOI21_X1 U10106 ( .B1(n8817), .B2(n9248), .A(n8706), .ZN(n8707) );
  OAI21_X1 U10107 ( .B1(n8804), .B2(n9282), .A(n8707), .ZN(n8708) );
  AOI21_X1 U10108 ( .B1(n9450), .B2(n8791), .A(n8708), .ZN(n8709) );
  OAI21_X1 U10109 ( .B1(n8710), .B2(n8773), .A(n8709), .ZN(P1_U3212) );
  NOR2_X1 U10110 ( .A1(n8711), .A2(n4521), .ZN(n8713) );
  XNOR2_X1 U10111 ( .A(n8713), .B(n8712), .ZN(n8718) );
  NOR2_X1 U10112 ( .A1(n8804), .A2(n9342), .ZN(n8716) );
  AOI22_X1 U10113 ( .A1(n8817), .A2(n9349), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8714) );
  OAI21_X1 U10114 ( .B1(n9371), .B2(n8819), .A(n8714), .ZN(n8715) );
  AOI211_X1 U10115 ( .C1(n9469), .C2(n8791), .A(n8716), .B(n8715), .ZN(n8717)
         );
  OAI21_X1 U10116 ( .B1(n8718), .B2(n8773), .A(n8717), .ZN(P1_U3214) );
  INV_X1 U10117 ( .A(n8719), .ZN(n8800) );
  NAND2_X1 U10118 ( .A1(n8721), .A2(n8720), .ZN(n8798) );
  NOR2_X1 U10119 ( .A1(n8721), .A2(n8720), .ZN(n8797) );
  AOI21_X1 U10120 ( .B1(n8800), .B2(n8798), .A(n8797), .ZN(n8725) );
  NAND2_X1 U10121 ( .A1(n8723), .A2(n8722), .ZN(n8724) );
  XNOR2_X1 U10122 ( .A(n8725), .B(n8724), .ZN(n8730) );
  NOR2_X1 U10123 ( .A1(n8804), .A2(n9401), .ZN(n8728) );
  NAND2_X1 U10124 ( .A1(n8817), .A2(n9206), .ZN(n8726) );
  NAND2_X1 U10125 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9165) );
  OAI211_X1 U10126 ( .C1(n9411), .C2(n8819), .A(n8726), .B(n9165), .ZN(n8727)
         );
  AOI211_X1 U10127 ( .C1(n9491), .C2(n8791), .A(n8728), .B(n8727), .ZN(n8729)
         );
  OAI21_X1 U10128 ( .B1(n8730), .B2(n8773), .A(n8729), .ZN(P1_U3217) );
  XOR2_X1 U10129 ( .A(n8732), .B(n8731), .Z(n8737) );
  NOR2_X1 U10130 ( .A1(n8804), .A2(n9373), .ZN(n8735) );
  INV_X1 U10131 ( .A(n9206), .ZN(n9410) );
  INV_X1 U10132 ( .A(n9371), .ZN(n9348) );
  AOI22_X1 U10133 ( .A1(n8817), .A2(n9348), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8733) );
  OAI21_X1 U10134 ( .B1(n9410), .B2(n8819), .A(n8733), .ZN(n8734) );
  AOI211_X1 U10135 ( .C1(n9481), .C2(n8791), .A(n8735), .B(n8734), .ZN(n8736)
         );
  OAI21_X1 U10136 ( .B1(n8737), .B2(n8773), .A(n8736), .ZN(P1_U3221) );
  XOR2_X1 U10137 ( .A(n8739), .B(n8738), .Z(n8744) );
  AND2_X1 U10138 ( .A1(n9305), .A2(n9524), .ZN(n9460) );
  NOR2_X1 U10139 ( .A1(n8804), .A2(n9307), .ZN(n8742) );
  INV_X1 U10140 ( .A(n9349), .ZN(n9316) );
  AOI22_X1 U10141 ( .A1(n8817), .A2(n9220), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8740) );
  OAI21_X1 U10142 ( .B1(n9316), .B2(n8819), .A(n8740), .ZN(n8741) );
  AOI211_X1 U10143 ( .C1(n9460), .C2(n8795), .A(n8742), .B(n8741), .ZN(n8743)
         );
  OAI21_X1 U10144 ( .B1(n8744), .B2(n8773), .A(n8743), .ZN(P1_U3223) );
  OAI21_X1 U10145 ( .B1(n8747), .B2(n8746), .A(n8745), .ZN(n8748) );
  NAND2_X1 U10146 ( .A1(n8748), .A2(n8812), .ZN(n8752) );
  NOR2_X1 U10147 ( .A1(n8804), .A2(n9415), .ZN(n8750) );
  NAND2_X1 U10148 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10142)
         );
  OAI21_X1 U10149 ( .B1(n8805), .B2(n9411), .A(n10142), .ZN(n8749) );
  AOI211_X1 U10150 ( .C1(n8808), .C2(n9421), .A(n8750), .B(n8749), .ZN(n8751)
         );
  OAI211_X1 U10151 ( .C1(n9418), .C2(n8824), .A(n8752), .B(n8751), .ZN(
        P1_U3226) );
  OAI21_X1 U10152 ( .B1(n8755), .B2(n8754), .A(n8753), .ZN(n8756) );
  NAND2_X1 U10153 ( .A1(n8756), .A2(n8812), .ZN(n8762) );
  INV_X1 U10154 ( .A(n9330), .ZN(n9335) );
  NOR2_X1 U10155 ( .A1(n9335), .A2(n10304), .ZN(n9464) );
  INV_X1 U10156 ( .A(n9218), .ZN(n9327) );
  AOI22_X1 U10157 ( .A1(n8817), .A2(n9327), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8759) );
  INV_X1 U10158 ( .A(n8757), .ZN(n9331) );
  NAND2_X1 U10159 ( .A1(n8821), .A2(n9331), .ZN(n8758) );
  OAI211_X1 U10160 ( .C1(n8836), .C2(n8819), .A(n8759), .B(n8758), .ZN(n8760)
         );
  AOI21_X1 U10161 ( .B1(n9464), .B2(n8795), .A(n8760), .ZN(n8761) );
  NAND2_X1 U10162 ( .A1(n8762), .A2(n8761), .ZN(P1_U3227) );
  INV_X1 U10163 ( .A(n8763), .ZN(n8768) );
  AOI21_X1 U10164 ( .B1(n8765), .B2(n8767), .A(n8764), .ZN(n8766) );
  AOI21_X1 U10165 ( .B1(n8768), .B2(n8767), .A(n8766), .ZN(n8774) );
  NOR2_X1 U10166 ( .A1(n8804), .A2(n9388), .ZN(n8771) );
  INV_X1 U10167 ( .A(n9203), .ZN(n9384) );
  AOI22_X1 U10168 ( .A1(n8817), .A2(n9361), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8769) );
  OAI21_X1 U10169 ( .B1(n9384), .B2(n8819), .A(n8769), .ZN(n8770) );
  AOI211_X1 U10170 ( .C1(n9486), .C2(n8791), .A(n8771), .B(n8770), .ZN(n8772)
         );
  OAI21_X1 U10171 ( .B1(n8774), .B2(n8773), .A(n8772), .ZN(P1_U3231) );
  INV_X1 U10172 ( .A(n8778), .ZN(n8775) );
  NOR2_X1 U10173 ( .A1(n8776), .A2(n8775), .ZN(n8781) );
  AOI21_X1 U10174 ( .B1(n8779), .B2(n8778), .A(n8777), .ZN(n8780) );
  OAI21_X1 U10175 ( .B1(n8781), .B2(n8780), .A(n8812), .ZN(n8785) );
  AOI22_X1 U10176 ( .A1(n8817), .A2(n9362), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8782) );
  OAI21_X1 U10177 ( .B1(n9385), .B2(n8819), .A(n8782), .ZN(n8783) );
  AOI21_X1 U10178 ( .B1(n9356), .B2(n8821), .A(n8783), .ZN(n8784) );
  OAI211_X1 U10179 ( .C1(n9358), .C2(n8824), .A(n8785), .B(n8784), .ZN(
        P1_U3233) );
  OAI21_X1 U10180 ( .B1(n8788), .B2(n8787), .A(n8786), .ZN(n8789) );
  NAND2_X1 U10181 ( .A1(n8789), .A2(n8812), .ZN(n8794) );
  AOI22_X1 U10182 ( .A1(n8808), .A2(n6920), .B1(n8817), .B2(n10225), .ZN(n8793) );
  AOI22_X1 U10183 ( .A1(n8791), .A2(n7018), .B1(n8790), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n8792) );
  NAND3_X1 U10184 ( .A1(n8794), .A2(n8793), .A3(n8792), .ZN(P1_U3235) );
  INV_X1 U10185 ( .A(n8795), .ZN(n8811) );
  NAND2_X1 U10186 ( .A1(n8796), .A2(n9524), .ZN(n9497) );
  INV_X1 U10187 ( .A(n8797), .ZN(n8799) );
  NAND2_X1 U10188 ( .A1(n8799), .A2(n8798), .ZN(n8801) );
  XNOR2_X1 U10189 ( .A(n8801), .B(n8800), .ZN(n8802) );
  NAND2_X1 U10190 ( .A1(n8802), .A2(n8812), .ZN(n8810) );
  NOR2_X1 U10191 ( .A1(n8804), .A2(n8803), .ZN(n8807) );
  NAND2_X1 U10192 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10160)
         );
  OAI21_X1 U10193 ( .B1(n8805), .B2(n9384), .A(n10160), .ZN(n8806) );
  AOI211_X1 U10194 ( .C1(n8808), .C2(n9130), .A(n8807), .B(n8806), .ZN(n8809)
         );
  OAI211_X1 U10195 ( .C1(n8811), .C2(n9497), .A(n8810), .B(n8809), .ZN(
        P1_U3236) );
  OAI211_X1 U10196 ( .C1(n8815), .C2(n8814), .A(n8813), .B(n8812), .ZN(n8823)
         );
  INV_X1 U10197 ( .A(n8816), .ZN(n9291) );
  INV_X1 U10198 ( .A(n9259), .ZN(n9298) );
  AOI22_X1 U10199 ( .A1(n8817), .A2(n9298), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8818) );
  OAI21_X1 U10200 ( .B1(n9218), .B2(n8819), .A(n8818), .ZN(n8820) );
  AOI21_X1 U10201 ( .B1(n9291), .B2(n8821), .A(n8820), .ZN(n8822) );
  OAI211_X1 U10202 ( .C1(n9293), .C2(n8824), .A(n8823), .B(n8822), .ZN(
        P1_U3238) );
  NAND2_X1 U10203 ( .A1(n8825), .A2(n8866), .ZN(n8827) );
  OR2_X1 U10204 ( .A1(n4485), .A2(n9737), .ZN(n8826) );
  INV_X1 U10205 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8831) );
  NAND2_X1 U10206 ( .A1(n8828), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8830) );
  NAND2_X1 U10207 ( .A1(n5325), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8829) );
  OAI211_X1 U10208 ( .C1(n8832), .C2(n8831), .A(n8830), .B(n8829), .ZN(n9247)
         );
  INV_X1 U10209 ( .A(n9247), .ZN(n8870) );
  OR2_X1 U10210 ( .A1(n9197), .A2(n8870), .ZN(n9111) );
  INV_X1 U10211 ( .A(n9111), .ZN(n8864) );
  NAND2_X1 U10212 ( .A1(n9444), .A2(n9275), .ZN(n9048) );
  NAND2_X1 U10213 ( .A1(n8833), .A2(n8866), .ZN(n8835) );
  OR2_X1 U10214 ( .A1(n4485), .A2(n9718), .ZN(n8834) );
  NAND2_X1 U10215 ( .A1(n9251), .A2(n9258), .ZN(n8928) );
  NAND2_X1 U10216 ( .A1(n9450), .A2(n9259), .ZN(n9044) );
  NAND2_X1 U10217 ( .A1(n9305), .A2(n9218), .ZN(n9030) );
  NAND2_X1 U10218 ( .A1(n9469), .A2(n8836), .ZN(n9104) );
  NAND2_X1 U10219 ( .A1(n9237), .A2(n9104), .ZN(n9347) );
  INV_X1 U10220 ( .A(n9347), .ZN(n8860) );
  NAND2_X1 U10221 ( .A1(n9481), .A2(n9385), .ZN(n9013) );
  NAND2_X1 U10222 ( .A1(n8879), .A2(n9013), .ZN(n9368) );
  INV_X1 U10223 ( .A(n9368), .ZN(n9234) );
  NAND2_X1 U10224 ( .A1(n9474), .A2(n9371), .ZN(n9235) );
  INV_X1 U10225 ( .A(n9235), .ZN(n8837) );
  NOR2_X1 U10226 ( .A1(n9236), .A2(n8837), .ZN(n9359) );
  INV_X1 U10227 ( .A(n9486), .ZN(n9392) );
  NAND2_X1 U10228 ( .A1(n9486), .A2(n9410), .ZN(n9232) );
  INV_X1 U10229 ( .A(n9232), .ZN(n8878) );
  OR2_X1 U10230 ( .A1(n9491), .A2(n9384), .ZN(n9008) );
  NAND2_X1 U10231 ( .A1(n9491), .A2(n9384), .ZN(n9011) );
  NAND2_X1 U10232 ( .A1(n9008), .A2(n9011), .ZN(n9407) );
  NOR2_X1 U10233 ( .A1(n10178), .A2(n10229), .ZN(n8840) );
  NAND4_X1 U10234 ( .A1(n8841), .A2(n8840), .A3(n8839), .A4(n8838), .ZN(n8844)
         );
  NAND2_X1 U10235 ( .A1(n7023), .A2(n10208), .ZN(n8842) );
  NOR3_X1 U10236 ( .A1(n8844), .A2(n8843), .A3(n8842), .ZN(n8849) );
  INV_X1 U10237 ( .A(n8845), .ZN(n8847) );
  AND4_X1 U10238 ( .A1(n8849), .A2(n8848), .A3(n8847), .A4(n8846), .ZN(n8851)
         );
  NAND4_X1 U10239 ( .A1(n8851), .A2(n8850), .A3(n10012), .A4(n8971), .ZN(n8852) );
  NOR3_X1 U10240 ( .A1(n8985), .A2(n8853), .A3(n8852), .ZN(n8854) );
  NAND3_X1 U10241 ( .A1(n9419), .A2(n8855), .A3(n8854), .ZN(n8857) );
  OR3_X1 U10242 ( .A1(n9407), .A2(n8857), .A3(n8856), .ZN(n8858) );
  NOR2_X1 U10243 ( .A1(n9381), .A2(n8858), .ZN(n8859) );
  NAND4_X1 U10244 ( .A1(n8860), .A2(n9234), .A3(n9359), .A4(n8859), .ZN(n8861)
         );
  OR2_X1 U10245 ( .A1(n9330), .A2(n9316), .ZN(n9020) );
  NAND2_X1 U10246 ( .A1(n9330), .A2(n9316), .ZN(n9311) );
  NAND2_X1 U10247 ( .A1(n9020), .A2(n9311), .ZN(n9322) );
  NOR2_X1 U10248 ( .A1(n8861), .A2(n9322), .ZN(n8862) );
  XNOR2_X1 U10249 ( .A(n9454), .B(n9220), .ZN(n9296) );
  NAND4_X1 U10250 ( .A1(n9222), .A2(n9313), .A3(n8862), .A4(n9296), .ZN(n8863)
         );
  NOR4_X1 U10251 ( .A1(n8864), .A2(n9267), .A3(n9244), .A4(n8863), .ZN(n8869)
         );
  NOR2_X1 U10252 ( .A1(n4484), .A2(n6563), .ZN(n8865) );
  INV_X1 U10253 ( .A(n9431), .ZN(n8868) );
  INV_X1 U10254 ( .A(n9194), .ZN(n8867) );
  NAND2_X1 U10255 ( .A1(n8868), .A2(n8867), .ZN(n9114) );
  NAND2_X1 U10256 ( .A1(n8869), .A2(n9114), .ZN(n8873) );
  AND2_X1 U10257 ( .A1(n9431), .A2(n9194), .ZN(n9071) );
  INV_X1 U10258 ( .A(n9071), .ZN(n8872) );
  NAND2_X1 U10259 ( .A1(n9197), .A2(n8870), .ZN(n8871) );
  NAND2_X1 U10260 ( .A1(n8872), .A2(n8871), .ZN(n9113) );
  OAI21_X1 U10261 ( .B1(n8873), .B2(n9113), .A(n9076), .ZN(n9066) );
  INV_X1 U10262 ( .A(n9066), .ZN(n8933) );
  AOI21_X1 U10263 ( .B1(n9194), .B2(n9111), .A(n9431), .ZN(n9051) );
  INV_X1 U10264 ( .A(n9051), .ZN(n9055) );
  AND2_X1 U10265 ( .A1(n9009), .A2(n8874), .ZN(n9227) );
  AND2_X1 U10266 ( .A1(n9011), .A2(n9226), .ZN(n8999) );
  INV_X1 U10267 ( .A(n8999), .ZN(n8877) );
  INV_X1 U10268 ( .A(n8879), .ZN(n8875) );
  OR2_X1 U10269 ( .A1(n9236), .A2(n8875), .ZN(n9015) );
  INV_X1 U10270 ( .A(n9015), .ZN(n9000) );
  INV_X1 U10271 ( .A(n9008), .ZN(n8876) );
  NOR2_X1 U10272 ( .A1(n9231), .A2(n8876), .ZN(n9001) );
  OAI211_X1 U10273 ( .C1(n9227), .C2(n8877), .A(n9000), .B(n9001), .ZN(n8882)
         );
  NAND2_X1 U10274 ( .A1(n8879), .A2(n8878), .ZN(n8880) );
  AND2_X1 U10275 ( .A1(n8880), .A2(n9013), .ZN(n8881) );
  AND2_X1 U10276 ( .A1(n8881), .A2(n9235), .ZN(n8917) );
  OR2_X1 U10277 ( .A1(n8917), .A2(n9236), .ZN(n9003) );
  AND2_X1 U10278 ( .A1(n8882), .A2(n9003), .ZN(n9075) );
  NAND2_X1 U10279 ( .A1(n9226), .A2(n8883), .ZN(n9229) );
  INV_X1 U10280 ( .A(n8884), .ZN(n8951) );
  NAND2_X1 U10281 ( .A1(n8950), .A2(n8949), .ZN(n8885) );
  NAND2_X1 U10282 ( .A1(n8885), .A2(n8953), .ZN(n8886) );
  AND3_X1 U10283 ( .A1(n8961), .A2(n8960), .A3(n8886), .ZN(n8887) );
  NAND2_X1 U10284 ( .A1(n8965), .A2(n8887), .ZN(n8912) );
  INV_X1 U10285 ( .A(n8912), .ZN(n8888) );
  OAI21_X1 U10286 ( .B1(n8889), .B2(n8951), .A(n8888), .ZN(n8896) );
  INV_X1 U10287 ( .A(n8890), .ZN(n8891) );
  NAND2_X1 U10288 ( .A1(n8962), .A2(n8891), .ZN(n8892) );
  NAND2_X1 U10289 ( .A1(n8892), .A2(n8961), .ZN(n8893) );
  NAND2_X1 U10290 ( .A1(n8894), .A2(n8893), .ZN(n8959) );
  NAND2_X1 U10291 ( .A1(n8959), .A2(n8965), .ZN(n8895) );
  AND3_X1 U10292 ( .A1(n8896), .A2(n8969), .A3(n8895), .ZN(n8899) );
  NAND2_X1 U10293 ( .A1(n8897), .A2(n8976), .ZN(n8967) );
  NAND2_X1 U10294 ( .A1(n8898), .A2(n8967), .ZN(n8915) );
  OAI211_X1 U10295 ( .C1(n8899), .C2(n8915), .A(n7708), .B(n8992), .ZN(n8900)
         );
  NAND2_X1 U10296 ( .A1(n8900), .A2(n8993), .ZN(n8901) );
  NOR2_X1 U10297 ( .A1(n9229), .A2(n8901), .ZN(n9094) );
  INV_X1 U10298 ( .A(n7221), .ZN(n8911) );
  AND2_X1 U10299 ( .A1(n10227), .A2(n8902), .ZN(n8903) );
  NAND2_X1 U10300 ( .A1(n9088), .A2(n8903), .ZN(n9085) );
  INV_X1 U10301 ( .A(n8904), .ZN(n8905) );
  AND2_X1 U10302 ( .A1(n8905), .A2(n10227), .ZN(n10175) );
  INV_X1 U10303 ( .A(n10175), .ZN(n8906) );
  AOI21_X1 U10304 ( .B1(n8907), .B2(n9083), .A(n8906), .ZN(n8909) );
  OAI21_X1 U10305 ( .B1(n8909), .B2(n9089), .A(n8908), .ZN(n8910) );
  OAI21_X1 U10306 ( .B1(n8911), .B2(n9085), .A(n8910), .ZN(n8934) );
  INV_X1 U10307 ( .A(n8940), .ZN(n8914) );
  INV_X1 U10308 ( .A(n8936), .ZN(n8913) );
  OR4_X1 U10309 ( .A1(n8915), .A2(n8914), .A3(n8913), .A4(n8912), .ZN(n8916)
         );
  OR3_X1 U10310 ( .A1(n9229), .A2(n4826), .A3(n8916), .ZN(n9097) );
  AOI21_X1 U10311 ( .B1(n8935), .B2(n8934), .A(n9097), .ZN(n8919) );
  INV_X1 U10312 ( .A(n8917), .ZN(n8918) );
  INV_X1 U10313 ( .A(n9011), .ZN(n9230) );
  NOR2_X1 U10314 ( .A1(n8918), .A2(n9230), .ZN(n9099) );
  OAI21_X1 U10315 ( .B1(n9094), .B2(n8919), .A(n9099), .ZN(n8920) );
  INV_X1 U10316 ( .A(n8920), .ZN(n8921) );
  OAI21_X1 U10317 ( .B1(n9075), .B2(n8921), .A(n9104), .ZN(n8922) );
  AND2_X1 U10318 ( .A1(n9020), .A2(n9237), .ZN(n9102) );
  NAND2_X1 U10319 ( .A1(n9030), .A2(n9311), .ZN(n9238) );
  AOI21_X1 U10320 ( .B1(n8922), .B2(n9102), .A(n9238), .ZN(n8930) );
  NAND2_X1 U10321 ( .A1(n9058), .A2(n9242), .ZN(n8927) );
  INV_X1 U10322 ( .A(n9043), .ZN(n9241) );
  OR2_X1 U10323 ( .A1(n9454), .A2(n9317), .ZN(n8923) );
  NAND2_X1 U10324 ( .A1(n8923), .A2(n9031), .ZN(n9240) );
  OR3_X1 U10325 ( .A1(n8927), .A2(n9241), .A3(n9240), .ZN(n9108) );
  NAND2_X1 U10326 ( .A1(n9247), .A2(n9194), .ZN(n8924) );
  AND2_X1 U10327 ( .A1(n9197), .A2(n8924), .ZN(n9059) );
  INV_X1 U10328 ( .A(n9059), .ZN(n9057) );
  NAND2_X1 U10329 ( .A1(n9454), .A2(n9317), .ZN(n9239) );
  OAI211_X1 U10330 ( .C1(n9241), .C2(n9239), .A(n9048), .B(n9044), .ZN(n8925)
         );
  INV_X1 U10331 ( .A(n8925), .ZN(n8926) );
  OR2_X1 U10332 ( .A1(n8927), .A2(n8926), .ZN(n8929) );
  AND2_X1 U10333 ( .A1(n8929), .A2(n8928), .ZN(n9107) );
  OAI211_X1 U10334 ( .C1(n8930), .C2(n9108), .A(n9057), .B(n9107), .ZN(n8931)
         );
  AOI211_X1 U10335 ( .C1(n9055), .C2(n8931), .A(n9076), .B(n9071), .ZN(n8932)
         );
  NOR2_X1 U10336 ( .A1(n8933), .A2(n8932), .ZN(n9069) );
  INV_X1 U10337 ( .A(n8934), .ZN(n8937) );
  INV_X1 U10338 ( .A(n8935), .ZN(n9091) );
  AOI21_X1 U10339 ( .B1(n8937), .B2(n8936), .A(n9091), .ZN(n8939) );
  AND2_X1 U10340 ( .A1(n8938), .A2(n10206), .ZN(n9438) );
  MUX2_X1 U10341 ( .A(n7232), .B(n8939), .S(n9438), .Z(n8947) );
  NAND2_X1 U10342 ( .A1(n8940), .A2(n8949), .ZN(n8948) );
  INV_X1 U10343 ( .A(n8948), .ZN(n8941) );
  OAI21_X1 U10344 ( .B1(n8947), .B2(n8942), .A(n8941), .ZN(n8946) );
  AND2_X1 U10345 ( .A1(n8953), .A2(n8943), .ZN(n8945) );
  NAND2_X1 U10346 ( .A1(n8961), .A2(n8950), .ZN(n8944) );
  AOI21_X1 U10347 ( .B1(n8946), .B2(n8945), .A(n8944), .ZN(n8958) );
  INV_X1 U10348 ( .A(n8947), .ZN(n8956) );
  NOR2_X1 U10349 ( .A1(n4639), .A2(n8948), .ZN(n8955) );
  NAND3_X1 U10350 ( .A1(n8951), .A2(n8950), .A3(n8949), .ZN(n8952) );
  NAND3_X1 U10351 ( .A1(n8962), .A2(n8953), .A3(n8952), .ZN(n8954) );
  AOI21_X1 U10352 ( .B1(n8956), .B2(n8955), .A(n8954), .ZN(n8957) );
  MUX2_X1 U10353 ( .A(n8958), .B(n8957), .S(n9438), .Z(n8972) );
  INV_X1 U10354 ( .A(n9438), .ZN(n9064) );
  NAND2_X1 U10355 ( .A1(n8959), .A2(n9064), .ZN(n8968) );
  NAND2_X1 U10356 ( .A1(n8961), .A2(n8960), .ZN(n8963) );
  NAND3_X1 U10357 ( .A1(n8963), .A2(n9438), .A3(n8962), .ZN(n8964) );
  AND2_X1 U10358 ( .A1(n8965), .A2(n8964), .ZN(n8966) );
  NAND4_X1 U10359 ( .A1(n8969), .A2(n8968), .A3(n8967), .A4(n8966), .ZN(n8970)
         );
  AOI21_X1 U10360 ( .B1(n8972), .B2(n8971), .A(n8970), .ZN(n8991) );
  NOR2_X1 U10361 ( .A1(n10013), .A2(n9438), .ZN(n8977) );
  NOR2_X1 U10362 ( .A1(n9132), .A2(n9438), .ZN(n8973) );
  AOI21_X1 U10363 ( .B1(n9516), .B2(n8977), .A(n8973), .ZN(n8983) );
  NAND2_X1 U10364 ( .A1(n10013), .A2(n9438), .ZN(n8975) );
  OAI22_X1 U10365 ( .A1(n9516), .A2(n8975), .B1(n8976), .B2(n9064), .ZN(n8974)
         );
  NAND2_X1 U10366 ( .A1(n10029), .A2(n8974), .ZN(n8982) );
  NOR2_X1 U10367 ( .A1(n8976), .A2(n8975), .ZN(n8980) );
  NAND2_X1 U10368 ( .A1(n8977), .A2(n8976), .ZN(n8978) );
  NAND2_X1 U10369 ( .A1(n9516), .A2(n8978), .ZN(n8979) );
  OAI21_X1 U10370 ( .B1(n9516), .B2(n8980), .A(n8979), .ZN(n8981) );
  OAI211_X1 U10371 ( .C1(n10029), .C2(n8983), .A(n8982), .B(n8981), .ZN(n8984)
         );
  OR2_X1 U10372 ( .A1(n8985), .A2(n8984), .ZN(n8990) );
  MUX2_X1 U10373 ( .A(n7707), .B(n8986), .S(n9064), .Z(n8987) );
  NOR2_X1 U10374 ( .A1(n8988), .A2(n8987), .ZN(n8989) );
  OAI21_X1 U10375 ( .B1(n8991), .B2(n8990), .A(n8989), .ZN(n8995) );
  MUX2_X1 U10376 ( .A(n8993), .B(n8992), .S(n9438), .Z(n8994) );
  NAND3_X1 U10377 ( .A1(n8995), .A2(n9419), .A3(n8994), .ZN(n8998) );
  INV_X1 U10378 ( .A(n9229), .ZN(n8996) );
  MUX2_X1 U10379 ( .A(n9227), .B(n8996), .S(n9438), .Z(n8997) );
  NAND2_X1 U10380 ( .A1(n8998), .A2(n8997), .ZN(n9010) );
  NAND2_X1 U10381 ( .A1(n9010), .A2(n8999), .ZN(n9002) );
  NAND3_X1 U10382 ( .A1(n9002), .A2(n9001), .A3(n9000), .ZN(n9004) );
  NAND3_X1 U10383 ( .A1(n9004), .A2(n9104), .A3(n9003), .ZN(n9005) );
  NAND2_X1 U10384 ( .A1(n9005), .A2(n9237), .ZN(n9006) );
  OR2_X1 U10385 ( .A1(n9330), .A2(n9349), .ZN(n9215) );
  NAND2_X1 U10386 ( .A1(n9330), .A2(n9349), .ZN(n9216) );
  NAND2_X1 U10387 ( .A1(n9215), .A2(n9216), .ZN(n9017) );
  NAND2_X1 U10388 ( .A1(n9006), .A2(n9017), .ZN(n9007) );
  NAND3_X1 U10389 ( .A1(n9007), .A2(n9031), .A3(n9020), .ZN(n9025) );
  NAND3_X1 U10390 ( .A1(n9010), .A2(n9009), .A3(n9008), .ZN(n9012) );
  NAND3_X1 U10391 ( .A1(n9012), .A2(n9232), .A3(n9011), .ZN(n9014) );
  INV_X1 U10392 ( .A(n9013), .ZN(n9233) );
  AOI21_X1 U10393 ( .B1(n9014), .B2(n4662), .A(n9233), .ZN(n9016) );
  OAI21_X1 U10394 ( .B1(n9016), .B2(n9015), .A(n9235), .ZN(n9018) );
  NAND3_X1 U10395 ( .A1(n9018), .A2(n9237), .A3(n9017), .ZN(n9023) );
  INV_X1 U10396 ( .A(n9238), .ZN(n9022) );
  INV_X1 U10397 ( .A(n9104), .ZN(n9019) );
  NAND2_X1 U10398 ( .A1(n9020), .A2(n9019), .ZN(n9021) );
  NAND3_X1 U10399 ( .A1(n9023), .A2(n9022), .A3(n9021), .ZN(n9024) );
  MUX2_X1 U10400 ( .A(n9025), .B(n9024), .S(n9438), .Z(n9035) );
  NAND2_X1 U10401 ( .A1(n9030), .A2(n9220), .ZN(n9026) );
  NAND2_X1 U10402 ( .A1(n9043), .A2(n9026), .ZN(n9028) );
  INV_X1 U10403 ( .A(n9031), .ZN(n9294) );
  OAI21_X1 U10404 ( .B1(n9293), .B2(n9294), .A(n9044), .ZN(n9027) );
  MUX2_X1 U10405 ( .A(n9028), .B(n9027), .S(n9438), .Z(n9029) );
  OAI21_X1 U10406 ( .B1(n9035), .B2(n9274), .A(n9029), .ZN(n9042) );
  NAND2_X1 U10407 ( .A1(n9030), .A2(n9064), .ZN(n9033) );
  NOR2_X1 U10408 ( .A1(n9220), .A2(n9064), .ZN(n9036) );
  NAND2_X1 U10409 ( .A1(n9031), .A2(n9036), .ZN(n9032) );
  OAI21_X1 U10410 ( .B1(n9454), .B2(n9033), .A(n9032), .ZN(n9034) );
  NAND2_X1 U10411 ( .A1(n9035), .A2(n9034), .ZN(n9041) );
  AND2_X1 U10412 ( .A1(n9220), .A2(n9064), .ZN(n9039) );
  INV_X1 U10413 ( .A(n9036), .ZN(n9037) );
  NAND2_X1 U10414 ( .A1(n9454), .A2(n9037), .ZN(n9038) );
  OAI21_X1 U10415 ( .B1(n9454), .B2(n9039), .A(n9038), .ZN(n9040) );
  NAND3_X1 U10416 ( .A1(n9042), .A2(n9041), .A3(n9040), .ZN(n9047) );
  INV_X1 U10417 ( .A(n9267), .ZN(n9046) );
  MUX2_X1 U10418 ( .A(n9044), .B(n9043), .S(n9438), .Z(n9045) );
  NAND3_X1 U10419 ( .A1(n9047), .A2(n9046), .A3(n9045), .ZN(n9050) );
  MUX2_X1 U10420 ( .A(n9048), .B(n9242), .S(n9064), .Z(n9049) );
  NAND2_X1 U10421 ( .A1(n9050), .A2(n9049), .ZN(n9054) );
  NOR2_X1 U10422 ( .A1(n9054), .A2(n9258), .ZN(n9052) );
  AOI21_X1 U10423 ( .B1(n9052), .B2(n9057), .A(n9051), .ZN(n9065) );
  INV_X1 U10424 ( .A(n9054), .ZN(n9053) );
  INV_X1 U10425 ( .A(n9251), .ZN(n9440) );
  AOI211_X1 U10426 ( .C1(n9054), .C2(n9129), .A(n9438), .B(n9440), .ZN(n9056)
         );
  OAI21_X1 U10427 ( .B1(n5064), .B2(n9056), .A(n9055), .ZN(n9063) );
  NOR2_X1 U10428 ( .A1(n9057), .A2(n9438), .ZN(n9061) );
  NOR3_X1 U10429 ( .A1(n9059), .A2(n9058), .A3(n9064), .ZN(n9060) );
  AOI211_X1 U10430 ( .C1(n9061), .C2(n9114), .A(n9071), .B(n9060), .ZN(n9062)
         );
  OAI211_X1 U10431 ( .C1(n9065), .C2(n9064), .A(n9063), .B(n9062), .ZN(n9070)
         );
  OAI21_X1 U10432 ( .B1(n9070), .B2(n9067), .A(n9066), .ZN(n9068) );
  MUX2_X1 U10433 ( .A(n9069), .B(n9068), .S(n10206), .Z(n9074) );
  INV_X1 U10434 ( .A(n9070), .ZN(n9072) );
  NOR4_X1 U10435 ( .A1(n9072), .A2(n9125), .A3(n9071), .A4(n9076), .ZN(n9073)
         );
  NOR3_X1 U10436 ( .A1(n9074), .A2(n9073), .A3(n9437), .ZN(n9128) );
  INV_X1 U10437 ( .A(n9075), .ZN(n9101) );
  AOI21_X1 U10438 ( .B1(n6920), .B2(n10251), .A(n9076), .ZN(n9079) );
  INV_X1 U10439 ( .A(n9077), .ZN(n9078) );
  AND2_X1 U10440 ( .A1(n9079), .A2(n9078), .ZN(n9081) );
  NAND3_X1 U10441 ( .A1(n9084), .A2(n9083), .A3(n9082), .ZN(n9087) );
  INV_X1 U10442 ( .A(n9085), .ZN(n9086) );
  NAND2_X1 U10443 ( .A1(n9087), .A2(n9086), .ZN(n9093) );
  OAI21_X1 U10444 ( .B1(n9090), .B2(n9089), .A(n9088), .ZN(n9092) );
  AOI21_X1 U10445 ( .B1(n9093), .B2(n9092), .A(n9091), .ZN(n9096) );
  INV_X1 U10446 ( .A(n9094), .ZN(n9095) );
  OAI21_X1 U10447 ( .B1(n9097), .B2(n9096), .A(n9095), .ZN(n9098) );
  NAND2_X1 U10448 ( .A1(n9099), .A2(n9098), .ZN(n9100) );
  NAND2_X1 U10449 ( .A1(n9101), .A2(n9100), .ZN(n9105) );
  INV_X1 U10450 ( .A(n9102), .ZN(n9103) );
  AOI21_X1 U10451 ( .B1(n9105), .B2(n9104), .A(n9103), .ZN(n9106) );
  NOR2_X1 U10452 ( .A1(n9106), .A2(n9238), .ZN(n9109) );
  OAI21_X1 U10453 ( .B1(n9109), .B2(n9108), .A(n9107), .ZN(n9110) );
  AND2_X1 U10454 ( .A1(n9111), .A2(n9110), .ZN(n9112) );
  OR2_X1 U10455 ( .A1(n9113), .A2(n9112), .ZN(n9115) );
  INV_X1 U10456 ( .A(n9116), .ZN(n9119) );
  NAND3_X1 U10457 ( .A1(n9120), .A2(n10206), .A3(n9437), .ZN(n9118) );
  OAI211_X1 U10458 ( .C1(n9120), .C2(n9119), .A(n9118), .B(n9117), .ZN(n9127)
         );
  NAND4_X1 U10459 ( .A1(n9122), .A2(n10049), .A3(n9193), .A4(n9121), .ZN(n9123) );
  OAI211_X1 U10460 ( .C1(n9125), .C2(n9124), .A(n9123), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9126) );
  OAI21_X1 U10461 ( .B1(n9128), .B2(n9127), .A(n9126), .ZN(P1_U3240) );
  MUX2_X1 U10462 ( .A(n9247), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9138), .Z(
        P1_U3585) );
  MUX2_X1 U10463 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9129), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10464 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9248), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10465 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9298), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10466 ( .A(n9220), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9138), .Z(
        P1_U3581) );
  MUX2_X1 U10467 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9327), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10468 ( .A(n9349), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9138), .Z(
        P1_U3579) );
  MUX2_X1 U10469 ( .A(n9362), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9138), .Z(
        P1_U3578) );
  MUX2_X1 U10470 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9348), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10471 ( .A(n9361), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9138), .Z(
        P1_U3576) );
  MUX2_X1 U10472 ( .A(n9206), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9138), .Z(
        P1_U3575) );
  MUX2_X1 U10473 ( .A(n9203), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9138), .Z(
        P1_U3574) );
  INV_X1 U10474 ( .A(n9411), .ZN(n9422) );
  MUX2_X1 U10475 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9422), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10476 ( .A(n9130), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9138), .Z(
        P1_U3572) );
  MUX2_X1 U10477 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9421), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10478 ( .A(n9131), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9138), .Z(
        P1_U3570) );
  MUX2_X1 U10479 ( .A(n9132), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9138), .Z(
        P1_U3569) );
  MUX2_X1 U10480 ( .A(n10013), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9138), .Z(
        P1_U3568) );
  MUX2_X1 U10481 ( .A(n9133), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9138), .Z(
        P1_U3567) );
  MUX2_X1 U10482 ( .A(n10014), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9138), .Z(
        P1_U3566) );
  MUX2_X1 U10483 ( .A(n9134), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9138), .Z(
        P1_U3565) );
  MUX2_X1 U10484 ( .A(n9135), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9138), .Z(
        P1_U3564) );
  MUX2_X1 U10485 ( .A(n9136), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9138), .Z(
        P1_U3563) );
  MUX2_X1 U10486 ( .A(n10174), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9138), .Z(
        P1_U3562) );
  MUX2_X1 U10487 ( .A(n10204), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9138), .Z(
        P1_U3561) );
  MUX2_X1 U10488 ( .A(n10224), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9138), .Z(
        P1_U3560) );
  MUX2_X1 U10489 ( .A(n9137), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9138), .Z(
        P1_U3559) );
  MUX2_X1 U10490 ( .A(n10225), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9138), .Z(
        P1_U3558) );
  MUX2_X1 U10491 ( .A(n7020), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9138), .Z(
        P1_U3557) );
  MUX2_X1 U10492 ( .A(n6920), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9138), .Z(
        P1_U3556) );
  AOI211_X1 U10493 ( .C1(n9141), .C2(n9140), .A(n9139), .B(n10159), .ZN(n9142)
         );
  AOI21_X1 U10494 ( .B1(n10129), .B2(n9143), .A(n9142), .ZN(n9151) );
  NAND2_X1 U10495 ( .A1(n10079), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n9149) );
  NAND3_X1 U10496 ( .A1(n10056), .A2(n9145), .A3(n9144), .ZN(n9147) );
  NAND3_X1 U10497 ( .A1(n10147), .A2(n9147), .A3(n9146), .ZN(n9148) );
  NAND4_X1 U10498 ( .A1(n9151), .A2(n9150), .A3(n9149), .A4(n9148), .ZN(
        P1_U3244) );
  OAI21_X1 U10499 ( .B1(n9154), .B2(n9153), .A(n9152), .ZN(n9155) );
  AOI22_X1 U10500 ( .A1(n9156), .A2(n10129), .B1(n10086), .B2(n9155), .ZN(
        n9164) );
  INV_X1 U10501 ( .A(n9157), .ZN(n9163) );
  NAND2_X1 U10502 ( .A1(n10079), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n9162) );
  OAI211_X1 U10503 ( .C1(n9160), .C2(n9159), .A(n10147), .B(n9158), .ZN(n9161)
         );
  NAND4_X1 U10504 ( .A1(n9164), .A2(n9163), .A3(n9162), .A4(n9161), .ZN(
        P1_U3246) );
  NAND2_X1 U10505 ( .A1(n9166), .A2(n9179), .ZN(n9168) );
  NAND2_X1 U10506 ( .A1(n9168), .A2(n9167), .ZN(n9169) );
  NOR2_X1 U10507 ( .A1(n9180), .A2(n9169), .ZN(n9170) );
  XNOR2_X1 U10508 ( .A(n9169), .B(n9180), .ZN(n10114) );
  NOR2_X1 U10509 ( .A1(n7751), .A2(n10114), .ZN(n10113) );
  NAND2_X1 U10510 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n10128), .ZN(n9171) );
  OAI21_X1 U10511 ( .B1(n10128), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9171), .ZN(
        n10124) );
  NOR2_X1 U10512 ( .A1(n10125), .A2(n10124), .ZN(n10123) );
  AOI21_X1 U10513 ( .B1(n10128), .B2(P1_REG2_REG_16__SCAN_IN), .A(n10123), 
        .ZN(n10136) );
  OR2_X1 U10514 ( .A1(n9177), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9173) );
  NAND2_X1 U10515 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9177), .ZN(n9172) );
  NAND2_X1 U10516 ( .A1(n9173), .A2(n9172), .ZN(n10137) );
  NOR2_X1 U10517 ( .A1(n10136), .A2(n10137), .ZN(n10138) );
  MUX2_X1 U10518 ( .A(n9174), .B(P1_REG2_REG_18__SCAN_IN), .S(n9176), .Z(
        n10154) );
  NOR2_X1 U10519 ( .A1(n10153), .A2(n10154), .ZN(n10155) );
  AOI21_X1 U10520 ( .B1(n9176), .B2(P1_REG2_REG_18__SCAN_IN), .A(n10155), .ZN(
        n9175) );
  XNOR2_X1 U10521 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9175), .ZN(n9190) );
  XNOR2_X1 U10522 ( .A(n9176), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n10167) );
  INV_X1 U10523 ( .A(n9177), .ZN(n10144) );
  XNOR2_X1 U10524 ( .A(n10144), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n10149) );
  INV_X1 U10525 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9183) );
  XOR2_X1 U10526 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10128), .Z(n10131) );
  NAND2_X1 U10527 ( .A1(n10117), .A2(n9181), .ZN(n9182) );
  NAND2_X1 U10528 ( .A1(n10131), .A2(n10132), .ZN(n10130) );
  AOI21_X1 U10529 ( .B1(n10162), .B2(n9186), .A(n10165), .ZN(n9188) );
  INV_X1 U10530 ( .A(n9190), .ZN(n9192) );
  INV_X1 U10531 ( .A(n9491), .ZN(n9400) );
  NAND2_X1 U10532 ( .A1(n9396), .A2(n9400), .ZN(n9397) );
  NAND2_X1 U10533 ( .A1(n9250), .A2(n9436), .ZN(n9432) );
  XNOR2_X1 U10534 ( .A(n9432), .B(n9431), .ZN(n9429) );
  NAND2_X1 U10535 ( .A1(n9429), .A2(n10221), .ZN(n9196) );
  AOI21_X1 U10536 ( .B1(n9193), .B2(P1_B_REG_SCAN_IN), .A(n10183), .ZN(n9246)
         );
  NAND2_X1 U10537 ( .A1(n9194), .A2(n9246), .ZN(n9434) );
  NOR2_X1 U10538 ( .A1(n10215), .A2(n9434), .ZN(n9198) );
  AOI21_X1 U10539 ( .B1(P1_REG2_REG_31__SCAN_IN), .B2(n10215), .A(n9198), .ZN(
        n9195) );
  OAI211_X1 U10540 ( .C1(n9431), .C2(n10239), .A(n9196), .B(n9195), .ZN(
        P1_U3261) );
  NAND2_X1 U10541 ( .A1(n4735), .A2(n9197), .ZN(n9433) );
  NAND3_X1 U10542 ( .A1(n9433), .A2(n10221), .A3(n9432), .ZN(n9200) );
  AOI21_X1 U10543 ( .B1(n10215), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9198), .ZN(
        n9199) );
  OAI211_X1 U10544 ( .C1(n9436), .C2(n10239), .A(n9200), .B(n9199), .ZN(
        P1_U3262) );
  NAND2_X1 U10545 ( .A1(n9395), .A2(n9202), .ZN(n9205) );
  NAND2_X1 U10546 ( .A1(n9491), .A2(n9203), .ZN(n9204) );
  NAND2_X1 U10547 ( .A1(n9205), .A2(n9204), .ZN(n9380) );
  OAI21_X1 U10548 ( .B1(n9486), .B2(n9206), .A(n9380), .ZN(n9208) );
  NAND2_X1 U10549 ( .A1(n9486), .A2(n9206), .ZN(n9207) );
  NAND2_X1 U10550 ( .A1(n9208), .A2(n9207), .ZN(n9367) );
  NAND2_X1 U10551 ( .A1(n9367), .A2(n9368), .ZN(n9210) );
  NAND2_X1 U10552 ( .A1(n9481), .A2(n9361), .ZN(n9209) );
  NOR2_X1 U10553 ( .A1(n9358), .A2(n9371), .ZN(n9212) );
  NAND2_X1 U10554 ( .A1(n9358), .A2(n9371), .ZN(n9211) );
  NAND2_X1 U10555 ( .A1(n9469), .A2(n9362), .ZN(n9213) );
  NAND2_X1 U10556 ( .A1(n9306), .A2(n9218), .ZN(n9219) );
  NOR2_X1 U10557 ( .A1(n9454), .A2(n9220), .ZN(n9221) );
  NAND2_X1 U10558 ( .A1(n9268), .A2(n9267), .ZN(n9266) );
  NAND2_X1 U10559 ( .A1(n9266), .A2(n4554), .ZN(n9225) );
  XNOR2_X1 U10560 ( .A(n9225), .B(n9224), .ZN(n9439) );
  INV_X1 U10561 ( .A(n9439), .ZN(n9256) );
  AOI22_X1 U10562 ( .A1(n9251), .A2(n10187), .B1(P1_REG2_REG_29__SCAN_IN), 
        .B2(n10215), .ZN(n9255) );
  INV_X1 U10563 ( .A(n9226), .ZN(n9228) );
  NOR2_X1 U10564 ( .A1(n9346), .A2(n9347), .ZN(n9324) );
  INV_X1 U10565 ( .A(n9242), .ZN(n9243) );
  AOI22_X1 U10566 ( .A1(n10226), .A2(n9248), .B1(n9247), .B2(n9246), .ZN(n9249) );
  OAI22_X1 U10567 ( .A1(n9441), .A2(n10206), .B1(n10237), .B2(n9252), .ZN(
        n9253) );
  OAI21_X1 U10568 ( .B1(n9443), .B2(n9253), .A(n9403), .ZN(n9254) );
  OAI211_X1 U10569 ( .C1(n9256), .C2(n9428), .A(n9255), .B(n9254), .ZN(
        P1_U3355) );
  AOI211_X1 U10570 ( .C1(n4526), .C2(n9267), .A(n10228), .B(n9257), .ZN(n9261)
         );
  OAI22_X1 U10571 ( .A1(n9259), .A2(n10209), .B1(n9258), .B2(n10183), .ZN(
        n9260) );
  NOR2_X1 U10572 ( .A1(n9261), .A2(n9260), .ZN(n9447) );
  AOI21_X1 U10573 ( .B1(n9444), .B2(n9278), .A(n4540), .ZN(n9445) );
  NOR2_X1 U10574 ( .A1(n4738), .A2(n10239), .ZN(n9265) );
  OAI22_X1 U10575 ( .A1(n9403), .A2(n9263), .B1(n9262), .B2(n10237), .ZN(n9264) );
  AOI211_X1 U10576 ( .C1(n9445), .C2(n10221), .A(n9265), .B(n9264), .ZN(n9270)
         );
  OAI21_X1 U10577 ( .B1(n9268), .B2(n9267), .A(n9266), .ZN(n9448) );
  OR2_X1 U10578 ( .A1(n9448), .A2(n9428), .ZN(n9269) );
  OAI211_X1 U10579 ( .C1(n9447), .C2(n10215), .A(n9270), .B(n9269), .ZN(
        P1_U3263) );
  XNOR2_X1 U10580 ( .A(n9271), .B(n9274), .ZN(n9453) );
  AOI211_X1 U10581 ( .C1(n9274), .C2(n9273), .A(n10228), .B(n9272), .ZN(n9277)
         );
  OAI22_X1 U10582 ( .A1(n9317), .A2(n10209), .B1(n9275), .B2(n10183), .ZN(
        n9276) );
  NOR2_X1 U10583 ( .A1(n9277), .A2(n9276), .ZN(n9452) );
  INV_X1 U10584 ( .A(n9289), .ZN(n9280) );
  INV_X1 U10585 ( .A(n9278), .ZN(n9279) );
  AOI211_X1 U10586 ( .C1(n9450), .C2(n9280), .A(n10306), .B(n9279), .ZN(n9449)
         );
  NAND2_X1 U10587 ( .A1(n9449), .A2(n9332), .ZN(n9281) );
  OAI211_X1 U10588 ( .C1(n9282), .C2(n10237), .A(n9452), .B(n9281), .ZN(n9286)
         );
  OAI22_X1 U10589 ( .A1(n9284), .A2(n10239), .B1(n9283), .B2(n9403), .ZN(n9285) );
  AOI21_X1 U10590 ( .B1(n9286), .B2(n9403), .A(n9285), .ZN(n9287) );
  OAI21_X1 U10591 ( .B1(n9453), .B2(n9428), .A(n9287), .ZN(P1_U3264) );
  XNOR2_X1 U10592 ( .A(n9288), .B(n9296), .ZN(n9458) );
  INV_X1 U10593 ( .A(n9304), .ZN(n9290) );
  AOI21_X1 U10594 ( .B1(n9454), .B2(n9290), .A(n9289), .ZN(n9455) );
  AOI22_X1 U10595 ( .A1(n10215), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9291), 
        .B2(n10203), .ZN(n9292) );
  OAI21_X1 U10596 ( .B1(n9293), .B2(n10239), .A(n9292), .ZN(n9301) );
  NOR2_X1 U10597 ( .A1(n9295), .A2(n9294), .ZN(n9297) );
  XNOR2_X1 U10598 ( .A(n9297), .B(n9296), .ZN(n9299) );
  AOI222_X1 U10599 ( .A1(n9424), .A2(n9299), .B1(n9298), .B2(n10223), .C1(
        n9327), .C2(n10226), .ZN(n9457) );
  NOR2_X1 U10600 ( .A1(n9457), .A2(n10215), .ZN(n9300) );
  AOI211_X1 U10601 ( .C1(n10221), .C2(n9455), .A(n9301), .B(n9300), .ZN(n9302)
         );
  OAI21_X1 U10602 ( .B1(n9428), .B2(n9458), .A(n9302), .ZN(P1_U3265) );
  XOR2_X1 U10603 ( .A(n9313), .B(n9303), .Z(n9463) );
  AOI211_X1 U10604 ( .C1(n9305), .C2(n9329), .A(n10306), .B(n9304), .ZN(n9459)
         );
  NOR2_X1 U10605 ( .A1(n9306), .A2(n10239), .ZN(n9310) );
  OAI22_X1 U10606 ( .A1(n9403), .A2(n9308), .B1(n9307), .B2(n10237), .ZN(n9309) );
  AOI211_X1 U10607 ( .C1(n9459), .C2(n9406), .A(n9310), .B(n9309), .ZN(n9319)
         );
  INV_X1 U10608 ( .A(n9311), .ZN(n9312) );
  NOR2_X1 U10609 ( .A1(n9321), .A2(n9312), .ZN(n9314) );
  XNOR2_X1 U10610 ( .A(n9314), .B(n9313), .ZN(n9315) );
  OAI222_X1 U10611 ( .A1(n10183), .A2(n9317), .B1(n10209), .B2(n9316), .C1(
        n9315), .C2(n10228), .ZN(n9461) );
  NAND2_X1 U10612 ( .A1(n9461), .A2(n9403), .ZN(n9318) );
  OAI211_X1 U10613 ( .C1(n9463), .C2(n9428), .A(n9319), .B(n9318), .ZN(
        P1_U3266) );
  XNOR2_X1 U10614 ( .A(n9320), .B(n9322), .ZN(n9468) );
  INV_X1 U10615 ( .A(n9321), .ZN(n9326) );
  OAI21_X1 U10616 ( .B1(n9324), .B2(n9323), .A(n9322), .ZN(n9325) );
  NAND2_X1 U10617 ( .A1(n9326), .A2(n9325), .ZN(n9328) );
  AOI222_X1 U10618 ( .A1(n9424), .A2(n9328), .B1(n9327), .B2(n10223), .C1(
        n9362), .C2(n10226), .ZN(n9467) );
  AOI211_X1 U10619 ( .C1(n9330), .C2(n9340), .A(n10306), .B(n4749), .ZN(n9465)
         );
  AOI22_X1 U10620 ( .A1(n9465), .A2(n9332), .B1(n10203), .B2(n9331), .ZN(n9333) );
  AOI21_X1 U10621 ( .B1(n9467), .B2(n9333), .A(n10215), .ZN(n9337) );
  OAI22_X1 U10622 ( .A1(n9335), .A2(n10239), .B1(n9403), .B2(n9334), .ZN(n9336) );
  NOR2_X1 U10623 ( .A1(n9337), .A2(n9336), .ZN(n9338) );
  OAI21_X1 U10624 ( .B1(n9428), .B2(n9468), .A(n9338), .ZN(P1_U3267) );
  XOR2_X1 U10625 ( .A(n9339), .B(n9347), .Z(n9473) );
  INV_X1 U10626 ( .A(n9355), .ZN(n9341) );
  AOI21_X1 U10627 ( .B1(n9469), .B2(n9341), .A(n4750), .ZN(n9470) );
  INV_X1 U10628 ( .A(n9342), .ZN(n9343) );
  AOI22_X1 U10629 ( .A1(n10215), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9343), 
        .B2(n10203), .ZN(n9344) );
  OAI21_X1 U10630 ( .B1(n9345), .B2(n10239), .A(n9344), .ZN(n9352) );
  XOR2_X1 U10631 ( .A(n9347), .B(n9346), .Z(n9350) );
  AOI222_X1 U10632 ( .A1(n9424), .A2(n9350), .B1(n9349), .B2(n10223), .C1(
        n9348), .C2(n10226), .ZN(n9472) );
  NOR2_X1 U10633 ( .A1(n9472), .A2(n10215), .ZN(n9351) );
  AOI211_X1 U10634 ( .C1(n9470), .C2(n10221), .A(n9352), .B(n9351), .ZN(n9353)
         );
  OAI21_X1 U10635 ( .B1(n9473), .B2(n9428), .A(n9353), .ZN(P1_U3268) );
  XOR2_X1 U10636 ( .A(n9354), .B(n9359), .Z(n9478) );
  AOI21_X1 U10637 ( .B1(n9474), .B2(n9372), .A(n9355), .ZN(n9475) );
  AOI22_X1 U10638 ( .A1(n10215), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9356), 
        .B2(n10203), .ZN(n9357) );
  OAI21_X1 U10639 ( .B1(n9358), .B2(n10239), .A(n9357), .ZN(n9365) );
  XOR2_X1 U10640 ( .A(n9360), .B(n9359), .Z(n9363) );
  AOI222_X1 U10641 ( .A1(n9424), .A2(n9363), .B1(n9362), .B2(n10223), .C1(
        n9361), .C2(n10226), .ZN(n9477) );
  NOR2_X1 U10642 ( .A1(n9477), .A2(n10215), .ZN(n9364) );
  AOI211_X1 U10643 ( .C1(n9475), .C2(n10221), .A(n9365), .B(n9364), .ZN(n9366)
         );
  OAI21_X1 U10644 ( .B1(n9478), .B2(n9428), .A(n9366), .ZN(P1_U3269) );
  XNOR2_X1 U10645 ( .A(n9367), .B(n9368), .ZN(n9483) );
  XNOR2_X1 U10646 ( .A(n9369), .B(n9368), .ZN(n9370) );
  OAI222_X1 U10647 ( .A1(n10183), .A2(n9371), .B1(n10209), .B2(n9410), .C1(
        n10228), .C2(n9370), .ZN(n9479) );
  INV_X1 U10648 ( .A(n9481), .ZN(n9377) );
  AOI211_X1 U10649 ( .C1(n9481), .C2(n9386), .A(n10306), .B(n4754), .ZN(n9480)
         );
  NAND2_X1 U10650 ( .A1(n9480), .A2(n9406), .ZN(n9376) );
  INV_X1 U10651 ( .A(n9373), .ZN(n9374) );
  AOI22_X1 U10652 ( .A1(n10215), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9374), 
        .B2(n10203), .ZN(n9375) );
  OAI211_X1 U10653 ( .C1(n9377), .C2(n10239), .A(n9376), .B(n9375), .ZN(n9378)
         );
  AOI21_X1 U10654 ( .B1(n9479), .B2(n9403), .A(n9378), .ZN(n9379) );
  OAI21_X1 U10655 ( .B1(n9483), .B2(n9428), .A(n9379), .ZN(P1_U3270) );
  XNOR2_X1 U10656 ( .A(n9380), .B(n9381), .ZN(n9488) );
  XOR2_X1 U10657 ( .A(n9382), .B(n9381), .Z(n9383) );
  OAI222_X1 U10658 ( .A1(n10183), .A2(n9385), .B1(n10209), .B2(n9384), .C1(
        n9383), .C2(n10228), .ZN(n9484) );
  INV_X1 U10659 ( .A(n9386), .ZN(n9387) );
  AOI211_X1 U10660 ( .C1(n9486), .C2(n9397), .A(n10306), .B(n9387), .ZN(n9485)
         );
  NAND2_X1 U10661 ( .A1(n9485), .A2(n9406), .ZN(n9391) );
  INV_X1 U10662 ( .A(n9388), .ZN(n9389) );
  AOI22_X1 U10663 ( .A1(n10215), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9389), 
        .B2(n10203), .ZN(n9390) );
  OAI211_X1 U10664 ( .C1(n9392), .C2(n10239), .A(n9391), .B(n9390), .ZN(n9393)
         );
  AOI21_X1 U10665 ( .B1(n9484), .B2(n9403), .A(n9393), .ZN(n9394) );
  OAI21_X1 U10666 ( .B1(n9488), .B2(n9428), .A(n9394), .ZN(P1_U3271) );
  XNOR2_X1 U10667 ( .A(n9395), .B(n9407), .ZN(n9493) );
  INV_X1 U10668 ( .A(n9396), .ZN(n9399) );
  INV_X1 U10669 ( .A(n9397), .ZN(n9398) );
  AOI211_X1 U10670 ( .C1(n9491), .C2(n9399), .A(n10306), .B(n9398), .ZN(n9490)
         );
  NOR2_X1 U10671 ( .A1(n9400), .A2(n10239), .ZN(n9405) );
  OAI22_X1 U10672 ( .A1(n9403), .A2(n9402), .B1(n9401), .B2(n10237), .ZN(n9404) );
  AOI211_X1 U10673 ( .C1(n9490), .C2(n9406), .A(n9405), .B(n9404), .ZN(n9413)
         );
  AOI21_X1 U10674 ( .B1(n9408), .B2(n9407), .A(n4532), .ZN(n9409) );
  OAI222_X1 U10675 ( .A1(n10209), .A2(n9411), .B1(n10183), .B2(n9410), .C1(
        n10228), .C2(n9409), .ZN(n9489) );
  NAND2_X1 U10676 ( .A1(n9489), .A2(n9403), .ZN(n9412) );
  OAI211_X1 U10677 ( .C1(n9493), .C2(n9428), .A(n9413), .B(n9412), .ZN(
        P1_U3272) );
  XNOR2_X1 U10678 ( .A(n4564), .B(n9419), .ZN(n9504) );
  AOI21_X1 U10679 ( .B1(n9500), .B2(n9414), .A(n4559), .ZN(n9501) );
  INV_X1 U10680 ( .A(n9415), .ZN(n9416) );
  AOI22_X1 U10681 ( .A1(n10215), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9416), 
        .B2(n10203), .ZN(n9417) );
  OAI21_X1 U10682 ( .B1(n9418), .B2(n10239), .A(n9417), .ZN(n9426) );
  XNOR2_X1 U10683 ( .A(n9420), .B(n9419), .ZN(n9423) );
  AOI222_X1 U10684 ( .A1(n9424), .A2(n9423), .B1(n9422), .B2(n10223), .C1(
        n9421), .C2(n10226), .ZN(n9503) );
  NOR2_X1 U10685 ( .A1(n9503), .A2(n10215), .ZN(n9425) );
  AOI211_X1 U10686 ( .C1(n9501), .C2(n10221), .A(n9426), .B(n9425), .ZN(n9427)
         );
  OAI21_X1 U10687 ( .B1(n9504), .B2(n9428), .A(n9427), .ZN(P1_U3274) );
  NAND2_X1 U10688 ( .A1(n9429), .A2(n10198), .ZN(n9430) );
  OAI211_X1 U10689 ( .C1(n9431), .C2(n10304), .A(n9430), .B(n9434), .ZN(n9530)
         );
  MUX2_X1 U10690 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9530), .S(n10326), .Z(
        P1_U3554) );
  NAND3_X1 U10691 ( .A1(n9433), .A2(n10198), .A3(n9432), .ZN(n9435) );
  OAI211_X1 U10692 ( .C1(n9436), .C2(n10304), .A(n9435), .B(n9434), .ZN(n9531)
         );
  MUX2_X1 U10693 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9531), .S(n10326), .Z(
        P1_U3553) );
  AND2_X1 U10694 ( .A1(n9438), .A2(n9437), .ZN(n10309) );
  OR2_X1 U10695 ( .A1(n10309), .A2(n10184), .ZN(n10295) );
  AOI22_X1 U10696 ( .A1(n9445), .A2(n10198), .B1(n9524), .B2(n9444), .ZN(n9446) );
  OAI211_X1 U10697 ( .C1(n9448), .C2(n9520), .A(n9447), .B(n9446), .ZN(n9533)
         );
  MUX2_X1 U10698 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9533), .S(n10326), .Z(
        P1_U3551) );
  AOI21_X1 U10699 ( .B1(n9524), .B2(n9450), .A(n9449), .ZN(n9451) );
  OAI211_X1 U10700 ( .C1(n9453), .C2(n9520), .A(n9452), .B(n9451), .ZN(n9534)
         );
  MUX2_X1 U10701 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9534), .S(n10326), .Z(
        P1_U3550) );
  AOI22_X1 U10702 ( .A1(n9455), .A2(n10198), .B1(n9524), .B2(n9454), .ZN(n9456) );
  OAI211_X1 U10703 ( .C1(n9458), .C2(n9520), .A(n9457), .B(n9456), .ZN(n9535)
         );
  MUX2_X1 U10704 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9535), .S(n10326), .Z(
        P1_U3549) );
  NOR3_X1 U10705 ( .A1(n9461), .A2(n9460), .A3(n9459), .ZN(n9462) );
  OAI21_X1 U10706 ( .B1(n9463), .B2(n9520), .A(n9462), .ZN(n9536) );
  MUX2_X1 U10707 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9536), .S(n10326), .Z(
        P1_U3548) );
  NOR2_X1 U10708 ( .A1(n9465), .A2(n9464), .ZN(n9466) );
  OAI211_X1 U10709 ( .C1(n9468), .C2(n9520), .A(n9467), .B(n9466), .ZN(n9537)
         );
  MUX2_X1 U10710 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9537), .S(n10326), .Z(
        P1_U3547) );
  AOI22_X1 U10711 ( .A1(n9470), .A2(n10198), .B1(n9524), .B2(n9469), .ZN(n9471) );
  OAI211_X1 U10712 ( .C1(n9473), .C2(n9520), .A(n9472), .B(n9471), .ZN(n9538)
         );
  MUX2_X1 U10713 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9538), .S(n10326), .Z(
        P1_U3546) );
  AOI22_X1 U10714 ( .A1(n9475), .A2(n10198), .B1(n9524), .B2(n9474), .ZN(n9476) );
  OAI211_X1 U10715 ( .C1(n9478), .C2(n9520), .A(n9477), .B(n9476), .ZN(n9539)
         );
  MUX2_X1 U10716 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9539), .S(n10326), .Z(
        P1_U3545) );
  AOI211_X1 U10717 ( .C1(n9524), .C2(n9481), .A(n9480), .B(n9479), .ZN(n9482)
         );
  OAI21_X1 U10718 ( .B1(n9483), .B2(n9520), .A(n9482), .ZN(n9540) );
  MUX2_X1 U10719 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9540), .S(n10326), .Z(
        P1_U3544) );
  AOI211_X1 U10720 ( .C1(n9524), .C2(n9486), .A(n9485), .B(n9484), .ZN(n9487)
         );
  OAI21_X1 U10721 ( .B1(n9488), .B2(n9520), .A(n9487), .ZN(n9541) );
  MUX2_X1 U10722 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9541), .S(n10326), .Z(
        P1_U3543) );
  AOI211_X1 U10723 ( .C1(n9524), .C2(n9491), .A(n9490), .B(n9489), .ZN(n9492)
         );
  OAI21_X1 U10724 ( .B1(n9493), .B2(n9520), .A(n9492), .ZN(n9542) );
  MUX2_X1 U10725 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9542), .S(n10326), .Z(
        P1_U3542) );
  NAND3_X1 U10726 ( .A1(n9495), .A2(n9494), .A3(n10295), .ZN(n9499) );
  NAND4_X1 U10727 ( .A1(n9499), .A2(n9498), .A3(n9497), .A4(n9496), .ZN(n9543)
         );
  MUX2_X1 U10728 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9543), .S(n10326), .Z(
        P1_U3541) );
  AOI22_X1 U10729 ( .A1(n9501), .A2(n10198), .B1(n9524), .B2(n9500), .ZN(n9502) );
  OAI211_X1 U10730 ( .C1(n9504), .C2(n9520), .A(n9503), .B(n9502), .ZN(n9544)
         );
  MUX2_X1 U10731 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9544), .S(n10326), .Z(
        P1_U3540) );
  AOI211_X1 U10732 ( .C1(n9524), .C2(n9507), .A(n9506), .B(n9505), .ZN(n9508)
         );
  OAI21_X1 U10733 ( .B1(n9509), .B2(n9520), .A(n9508), .ZN(n9545) );
  MUX2_X1 U10734 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9545), .S(n10326), .Z(
        P1_U3539) );
  OAI22_X1 U10735 ( .A1(n9511), .A2(n10306), .B1(n9510), .B2(n10304), .ZN(
        n9513) );
  AOI211_X1 U10736 ( .C1(n10309), .C2(n9514), .A(n9513), .B(n9512), .ZN(n9546)
         );
  MUX2_X1 U10737 ( .A(n5588), .B(n9546), .S(n10326), .Z(n9515) );
  INV_X1 U10738 ( .A(n9515), .ZN(P1_U3538) );
  AOI22_X1 U10739 ( .A1(n9517), .A2(n10198), .B1(n9524), .B2(n9516), .ZN(n9518) );
  OAI211_X1 U10740 ( .C1(n9521), .C2(n9520), .A(n9519), .B(n9518), .ZN(n9549)
         );
  MUX2_X1 U10741 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9549), .S(n10326), .Z(
        P1_U3536) );
  INV_X1 U10742 ( .A(n10309), .ZN(n9529) );
  INV_X1 U10743 ( .A(n9522), .ZN(n9528) );
  AOI22_X1 U10744 ( .A1(n9525), .A2(n10198), .B1(n9524), .B2(n9523), .ZN(n9526) );
  OAI211_X1 U10745 ( .C1(n9529), .C2(n9528), .A(n9527), .B(n9526), .ZN(n9550)
         );
  MUX2_X1 U10746 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9550), .S(n10326), .Z(
        P1_U3534) );
  MUX2_X1 U10747 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9530), .S(n10315), .Z(
        P1_U3522) );
  MUX2_X1 U10748 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9531), .S(n10315), .Z(
        P1_U3521) );
  MUX2_X1 U10749 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9533), .S(n10315), .Z(
        P1_U3519) );
  MUX2_X1 U10750 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9534), .S(n10315), .Z(
        P1_U3518) );
  MUX2_X1 U10751 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9535), .S(n10315), .Z(
        P1_U3517) );
  MUX2_X1 U10752 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9536), .S(n10315), .Z(
        P1_U3516) );
  MUX2_X1 U10753 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9537), .S(n10315), .Z(
        P1_U3515) );
  MUX2_X1 U10754 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9538), .S(n10315), .Z(
        P1_U3514) );
  MUX2_X1 U10755 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9539), .S(n10315), .Z(
        P1_U3513) );
  MUX2_X1 U10756 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9540), .S(n10315), .Z(
        P1_U3512) );
  MUX2_X1 U10757 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9541), .S(n10315), .Z(
        P1_U3511) );
  MUX2_X1 U10758 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9542), .S(n10315), .Z(
        P1_U3510) );
  MUX2_X1 U10759 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9543), .S(n10315), .Z(
        P1_U3508) );
  MUX2_X1 U10760 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9544), .S(n10315), .Z(
        P1_U3505) );
  MUX2_X1 U10761 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9545), .S(n10315), .Z(
        P1_U3502) );
  INV_X1 U10762 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9547) );
  MUX2_X1 U10763 ( .A(n9547), .B(n9546), .S(n10315), .Z(n9548) );
  INV_X1 U10764 ( .A(n9548), .ZN(P1_U3499) );
  MUX2_X1 U10765 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9549), .S(n10315), .Z(
        P1_U3493) );
  MUX2_X1 U10766 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n9550), .S(n10315), .Z(
        P1_U3487) );
  MUX2_X1 U10767 ( .A(n9551), .B(P1_D_REG_0__SCAN_IN), .S(n10247), .Z(P1_U3440) );
  NAND3_X1 U10768 ( .A1(n9552), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n9554) );
  OAI22_X1 U10769 ( .A1(n9555), .A2(n9554), .B1(n6563), .B2(n9553), .ZN(n9556)
         );
  INV_X1 U10770 ( .A(n9556), .ZN(n9557) );
  OAI21_X1 U10771 ( .B1(n9558), .B2(n9560), .A(n9557), .ZN(P1_U3322) );
  OAI222_X1 U10772 ( .A1(n9562), .A2(n9718), .B1(P1_U3084), .B2(n9561), .C1(
        n9560), .C2(n9559), .ZN(P1_U3324) );
  MUX2_X1 U10773 ( .A(n9563), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U10774 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10517) );
  NOR2_X1 U10775 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9564) );
  AOI21_X1 U10776 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9564), .ZN(n10484) );
  NOR2_X1 U10777 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9565) );
  AOI21_X1 U10778 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9565), .ZN(n10487) );
  NOR2_X1 U10779 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9566) );
  AOI21_X1 U10780 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9566), .ZN(n10490) );
  NOR2_X1 U10781 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9567) );
  AOI21_X1 U10782 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9567), .ZN(n10493) );
  NOR2_X1 U10783 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9568) );
  AOI21_X1 U10784 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9568), .ZN(n10496) );
  NOR2_X1 U10785 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9575) );
  XNOR2_X1 U10786 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10524) );
  NAND2_X1 U10787 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9573) );
  XOR2_X1 U10788 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10522) );
  NAND2_X1 U10789 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9571) );
  XOR2_X1 U10790 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10511) );
  AOI21_X1 U10791 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10478) );
  INV_X1 U10792 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9569) );
  NAND3_X1 U10793 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10480) );
  OAI21_X1 U10794 ( .B1(n10478), .B2(n9569), .A(n10480), .ZN(n10510) );
  NAND2_X1 U10795 ( .A1(n10511), .A2(n10510), .ZN(n9570) );
  NAND2_X1 U10796 ( .A1(n9571), .A2(n9570), .ZN(n10521) );
  NAND2_X1 U10797 ( .A1(n10522), .A2(n10521), .ZN(n9572) );
  NAND2_X1 U10798 ( .A1(n9573), .A2(n9572), .ZN(n10523) );
  NOR2_X1 U10799 ( .A1(n10524), .A2(n10523), .ZN(n9574) );
  NOR2_X1 U10800 ( .A1(n9575), .A2(n9574), .ZN(n9576) );
  NOR2_X1 U10801 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9576), .ZN(n10513) );
  AND2_X1 U10802 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9576), .ZN(n10512) );
  NOR2_X1 U10803 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10512), .ZN(n9577) );
  NOR2_X1 U10804 ( .A1(n10513), .A2(n9577), .ZN(n9578) );
  NAND2_X1 U10805 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n9578), .ZN(n9580) );
  XOR2_X1 U10806 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n9578), .Z(n10520) );
  NAND2_X1 U10807 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10520), .ZN(n9579) );
  NAND2_X1 U10808 ( .A1(n9580), .A2(n9579), .ZN(n9581) );
  NAND2_X1 U10809 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9581), .ZN(n9583) );
  XOR2_X1 U10810 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9581), .Z(n10509) );
  NAND2_X1 U10811 ( .A1(n10509), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n9582) );
  NAND2_X1 U10812 ( .A1(n9583), .A2(n9582), .ZN(n9584) );
  NAND2_X1 U10813 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9584), .ZN(n9586) );
  XOR2_X1 U10814 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9584), .Z(n10519) );
  NAND2_X1 U10815 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10519), .ZN(n9585) );
  NAND2_X1 U10816 ( .A1(n9586), .A2(n9585), .ZN(n9587) );
  AND2_X1 U10817 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9587), .ZN(n9588) );
  XNOR2_X1 U10818 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9587), .ZN(n10508) );
  NAND2_X1 U10819 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9589) );
  OAI21_X1 U10820 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9589), .ZN(n10504) );
  NAND2_X1 U10821 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9590) );
  OAI21_X1 U10822 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9590), .ZN(n10501) );
  AOI21_X1 U10823 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10500), .ZN(n10499) );
  NOR2_X1 U10824 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9591) );
  AOI21_X1 U10825 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9591), .ZN(n10498) );
  NAND2_X1 U10826 ( .A1(n10499), .A2(n10498), .ZN(n10497) );
  OAI21_X1 U10827 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10497), .ZN(n10495) );
  NAND2_X1 U10828 ( .A1(n10496), .A2(n10495), .ZN(n10494) );
  OAI21_X1 U10829 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10494), .ZN(n10492) );
  NAND2_X1 U10830 ( .A1(n10493), .A2(n10492), .ZN(n10491) );
  OAI21_X1 U10831 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10491), .ZN(n10489) );
  NAND2_X1 U10832 ( .A1(n10490), .A2(n10489), .ZN(n10488) );
  OAI21_X1 U10833 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10488), .ZN(n10486) );
  NAND2_X1 U10834 ( .A1(n10487), .A2(n10486), .ZN(n10485) );
  OAI21_X1 U10835 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10485), .ZN(n10483) );
  NAND2_X1 U10836 ( .A1(n10484), .A2(n10483), .ZN(n10482) );
  OAI21_X1 U10837 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10482), .ZN(n10516) );
  NOR2_X1 U10838 ( .A1(n10517), .A2(n10516), .ZN(n9592) );
  NAND2_X1 U10839 ( .A1(n10517), .A2(n10516), .ZN(n10515) );
  OAI21_X1 U10840 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n9592), .A(n10515), .ZN(
        n9970) );
  OAI22_X1 U10841 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(keyinput_g105), .B1(SI_20_), .B2(keyinput_g12), .ZN(n9593) );
  AOI221_X1 U10842 ( .B1(P1_IR_REG_14__SCAN_IN), .B2(keyinput_g105), .C1(
        keyinput_g12), .C2(SI_20_), .A(n9593), .ZN(n9600) );
  OAI22_X1 U10843 ( .A1(SI_23_), .A2(keyinput_g9), .B1(SI_3_), .B2(
        keyinput_g29), .ZN(n9594) );
  AOI221_X1 U10844 ( .B1(SI_23_), .B2(keyinput_g9), .C1(keyinput_g29), .C2(
        SI_3_), .A(n9594), .ZN(n9599) );
  OAI22_X1 U10845 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(keyinput_g116), .B1(
        P2_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .ZN(n9595) );
  AOI221_X1 U10846 ( .B1(P1_IR_REG_25__SCAN_IN), .B2(keyinput_g116), .C1(
        keyinput_g55), .C2(P2_REG3_REG_20__SCAN_IN), .A(n9595), .ZN(n9598) );
  OAI22_X1 U10847 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput_g111), .B1(SI_26_), .B2(keyinput_g6), .ZN(n9596) );
  AOI221_X1 U10848 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput_g111), .C1(
        keyinput_g6), .C2(SI_26_), .A(n9596), .ZN(n9597) );
  NAND4_X1 U10849 ( .A1(n9600), .A2(n9599), .A3(n9598), .A4(n9597), .ZN(n9630)
         );
  OAI22_X1 U10850 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(keyinput_g74), .B1(
        keyinput_g56), .B2(P2_REG3_REG_13__SCAN_IN), .ZN(n9601) );
  AOI221_X1 U10851 ( .B1(P2_DATAO_REG_22__SCAN_IN), .B2(keyinput_g74), .C1(
        P2_REG3_REG_13__SCAN_IN), .C2(keyinput_g56), .A(n9601), .ZN(n9608) );
  OAI22_X1 U10852 ( .A1(SI_0_), .A2(keyinput_g32), .B1(keyinput_g34), .B2(
        P2_STATE_REG_SCAN_IN), .ZN(n9602) );
  AOI221_X1 U10853 ( .B1(SI_0_), .B2(keyinput_g32), .C1(P2_STATE_REG_SCAN_IN), 
        .C2(keyinput_g34), .A(n9602), .ZN(n9607) );
  OAI22_X1 U10854 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(keyinput_g102), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(keyinput_g69), .ZN(n9603) );
  AOI221_X1 U10855 ( .B1(P1_IR_REG_11__SCAN_IN), .B2(keyinput_g102), .C1(
        keyinput_g69), .C2(P2_DATAO_REG_27__SCAN_IN), .A(n9603), .ZN(n9606) );
  OAI22_X1 U10856 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(keyinput_g110), .B1(
        keyinput_g72), .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9604) );
  AOI221_X1 U10857 ( .B1(P1_IR_REG_19__SCAN_IN), .B2(keyinput_g110), .C1(
        P2_DATAO_REG_24__SCAN_IN), .C2(keyinput_g72), .A(n9604), .ZN(n9605) );
  NAND4_X1 U10858 ( .A1(n9608), .A2(n9607), .A3(n9606), .A4(n9605), .ZN(n9629)
         );
  OAI22_X1 U10859 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_g51), .B1(
        P2_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .ZN(n9609) );
  AOI221_X1 U10860 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_g51), .C1(
        keyinput_g61), .C2(P2_REG3_REG_6__SCAN_IN), .A(n9609), .ZN(n9616) );
  OAI22_X1 U10861 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(keyinput_g98), .B1(
        keyinput_g11), .B2(SI_21_), .ZN(n9610) );
  AOI221_X1 U10862 ( .B1(P1_IR_REG_7__SCAN_IN), .B2(keyinput_g98), .C1(SI_21_), 
        .C2(keyinput_g11), .A(n9610), .ZN(n9615) );
  OAI22_X1 U10863 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_g60), .B1(
        keyinput_g48), .B2(P2_REG3_REG_16__SCAN_IN), .ZN(n9611) );
  AOI221_X1 U10864 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .C1(
        P2_REG3_REG_16__SCAN_IN), .C2(keyinput_g48), .A(n9611), .ZN(n9614) );
  OAI22_X1 U10865 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput_g36), .B1(
        SI_30_), .B2(keyinput_g2), .ZN(n9612) );
  AOI221_X1 U10866 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .C1(
        keyinput_g2), .C2(SI_30_), .A(n9612), .ZN(n9613) );
  NAND4_X1 U10867 ( .A1(n9616), .A2(n9615), .A3(n9614), .A4(n9613), .ZN(n9628)
         );
  OAI22_X1 U10868 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(keyinput_g76), .B1(
        keyinput_g63), .B2(P2_REG3_REG_15__SCAN_IN), .ZN(n9617) );
  AOI221_X1 U10869 ( .B1(P2_DATAO_REG_20__SCAN_IN), .B2(keyinput_g76), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput_g63), .A(n9617), .ZN(n9626) );
  OAI22_X1 U10870 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(keyinput_g107), .B1(
        keyinput_g101), .B2(P1_IR_REG_10__SCAN_IN), .ZN(n9618) );
  AOI221_X1 U10871 ( .B1(P1_IR_REG_16__SCAN_IN), .B2(keyinput_g107), .C1(
        P1_IR_REG_10__SCAN_IN), .C2(keyinput_g101), .A(n9618), .ZN(n9625) );
  OAI22_X1 U10872 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(keyinput_g73), .B1(
        SI_12_), .B2(keyinput_g20), .ZN(n9619) );
  AOI221_X1 U10873 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(keyinput_g73), .C1(
        keyinput_g20), .C2(SI_12_), .A(n9619), .ZN(n9624) );
  XNOR2_X1 U10874 ( .A(n9620), .B(keyinput_g97), .ZN(n9622) );
  XNOR2_X1 U10875 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput_g113), .ZN(n9621)
         );
  NOR2_X1 U10876 ( .A1(n9622), .A2(n9621), .ZN(n9623) );
  NAND4_X1 U10877 ( .A1(n9626), .A2(n9625), .A3(n9624), .A4(n9623), .ZN(n9627)
         );
  NOR4_X1 U10878 ( .A1(n9630), .A2(n9629), .A3(n9628), .A4(n9627), .ZN(n9968)
         );
  OAI22_X1 U10879 ( .A1(SI_15_), .A2(keyinput_g17), .B1(keyinput_g26), .B2(
        SI_6_), .ZN(n9631) );
  AOI221_X1 U10880 ( .B1(SI_15_), .B2(keyinput_g17), .C1(SI_6_), .C2(
        keyinput_g26), .A(n9631), .ZN(n9638) );
  OAI22_X1 U10881 ( .A1(SI_16_), .A2(keyinput_g16), .B1(keyinput_g88), .B2(
        P2_DATAO_REG_8__SCAN_IN), .ZN(n9632) );
  AOI221_X1 U10882 ( .B1(SI_16_), .B2(keyinput_g16), .C1(
        P2_DATAO_REG_8__SCAN_IN), .C2(keyinput_g88), .A(n9632), .ZN(n9637) );
  OAI22_X1 U10883 ( .A1(SI_19_), .A2(keyinput_g13), .B1(keyinput_g37), .B2(
        P2_REG3_REG_14__SCAN_IN), .ZN(n9633) );
  AOI221_X1 U10884 ( .B1(SI_19_), .B2(keyinput_g13), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput_g37), .A(n9633), .ZN(n9636) );
  OAI22_X1 U10885 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(keyinput_g112), .B1(SI_24_), .B2(keyinput_g8), .ZN(n9634) );
  AOI221_X1 U10886 ( .B1(P1_IR_REG_21__SCAN_IN), .B2(keyinput_g112), .C1(
        keyinput_g8), .C2(SI_24_), .A(n9634), .ZN(n9635) );
  NAND4_X1 U10887 ( .A1(n9638), .A2(n9637), .A3(n9636), .A4(n9635), .ZN(n9767)
         );
  OAI22_X1 U10888 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput_g104), .B1(SI_8_), 
        .B2(keyinput_g24), .ZN(n9639) );
  AOI221_X1 U10889 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput_g104), .C1(
        keyinput_g24), .C2(SI_8_), .A(n9639), .ZN(n9664) );
  OAI22_X1 U10890 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(keyinput_g93), .B1(
        keyinput_g42), .B2(P2_REG3_REG_28__SCAN_IN), .ZN(n9640) );
  AOI221_X1 U10891 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(keyinput_g93), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_g42), .A(n9640), .ZN(n9643) );
  OAI22_X1 U10892 ( .A1(P1_D_REG_4__SCAN_IN), .A2(keyinput_g127), .B1(
        keyinput_g45), .B2(P2_REG3_REG_21__SCAN_IN), .ZN(n9641) );
  AOI221_X1 U10893 ( .B1(P1_D_REG_4__SCAN_IN), .B2(keyinput_g127), .C1(
        P2_REG3_REG_21__SCAN_IN), .C2(keyinput_g45), .A(n9641), .ZN(n9642) );
  OAI211_X1 U10894 ( .C1(n9842), .C2(keyinput_g43), .A(n9643), .B(n9642), .ZN(
        n9644) );
  AOI21_X1 U10895 ( .B1(n9842), .B2(keyinput_g43), .A(n9644), .ZN(n9663) );
  AOI22_X1 U10896 ( .A1(P2_B_REG_SCAN_IN), .A2(keyinput_g64), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(keyinput_g89), .ZN(n9645) );
  OAI221_X1 U10897 ( .B1(P2_B_REG_SCAN_IN), .B2(keyinput_g64), .C1(
        P2_DATAO_REG_7__SCAN_IN), .C2(keyinput_g89), .A(n9645), .ZN(n9652) );
  AOI22_X1 U10898 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_g57), .B1(SI_9_), .B2(keyinput_g23), .ZN(n9646) );
  OAI221_X1 U10899 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .C1(
        SI_9_), .C2(keyinput_g23), .A(n9646), .ZN(n9651) );
  AOI22_X1 U10900 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput_g65), .B1(
        SI_13_), .B2(keyinput_g19), .ZN(n9647) );
  OAI221_X1 U10901 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(keyinput_g65), .C1(
        SI_13_), .C2(keyinput_g19), .A(n9647), .ZN(n9650) );
  AOI22_X1 U10902 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput_g52), .B1(SI_25_), .B2(keyinput_g7), .ZN(n9648) );
  OAI221_X1 U10903 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput_g52), .C1(
        SI_25_), .C2(keyinput_g7), .A(n9648), .ZN(n9649) );
  NOR4_X1 U10904 ( .A1(n9652), .A2(n9651), .A3(n9650), .A4(n9649), .ZN(n9662)
         );
  AOI22_X1 U10905 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(keyinput_g68), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_g85), .ZN(n9653) );
  OAI221_X1 U10906 ( .B1(P2_DATAO_REG_28__SCAN_IN), .B2(keyinput_g68), .C1(
        P2_DATAO_REG_11__SCAN_IN), .C2(keyinput_g85), .A(n9653), .ZN(n9660) );
  AOI22_X1 U10907 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_g62), .B1(
        P1_IR_REG_23__SCAN_IN), .B2(keyinput_g114), .ZN(n9654) );
  OAI221_X1 U10908 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .C1(
        P1_IR_REG_23__SCAN_IN), .C2(keyinput_g114), .A(n9654), .ZN(n9659) );
  AOI22_X1 U10909 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput_g92), .B1(
        P1_IR_REG_17__SCAN_IN), .B2(keyinput_g108), .ZN(n9655) );
  OAI221_X1 U10910 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput_g92), .C1(
        P1_IR_REG_17__SCAN_IN), .C2(keyinput_g108), .A(n9655), .ZN(n9658) );
  AOI22_X1 U10911 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_g0), .B1(
        P2_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .ZN(n9656) );
  OAI221_X1 U10912 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_g0), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_g46), .A(n9656), .ZN(n9657) );
  NOR4_X1 U10913 ( .A1(n9660), .A2(n9659), .A3(n9658), .A4(n9657), .ZN(n9661)
         );
  NAND4_X1 U10914 ( .A1(n9664), .A2(n9663), .A3(n9662), .A4(n9661), .ZN(n9766)
         );
  INV_X1 U10915 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9666) );
  AOI22_X1 U10916 ( .A1(n5076), .A2(keyinput_g31), .B1(n9666), .B2(
        keyinput_g106), .ZN(n9665) );
  OAI221_X1 U10917 ( .B1(n5076), .B2(keyinput_g31), .C1(n9666), .C2(
        keyinput_g106), .A(n9665), .ZN(n9675) );
  INV_X1 U10918 ( .A(SI_11_), .ZN(n9847) );
  AOI22_X1 U10919 ( .A1(n6036), .A2(keyinput_g35), .B1(n9847), .B2(
        keyinput_g21), .ZN(n9667) );
  OAI221_X1 U10920 ( .B1(n6036), .B2(keyinput_g35), .C1(n9847), .C2(
        keyinput_g21), .A(n9667), .ZN(n9674) );
  AOI22_X1 U10921 ( .A1(n9669), .A2(keyinput_g22), .B1(n9899), .B2(
        keyinput_g81), .ZN(n9668) );
  OAI221_X1 U10922 ( .B1(n9669), .B2(keyinput_g22), .C1(n9899), .C2(
        keyinput_g81), .A(n9668), .ZN(n9673) );
  INV_X1 U10923 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9872) );
  XOR2_X1 U10924 ( .A(n9872), .B(keyinput_g115), .Z(n9671) );
  XNOR2_X1 U10925 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_g95), .ZN(n9670) );
  NAND2_X1 U10926 ( .A1(n9671), .A2(n9670), .ZN(n9672) );
  NOR4_X1 U10927 ( .A1(n9675), .A2(n9674), .A3(n9673), .A4(n9672), .ZN(n9713)
         );
  AOI22_X1 U10928 ( .A1(n6063), .A2(keyinput_g53), .B1(keyinput_g3), .B2(n9677), .ZN(n9676) );
  OAI221_X1 U10929 ( .B1(n6063), .B2(keyinput_g53), .C1(n9677), .C2(
        keyinput_g3), .A(n9676), .ZN(n9686) );
  AOI22_X1 U10930 ( .A1(n9908), .A2(keyinput_g91), .B1(n9932), .B2(
        keyinput_g96), .ZN(n9678) );
  OAI221_X1 U10931 ( .B1(n9908), .B2(keyinput_g91), .C1(n9932), .C2(
        keyinput_g96), .A(n9678), .ZN(n9685) );
  AOI22_X1 U10932 ( .A1(n9681), .A2(keyinput_g4), .B1(n9680), .B2(keyinput_g87), .ZN(n9679) );
  OAI221_X1 U10933 ( .B1(n9681), .B2(keyinput_g4), .C1(n9680), .C2(
        keyinput_g87), .A(n9679), .ZN(n9684) );
  INV_X1 U10934 ( .A(SI_18_), .ZN(n9943) );
  AOI22_X1 U10935 ( .A1(n9943), .A2(keyinput_g14), .B1(keyinput_g50), .B2(
        n9949), .ZN(n9682) );
  OAI221_X1 U10936 ( .B1(n9943), .B2(keyinput_g14), .C1(n9949), .C2(
        keyinput_g50), .A(n9682), .ZN(n9683) );
  NOR4_X1 U10937 ( .A1(n9686), .A2(n9685), .A3(n9684), .A4(n9683), .ZN(n9712)
         );
  AOI22_X1 U10938 ( .A1(n9688), .A2(keyinput_g123), .B1(keyinput_g10), .B2(
        n9915), .ZN(n9687) );
  OAI221_X1 U10939 ( .B1(n9688), .B2(keyinput_g123), .C1(n9915), .C2(
        keyinput_g10), .A(n9687), .ZN(n9698) );
  AOI22_X1 U10940 ( .A1(n5931), .A2(keyinput_g41), .B1(n9690), .B2(
        keyinput_g47), .ZN(n9689) );
  OAI221_X1 U10941 ( .B1(n5931), .B2(keyinput_g41), .C1(n9690), .C2(
        keyinput_g47), .A(n9689), .ZN(n9697) );
  AOI22_X1 U10942 ( .A1(n9692), .A2(keyinput_g39), .B1(n9859), .B2(
        keyinput_g71), .ZN(n9691) );
  OAI221_X1 U10943 ( .B1(n9692), .B2(keyinput_g39), .C1(n9859), .C2(
        keyinput_g71), .A(n9691), .ZN(n9696) );
  XOR2_X1 U10944 ( .A(n5332), .B(keyinput_g94), .Z(n9694) );
  XNOR2_X1 U10945 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_g99), .ZN(n9693) );
  NAND2_X1 U10946 ( .A1(n9694), .A2(n9693), .ZN(n9695) );
  NOR4_X1 U10947 ( .A1(n9698), .A2(n9697), .A3(n9696), .A4(n9695), .ZN(n9711)
         );
  INV_X1 U10948 ( .A(SI_7_), .ZN(n9855) );
  AOI22_X1 U10949 ( .A1(n9855), .A2(keyinput_g25), .B1(keyinput_g40), .B2(
        n10378), .ZN(n9699) );
  OAI221_X1 U10950 ( .B1(n9855), .B2(keyinput_g25), .C1(n10378), .C2(
        keyinput_g40), .A(n9699), .ZN(n9709) );
  INV_X1 U10951 ( .A(SI_4_), .ZN(n9917) );
  AOI22_X1 U10952 ( .A1(n6090), .A2(keyinput_g58), .B1(n9917), .B2(
        keyinput_g28), .ZN(n9700) );
  OAI221_X1 U10953 ( .B1(n6090), .B2(keyinput_g58), .C1(n9917), .C2(
        keyinput_g28), .A(n9700), .ZN(n9708) );
  AOI22_X1 U10954 ( .A1(n9703), .A2(keyinput_g82), .B1(n9702), .B2(
        keyinput_g75), .ZN(n9701) );
  OAI221_X1 U10955 ( .B1(n9703), .B2(keyinput_g82), .C1(n9702), .C2(
        keyinput_g75), .A(n9701), .ZN(n9707) );
  XNOR2_X1 U10956 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_g118), .ZN(n9705)
         );
  XNOR2_X1 U10957 ( .A(SI_5_), .B(keyinput_g27), .ZN(n9704) );
  NAND2_X1 U10958 ( .A1(n9705), .A2(n9704), .ZN(n9706) );
  NOR4_X1 U10959 ( .A1(n9709), .A2(n9708), .A3(n9707), .A4(n9706), .ZN(n9710)
         );
  NAND4_X1 U10960 ( .A1(n9713), .A2(n9712), .A3(n9711), .A4(n9710), .ZN(n9765)
         );
  AOI22_X1 U10961 ( .A1(n9854), .A2(keyinput_g124), .B1(keyinput_g121), .B2(
        n9552), .ZN(n9714) );
  OAI221_X1 U10962 ( .B1(n9854), .B2(keyinput_g124), .C1(n9552), .C2(
        keyinput_g121), .A(n9714), .ZN(n9724) );
  INV_X1 U10963 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9716) );
  AOI22_X1 U10964 ( .A1(n5220), .A2(keyinput_g120), .B1(n9716), .B2(
        keyinput_g109), .ZN(n9715) );
  OAI221_X1 U10965 ( .B1(n5220), .B2(keyinput_g120), .C1(n9716), .C2(
        keyinput_g109), .A(n9715), .ZN(n9723) );
  AOI22_X1 U10966 ( .A1(n9940), .A2(keyinput_g70), .B1(keyinput_g67), .B2(
        n9718), .ZN(n9717) );
  OAI221_X1 U10967 ( .B1(n9940), .B2(keyinput_g70), .C1(n9718), .C2(
        keyinput_g67), .A(n9717), .ZN(n9722) );
  XNOR2_X1 U10968 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_g103), .ZN(n9720)
         );
  XNOR2_X1 U10969 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_g33), .ZN(n9719) );
  NAND2_X1 U10970 ( .A1(n9720), .A2(n9719), .ZN(n9721) );
  NOR4_X1 U10971 ( .A1(n9724), .A2(n9723), .A3(n9722), .A4(n9721), .ZN(n9763)
         );
  AOI22_X1 U10972 ( .A1(n9726), .A2(keyinput_g80), .B1(n5212), .B2(
        keyinput_g117), .ZN(n9725) );
  OAI221_X1 U10973 ( .B1(n9726), .B2(keyinput_g80), .C1(n5212), .C2(
        keyinput_g117), .A(n9725), .ZN(n9735) );
  AOI22_X1 U10974 ( .A1(n9728), .A2(keyinput_g84), .B1(n5479), .B2(
        keyinput_g100), .ZN(n9727) );
  OAI221_X1 U10975 ( .B1(n9728), .B2(keyinput_g84), .C1(n5479), .C2(
        keyinput_g100), .A(n9727), .ZN(n9734) );
  XNOR2_X1 U10976 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_g79), .ZN(n9732)
         );
  XNOR2_X1 U10977 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_g122), .ZN(n9731)
         );
  XNOR2_X1 U10978 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_g119), .ZN(n9730)
         );
  XNOR2_X1 U10979 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_g78), .ZN(n9729)
         );
  NAND4_X1 U10980 ( .A1(n9732), .A2(n9731), .A3(n9730), .A4(n9729), .ZN(n9733)
         );
  NOR3_X1 U10981 ( .A1(n9735), .A2(n9734), .A3(n9733), .ZN(n9762) );
  AOI22_X1 U10982 ( .A1(n9738), .A2(keyinput_g83), .B1(keyinput_g66), .B2(
        n9737), .ZN(n9736) );
  OAI221_X1 U10983 ( .B1(n9738), .B2(keyinput_g83), .C1(n9737), .C2(
        keyinput_g66), .A(n9736), .ZN(n9746) );
  INV_X1 U10984 ( .A(SI_14_), .ZN(n9925) );
  AOI22_X1 U10985 ( .A1(n9925), .A2(keyinput_g18), .B1(keyinput_g49), .B2(
        n6914), .ZN(n9739) );
  OAI221_X1 U10986 ( .B1(n9925), .B2(keyinput_g18), .C1(n6914), .C2(
        keyinput_g49), .A(n9739), .ZN(n9745) );
  INV_X1 U10987 ( .A(SI_17_), .ZN(n9931) );
  AOI22_X1 U10988 ( .A1(n9903), .A2(keyinput_g38), .B1(n9931), .B2(
        keyinput_g15), .ZN(n9740) );
  OAI221_X1 U10989 ( .B1(n9903), .B2(keyinput_g38), .C1(n9931), .C2(
        keyinput_g15), .A(n9740), .ZN(n9744) );
  INV_X1 U10990 ( .A(SI_31_), .ZN(n9742) );
  AOI22_X1 U10991 ( .A1(n9860), .A2(keyinput_g59), .B1(keyinput_g1), .B2(n9742), .ZN(n9741) );
  OAI221_X1 U10992 ( .B1(n9860), .B2(keyinput_g59), .C1(n9742), .C2(
        keyinput_g1), .A(n9741), .ZN(n9743) );
  NOR4_X1 U10993 ( .A1(n9746), .A2(n9745), .A3(n9744), .A4(n9743), .ZN(n9761)
         );
  INV_X1 U10994 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10245) );
  AOI22_X1 U10995 ( .A1(n9748), .A2(keyinput_g77), .B1(n10245), .B2(
        keyinput_g126), .ZN(n9747) );
  OAI221_X1 U10996 ( .B1(n9748), .B2(keyinput_g77), .C1(n10245), .C2(
        keyinput_g126), .A(n9747), .ZN(n9759) );
  INV_X1 U10997 ( .A(SI_2_), .ZN(n9947) );
  AOI22_X1 U10998 ( .A1(n9947), .A2(keyinput_g30), .B1(n9750), .B2(
        keyinput_g86), .ZN(n9749) );
  OAI221_X1 U10999 ( .B1(n9947), .B2(keyinput_g30), .C1(n9750), .C2(
        keyinput_g86), .A(n9749), .ZN(n9758) );
  AOI22_X1 U11000 ( .A1(n9753), .A2(keyinput_g5), .B1(keyinput_g54), .B2(n9752), .ZN(n9751) );
  OAI221_X1 U11001 ( .B1(n9753), .B2(keyinput_g5), .C1(n9752), .C2(
        keyinput_g54), .A(n9751), .ZN(n9757) );
  AOI22_X1 U11002 ( .A1(n9755), .A2(keyinput_g90), .B1(keyinput_g44), .B2(
        n9841), .ZN(n9754) );
  OAI221_X1 U11003 ( .B1(n9755), .B2(keyinput_g90), .C1(n9841), .C2(
        keyinput_g44), .A(n9754), .ZN(n9756) );
  NOR4_X1 U11004 ( .A1(n9759), .A2(n9758), .A3(n9757), .A4(n9756), .ZN(n9760)
         );
  NAND4_X1 U11005 ( .A1(n9763), .A2(n9762), .A3(n9761), .A4(n9760), .ZN(n9764)
         );
  NOR4_X1 U11006 ( .A1(n9767), .A2(n9766), .A3(n9765), .A4(n9764), .ZN(n9967)
         );
  XOR2_X1 U11007 ( .A(SI_27_), .B(keyinput_f5), .Z(n9774) );
  AOI22_X1 U11008 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_f47), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(keyinput_f83), .ZN(n9768) );
  OAI221_X1 U11009 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .C1(
        P2_DATAO_REG_13__SCAN_IN), .C2(keyinput_f83), .A(n9768), .ZN(n9773) );
  AOI22_X1 U11010 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput_f87), .B1(
        P1_IR_REG_20__SCAN_IN), .B2(keyinput_f111), .ZN(n9769) );
  OAI221_X1 U11011 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput_f87), .C1(
        P1_IR_REG_20__SCAN_IN), .C2(keyinput_f111), .A(n9769), .ZN(n9772) );
  AOI22_X1 U11012 ( .A1(SI_28_), .A2(keyinput_f4), .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_f88), .ZN(n9770) );
  OAI221_X1 U11013 ( .B1(SI_28_), .B2(keyinput_f4), .C1(
        P2_DATAO_REG_8__SCAN_IN), .C2(keyinput_f88), .A(n9770), .ZN(n9771) );
  NOR4_X1 U11014 ( .A1(n9774), .A2(n9773), .A3(n9772), .A4(n9771), .ZN(n9802)
         );
  AOI22_X1 U11015 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput_f33), .B1(
        P1_IR_REG_10__SCAN_IN), .B2(keyinput_f101), .ZN(n9775) );
  OAI221_X1 U11016 ( .B1(P2_RD_REG_SCAN_IN), .B2(keyinput_f33), .C1(
        P1_IR_REG_10__SCAN_IN), .C2(keyinput_f101), .A(n9775), .ZN(n9782) );
  AOI22_X1 U11017 ( .A1(SI_3_), .A2(keyinput_f29), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(keyinput_f84), .ZN(n9776) );
  OAI221_X1 U11018 ( .B1(SI_3_), .B2(keyinput_f29), .C1(
        P2_DATAO_REG_12__SCAN_IN), .C2(keyinput_f84), .A(n9776), .ZN(n9781) );
  AOI22_X1 U11019 ( .A1(SI_29_), .A2(keyinput_f3), .B1(SI_0_), .B2(
        keyinput_f32), .ZN(n9777) );
  OAI221_X1 U11020 ( .B1(SI_29_), .B2(keyinput_f3), .C1(SI_0_), .C2(
        keyinput_f32), .A(n9777), .ZN(n9780) );
  AOI22_X1 U11021 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(keyinput_f77), .B1(
        SI_20_), .B2(keyinput_f12), .ZN(n9778) );
  OAI221_X1 U11022 ( .B1(P2_DATAO_REG_19__SCAN_IN), .B2(keyinput_f77), .C1(
        SI_20_), .C2(keyinput_f12), .A(n9778), .ZN(n9779) );
  NOR4_X1 U11023 ( .A1(n9782), .A2(n9781), .A3(n9780), .A4(n9779), .ZN(n9801)
         );
  AOI22_X1 U11024 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput_f63), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .ZN(n9783) );
  OAI221_X1 U11025 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_f62), .A(n9783), .ZN(n9790) );
  AOI22_X1 U11026 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(keyinput_f86), .B1(
        SI_13_), .B2(keyinput_f19), .ZN(n9784) );
  OAI221_X1 U11027 ( .B1(P2_DATAO_REG_10__SCAN_IN), .B2(keyinput_f86), .C1(
        SI_13_), .C2(keyinput_f19), .A(n9784), .ZN(n9789) );
  AOI22_X1 U11028 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput_f104), .B1(
        P1_IR_REG_18__SCAN_IN), .B2(keyinput_f109), .ZN(n9785) );
  OAI221_X1 U11029 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput_f104), .C1(
        P1_IR_REG_18__SCAN_IN), .C2(keyinput_f109), .A(n9785), .ZN(n9788) );
  AOI22_X1 U11030 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(keyinput_f73), .B1(
        P1_IR_REG_27__SCAN_IN), .B2(keyinput_f118), .ZN(n9786) );
  OAI221_X1 U11031 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(keyinput_f73), .C1(
        P1_IR_REG_27__SCAN_IN), .C2(keyinput_f118), .A(n9786), .ZN(n9787) );
  NOR4_X1 U11032 ( .A1(n9790), .A2(n9789), .A3(n9788), .A4(n9787), .ZN(n9800)
         );
  AOI22_X1 U11033 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(keyinput_f76), .B1(
        P1_IR_REG_12__SCAN_IN), .B2(keyinput_f103), .ZN(n9791) );
  OAI221_X1 U11034 ( .B1(P2_DATAO_REG_20__SCAN_IN), .B2(keyinput_f76), .C1(
        P1_IR_REG_12__SCAN_IN), .C2(keyinput_f103), .A(n9791), .ZN(n9798) );
  AOI22_X1 U11035 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(keyinput_f93), .B1(
        P1_IR_REG_16__SCAN_IN), .B2(keyinput_f107), .ZN(n9792) );
  OAI221_X1 U11036 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(keyinput_f93), .C1(
        P1_IR_REG_16__SCAN_IN), .C2(keyinput_f107), .A(n9792), .ZN(n9797) );
  AOI22_X1 U11037 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(keyinput_f120), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_f79), .ZN(n9793) );
  OAI221_X1 U11038 ( .B1(P1_IR_REG_29__SCAN_IN), .B2(keyinput_f120), .C1(
        P2_DATAO_REG_17__SCAN_IN), .C2(keyinput_f79), .A(n9793), .ZN(n9796) );
  AOI22_X1 U11039 ( .A1(SI_10_), .A2(keyinput_f22), .B1(P1_D_REG_0__SCAN_IN), 
        .B2(keyinput_f123), .ZN(n9794) );
  OAI221_X1 U11040 ( .B1(SI_10_), .B2(keyinput_f22), .C1(P1_D_REG_0__SCAN_IN), 
        .C2(keyinput_f123), .A(n9794), .ZN(n9795) );
  NOR4_X1 U11041 ( .A1(n9798), .A2(n9797), .A3(n9796), .A4(n9795), .ZN(n9799)
         );
  NAND4_X1 U11042 ( .A1(n9802), .A2(n9801), .A3(n9800), .A4(n9799), .ZN(n9961)
         );
  AOI22_X1 U11043 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_f45), .B1(
        P2_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .ZN(n9803) );
  OAI221_X1 U11044 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_f45), .C1(
        P2_REG3_REG_24__SCAN_IN), .C2(keyinput_f51), .A(n9803), .ZN(n9810) );
  AOI22_X1 U11045 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(keyinput_f67), .B1(
        P2_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .ZN(n9804) );
  OAI221_X1 U11046 ( .B1(P2_DATAO_REG_29__SCAN_IN), .B2(keyinput_f67), .C1(
        P2_REG3_REG_10__SCAN_IN), .C2(keyinput_f39), .A(n9804), .ZN(n9809) );
  AOI22_X1 U11047 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_f42), .B1(
        SI_26_), .B2(keyinput_f6), .ZN(n9805) );
  OAI221_X1 U11048 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .C1(
        SI_26_), .C2(keyinput_f6), .A(n9805), .ZN(n9808) );
  AOI22_X1 U11049 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_f46), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .ZN(n9806) );
  OAI221_X1 U11050 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n9806), .ZN(n9807) );
  NOR4_X1 U11051 ( .A1(n9810), .A2(n9809), .A3(n9808), .A4(n9807), .ZN(n9838)
         );
  AOI22_X1 U11052 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput_f65), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(keyinput_f80), .ZN(n9811) );
  OAI221_X1 U11053 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(keyinput_f65), .C1(
        P2_DATAO_REG_16__SCAN_IN), .C2(keyinput_f80), .A(n9811), .ZN(n9818) );
  AOI22_X1 U11054 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_f58), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(keyinput_f78), .ZN(n9812) );
  OAI221_X1 U11055 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .C1(
        P2_DATAO_REG_18__SCAN_IN), .C2(keyinput_f78), .A(n9812), .ZN(n9817) );
  AOI22_X1 U11056 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(keyinput_f82), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_f75), .ZN(n9813) );
  OAI221_X1 U11057 ( .B1(P2_DATAO_REG_14__SCAN_IN), .B2(keyinput_f82), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput_f75), .A(n9813), .ZN(n9816) );
  AOI22_X1 U11058 ( .A1(SI_6_), .A2(keyinput_f26), .B1(P1_IR_REG_9__SCAN_IN), 
        .B2(keyinput_f100), .ZN(n9814) );
  OAI221_X1 U11059 ( .B1(SI_6_), .B2(keyinput_f26), .C1(P1_IR_REG_9__SCAN_IN), 
        .C2(keyinput_f100), .A(n9814), .ZN(n9815) );
  NOR4_X1 U11060 ( .A1(n9818), .A2(n9817), .A3(n9816), .A4(n9815), .ZN(n9837)
         );
  AOI22_X1 U11061 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(keyinput_f74), .B1(
        P1_IR_REG_7__SCAN_IN), .B2(keyinput_f98), .ZN(n9819) );
  OAI221_X1 U11062 ( .B1(P2_DATAO_REG_22__SCAN_IN), .B2(keyinput_f74), .C1(
        P1_IR_REG_7__SCAN_IN), .C2(keyinput_f98), .A(n9819), .ZN(n9826) );
  AOI22_X1 U11063 ( .A1(SI_19_), .A2(keyinput_f13), .B1(P1_IR_REG_1__SCAN_IN), 
        .B2(keyinput_f92), .ZN(n9820) );
  OAI221_X1 U11064 ( .B1(SI_19_), .B2(keyinput_f13), .C1(P1_IR_REG_1__SCAN_IN), 
        .C2(keyinput_f92), .A(n9820), .ZN(n9825) );
  AOI22_X1 U11065 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(keyinput_f121), .B1(
        P1_IR_REG_14__SCAN_IN), .B2(keyinput_f105), .ZN(n9821) );
  OAI221_X1 U11066 ( .B1(P1_IR_REG_30__SCAN_IN), .B2(keyinput_f121), .C1(
        P1_IR_REG_14__SCAN_IN), .C2(keyinput_f105), .A(n9821), .ZN(n9824) );
  AOI22_X1 U11067 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(keyinput_f66), .B1(
        P1_IR_REG_4__SCAN_IN), .B2(keyinput_f95), .ZN(n9822) );
  OAI221_X1 U11068 ( .B1(P2_DATAO_REG_30__SCAN_IN), .B2(keyinput_f66), .C1(
        P1_IR_REG_4__SCAN_IN), .C2(keyinput_f95), .A(n9822), .ZN(n9823) );
  NOR4_X1 U11069 ( .A1(n9826), .A2(n9825), .A3(n9824), .A4(n9823), .ZN(n9836)
         );
  AOI22_X1 U11070 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(keyinput_f89), .B1(
        P1_IR_REG_11__SCAN_IN), .B2(keyinput_f102), .ZN(n9827) );
  OAI221_X1 U11071 ( .B1(P2_DATAO_REG_7__SCAN_IN), .B2(keyinput_f89), .C1(
        P1_IR_REG_11__SCAN_IN), .C2(keyinput_f102), .A(n9827), .ZN(n9834) );
  AOI22_X1 U11072 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_f54), .B1(
        P2_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .ZN(n9828) );
  OAI221_X1 U11073 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_f54), .C1(
        P2_REG3_REG_9__SCAN_IN), .C2(keyinput_f53), .A(n9828), .ZN(n9833) );
  AOI22_X1 U11074 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(keyinput_f35), .B1(
        P1_IR_REG_15__SCAN_IN), .B2(keyinput_f106), .ZN(n9829) );
  OAI221_X1 U11075 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_f35), .C1(
        P1_IR_REG_15__SCAN_IN), .C2(keyinput_f106), .A(n9829), .ZN(n9832) );
  AOI22_X1 U11076 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(keyinput_f113), .B1(n6121), 
        .B2(keyinput_f56), .ZN(n9830) );
  OAI221_X1 U11077 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(keyinput_f113), .C1(n6121), .C2(keyinput_f56), .A(n9830), .ZN(n9831) );
  NOR4_X1 U11078 ( .A1(n9834), .A2(n9833), .A3(n9832), .A4(n9831), .ZN(n9835)
         );
  NAND4_X1 U11079 ( .A1(n9838), .A2(n9837), .A3(n9836), .A4(n9835), .ZN(n9960)
         );
  AOI22_X1 U11080 ( .A1(n5931), .A2(keyinput_f41), .B1(n5076), .B2(
        keyinput_f31), .ZN(n9839) );
  OAI221_X1 U11081 ( .B1(n5931), .B2(keyinput_f41), .C1(n5076), .C2(
        keyinput_f31), .A(n9839), .ZN(n9852) );
  AOI22_X1 U11082 ( .A1(n9842), .A2(keyinput_f43), .B1(keyinput_f44), .B2(
        n9841), .ZN(n9840) );
  OAI221_X1 U11083 ( .B1(n9842), .B2(keyinput_f43), .C1(n9841), .C2(
        keyinput_f44), .A(n9840), .ZN(n9851) );
  INV_X1 U11084 ( .A(SI_30_), .ZN(n9845) );
  AOI22_X1 U11085 ( .A1(n9845), .A2(keyinput_f2), .B1(n9844), .B2(keyinput_f24), .ZN(n9843) );
  OAI221_X1 U11086 ( .B1(n9845), .B2(keyinput_f2), .C1(n9844), .C2(
        keyinput_f24), .A(n9843), .ZN(n9850) );
  AOI22_X1 U11087 ( .A1(n9848), .A2(keyinput_f61), .B1(n9847), .B2(
        keyinput_f21), .ZN(n9846) );
  OAI221_X1 U11088 ( .B1(n9848), .B2(keyinput_f61), .C1(n9847), .C2(
        keyinput_f21), .A(n9846), .ZN(n9849) );
  NOR4_X1 U11089 ( .A1(n9852), .A2(n9851), .A3(n9850), .A4(n9849), .ZN(n9897)
         );
  AOI22_X1 U11090 ( .A1(n9855), .A2(keyinput_f25), .B1(n9854), .B2(
        keyinput_f124), .ZN(n9853) );
  OAI221_X1 U11091 ( .B1(n9855), .B2(keyinput_f25), .C1(n9854), .C2(
        keyinput_f124), .A(n9853), .ZN(n9866) );
  AOI22_X1 U11092 ( .A1(n5240), .A2(keyinput_f110), .B1(keyinput_f7), .B2(
        n9857), .ZN(n9856) );
  OAI221_X1 U11093 ( .B1(n5240), .B2(keyinput_f110), .C1(n9857), .C2(
        keyinput_f7), .A(n9856), .ZN(n9865) );
  AOI22_X1 U11094 ( .A1(n9860), .A2(keyinput_f59), .B1(n9859), .B2(
        keyinput_f71), .ZN(n9858) );
  OAI221_X1 U11095 ( .B1(n9860), .B2(keyinput_f59), .C1(n9859), .C2(
        keyinput_f71), .A(n9858), .ZN(n9864) );
  XNOR2_X1 U11096 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_f97), .ZN(n9862) );
  XNOR2_X1 U11097 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput_f34), .ZN(n9861) );
  NAND2_X1 U11098 ( .A1(n9862), .A2(n9861), .ZN(n9863) );
  NOR4_X1 U11099 ( .A1(n9866), .A2(n9865), .A3(n9864), .A4(n9863), .ZN(n9896)
         );
  AOI22_X1 U11100 ( .A1(n9869), .A2(keyinput_f64), .B1(n9868), .B2(
        keyinput_f20), .ZN(n9867) );
  OAI221_X1 U11101 ( .B1(n9869), .B2(keyinput_f64), .C1(n9868), .C2(
        keyinput_f20), .A(n9867), .ZN(n9882) );
  AOI22_X1 U11102 ( .A1(n9872), .A2(keyinput_f115), .B1(keyinput_f60), .B2(
        n9871), .ZN(n9870) );
  OAI221_X1 U11103 ( .B1(n9872), .B2(keyinput_f115), .C1(n9871), .C2(
        keyinput_f60), .A(n9870), .ZN(n9881) );
  INV_X1 U11104 ( .A(P2_WR_REG_SCAN_IN), .ZN(n9874) );
  AOI22_X1 U11105 ( .A1(n9875), .A2(keyinput_f16), .B1(keyinput_f0), .B2(n9874), .ZN(n9873) );
  OAI221_X1 U11106 ( .B1(n9875), .B2(keyinput_f16), .C1(n9874), .C2(
        keyinput_f0), .A(n9873), .ZN(n9880) );
  AOI22_X1 U11107 ( .A1(n9878), .A2(keyinput_f68), .B1(n9877), .B2(
        keyinput_f11), .ZN(n9876) );
  OAI221_X1 U11108 ( .B1(n9878), .B2(keyinput_f68), .C1(n9877), .C2(
        keyinput_f11), .A(n9876), .ZN(n9879) );
  NOR4_X1 U11109 ( .A1(n9882), .A2(n9881), .A3(n9880), .A4(n9879), .ZN(n9895)
         );
  AOI22_X1 U11110 ( .A1(n9884), .A2(keyinput_f9), .B1(n5839), .B2(
        keyinput_f114), .ZN(n9883) );
  OAI221_X1 U11111 ( .B1(n9884), .B2(keyinput_f9), .C1(n5839), .C2(
        keyinput_f114), .A(n9883), .ZN(n9893) );
  XNOR2_X1 U11112 ( .A(n9885), .B(keyinput_f119), .ZN(n9892) );
  XNOR2_X1 U11113 ( .A(keyinput_f117), .B(n5212), .ZN(n9891) );
  XNOR2_X1 U11114 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_f57), .ZN(n9889)
         );
  XNOR2_X1 U11115 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_f99), .ZN(n9888) );
  XNOR2_X1 U11116 ( .A(SI_31_), .B(keyinput_f1), .ZN(n9887) );
  XNOR2_X1 U11117 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_f122), .ZN(n9886)
         );
  NAND4_X1 U11118 ( .A1(n9889), .A2(n9888), .A3(n9887), .A4(n9886), .ZN(n9890)
         );
  NOR4_X1 U11119 ( .A1(n9893), .A2(n9892), .A3(n9891), .A4(n9890), .ZN(n9894)
         );
  NAND4_X1 U11120 ( .A1(n9897), .A2(n9896), .A3(n9895), .A4(n9894), .ZN(n9959)
         );
  AOI22_X1 U11121 ( .A1(n9900), .A2(keyinput_f55), .B1(n9899), .B2(
        keyinput_f81), .ZN(n9898) );
  OAI221_X1 U11122 ( .B1(n9900), .B2(keyinput_f55), .C1(n9899), .C2(
        keyinput_f81), .A(n9898), .ZN(n9912) );
  AOI22_X1 U11123 ( .A1(n9903), .A2(keyinput_f38), .B1(keyinput_f52), .B2(
        n9902), .ZN(n9901) );
  OAI221_X1 U11124 ( .B1(n9903), .B2(keyinput_f38), .C1(n9902), .C2(
        keyinput_f52), .A(n9901), .ZN(n9911) );
  AOI22_X1 U11125 ( .A1(n6914), .A2(keyinput_f49), .B1(n9905), .B2(
        keyinput_f23), .ZN(n9904) );
  OAI221_X1 U11126 ( .B1(n6914), .B2(keyinput_f49), .C1(n9905), .C2(
        keyinput_f23), .A(n9904), .ZN(n9910) );
  AOI22_X1 U11127 ( .A1(n9908), .A2(keyinput_f91), .B1(n9907), .B2(
        keyinput_f108), .ZN(n9906) );
  OAI221_X1 U11128 ( .B1(n9908), .B2(keyinput_f91), .C1(n9907), .C2(
        keyinput_f108), .A(n9906), .ZN(n9909) );
  NOR4_X1 U11129 ( .A1(n9912), .A2(n9911), .A3(n9910), .A4(n9909), .ZN(n9957)
         );
  INV_X1 U11130 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10244) );
  AOI22_X1 U11131 ( .A1(n10244), .A2(keyinput_f127), .B1(keyinput_f40), .B2(
        n10378), .ZN(n9913) );
  OAI221_X1 U11132 ( .B1(n10244), .B2(keyinput_f127), .C1(n10378), .C2(
        keyinput_f40), .A(n9913), .ZN(n9923) );
  AOI22_X1 U11133 ( .A1(n10245), .A2(keyinput_f126), .B1(keyinput_f10), .B2(
        n9915), .ZN(n9914) );
  OAI221_X1 U11134 ( .B1(n10245), .B2(keyinput_f126), .C1(n9915), .C2(
        keyinput_f10), .A(n9914), .ZN(n9922) );
  AOI22_X1 U11135 ( .A1(n5167), .A2(keyinput_f8), .B1(keyinput_f28), .B2(n9917), .ZN(n9916) );
  OAI221_X1 U11136 ( .B1(n5167), .B2(keyinput_f8), .C1(n9917), .C2(
        keyinput_f28), .A(n9916), .ZN(n9921) );
  XNOR2_X1 U11137 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_f116), .ZN(n9919)
         );
  XNOR2_X1 U11138 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput_f90), .ZN(n9918)
         );
  NAND2_X1 U11139 ( .A1(n9919), .A2(n9918), .ZN(n9920) );
  NOR4_X1 U11140 ( .A1(n9923), .A2(n9922), .A3(n9921), .A4(n9920), .ZN(n9956)
         );
  AOI22_X1 U11141 ( .A1(n9926), .A2(keyinput_f48), .B1(n9925), .B2(
        keyinput_f18), .ZN(n9924) );
  OAI221_X1 U11142 ( .B1(n9926), .B2(keyinput_f48), .C1(n9925), .C2(
        keyinput_f18), .A(n9924), .ZN(n9938) );
  AOI22_X1 U11143 ( .A1(n9929), .A2(keyinput_f37), .B1(n9928), .B2(
        keyinput_f72), .ZN(n9927) );
  OAI221_X1 U11144 ( .B1(n9929), .B2(keyinput_f37), .C1(n9928), .C2(
        keyinput_f72), .A(n9927), .ZN(n9937) );
  AOI22_X1 U11145 ( .A1(n9932), .A2(keyinput_f96), .B1(keyinput_f15), .B2(
        n9931), .ZN(n9930) );
  OAI221_X1 U11146 ( .B1(n9932), .B2(keyinput_f96), .C1(n9931), .C2(
        keyinput_f15), .A(n9930), .ZN(n9936) );
  AOI22_X1 U11147 ( .A1(n5332), .A2(keyinput_f94), .B1(keyinput_f85), .B2(
        n9934), .ZN(n9933) );
  OAI221_X1 U11148 ( .B1(n5332), .B2(keyinput_f94), .C1(n9934), .C2(
        keyinput_f85), .A(n9933), .ZN(n9935) );
  NOR4_X1 U11149 ( .A1(n9938), .A2(n9937), .A3(n9936), .A4(n9935), .ZN(n9955)
         );
  AOI22_X1 U11150 ( .A1(n9941), .A2(keyinput_f17), .B1(n9940), .B2(
        keyinput_f70), .ZN(n9939) );
  OAI221_X1 U11151 ( .B1(n9941), .B2(keyinput_f17), .C1(n9940), .C2(
        keyinput_f70), .A(n9939), .ZN(n9953) );
  AOI22_X1 U11152 ( .A1(n9944), .A2(keyinput_f27), .B1(n9943), .B2(
        keyinput_f14), .ZN(n9942) );
  OAI221_X1 U11153 ( .B1(n9944), .B2(keyinput_f27), .C1(n9943), .C2(
        keyinput_f14), .A(n9942), .ZN(n9952) );
  AOI22_X1 U11154 ( .A1(n9947), .A2(keyinput_f30), .B1(n9946), .B2(
        keyinput_f69), .ZN(n9945) );
  OAI221_X1 U11155 ( .B1(n9947), .B2(keyinput_f30), .C1(n9946), .C2(
        keyinput_f69), .A(n9945), .ZN(n9951) );
  AOI22_X1 U11156 ( .A1(n5232), .A2(keyinput_f112), .B1(keyinput_f50), .B2(
        n9949), .ZN(n9948) );
  OAI221_X1 U11157 ( .B1(n5232), .B2(keyinput_f112), .C1(n9949), .C2(
        keyinput_f50), .A(n9948), .ZN(n9950) );
  NOR4_X1 U11158 ( .A1(n9953), .A2(n9952), .A3(n9951), .A4(n9950), .ZN(n9954)
         );
  NAND4_X1 U11159 ( .A1(n9957), .A2(n9956), .A3(n9955), .A4(n9954), .ZN(n9958)
         );
  OR4_X1 U11160 ( .A1(n9961), .A2(n9960), .A3(n9959), .A4(n9958), .ZN(n9963)
         );
  AOI21_X1 U11161 ( .B1(keyinput_f125), .B2(n9963), .A(keyinput_g125), .ZN(
        n9965) );
  INV_X1 U11162 ( .A(keyinput_f125), .ZN(n9962) );
  AOI21_X1 U11163 ( .B1(n9963), .B2(n9962), .A(P1_D_REG_2__SCAN_IN), .ZN(n9964) );
  AOI22_X1 U11164 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9965), .B1(keyinput_g125), 
        .B2(n9964), .ZN(n9966) );
  AOI21_X1 U11165 ( .B1(n9968), .B2(n9967), .A(n9966), .ZN(n9969) );
  XNOR2_X1 U11166 ( .A(n9970), .B(n9969), .ZN(n9974) );
  NOR2_X1 U11167 ( .A1(n9972), .A2(n9971), .ZN(n9973) );
  XOR2_X1 U11168 ( .A(n9974), .B(n9973), .Z(ADD_1071_U4) );
  NAND2_X1 U11169 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9976) );
  AOI21_X1 U11170 ( .B1(n9977), .B2(n9976), .A(n9975), .ZN(n9978) );
  NAND2_X1 U11171 ( .A1(n10331), .A2(n9978), .ZN(n9980) );
  AOI22_X1 U11172 ( .A1(n10333), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n9979) );
  OAI211_X1 U11173 ( .C1(n10327), .C2(n9981), .A(n9980), .B(n9979), .ZN(n9982)
         );
  INV_X1 U11174 ( .A(n9982), .ZN(n9987) );
  NOR2_X1 U11175 ( .A1(n10335), .A2(n5952), .ZN(n9985) );
  OAI211_X1 U11176 ( .C1(n9985), .C2(n9984), .A(n10330), .B(n9983), .ZN(n9986)
         );
  NAND2_X1 U11177 ( .A1(n9987), .A2(n9986), .ZN(P2_U3246) );
  AOI22_X1 U11178 ( .A1(n10333), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n10000) );
  AOI211_X1 U11179 ( .C1(n9991), .C2(n9990), .A(n9989), .B(n9988), .ZN(n9992)
         );
  AOI21_X1 U11180 ( .B1(n9994), .B2(n9993), .A(n9992), .ZN(n9999) );
  OAI211_X1 U11181 ( .C1(n9997), .C2(n9996), .A(n10330), .B(n9995), .ZN(n9998)
         );
  NAND3_X1 U11182 ( .A1(n10000), .A2(n9999), .A3(n9998), .ZN(P2_U3247) );
  OAI21_X1 U11183 ( .B1(n10002), .B2(n10304), .A(n10001), .ZN(n10003) );
  AOI21_X1 U11184 ( .B1(n10004), .B2(n10309), .A(n10003), .ZN(n10005) );
  AND2_X1 U11185 ( .A1(n10006), .A2(n10005), .ZN(n10008) );
  INV_X1 U11186 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10007) );
  AOI22_X1 U11187 ( .A1(n10315), .A2(n10008), .B1(n10007), .B2(n10313), .ZN(
        P1_U3484) );
  AOI22_X1 U11188 ( .A1(n10326), .A2(n10008), .B1(n6831), .B2(n10324), .ZN(
        P1_U3533) );
  AOI21_X1 U11189 ( .B1(n10012), .B2(n10010), .A(n10009), .ZN(n10037) );
  XOR2_X1 U11190 ( .A(n10012), .B(n10011), .Z(n10016) );
  AOI22_X1 U11191 ( .A1(n10014), .A2(n10226), .B1(n10223), .B2(n10013), .ZN(
        n10015) );
  OAI21_X1 U11192 ( .B1(n10016), .B2(n10228), .A(n10015), .ZN(n10017) );
  AOI21_X1 U11193 ( .B1(n10037), .B2(n10184), .A(n10017), .ZN(n10034) );
  INV_X1 U11194 ( .A(n10018), .ZN(n10019) );
  AOI222_X1 U11195 ( .A1(n10020), .A2(n10187), .B1(n10019), .B2(n10203), .C1(
        P1_REG2_REG_12__SCAN_IN), .C2(n10215), .ZN(n10026) );
  OAI211_X1 U11196 ( .C1(n10022), .C2(n10033), .A(n10198), .B(n10021), .ZN(
        n10032) );
  INV_X1 U11197 ( .A(n10032), .ZN(n10023) );
  AOI22_X1 U11198 ( .A1(n10037), .A2(n10222), .B1(n10024), .B2(n10023), .ZN(
        n10025) );
  OAI211_X1 U11199 ( .C1(n10215), .C2(n10034), .A(n10026), .B(n10025), .ZN(
        P1_U3279) );
  OAI211_X1 U11200 ( .C1(n10029), .C2(n10304), .A(n10028), .B(n10027), .ZN(
        n10030) );
  AOI21_X1 U11201 ( .B1(n10031), .B2(n10295), .A(n10030), .ZN(n10039) );
  AOI22_X1 U11202 ( .A1(n10326), .A2(n10039), .B1(n5570), .B2(n10324), .ZN(
        P1_U3537) );
  OAI21_X1 U11203 ( .B1(n10033), .B2(n10304), .A(n10032), .ZN(n10036) );
  INV_X1 U11204 ( .A(n10034), .ZN(n10035) );
  AOI211_X1 U11205 ( .C1(n10309), .C2(n10037), .A(n10036), .B(n10035), .ZN(
        n10041) );
  AOI22_X1 U11206 ( .A1(n10326), .A2(n10041), .B1(n5529), .B2(n10324), .ZN(
        P1_U3535) );
  INV_X1 U11207 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10038) );
  AOI22_X1 U11208 ( .A1(n10315), .A2(n10039), .B1(n10038), .B2(n10313), .ZN(
        P1_U3496) );
  INV_X1 U11209 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10040) );
  AOI22_X1 U11210 ( .A1(n10315), .A2(n10041), .B1(n10040), .B2(n10313), .ZN(
        P1_U3490) );
  XNOR2_X1 U11211 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X1 U11212 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10064) );
  INV_X1 U11213 ( .A(n10042), .ZN(n10045) );
  AOI211_X1 U11214 ( .C1(n10045), .C2(n10044), .A(n10043), .B(n10159), .ZN(
        n10061) );
  INV_X1 U11215 ( .A(n10046), .ZN(n10047) );
  MUX2_X1 U11216 ( .A(n10048), .B(n10047), .S(n6468), .Z(n10050) );
  NAND2_X1 U11217 ( .A1(n10050), .A2(n10049), .ZN(n10051) );
  OAI211_X1 U11218 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n10052), .A(n10051), .B(
        P1_U4006), .ZN(n10076) );
  MUX2_X1 U11219 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10054), .S(n10053), .Z(
        n10057) );
  OAI211_X1 U11220 ( .C1(n10057), .C2(n4580), .A(n10147), .B(n10056), .ZN(
        n10058) );
  OAI211_X1 U11221 ( .C1(n10163), .C2(n10059), .A(n10076), .B(n10058), .ZN(
        n10060) );
  AOI211_X1 U11222 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(P1_U3084), .A(n10061), 
        .B(n10060), .ZN(n10063) );
  OAI21_X1 U11223 ( .B1(n10172), .B2(n10064), .A(n10063), .ZN(P1_U3243) );
  OAI21_X1 U11224 ( .B1(n10067), .B2(n4724), .A(n10066), .ZN(n10068) );
  AOI22_X1 U11225 ( .A1(n10069), .A2(n10129), .B1(n10086), .B2(n10068), .ZN(
        n10078) );
  AOI21_X1 U11226 ( .B1(n10072), .B2(n10071), .A(n10070), .ZN(n10073) );
  NOR2_X1 U11227 ( .A1(n10169), .A2(n10073), .ZN(n10074) );
  AOI211_X1 U11228 ( .C1(P1_ADDR_REG_4__SCAN_IN), .C2(n10079), .A(n10075), .B(
        n10074), .ZN(n10077) );
  NAND3_X1 U11229 ( .A1(n10078), .A2(n10077), .A3(n10076), .ZN(P1_U3245) );
  AOI22_X1 U11230 ( .A1(n10129), .A2(n10080), .B1(n10079), .B2(
        P1_ADDR_REG_8__SCAN_IN), .ZN(n10093) );
  INV_X1 U11231 ( .A(n10081), .ZN(n10092) );
  OAI21_X1 U11232 ( .B1(n10084), .B2(n10083), .A(n10082), .ZN(n10085) );
  NAND2_X1 U11233 ( .A1(n10086), .A2(n10085), .ZN(n10091) );
  OAI211_X1 U11234 ( .C1(n10089), .C2(n10088), .A(n10147), .B(n10087), .ZN(
        n10090) );
  NAND4_X1 U11235 ( .A1(n10093), .A2(n10092), .A3(n10091), .A4(n10090), .ZN(
        P1_U3249) );
  INV_X1 U11236 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10112) );
  INV_X1 U11237 ( .A(n10094), .ZN(n10097) );
  INV_X1 U11238 ( .A(n10095), .ZN(n10096) );
  NAND2_X1 U11239 ( .A1(n10097), .A2(n10096), .ZN(n10098) );
  NAND2_X1 U11240 ( .A1(n10099), .A2(n10098), .ZN(n10100) );
  OR2_X1 U11241 ( .A1(n10159), .A2(n10100), .ZN(n10103) );
  INV_X1 U11242 ( .A(n10101), .ZN(n10102) );
  OAI211_X1 U11243 ( .C1(n10163), .C2(n10104), .A(n10103), .B(n10102), .ZN(
        n10105) );
  INV_X1 U11244 ( .A(n10105), .ZN(n10111) );
  AOI21_X1 U11245 ( .B1(n10108), .B2(n10107), .A(n10106), .ZN(n10109) );
  OR2_X1 U11246 ( .A1(n10109), .A2(n10169), .ZN(n10110) );
  OAI211_X1 U11247 ( .C1(n10112), .C2(n10172), .A(n10111), .B(n10110), .ZN(
        P1_U3254) );
  INV_X1 U11248 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10122) );
  AOI211_X1 U11249 ( .C1(n10114), .C2(n7751), .A(n10113), .B(n10159), .ZN(
        n10115) );
  AOI211_X1 U11250 ( .C1(n10129), .C2(n10117), .A(n10116), .B(n10115), .ZN(
        n10121) );
  OAI211_X1 U11251 ( .C1(n10119), .C2(P1_REG1_REG_15__SCAN_IN), .A(n10147), 
        .B(n10118), .ZN(n10120) );
  OAI211_X1 U11252 ( .C1(n10122), .C2(n10172), .A(n10121), .B(n10120), .ZN(
        P1_U3256) );
  INV_X1 U11253 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10135) );
  AOI211_X1 U11254 ( .C1(n10125), .C2(n10124), .A(n10123), .B(n10159), .ZN(
        n10126) );
  AOI211_X1 U11255 ( .C1(n10129), .C2(n10128), .A(n10127), .B(n10126), .ZN(
        n10134) );
  OAI211_X1 U11256 ( .C1(n10132), .C2(n10131), .A(n10147), .B(n10130), .ZN(
        n10133) );
  OAI211_X1 U11257 ( .C1(n10135), .C2(n10172), .A(n10134), .B(n10133), .ZN(
        P1_U3257) );
  INV_X1 U11258 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10152) );
  NAND2_X1 U11259 ( .A1(n10137), .A2(n10136), .ZN(n10140) );
  INV_X1 U11260 ( .A(n10138), .ZN(n10139) );
  NAND2_X1 U11261 ( .A1(n10140), .A2(n10139), .ZN(n10141) );
  OAI211_X1 U11262 ( .C1(n10163), .C2(n10144), .A(n10143), .B(n10142), .ZN(
        n10145) );
  INV_X1 U11263 ( .A(n10145), .ZN(n10151) );
  OAI211_X1 U11264 ( .C1(n10149), .C2(n10148), .A(n10147), .B(n10146), .ZN(
        n10150) );
  OAI211_X1 U11265 ( .C1(n10152), .C2(n10172), .A(n10151), .B(n10150), .ZN(
        P1_U3258) );
  NAND2_X1 U11266 ( .A1(n10154), .A2(n10153), .ZN(n10157) );
  INV_X1 U11267 ( .A(n10155), .ZN(n10156) );
  NAND2_X1 U11268 ( .A1(n10157), .A2(n10156), .ZN(n10158) );
  OAI211_X1 U11269 ( .C1(n10163), .C2(n10162), .A(n10161), .B(n10160), .ZN(
        n10164) );
  INV_X1 U11270 ( .A(n10164), .ZN(n10171) );
  AOI21_X1 U11271 ( .B1(n10167), .B2(n10166), .A(n10165), .ZN(n10168) );
  OR2_X1 U11272 ( .A1(n10169), .A2(n10168), .ZN(n10170) );
  OAI211_X1 U11273 ( .C1(n10517), .C2(n10172), .A(n10171), .B(n10170), .ZN(
        P1_U3259) );
  OAI21_X1 U11274 ( .B1(n4573), .B2(n10178), .A(n10173), .ZN(n10288) );
  INV_X1 U11275 ( .A(n10174), .ZN(n10182) );
  NAND2_X1 U11276 ( .A1(n10232), .A2(n10175), .ZN(n10177) );
  NAND2_X1 U11277 ( .A1(n10177), .A2(n10176), .ZN(n10179) );
  XNOR2_X1 U11278 ( .A(n10179), .B(n10178), .ZN(n10180) );
  OAI222_X1 U11279 ( .A1(n10183), .A2(n10182), .B1(n10209), .B2(n10181), .C1(
        n10180), .C2(n10228), .ZN(n10286) );
  AOI21_X1 U11280 ( .B1(n10184), .B2(n10288), .A(n10286), .ZN(n10195) );
  INV_X1 U11281 ( .A(n10185), .ZN(n10186) );
  AOI222_X1 U11282 ( .A1(n10188), .A2(n10187), .B1(P1_REG2_REG_6__SCAN_IN), 
        .B2(n10215), .C1(n10186), .C2(n10203), .ZN(n10194) );
  NOR2_X1 U11283 ( .A1(n10197), .A2(n10189), .ZN(n10190) );
  OR2_X1 U11284 ( .A1(n10191), .A2(n10190), .ZN(n10285) );
  INV_X1 U11285 ( .A(n10285), .ZN(n10192) );
  AOI22_X1 U11286 ( .A1(n10288), .A2(n10222), .B1(n10221), .B2(n10192), .ZN(
        n10193) );
  OAI211_X1 U11287 ( .C1(n10215), .C2(n10195), .A(n10194), .B(n10193), .ZN(
        P1_U3285) );
  XOR2_X1 U11288 ( .A(n10208), .B(n10196), .Z(n10281) );
  INV_X1 U11289 ( .A(n10197), .ZN(n10199) );
  OAI211_X1 U11290 ( .C1(n10278), .C2(n4747), .A(n10199), .B(n10198), .ZN(
        n10277) );
  AOI22_X1 U11291 ( .A1(n10203), .A2(n10202), .B1(n10201), .B2(n10200), .ZN(
        n10205) );
  NAND2_X1 U11292 ( .A1(n10204), .A2(n10223), .ZN(n10276) );
  OAI211_X1 U11293 ( .C1(n10277), .C2(n10206), .A(n10205), .B(n10276), .ZN(
        n10212) );
  XNOR2_X1 U11294 ( .A(n10207), .B(n10208), .ZN(n10211) );
  OAI22_X1 U11295 ( .A1(n10211), .A2(n10228), .B1(n10210), .B2(n10209), .ZN(
        n10279) );
  AOI211_X1 U11296 ( .C1(n10213), .C2(n10281), .A(n10212), .B(n10279), .ZN(
        n10214) );
  AOI22_X1 U11297 ( .A1(n10215), .A2(n5383), .B1(n10214), .B2(n9403), .ZN(
        P1_U3286) );
  XOR2_X1 U11298 ( .A(n10216), .B(n10229), .Z(n10236) );
  INV_X1 U11299 ( .A(n10236), .ZN(n10274) );
  INV_X1 U11300 ( .A(n10217), .ZN(n10219) );
  OAI21_X1 U11301 ( .B1(n10219), .B2(n10270), .A(n10218), .ZN(n10271) );
  INV_X1 U11302 ( .A(n10271), .ZN(n10220) );
  AOI22_X1 U11303 ( .A1(n10274), .A2(n10222), .B1(n10221), .B2(n10220), .ZN(
        n10243) );
  AOI22_X1 U11304 ( .A1(n10226), .A2(n10225), .B1(n10224), .B2(n10223), .ZN(
        n10234) );
  AOI21_X1 U11305 ( .B1(n10230), .B2(n10229), .A(n10228), .ZN(n10231) );
  OAI21_X1 U11306 ( .B1(n10232), .B2(n4652), .A(n10231), .ZN(n10233) );
  OAI211_X1 U11307 ( .C1(n10236), .C2(n10235), .A(n10234), .B(n10233), .ZN(
        n10272) );
  MUX2_X1 U11308 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10272), .S(n9403), .Z(
        n10241) );
  OAI22_X1 U11309 ( .A1(n10239), .A2(n10270), .B1(n10238), .B2(n10237), .ZN(
        n10240) );
  NOR2_X1 U11310 ( .A1(n10241), .A2(n10240), .ZN(n10242) );
  NAND2_X1 U11311 ( .A1(n10243), .A2(n10242), .ZN(P1_U3287) );
  AND2_X1 U11312 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10247), .ZN(P1_U3292) );
  AND2_X1 U11313 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10247), .ZN(P1_U3293) );
  AND2_X1 U11314 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10247), .ZN(P1_U3294) );
  AND2_X1 U11315 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10247), .ZN(P1_U3295) );
  AND2_X1 U11316 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10247), .ZN(P1_U3296) );
  AND2_X1 U11317 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10247), .ZN(P1_U3297) );
  AND2_X1 U11318 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10247), .ZN(P1_U3298) );
  AND2_X1 U11319 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10247), .ZN(P1_U3299) );
  AND2_X1 U11320 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10247), .ZN(P1_U3300) );
  AND2_X1 U11321 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10247), .ZN(P1_U3301) );
  AND2_X1 U11322 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10247), .ZN(P1_U3302) );
  AND2_X1 U11323 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10247), .ZN(P1_U3303) );
  AND2_X1 U11324 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10247), .ZN(P1_U3304) );
  AND2_X1 U11325 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10247), .ZN(P1_U3305) );
  AND2_X1 U11326 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10247), .ZN(P1_U3306) );
  AND2_X1 U11327 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10247), .ZN(P1_U3307) );
  AND2_X1 U11328 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10247), .ZN(P1_U3308) );
  AND2_X1 U11329 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10247), .ZN(P1_U3309) );
  AND2_X1 U11330 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10247), .ZN(P1_U3310) );
  AND2_X1 U11331 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10247), .ZN(P1_U3311) );
  AND2_X1 U11332 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10247), .ZN(P1_U3312) );
  AND2_X1 U11333 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10247), .ZN(P1_U3313) );
  AND2_X1 U11334 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10247), .ZN(P1_U3314) );
  AND2_X1 U11335 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10247), .ZN(P1_U3315) );
  AND2_X1 U11336 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10247), .ZN(P1_U3316) );
  AND2_X1 U11337 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10247), .ZN(P1_U3317) );
  AND2_X1 U11338 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10247), .ZN(P1_U3318) );
  INV_X1 U11339 ( .A(n10247), .ZN(n10246) );
  NOR2_X1 U11340 ( .A1(n10246), .A2(n10244), .ZN(P1_U3319) );
  NOR2_X1 U11341 ( .A1(n10246), .A2(n10245), .ZN(P1_U3320) );
  AND2_X1 U11342 ( .A1(n10247), .A2(P1_D_REG_2__SCAN_IN), .ZN(P1_U3321) );
  INV_X1 U11343 ( .A(n10248), .ZN(n10254) );
  INV_X1 U11344 ( .A(n10249), .ZN(n10250) );
  OAI21_X1 U11345 ( .B1(n10251), .B2(n10304), .A(n10250), .ZN(n10253) );
  AOI211_X1 U11346 ( .C1(n10309), .C2(n10254), .A(n10253), .B(n10252), .ZN(
        n10316) );
  INV_X1 U11347 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10255) );
  AOI22_X1 U11348 ( .A1(n10315), .A2(n10316), .B1(n10255), .B2(n10313), .ZN(
        P1_U3457) );
  INV_X1 U11349 ( .A(n10256), .ZN(n10261) );
  OAI22_X1 U11350 ( .A1(n10258), .A2(n10306), .B1(n10257), .B2(n10304), .ZN(
        n10260) );
  AOI211_X1 U11351 ( .C1(n10309), .C2(n10261), .A(n10260), .B(n10259), .ZN(
        n10317) );
  INV_X1 U11352 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10262) );
  AOI22_X1 U11353 ( .A1(n10315), .A2(n10317), .B1(n10262), .B2(n10313), .ZN(
        P1_U3460) );
  INV_X1 U11354 ( .A(n10263), .ZN(n10268) );
  OAI22_X1 U11355 ( .A1(n10265), .A2(n10306), .B1(n10264), .B2(n10304), .ZN(
        n10267) );
  AOI211_X1 U11356 ( .C1(n10309), .C2(n10268), .A(n10267), .B(n10266), .ZN(
        n10318) );
  INV_X1 U11357 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10269) );
  AOI22_X1 U11358 ( .A1(n10315), .A2(n10318), .B1(n10269), .B2(n10313), .ZN(
        P1_U3463) );
  OAI22_X1 U11359 ( .A1(n10271), .A2(n10306), .B1(n10270), .B2(n10304), .ZN(
        n10273) );
  AOI211_X1 U11360 ( .C1(n10309), .C2(n10274), .A(n10273), .B(n10272), .ZN(
        n10319) );
  INV_X1 U11361 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10275) );
  AOI22_X1 U11362 ( .A1(n10315), .A2(n10319), .B1(n10275), .B2(n10313), .ZN(
        P1_U3466) );
  OAI211_X1 U11363 ( .C1(n10278), .C2(n10304), .A(n10277), .B(n10276), .ZN(
        n10280) );
  AOI211_X1 U11364 ( .C1(n10281), .C2(n10295), .A(n10280), .B(n10279), .ZN(
        n10320) );
  INV_X1 U11365 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10282) );
  AOI22_X1 U11366 ( .A1(n10315), .A2(n10320), .B1(n10282), .B2(n10313), .ZN(
        P1_U3469) );
  INV_X1 U11367 ( .A(n10283), .ZN(n10284) );
  OAI21_X1 U11368 ( .B1(n10285), .B2(n10306), .A(n10284), .ZN(n10287) );
  AOI211_X1 U11369 ( .C1(n10295), .C2(n10288), .A(n10287), .B(n10286), .ZN(
        n10321) );
  INV_X1 U11370 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U11371 ( .A1(n10315), .A2(n10321), .B1(n10289), .B2(n10313), .ZN(
        P1_U3472) );
  OAI211_X1 U11372 ( .C1(n10292), .C2(n10304), .A(n10291), .B(n10290), .ZN(
        n10293) );
  AOI21_X1 U11373 ( .B1(n10295), .B2(n10294), .A(n10293), .ZN(n10322) );
  INV_X1 U11374 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10296) );
  AOI22_X1 U11375 ( .A1(n10315), .A2(n10322), .B1(n10296), .B2(n10313), .ZN(
        P1_U3475) );
  INV_X1 U11376 ( .A(n10297), .ZN(n10302) );
  OAI21_X1 U11377 ( .B1(n10299), .B2(n10306), .A(n10298), .ZN(n10301) );
  AOI211_X1 U11378 ( .C1(n10309), .C2(n10302), .A(n10301), .B(n10300), .ZN(
        n10323) );
  INV_X1 U11379 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10303) );
  AOI22_X1 U11380 ( .A1(n10315), .A2(n10323), .B1(n10303), .B2(n10313), .ZN(
        P1_U3478) );
  OAI22_X1 U11381 ( .A1(n10307), .A2(n10306), .B1(n10305), .B2(n10304), .ZN(
        n10308) );
  AOI21_X1 U11382 ( .B1(n10310), .B2(n10309), .A(n10308), .ZN(n10311) );
  AND2_X1 U11383 ( .A1(n10312), .A2(n10311), .ZN(n10325) );
  INV_X1 U11384 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10314) );
  AOI22_X1 U11385 ( .A1(n10315), .A2(n10325), .B1(n10314), .B2(n10313), .ZN(
        P1_U3481) );
  AOI22_X1 U11386 ( .A1(n10326), .A2(n10316), .B1(n6590), .B2(n10324), .ZN(
        P1_U3524) );
  AOI22_X1 U11387 ( .A1(n10326), .A2(n10317), .B1(n10054), .B2(n10324), .ZN(
        P1_U3525) );
  AOI22_X1 U11388 ( .A1(n10326), .A2(n10318), .B1(n6476), .B2(n10324), .ZN(
        P1_U3526) );
  AOI22_X1 U11389 ( .A1(n10326), .A2(n10319), .B1(n5344), .B2(n10324), .ZN(
        P1_U3527) );
  AOI22_X1 U11390 ( .A1(n10326), .A2(n10320), .B1(n6472), .B2(n10324), .ZN(
        P1_U3528) );
  AOI22_X1 U11391 ( .A1(n10326), .A2(n10321), .B1(n6480), .B2(n10324), .ZN(
        P1_U3529) );
  AOI22_X1 U11392 ( .A1(n10326), .A2(n10322), .B1(n6481), .B2(n10324), .ZN(
        P1_U3530) );
  AOI22_X1 U11393 ( .A1(n10326), .A2(n10323), .B1(n6471), .B2(n10324), .ZN(
        P1_U3531) );
  AOI22_X1 U11394 ( .A1(n10326), .A2(n10325), .B1(n5454), .B2(n10324), .ZN(
        P1_U3532) );
  OAI211_X1 U11395 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n10328), .A(n10327), .B(
        P2_IR_REG_0__SCAN_IN), .ZN(n10329) );
  AOI21_X1 U11396 ( .B1(n10331), .B2(n5953), .A(n10329), .ZN(n10337) );
  AOI22_X1 U11397 ( .A1(n10331), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10330), .ZN(n10336) );
  AOI22_X1 U11398 ( .A1(n10333), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10334) );
  OAI221_X1 U11399 ( .B1(n10337), .B2(n10336), .C1(n10337), .C2(n10335), .A(
        n10334), .ZN(P2_U3245) );
  XNOR2_X1 U11400 ( .A(n10338), .B(n10345), .ZN(n10340) );
  AOI21_X1 U11401 ( .B1(n10340), .B2(n10369), .A(n10339), .ZN(n10443) );
  AOI222_X1 U11402 ( .A1(n10347), .A2(n10381), .B1(P2_REG2_REG_6__SCAN_IN), 
        .B2(n10389), .C1(n10379), .C2(n10341), .ZN(n10354) );
  NAND2_X1 U11403 ( .A1(n10356), .A2(n10342), .ZN(n10343) );
  AND2_X1 U11404 ( .A1(n10344), .A2(n10343), .ZN(n10346) );
  XNOR2_X1 U11405 ( .A(n10346), .B(n10345), .ZN(n10446) );
  NAND2_X1 U11406 ( .A1(n10359), .A2(n10347), .ZN(n10348) );
  NAND2_X1 U11407 ( .A1(n10348), .A2(n10360), .ZN(n10350) );
  OR2_X1 U11408 ( .A1(n10350), .A2(n10349), .ZN(n10442) );
  INV_X1 U11409 ( .A(n10442), .ZN(n10351) );
  AOI22_X1 U11410 ( .A1(n10446), .A2(n10352), .B1(n10383), .B2(n10351), .ZN(
        n10353) );
  OAI211_X1 U11411 ( .C1(n10389), .C2(n10443), .A(n10354), .B(n10353), .ZN(
        P2_U3290) );
  NAND2_X1 U11412 ( .A1(n10356), .A2(n10355), .ZN(n10357) );
  XNOR2_X1 U11413 ( .A(n6332), .B(n10357), .ZN(n10440) );
  INV_X1 U11414 ( .A(n10358), .ZN(n10361) );
  OAI211_X1 U11415 ( .C1(n10361), .C2(n10437), .A(n10360), .B(n10359), .ZN(
        n10436) );
  INV_X1 U11416 ( .A(n10362), .ZN(n10365) );
  AOI22_X1 U11417 ( .A1(n10379), .A2(n10365), .B1(n10364), .B2(n10363), .ZN(
        n10366) );
  OAI21_X1 U11418 ( .B1(n10436), .B2(n10367), .A(n10366), .ZN(n10374) );
  OAI211_X1 U11419 ( .C1(n10371), .C2(n10370), .A(n10368), .B(n10369), .ZN(
        n10373) );
  NAND2_X1 U11420 ( .A1(n10373), .A2(n10372), .ZN(n10438) );
  AOI211_X1 U11421 ( .C1(n10440), .C2(n10375), .A(n10374), .B(n10438), .ZN(
        n10377) );
  AOI22_X1 U11422 ( .A1(n10389), .A2(n5990), .B1(n10377), .B2(n10376), .ZN(
        P2_U3291) );
  AOI22_X1 U11423 ( .A1(n10379), .A2(n10378), .B1(P2_REG2_REG_3__SCAN_IN), 
        .B2(n10389), .ZN(n10387) );
  INV_X1 U11424 ( .A(n10380), .ZN(n10384) );
  AOI222_X1 U11425 ( .A1(n10385), .A2(n10384), .B1(n10383), .B2(n10382), .C1(
        n5984), .C2(n10381), .ZN(n10386) );
  OAI211_X1 U11426 ( .C1(n10389), .C2(n10388), .A(n10387), .B(n10386), .ZN(
        P2_U3293) );
  NOR2_X1 U11427 ( .A1(n10391), .A2(n10390), .ZN(n10406) );
  INV_X1 U11428 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n10392) );
  NOR2_X1 U11429 ( .A1(n10427), .A2(n10392), .ZN(P2_U3297) );
  INV_X1 U11430 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n10393) );
  NOR2_X1 U11431 ( .A1(n10427), .A2(n10393), .ZN(P2_U3298) );
  INV_X1 U11432 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n10394) );
  NOR2_X1 U11433 ( .A1(n10427), .A2(n10394), .ZN(P2_U3299) );
  INV_X1 U11434 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n10395) );
  NOR2_X1 U11435 ( .A1(n10427), .A2(n10395), .ZN(P2_U3300) );
  INV_X1 U11436 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n10396) );
  NOR2_X1 U11437 ( .A1(n10406), .A2(n10396), .ZN(P2_U3301) );
  INV_X1 U11438 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n10397) );
  NOR2_X1 U11439 ( .A1(n10406), .A2(n10397), .ZN(P2_U3302) );
  INV_X1 U11440 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n10398) );
  NOR2_X1 U11441 ( .A1(n10406), .A2(n10398), .ZN(P2_U3303) );
  INV_X1 U11442 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n10399) );
  NOR2_X1 U11443 ( .A1(n10406), .A2(n10399), .ZN(P2_U3304) );
  INV_X1 U11444 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10400) );
  NOR2_X1 U11445 ( .A1(n10406), .A2(n10400), .ZN(P2_U3305) );
  INV_X1 U11446 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n10401) );
  NOR2_X1 U11447 ( .A1(n10406), .A2(n10401), .ZN(P2_U3306) );
  INV_X1 U11448 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n10402) );
  NOR2_X1 U11449 ( .A1(n10406), .A2(n10402), .ZN(P2_U3307) );
  INV_X1 U11450 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n10403) );
  NOR2_X1 U11451 ( .A1(n10406), .A2(n10403), .ZN(P2_U3308) );
  INV_X1 U11452 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n10404) );
  NOR2_X1 U11453 ( .A1(n10406), .A2(n10404), .ZN(P2_U3309) );
  INV_X1 U11454 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n10405) );
  NOR2_X1 U11455 ( .A1(n10406), .A2(n10405), .ZN(P2_U3310) );
  INV_X1 U11456 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n10407) );
  NOR2_X1 U11457 ( .A1(n10427), .A2(n10407), .ZN(P2_U3311) );
  INV_X1 U11458 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n10408) );
  NOR2_X1 U11459 ( .A1(n10427), .A2(n10408), .ZN(P2_U3312) );
  INV_X1 U11460 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10409) );
  NOR2_X1 U11461 ( .A1(n10427), .A2(n10409), .ZN(P2_U3313) );
  INV_X1 U11462 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n10410) );
  NOR2_X1 U11463 ( .A1(n10427), .A2(n10410), .ZN(P2_U3314) );
  INV_X1 U11464 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n10411) );
  NOR2_X1 U11465 ( .A1(n10427), .A2(n10411), .ZN(P2_U3315) );
  INV_X1 U11466 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10412) );
  NOR2_X1 U11467 ( .A1(n10427), .A2(n10412), .ZN(P2_U3316) );
  INV_X1 U11468 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n10413) );
  NOR2_X1 U11469 ( .A1(n10427), .A2(n10413), .ZN(P2_U3317) );
  INV_X1 U11470 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10414) );
  NOR2_X1 U11471 ( .A1(n10427), .A2(n10414), .ZN(P2_U3318) );
  INV_X1 U11472 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10415) );
  NOR2_X1 U11473 ( .A1(n10427), .A2(n10415), .ZN(P2_U3319) );
  INV_X1 U11474 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n10416) );
  NOR2_X1 U11475 ( .A1(n10427), .A2(n10416), .ZN(P2_U3320) );
  INV_X1 U11476 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10417) );
  NOR2_X1 U11477 ( .A1(n10427), .A2(n10417), .ZN(P2_U3321) );
  INV_X1 U11478 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n10418) );
  NOR2_X1 U11479 ( .A1(n10427), .A2(n10418), .ZN(P2_U3322) );
  NOR2_X1 U11480 ( .A1(n10427), .A2(n10419), .ZN(P2_U3323) );
  NOR2_X1 U11481 ( .A1(n10427), .A2(n10420), .ZN(P2_U3324) );
  NOR2_X1 U11482 ( .A1(n10427), .A2(n10421), .ZN(P2_U3325) );
  NOR2_X1 U11483 ( .A1(n10427), .A2(n10422), .ZN(P2_U3326) );
  OAI22_X1 U11484 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n10427), .B1(n10423), .B2(
        n10425), .ZN(n10424) );
  INV_X1 U11485 ( .A(n10424), .ZN(P2_U3437) );
  OAI22_X1 U11486 ( .A1(P2_D_REG_1__SCAN_IN), .A2(n10427), .B1(n10426), .B2(
        n10425), .ZN(n10428) );
  INV_X1 U11487 ( .A(n10428), .ZN(P2_U3438) );
  INV_X1 U11488 ( .A(n10429), .ZN(n10435) );
  OAI22_X1 U11489 ( .A1(n10433), .A2(n10432), .B1(n10431), .B2(n10430), .ZN(
        n10434) );
  NOR2_X1 U11490 ( .A1(n10435), .A2(n10434), .ZN(n10470) );
  AOI22_X1 U11491 ( .A1(n10469), .A2(n10470), .B1(n5951), .B2(n10468), .ZN(
        P2_U3451) );
  OAI21_X1 U11492 ( .B1(n10437), .B2(n10460), .A(n10436), .ZN(n10439) );
  AOI211_X1 U11493 ( .C1(n10440), .C2(n10466), .A(n10439), .B(n10438), .ZN(
        n10471) );
  INV_X1 U11494 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10441) );
  AOI22_X1 U11495 ( .A1(n10469), .A2(n10471), .B1(n10441), .B2(n10468), .ZN(
        P2_U3466) );
  OAI211_X1 U11496 ( .C1(n10444), .C2(n10460), .A(n10443), .B(n10442), .ZN(
        n10445) );
  AOI21_X1 U11497 ( .B1(n10446), .B2(n10466), .A(n10445), .ZN(n10472) );
  AOI22_X1 U11498 ( .A1(n10469), .A2(n10472), .B1(n6008), .B2(n10468), .ZN(
        P2_U3469) );
  INV_X1 U11499 ( .A(n10447), .ZN(n10452) );
  OAI22_X1 U11500 ( .A1(n10449), .A2(n10462), .B1(n10448), .B2(n10460), .ZN(
        n10451) );
  AOI211_X1 U11501 ( .C1(n10453), .C2(n10452), .A(n10451), .B(n10450), .ZN(
        n10473) );
  AOI22_X1 U11502 ( .A1(n10469), .A2(n10473), .B1(n6051), .B2(n10468), .ZN(
        P2_U3475) );
  OAI22_X1 U11503 ( .A1(n10455), .A2(n10462), .B1(n10454), .B2(n10460), .ZN(
        n10456) );
  AOI211_X1 U11504 ( .C1(n10458), .C2(n10466), .A(n10457), .B(n10456), .ZN(
        n10474) );
  INV_X1 U11505 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10459) );
  AOI22_X1 U11506 ( .A1(n10469), .A2(n10474), .B1(n10459), .B2(n10468), .ZN(
        P2_U3481) );
  OAI22_X1 U11507 ( .A1(n10463), .A2(n10462), .B1(n10461), .B2(n10460), .ZN(
        n10465) );
  AOI211_X1 U11508 ( .C1(n10467), .C2(n10466), .A(n10465), .B(n10464), .ZN(
        n10476) );
  AOI22_X1 U11509 ( .A1(n10469), .A2(n10476), .B1(n6107), .B2(n10468), .ZN(
        P2_U3487) );
  AOI22_X1 U11510 ( .A1(n10477), .A2(n10470), .B1(n5952), .B2(n10475), .ZN(
        P2_U3520) );
  AOI22_X1 U11511 ( .A1(n10477), .A2(n10471), .B1(n5989), .B2(n10475), .ZN(
        P2_U3525) );
  AOI22_X1 U11512 ( .A1(n10477), .A2(n10472), .B1(n6659), .B2(n10475), .ZN(
        P2_U3526) );
  AOI22_X1 U11513 ( .A1(n10477), .A2(n10473), .B1(n6990), .B2(n10475), .ZN(
        P2_U3528) );
  AOI22_X1 U11514 ( .A1(n10477), .A2(n10474), .B1(n6992), .B2(n10475), .ZN(
        P2_U3530) );
  AOI22_X1 U11515 ( .A1(n10477), .A2(n10476), .B1(n6111), .B2(n10475), .ZN(
        P2_U3532) );
  INV_X1 U11516 ( .A(n10478), .ZN(n10479) );
  NAND2_X1 U11517 ( .A1(n10480), .A2(n10479), .ZN(n10481) );
  XNOR2_X1 U11518 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10481), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11519 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11520 ( .B1(n10484), .B2(n10483), .A(n10482), .ZN(ADD_1071_U56) );
  OAI21_X1 U11521 ( .B1(n10487), .B2(n10486), .A(n10485), .ZN(ADD_1071_U57) );
  OAI21_X1 U11522 ( .B1(n10490), .B2(n10489), .A(n10488), .ZN(ADD_1071_U58) );
  OAI21_X1 U11523 ( .B1(n10493), .B2(n10492), .A(n10491), .ZN(ADD_1071_U59) );
  OAI21_X1 U11524 ( .B1(n10496), .B2(n10495), .A(n10494), .ZN(ADD_1071_U60) );
  OAI21_X1 U11525 ( .B1(n10499), .B2(n10498), .A(n10497), .ZN(ADD_1071_U61) );
  AOI21_X1 U11526 ( .B1(n10502), .B2(n10501), .A(n10500), .ZN(ADD_1071_U62) );
  AOI21_X1 U11527 ( .B1(n10505), .B2(n10504), .A(n10503), .ZN(ADD_1071_U63) );
  AOI21_X1 U11528 ( .B1(n10508), .B2(n10507), .A(n10506), .ZN(ADD_1071_U47) );
  XOR2_X1 U11529 ( .A(n10509), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U11530 ( .A(n10511), .B(n10510), .Z(ADD_1071_U54) );
  NOR2_X1 U11531 ( .A1(n10513), .A2(n10512), .ZN(n10514) );
  XOR2_X1 U11532 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10514), .Z(ADD_1071_U51) );
  OAI21_X1 U11533 ( .B1(n10517), .B2(n10516), .A(n10515), .ZN(n10518) );
  XNOR2_X1 U11534 ( .A(n10518), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11535 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10519), .Z(ADD_1071_U48) );
  XOR2_X1 U11536 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10520), .Z(ADD_1071_U50) );
  XOR2_X1 U11537 ( .A(n10522), .B(n10521), .Z(ADD_1071_U53) );
  XNOR2_X1 U11538 ( .A(n10524), .B(n10523), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U5537 ( .A(n5285), .Z(n5817) );
endmodule

