

module b14_C_SARLock_k_64_8 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, U3352, U3351, U3350, U3349, U3348, U3347, 
        U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, 
        U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, 
        U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, 
        U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, 
        U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, 
        U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, 
        U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, 
        U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, 
        U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, 
        U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, 
        U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, 
        U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, 
        U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, 
        U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, 
        U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, 
        U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, 
        U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, 
        U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, 
        U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, 
        U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, 
        U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, 
        U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, 
        U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, 
        U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621;

  INV_X4 U2265 ( .A(n2496), .ZN(n2456) );
  INV_X1 U2266 ( .A(n2437), .ZN(n3609) );
  AND3_X1 U2268 ( .A1(n2162), .A2(n2028), .A3(n2160), .ZN(n2305) );
  OR2_X1 U2269 ( .A1(n2308), .A2(IR_REG_27__SCAN_IN), .ZN(n2282) );
  NOR2_X1 U2270 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2247)
         );
  NAND2_X1 U2271 ( .A1(n3555), .A2(n3553), .ZN(n2073) );
  AND2_X1 U2272 ( .A1(n2305), .A2(n2276), .ZN(n2295) );
  NAND2_X1 U2274 ( .A1(n4335), .A2(n4336), .ZN(n2024) );
  AOI21_X1 U2275 ( .B1(n4026), .B2(n4032), .A(n3803), .ZN(n4004) );
  CLKBUF_X2 U2276 ( .A(n2454), .Z(n3349) );
  INV_X2 U2277 ( .A(n2692), .ZN(n2397) );
  NAND4_X1 U2279 ( .A1(n2375), .A2(n2374), .A3(n2373), .A4(n2372), .ZN(n3056)
         );
  INV_X1 U2280 ( .A(n4521), .ZN(n4061) );
  OR2_X1 U2281 ( .A1(n4466), .A2(n3257), .ZN(n3265) );
  AND2_X1 U2282 ( .A1(n2034), .A2(n2162), .ZN(n2150) );
  AND2_X1 U2283 ( .A1(n2290), .A2(n2289), .ZN(n3687) );
  AND2_X2 U2284 ( .A1(n2146), .A2(n2043), .ZN(n2022) );
  NOR2_X2 U2285 ( .A1(n3138), .A2(n3137), .ZN(n3140) );
  OAI22_X2 U2286 ( .A1(n3272), .A2(n2144), .B1(n3273), .B2(n2143), .ZN(n2626)
         );
  OAI21_X2 U2287 ( .B1(n3238), .B2(n3239), .A(n3240), .ZN(n3272) );
  NAND2_X1 U2288 ( .A1(n4335), .A2(n4336), .ZN(n2023) );
  INV_X1 U2289 ( .A(n2024), .ZN(n2025) );
  AOI21_X1 U2290 ( .B1(n3421), .B2(n3422), .A(n3424), .ZN(n3510) );
  NOR3_X1 U2291 ( .A1(n2022), .A2(n3396), .A3(n3395), .ZN(n3394) );
  CLKBUF_X1 U2293 ( .A(n2439), .Z(n2792) );
  AND4_X1 U2294 ( .A1(n2453), .A2(n2452), .A3(n2451), .A4(n2450), .ZN(n2990)
         );
  NAND2_X1 U2295 ( .A1(n2845), .A2(n3687), .ZN(n3033) );
  INV_X1 U2296 ( .A(n2252), .ZN(n2162) );
  NAND4_X1 U2297 ( .A1(n2250), .A2(n2249), .A3(n2248), .A4(n2247), .ZN(n2252)
         );
  AND3_X1 U2298 ( .A1(n2246), .A2(n2245), .A3(n2244), .ZN(n2250) );
  NOR2_X1 U2299 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2303)
         );
  OAI21_X1 U2300 ( .B1(n2022), .B2(n2740), .A(n2739), .ZN(n3452) );
  AND2_X1 U2301 ( .A1(n3848), .A2(n3857), .ZN(n3850) );
  AND2_X1 U2302 ( .A1(n3908), .A2(n3785), .ZN(n3891) );
  OAI21_X1 U2303 ( .B1(n3987), .B2(n3779), .A(n3781), .ZN(n3971) );
  NAND2_X1 U2304 ( .A1(n3777), .A2(n3776), .ZN(n4045) );
  OR2_X1 U2305 ( .A1(n3809), .A2(n2055), .ZN(n2051) );
  NAND2_X1 U2306 ( .A1(n3879), .A2(n2167), .ZN(n3839) );
  NAND2_X1 U2307 ( .A1(n3660), .A2(n3288), .ZN(n3322) );
  NAND2_X1 U2308 ( .A1(n2065), .A2(n3802), .ZN(n4026) );
  NAND2_X1 U2309 ( .A1(n2064), .A2(n2044), .ZN(n2065) );
  NOR3_X2 U2310 ( .A1(n3265), .A2(n3295), .A3(n2164), .ZN(n2163) );
  OAI22_X1 U2311 ( .A1(n4371), .A2(n2099), .B1(n2490), .B2(n4554), .ZN(n2321)
         );
  OAI21_X1 U2312 ( .B1(n3036), .B2(n3002), .A(n3563), .ZN(n3133) );
  AND2_X1 U2313 ( .A1(n2976), .A2(n2133), .ZN(n2132) );
  NOR2_X1 U2314 ( .A1(n2975), .A2(n2136), .ZN(n2135) );
  NAND2_X1 U2315 ( .A1(n2995), .A2(n2069), .ZN(n2068) );
  NOR2_X1 U2316 ( .A1(n4359), .A2(n4360), .ZN(n4358) );
  INV_X1 U2317 ( .A(n2990), .ZN(n4491) );
  AND2_X2 U2318 ( .A1(n2840), .A2(n3033), .ZN(n2793) );
  XNOR2_X1 U2319 ( .A(n2297), .B(n2296), .ZN(n2884) );
  NAND3_X2 U2320 ( .A1(n2282), .A2(n2281), .A3(n2280), .ZN(n2454) );
  XNOR2_X1 U2321 ( .A(n2366), .B(n3346), .ZN(n2370) );
  OAI21_X1 U2322 ( .B1(n2298), .B2(IR_REG_25__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2299) );
  NAND2_X1 U2323 ( .A1(n2388), .A2(n2027), .ZN(n2123) );
  NAND2_X1 U2324 ( .A1(n2152), .A2(IR_REG_31__SCAN_IN), .ZN(n2366) );
  MUX2_X1 U2325 ( .A(IR_REG_31__SCAN_IN), .B(n2288), .S(IR_REG_21__SCAN_IN), 
        .Z(n2290) );
  AND3_X1 U2326 ( .A1(n2087), .A2(n2303), .A3(n2304), .ZN(n2362) );
  AND2_X1 U2327 ( .A1(n2273), .A2(n2272), .ZN(n2376) );
  AND3_X1 U2328 ( .A1(n2157), .A2(n2156), .A3(n2155), .ZN(n2273) );
  AND2_X1 U2329 ( .A1(n2302), .A2(n2276), .ZN(n2087) );
  NAND2_X1 U2330 ( .A1(n2365), .A2(n2382), .ZN(n2124) );
  AND2_X1 U2331 ( .A1(n2089), .A2(n2090), .ZN(n2088) );
  AND3_X1 U2332 ( .A1(n2200), .A2(n2199), .A3(n2190), .ZN(n2201) );
  INV_X1 U2333 ( .A(IR_REG_27__SCAN_IN), .ZN(n2302) );
  NOR2_X1 U2334 ( .A1(IR_REG_26__SCAN_IN), .A2(IR_REG_25__SCAN_IN), .ZN(n2304)
         );
  NOR2_X1 U2335 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2274)
         );
  NOR2_X1 U2336 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2249)
         );
  NOR2_X1 U2337 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2248)
         );
  AOI21_X2 U2338 ( .B1(n3984), .B2(n3807), .A(n3806), .ZN(n3925) );
  NAND2_X1 U2339 ( .A1(n2393), .A2(n3018), .ZN(n2498) );
  INV_X4 U2340 ( .A(n2439), .ZN(n2393) );
  NOR2_X2 U2341 ( .A1(n4018), .A2(n3632), .ZN(n2169) );
  NOR2_X2 U2342 ( .A1(n3206), .A2(n3205), .ZN(n4468) );
  XNOR2_X2 U2343 ( .A(n2294), .B(n2293), .ZN(n2799) );
  INV_X1 U2344 ( .A(IR_REG_1__SCAN_IN), .ZN(n2089) );
  NAND2_X1 U2345 ( .A1(n3895), .A2(n3881), .ZN(n3818) );
  NOR2_X1 U2346 ( .A1(n2251), .A2(IR_REG_21__SCAN_IN), .ZN(n2159) );
  AND2_X1 U2347 ( .A1(n2644), .A2(n2643), .ZN(n2645) );
  INV_X1 U2348 ( .A(n3033), .ZN(n2383) );
  NOR2_X1 U2349 ( .A1(n2102), .A2(REG2_REG_16__SCAN_IN), .ZN(n2101) );
  INV_X1 U2350 ( .A(n2106), .ZN(n2102) );
  NAND2_X1 U2351 ( .A1(n3738), .A2(n2315), .ZN(n2316) );
  OR2_X1 U2352 ( .A1(n2910), .A2(n4612), .ZN(n2096) );
  NAND2_X1 U2353 ( .A1(n2117), .A2(n2116), .ZN(n4393) );
  OR2_X1 U2354 ( .A1(n4385), .A2(n2119), .ZN(n2116) );
  INV_X1 U2355 ( .A(n4394), .ZN(n2118) );
  NAND2_X1 U2356 ( .A1(n3888), .A2(n2052), .ZN(n3816) );
  NAND2_X1 U2357 ( .A1(n3817), .A2(n3894), .ZN(n2052) );
  OR2_X1 U2358 ( .A1(n3436), .A2(n3525), .ZN(n3318) );
  NAND2_X1 U2359 ( .A1(n3436), .A2(n3525), .ZN(n3316) );
  NAND2_X1 U2360 ( .A1(n2068), .A2(n2066), .ZN(n3148) );
  NOR2_X1 U2361 ( .A1(n2036), .A2(n2067), .ZN(n2066) );
  INV_X1 U2362 ( .A(n2071), .ZN(n2067) );
  NOR2_X2 U2363 ( .A1(n3839), .A2(n3824), .ZN(n4067) );
  XNOR2_X1 U2364 ( .A(n2368), .B(n2151), .ZN(n2369) );
  AND2_X1 U2365 ( .A1(n2376), .A2(n2362), .ZN(n2086) );
  INV_X1 U2366 ( .A(n2251), .ZN(n2160) );
  AND2_X1 U2367 ( .A1(n2272), .A2(n2271), .ZN(n2161) );
  NAND2_X1 U2368 ( .A1(n4491), .A2(n3062), .ZN(n3555) );
  NAND2_X1 U2369 ( .A1(n2308), .A2(IR_REG_28__SCAN_IN), .ZN(n2281) );
  OR2_X1 U2370 ( .A1(n2913), .A2(n2193), .ZN(n2197) );
  OAI22_X1 U2371 ( .A1(n3341), .A2(n2122), .B1(n2255), .B2(n3268), .ZN(n2258)
         );
  NOR2_X1 U2372 ( .A1(n4337), .A2(REG2_REG_13__SCAN_IN), .ZN(n2122) );
  NOR2_X1 U2373 ( .A1(n2608), .A2(n3529), .ZN(n2635) );
  NAND2_X1 U2374 ( .A1(n3203), .A2(n2040), .ZN(n2062) );
  NAND2_X1 U2375 ( .A1(n3072), .A2(n3559), .ZN(n3036) );
  INV_X1 U2376 ( .A(n3000), .ZN(n2078) );
  INV_X1 U2377 ( .A(IR_REG_17__SCAN_IN), .ZN(n2272) );
  INV_X1 U2378 ( .A(IR_REG_16__SCAN_IN), .ZN(n2155) );
  XNOR2_X1 U2379 ( .A(n2604), .B(n2793), .ZN(n3273) );
  NAND2_X1 U2380 ( .A1(n2140), .A2(n2142), .ZN(n2139) );
  INV_X1 U2381 ( .A(n2178), .ZN(n2140) );
  XNOR2_X1 U2382 ( .A(n2419), .B(n2778), .ZN(n2472) );
  NOR2_X1 U2383 ( .A1(n2738), .A2(n2737), .ZN(n2739) );
  NAND2_X1 U2384 ( .A1(n2736), .A2(n2735), .ZN(n2740) );
  OAI211_X1 U2385 ( .C1(n2134), .C2(n2130), .A(n3362), .B(n2127), .ZN(n2520)
         );
  NAND2_X1 U2386 ( .A1(n2129), .A2(n2128), .ZN(n2127) );
  OAI211_X1 U2387 ( .C1(n2384), .C2(n2432), .A(n2431), .B(n2433), .ZN(n2886)
         );
  NAND2_X1 U2388 ( .A1(n3412), .A2(n2704), .ZN(n2147) );
  NAND2_X1 U2389 ( .A1(n3474), .A2(n2148), .ZN(n2146) );
  NOR2_X1 U2390 ( .A1(n2705), .A2(n2149), .ZN(n2148) );
  OR2_X1 U2391 ( .A1(n2628), .A2(n2627), .ZN(n2629) );
  NAND2_X1 U2392 ( .A1(n2311), .A2(REG2_REG_1__SCAN_IN), .ZN(n2184) );
  XNOR2_X1 U2393 ( .A(n2197), .B(n3751), .ZN(n3744) );
  NAND2_X1 U2394 ( .A1(n2096), .A2(n2037), .ZN(n2317) );
  OAI21_X1 U2395 ( .B1(n3744), .B2(n2114), .A(n2112), .ZN(n2115) );
  INV_X1 U2396 ( .A(n2198), .ZN(n2114) );
  AOI21_X1 U2397 ( .B1(n2198), .B2(n2113), .A(n2921), .ZN(n2112) );
  NAND2_X1 U2398 ( .A1(n3744), .A2(REG2_REG_4__SCAN_IN), .ZN(n3747) );
  NOR2_X1 U2399 ( .A1(n4368), .A2(REG1_REG_7__SCAN_IN), .ZN(n2099) );
  NOR2_X1 U2400 ( .A1(n4393), .A2(n2180), .ZN(n2237) );
  NAND2_X1 U2401 ( .A1(n4398), .A2(n2326), .ZN(n2327) );
  NAND2_X1 U2402 ( .A1(n2557), .A2(REG1_REG_11__SCAN_IN), .ZN(n2326) );
  NAND2_X1 U2403 ( .A1(n2330), .A2(n2172), .ZN(n2331) );
  NAND2_X1 U2404 ( .A1(n3336), .A2(n2329), .ZN(n2330) );
  INV_X1 U2405 ( .A(n3335), .ZN(n2329) );
  AND2_X1 U2406 ( .A1(n2108), .A2(n2031), .ZN(n2270) );
  NOR2_X1 U2407 ( .A1(n2270), .A2(n2269), .ZN(n2354) );
  AND2_X1 U2408 ( .A1(n3828), .A2(n3644), .ZN(n3857) );
  NAND2_X1 U2409 ( .A1(n2051), .A2(n2050), .ZN(n2053) );
  AND2_X1 U2410 ( .A1(n3815), .A2(n2054), .ZN(n2050) );
  INV_X1 U2411 ( .A(n3852), .ZN(n3895) );
  NAND2_X1 U2412 ( .A1(n3799), .A2(n3798), .ZN(n2064) );
  AND2_X1 U2413 ( .A1(n3532), .A2(n3302), .ZN(n3303) );
  OR3_X1 U2414 ( .A1(n2597), .A2(n2596), .A3(n2595), .ZN(n2608) );
  OAI22_X1 U2415 ( .A1(n2060), .A2(n2062), .B1(n3260), .B2(n4457), .ZN(n2059)
         );
  INV_X1 U2416 ( .A(n3204), .ZN(n2060) );
  NAND2_X1 U2417 ( .A1(n4450), .A2(n2061), .ZN(n2058) );
  INV_X1 U2418 ( .A(n2062), .ZN(n2061) );
  NAND2_X1 U2419 ( .A1(n2565), .A2(REG3_REG_12__SCAN_IN), .ZN(n2597) );
  INV_X1 U2420 ( .A(n2566), .ZN(n2565) );
  NAND2_X1 U2421 ( .A1(n2085), .A2(n3541), .ZN(n4455) );
  NAND2_X1 U2422 ( .A1(n2084), .A2(n2082), .ZN(n2085) );
  AOI21_X1 U2423 ( .B1(n3581), .B2(n3188), .A(n2083), .ZN(n2082) );
  OAI21_X1 U2424 ( .B1(n3153), .B2(n3152), .A(n3574), .ZN(n3167) );
  NOR2_X1 U2425 ( .A1(n2996), .A2(n2070), .ZN(n2069) );
  INV_X1 U2426 ( .A(n2994), .ZN(n2070) );
  AND3_X1 U2427 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2475) );
  INV_X1 U2428 ( .A(n3014), .ZN(n3029) );
  NOR2_X1 U2429 ( .A1(n3851), .A2(n3841), .ZN(n2167) );
  NAND2_X1 U2430 ( .A1(n2798), .A2(n2801), .ZN(n2881) );
  NAND2_X1 U2431 ( .A1(n2381), .A2(n2380), .ZN(n2388) );
  INV_X1 U2432 ( .A(IR_REG_4__SCAN_IN), .ZN(n2199) );
  INV_X1 U2433 ( .A(n2088), .ZN(n2074) );
  INV_X1 U2434 ( .A(n3768), .ZN(n3763) );
  NAND2_X1 U2435 ( .A1(n2098), .A2(n2097), .ZN(n3740) );
  NAND2_X1 U2436 ( .A1(n2188), .A2(n4610), .ZN(n2097) );
  OR2_X1 U2437 ( .A1(n2188), .A2(n4610), .ZN(n2098) );
  XNOR2_X1 U2438 ( .A(n2317), .B(n3751), .ZN(n3754) );
  NAND2_X1 U2439 ( .A1(n3754), .A2(REG1_REG_4__SCAN_IN), .ZN(n3753) );
  XNOR2_X1 U2440 ( .A(n2324), .B(n2095), .ZN(n4390) );
  NAND2_X1 U2441 ( .A1(n4390), .A2(REG1_REG_10__SCAN_IN), .ZN(n4389) );
  NAND2_X1 U2442 ( .A1(n4399), .A2(n4400), .ZN(n4398) );
  XNOR2_X1 U2443 ( .A(n2327), .B(n4547), .ZN(n4409) );
  NAND2_X1 U2444 ( .A1(n4409), .A2(REG1_REG_12__SCAN_IN), .ZN(n4408) );
  XNOR2_X1 U2445 ( .A(n2331), .B(n2257), .ZN(n4418) );
  NAND2_X1 U2446 ( .A1(n4418), .A2(REG1_REG_14__SCAN_IN), .ZN(n4417) );
  NAND2_X1 U2447 ( .A1(n4423), .A2(n4424), .ZN(n4421) );
  NOR2_X1 U2448 ( .A1(n4436), .A2(n2334), .ZN(n2336) );
  AOI21_X1 U2449 ( .B1(n4435), .B2(ADDR_REG_17__SCAN_IN), .A(n3446), .ZN(n2340) );
  AOI21_X1 U2450 ( .B1(n3838), .B2(n3836), .A(n2174), .ZN(n3823) );
  AND2_X1 U2451 ( .A1(n4041), .A2(n4596), .ZN(n4504) );
  INV_X1 U2452 ( .A(n3395), .ZN(n2736) );
  NAND2_X1 U2453 ( .A1(n2503), .A2(n2131), .ZN(n2130) );
  INV_X1 U2454 ( .A(n3363), .ZN(n2131) );
  INV_X1 U2455 ( .A(n2130), .ZN(n2128) );
  NOR2_X1 U2456 ( .A1(n3274), .A2(n2607), .ZN(n2144) );
  INV_X1 U2457 ( .A(n3274), .ZN(n2143) );
  AND2_X1 U2458 ( .A1(n3907), .A2(n3636), .ZN(n3785) );
  OR2_X1 U2459 ( .A1(n4394), .A2(n4386), .ZN(n2119) );
  NAND2_X1 U2460 ( .A1(n4421), .A2(n2173), .ZN(n2333) );
  INV_X1 U2461 ( .A(n2334), .ZN(n2093) );
  AOI21_X1 U2462 ( .B1(n3891), .B2(n3787), .A(n3786), .ZN(n3848) );
  NOR2_X1 U2463 ( .A1(n2676), .A2(n2675), .ZN(n2693) );
  OR2_X1 U2464 ( .A1(n4045), .A2(n3778), .ZN(n3987) );
  AND2_X1 U2465 ( .A1(n2635), .A2(n2634), .ZN(n2647) );
  NAND2_X1 U2466 ( .A1(n2081), .A2(n3548), .ZN(n3660) );
  NAND2_X1 U2467 ( .A1(n3190), .A2(n2079), .ZN(n3287) );
  NOR2_X1 U2468 ( .A1(n3547), .A2(n2080), .ZN(n2079) );
  INV_X1 U2469 ( .A(n3542), .ZN(n2083) );
  INV_X1 U2470 ( .A(n2075), .ZN(n3070) );
  AOI21_X1 U2471 ( .B1(n4486), .B2(n3000), .A(n2073), .ZN(n2075) );
  AND2_X1 U2472 ( .A1(n3900), .A2(n3881), .ZN(n3879) );
  NAND2_X1 U2473 ( .A1(n2168), .A2(n3195), .ZN(n3206) );
  NOR2_X1 U2474 ( .A1(n3159), .A2(n3367), .ZN(n2168) );
  NAND2_X1 U2475 ( .A1(n4565), .A2(n3077), .ZN(n3076) );
  INV_X1 U2476 ( .A(IR_REG_18__SCAN_IN), .ZN(n2377) );
  OR2_X1 U2477 ( .A1(n2242), .A2(IR_REG_10__SCAN_IN), .ZN(n2232) );
  INV_X1 U2478 ( .A(IR_REG_11__SCAN_IN), .ZN(n2240) );
  NAND2_X1 U2479 ( .A1(n2088), .A2(n2190), .ZN(n2191) );
  INV_X1 U2480 ( .A(n2473), .ZN(n2136) );
  OAI22_X1 U2481 ( .A1(n2948), .A2(n2496), .B1(n2439), .B2(n2970), .ZN(n2403)
         );
  INV_X1 U2482 ( .A(n3122), .ZN(n2528) );
  OR2_X1 U2483 ( .A1(n3462), .A2(n3464), .ZN(n3084) );
  INV_X1 U2484 ( .A(n3995), .ZN(n3632) );
  AND2_X1 U2485 ( .A1(n2560), .A2(n2559), .ZN(n2562) );
  NAND2_X1 U2486 ( .A1(n2154), .A2(n2153), .ZN(n3216) );
  AOI21_X1 U2487 ( .B1(n3464), .B2(n2545), .A(n2033), .ZN(n2153) );
  NAND2_X1 U2488 ( .A1(n3462), .A2(n2545), .ZN(n2154) );
  INV_X1 U2489 ( .A(n3871), .ZN(n3881) );
  AND2_X1 U2490 ( .A1(n3020), .A2(n2817), .ZN(n2849) );
  INV_X1 U2491 ( .A(n2839), .ZN(n2786) );
  NAND2_X1 U2492 ( .A1(n2692), .A2(REG1_REG_1__SCAN_IN), .ZN(n2893) );
  XNOR2_X1 U2493 ( .A(n2192), .B(n2858), .ZN(n2914) );
  XNOR2_X1 U2494 ( .A(n2217), .B(n4552), .ZN(n4375) );
  OAI21_X1 U2495 ( .B1(n4353), .B2(n2110), .A(n2109), .ZN(n2217) );
  NAND2_X1 U2496 ( .A1(n4364), .A2(n2212), .ZN(n2109) );
  NAND2_X1 U2497 ( .A1(n2111), .A2(n2212), .ZN(n2110) );
  INV_X1 U2498 ( .A(n2209), .ZN(n2111) );
  OR2_X1 U2499 ( .A1(n3118), .A2(n3117), .ZN(n3115) );
  NAND2_X1 U2500 ( .A1(n3115), .A2(n2227), .ZN(n2229) );
  OR2_X1 U2501 ( .A1(n4385), .A2(n4386), .ZN(n2121) );
  NOR2_X1 U2502 ( .A1(n2238), .A2(n4403), .ZN(n3341) );
  XNOR2_X1 U2503 ( .A(n2258), .B(n2257), .ZN(n4413) );
  NAND2_X1 U2504 ( .A1(n2104), .A2(n4541), .ZN(n2103) );
  INV_X1 U2505 ( .A(n4425), .ZN(n2104) );
  NAND2_X1 U2506 ( .A1(n4425), .A2(n2105), .ZN(n2100) );
  OAI21_X1 U2507 ( .B1(n4436), .B2(n2092), .A(n2091), .ZN(n2348) );
  NAND2_X1 U2508 ( .A1(n2335), .A2(n2094), .ZN(n2091) );
  NAND2_X1 U2509 ( .A1(n2093), .A2(n2094), .ZN(n2092) );
  NAND2_X1 U2510 ( .A1(n4540), .A2(n4123), .ZN(n2094) );
  NOR2_X1 U2511 ( .A1(n2641), .A2(REG2_REG_17__SCAN_IN), .ZN(n2353) );
  NAND2_X1 U2512 ( .A1(n2348), .A2(n2347), .ZN(n3761) );
  NAND2_X1 U2513 ( .A1(n3831), .A2(n3851), .ZN(n3820) );
  NOR2_X1 U2514 ( .A1(n3831), .A2(n3851), .ZN(n2072) );
  OR2_X1 U2515 ( .A1(n2772), .A2(n3377), .ZN(n2784) );
  AND2_X1 U2516 ( .A1(n2791), .A2(n2790), .ZN(n3854) );
  OR2_X1 U2517 ( .A1(n3843), .A2(n2023), .ZN(n2791) );
  INV_X1 U2518 ( .A(n2744), .ZN(n2743) );
  INV_X1 U2519 ( .A(n3812), .ZN(n2054) );
  NAND2_X1 U2520 ( .A1(n2707), .A2(REG3_REG_22__SCAN_IN), .ZN(n2717) );
  AND2_X1 U2521 ( .A1(n3934), .A2(n3622), .ZN(n3952) );
  NOR2_X1 U2522 ( .A1(n3700), .A2(n4033), .ZN(n3803) );
  INV_X1 U2523 ( .A(n4019), .ZN(n4014) );
  NAND2_X1 U2524 ( .A1(n2647), .A2(REG3_REG_18__SCAN_IN), .ZN(n2663) );
  INV_X1 U2525 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2596) );
  NAND2_X1 U2526 ( .A1(n2063), .A2(n3282), .ZN(n3304) );
  NAND2_X1 U2527 ( .A1(n2058), .A2(n2057), .ZN(n2063) );
  NOR2_X1 U2528 ( .A1(n2059), .A2(n3283), .ZN(n2057) );
  INV_X1 U2529 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2595) );
  NOR2_X1 U2530 ( .A1(n3265), .A2(n3281), .ZN(n3294) );
  NAND2_X1 U2531 ( .A1(n3190), .A2(n3545), .ZN(n3259) );
  INV_X1 U2532 ( .A(n3212), .ZN(n4467) );
  INV_X1 U2533 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3089) );
  OR2_X1 U2534 ( .A1(n2532), .A2(n3089), .ZN(n2550) );
  NOR2_X1 U2535 ( .A1(n2507), .A2(n2506), .ZN(n2522) );
  NAND2_X1 U2536 ( .A1(n3167), .A2(n3580), .ZN(n3155) );
  INV_X1 U2537 ( .A(n3387), .ZN(n3099) );
  NAND2_X1 U2538 ( .A1(n3095), .A2(n3565), .ZN(n3153) );
  AND4_X1 U2539 ( .A1(n2495), .A2(n2494), .A3(n2493), .A4(n2492), .ZN(n3369)
         );
  INV_X1 U2540 ( .A(n3105), .ZN(n3016) );
  OAI21_X1 U2541 ( .B1(n3133), .B2(n3131), .A(n3569), .ZN(n3094) );
  OR2_X1 U2542 ( .A1(n3076), .A2(n3043), .ZN(n3138) );
  NAND2_X1 U2543 ( .A1(n3052), .A2(n2991), .ZN(n3068) );
  OAI21_X1 U2544 ( .B1(n4486), .B2(n2073), .A(n2076), .ZN(n3001) );
  INV_X1 U2545 ( .A(n3553), .ZN(n2077) );
  INV_X1 U2546 ( .A(n3558), .ZN(n3077) );
  INV_X1 U2547 ( .A(n4493), .ZN(n4460) );
  AND2_X1 U2548 ( .A1(n3006), .A2(n3005), .ZN(n4462) );
  OR2_X1 U2549 ( .A1(n2998), .A2(n3647), .ZN(n4486) );
  OR2_X1 U2550 ( .A1(n4341), .A2(n3007), .ZN(n4493) );
  NAND2_X1 U2551 ( .A1(n4509), .A2(n4502), .ZN(n4501) );
  INV_X1 U2552 ( .A(n4462), .ZN(n4511) );
  INV_X1 U2553 ( .A(n4497), .ZN(n4512) );
  INV_X1 U2554 ( .A(n4489), .ZN(n4456) );
  NAND2_X1 U2555 ( .A1(n3879), .A2(n3860), .ZN(n3859) );
  NOR2_X1 U2556 ( .A1(n3916), .A2(n3899), .ZN(n3900) );
  OR2_X1 U2557 ( .A1(n3943), .A2(n3813), .ZN(n3916) );
  NOR2_X1 U2558 ( .A1(n3976), .A2(n3963), .ZN(n3962) );
  NAND2_X1 U2559 ( .A1(n3962), .A2(n3941), .ZN(n3943) );
  INV_X1 U2560 ( .A(n3808), .ZN(n3941) );
  NAND2_X1 U2561 ( .A1(n2169), .A2(n3977), .ZN(n3976) );
  AND2_X1 U2562 ( .A1(n4053), .A2(n4029), .ZN(n4027) );
  NOR2_X1 U2563 ( .A1(n4052), .A2(n3801), .ZN(n4053) );
  NAND2_X1 U2564 ( .A1(n3525), .A2(n2165), .ZN(n2164) );
  NOR3_X1 U2565 ( .A1(n3265), .A2(n3295), .A3(n3281), .ZN(n3309) );
  NAND2_X1 U2566 ( .A1(n4468), .A2(n4467), .ZN(n4466) );
  INV_X1 U2567 ( .A(n2168), .ZN(n3164) );
  AND2_X1 U2568 ( .A1(n3140), .A2(n3016), .ZN(n3100) );
  AND3_X1 U2569 ( .A1(n4509), .A2(n4502), .A3(n3062), .ZN(n4565) );
  INV_X1 U2570 ( .A(n3020), .ZN(n3031) );
  NOR2_X1 U2571 ( .A1(n3015), .A2(n3029), .ZN(n3021) );
  OR2_X1 U2572 ( .A1(n3013), .A2(n3027), .ZN(n3015) );
  AND2_X1 U2573 ( .A1(n2277), .A2(n2276), .ZN(n2278) );
  XNOR2_X1 U2574 ( .A(n2286), .B(n2276), .ZN(n2828) );
  AND2_X1 U2575 ( .A1(n2376), .A2(n2275), .ZN(n2364) );
  AND2_X1 U2576 ( .A1(n2221), .A2(n2220), .ZN(n2223) );
  INV_X1 U2577 ( .A(IR_REG_5__SCAN_IN), .ZN(n2246) );
  XNOR2_X1 U2578 ( .A(n2194), .B(IR_REG_3__SCAN_IN), .ZN(n2858) );
  MUX2_X1 U2579 ( .A(IR_REG_31__SCAN_IN), .B(n2181), .S(IR_REG_1__SCAN_IN), 
        .Z(n2182) );
  AOI21_X1 U2580 ( .B1(n3510), .B2(n3507), .A(n3506), .ZN(n3376) );
  NAND2_X1 U2581 ( .A1(n3084), .A2(n2545), .ZN(n3086) );
  OR2_X1 U2582 ( .A1(n2030), .A2(n3494), .ZN(n2137) );
  OR2_X1 U2583 ( .A1(n3441), .A2(n2139), .ZN(n2138) );
  AND2_X1 U2584 ( .A1(n2827), .A2(n2176), .ZN(n2825) );
  NAND2_X1 U2585 ( .A1(n2126), .A2(n2503), .ZN(n3365) );
  NAND2_X1 U2586 ( .A1(n2134), .A2(n2132), .ZN(n2126) );
  AND4_X1 U2587 ( .A1(n2713), .A2(n2712), .A3(n2711), .A4(n2710), .ZN(n3972)
         );
  NAND2_X1 U2588 ( .A1(n3474), .A2(n3477), .ZN(n3414) );
  NAND2_X1 U2589 ( .A1(n3215), .A2(n3219), .ZN(n3182) );
  INV_X1 U2590 ( .A(n3531), .ZN(n3498) );
  INV_X1 U2591 ( .A(n2999), .ZN(n4509) );
  INV_X1 U2592 ( .A(n3486), .ZN(n2145) );
  NAND2_X1 U2593 ( .A1(n2146), .A2(n2147), .ZN(n3485) );
  NAND2_X1 U2594 ( .A1(n2460), .A2(n2459), .ZN(n2463) );
  OR2_X1 U2595 ( .A1(n3441), .A2(n2178), .ZN(n2141) );
  INV_X1 U2596 ( .A(n3514), .ZN(n3538) );
  AND4_X1 U2597 ( .A1(n2602), .A2(n2601), .A3(n2600), .A4(n2599), .ZN(n3532)
         );
  INV_X1 U2598 ( .A(n3517), .ZN(n3523) );
  OR2_X1 U2599 ( .A1(n3882), .A2(n2024), .ZN(n2763) );
  INV_X1 U2600 ( .A(n3814), .ZN(n3938) );
  NAND4_X1 U2601 ( .A1(n2681), .A2(n2680), .A3(n2679), .A4(n2678), .ZN(n4015)
         );
  NAND4_X1 U2602 ( .A1(n2571), .A2(n2570), .A3(n2569), .A4(n2568), .ZN(n3703)
         );
  NAND4_X1 U2603 ( .A1(n2416), .A2(n2415), .A3(n2414), .A4(n2413), .ZN(n3708)
         );
  NAND4_X1 U2604 ( .A1(n2426), .A2(n2425), .A3(n2424), .A4(n2423), .ZN(n3711)
         );
  OR2_X1 U2605 ( .A1(n2384), .A2(n2883), .ZN(n3726) );
  NAND2_X1 U2606 ( .A1(n2313), .A2(n2312), .ZN(n3714) );
  NAND2_X1 U2607 ( .A1(n2311), .A2(REG1_REG_1__SCAN_IN), .ZN(n2312) );
  OR2_X1 U2608 ( .A1(n2311), .A2(REG1_REG_1__SCAN_IN), .ZN(n2313) );
  NAND2_X1 U2609 ( .A1(n3740), .A2(n3739), .ZN(n3738) );
  XNOR2_X1 U2610 ( .A(n2316), .B(n2858), .ZN(n2910) );
  INV_X1 U2611 ( .A(n2096), .ZN(n2909) );
  AND2_X1 U2612 ( .A1(n3753), .A2(n2318), .ZN(n2925) );
  AND2_X1 U2613 ( .A1(n3747), .A2(n2198), .ZN(n2922) );
  NOR2_X1 U2614 ( .A1(n4353), .A2(n2209), .ZN(n4365) );
  AND2_X1 U2615 ( .A1(n2320), .A2(n2179), .ZN(n4371) );
  XNOR2_X1 U2616 ( .A(n2321), .B(n4552), .ZN(n4381) );
  XNOR2_X1 U2617 ( .A(n2229), .B(n2539), .ZN(n4385) );
  NAND2_X1 U2618 ( .A1(n4389), .A2(n2325), .ZN(n4399) );
  NOR2_X1 U2619 ( .A1(n4405), .A2(n4404), .ZN(n4403) );
  NAND2_X1 U2620 ( .A1(n4408), .A2(n2328), .ZN(n3336) );
  NAND2_X1 U2621 ( .A1(n4417), .A2(n2332), .ZN(n4423) );
  INV_X1 U2622 ( .A(n4426), .ZN(n4440) );
  INV_X1 U2623 ( .A(n4442), .ZN(n4422) );
  INV_X1 U2624 ( .A(n3819), .ZN(n3858) );
  AND2_X1 U2625 ( .A1(n2064), .A2(n2041), .ZN(n4044) );
  NAND2_X1 U2626 ( .A1(n2058), .A2(n2056), .ZN(n3284) );
  INV_X1 U2627 ( .A(n2059), .ZN(n2056) );
  INV_X1 U2628 ( .A(n4504), .ZN(n4056) );
  NAND2_X1 U2629 ( .A1(n4495), .A2(n2989), .ZN(n3050) );
  INV_X1 U2630 ( .A(n4621), .ZN(n4618) );
  AND2_X2 U2631 ( .A1(n3021), .A2(n3020), .ZN(n4621) );
  AOI21_X1 U2632 ( .B1(n4596), .B2(n4074), .A(n4073), .ZN(n4075) );
  AND2_X1 U2633 ( .A1(n4606), .A2(n4596), .ZN(n4148) );
  AND2_X2 U2634 ( .A1(n3021), .A2(n3031), .ZN(n4606) );
  NAND2_X1 U2635 ( .A1(n2882), .A2(n2881), .ZN(n4530) );
  AND2_X1 U2636 ( .A1(n2159), .A2(n2038), .ZN(n2049) );
  INV_X1 U2637 ( .A(n2370), .ZN(n4335) );
  INV_X1 U2638 ( .A(n2369), .ZN(n4336) );
  NAND2_X1 U2639 ( .A1(n2389), .A2(n2388), .ZN(n3768) );
  NAND2_X1 U2640 ( .A1(n2074), .A2(IR_REG_31__SCAN_IN), .ZN(n2187) );
  INV_X1 U2641 ( .A(n2310), .ZN(n2344) );
  AOI22_X1 U2642 ( .A1(n4343), .A2(n4504), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4521), .ZN(n4344) );
  XNOR2_X1 U2643 ( .A(n2187), .B(IR_REG_2__SCAN_IN), .ZN(n2188) );
  AND2_X1 U2644 ( .A1(n2115), .A2(n2042), .ZN(n2026) );
  AND2_X1 U2645 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2027)
         );
  AND3_X1 U2646 ( .A1(n2275), .A2(n2273), .A3(n2161), .ZN(n2028) );
  INV_X1 U2647 ( .A(n3281), .ZN(n2165) );
  NAND4_X1 U2648 ( .A1(n2750), .A2(n2749), .A3(n2748), .A4(n2747), .ZN(n3913)
         );
  INV_X1 U2649 ( .A(n3913), .ZN(n3817) );
  OR2_X1 U2650 ( .A1(n4036), .A2(n4055), .ZN(n2029) );
  AND2_X1 U2651 ( .A1(n2039), .A2(n3493), .ZN(n2030) );
  NAND2_X1 U2652 ( .A1(n2384), .A2(n3033), .ZN(n2439) );
  OR2_X1 U2653 ( .A1(n4541), .A2(n2266), .ZN(n2031) );
  NAND2_X1 U2654 ( .A1(n4335), .A2(n2369), .ZN(n2746) );
  AND2_X1 U2655 ( .A1(n2051), .A2(n2054), .ZN(n2032) );
  INV_X1 U2656 ( .A(IR_REG_3__SCAN_IN), .ZN(n2200) );
  INV_X1 U2657 ( .A(IR_REG_2__SCAN_IN), .ZN(n2190) );
  AND2_X1 U2658 ( .A1(n2548), .A2(n2547), .ZN(n2033) );
  AND2_X1 U2659 ( .A1(n2275), .A2(n2363), .ZN(n2034) );
  NAND2_X1 U2660 ( .A1(n2182), .A2(n2074), .ZN(n2311) );
  INV_X1 U2661 ( .A(n2311), .ZN(n4339) );
  NOR2_X1 U2662 ( .A1(n2336), .A2(n2335), .ZN(n2035) );
  NOR2_X1 U2663 ( .A1(n3707), .A2(n3105), .ZN(n2036) );
  NAND2_X1 U2664 ( .A1(n2316), .A2(n2858), .ZN(n2037) );
  INV_X1 U2665 ( .A(IR_REG_21__SCAN_IN), .ZN(n2271) );
  AND3_X1 U2666 ( .A1(n2376), .A2(n2151), .A3(n2362), .ZN(n2038) );
  NAND2_X1 U2667 ( .A1(n2088), .A2(n2201), .ZN(n2251) );
  INV_X1 U2668 ( .A(IR_REG_31__SCAN_IN), .ZN(n2365) );
  INV_X1 U2669 ( .A(n3295), .ZN(n3302) );
  NAND2_X1 U2670 ( .A1(n2646), .A2(n3442), .ZN(n2039) );
  NAND2_X1 U2671 ( .A1(n2370), .A2(n2369), .ZN(n2437) );
  INV_X1 U2672 ( .A(IR_REG_28__SCAN_IN), .ZN(n2363) );
  XNOR2_X1 U2673 ( .A(n2299), .B(IR_REG_26__SCAN_IN), .ZN(n2798) );
  NAND2_X1 U2674 ( .A1(n2138), .A2(n2137), .ZN(n3404) );
  AOI22_X1 U2675 ( .A1(n4004), .A2(n3805), .B1(n4014), .B2(n4034), .ZN(n3984)
         );
  INV_X1 U2676 ( .A(IR_REG_29__SCAN_IN), .ZN(n2151) );
  OR2_X1 U2677 ( .A1(n3703), .A2(n3257), .ZN(n2040) );
  INV_X1 U2678 ( .A(IR_REG_9__SCAN_IN), .ZN(n2244) );
  INV_X1 U2679 ( .A(n2169), .ZN(n3994) );
  OR2_X1 U2680 ( .A1(n3528), .A2(n3329), .ZN(n2041) );
  OR2_X1 U2681 ( .A1(n2207), .A2(n2205), .ZN(n2042) );
  AND2_X1 U2682 ( .A1(n2147), .A2(n2145), .ZN(n2043) );
  AND2_X1 U2683 ( .A1(n2041), .A2(n2029), .ZN(n2044) );
  AND2_X1 U2684 ( .A1(n2141), .A2(n2039), .ZN(n2045) );
  NAND2_X1 U2685 ( .A1(n3814), .A2(n3917), .ZN(n2046) );
  INV_X1 U2686 ( .A(n3494), .ZN(n2142) );
  AND2_X1 U2687 ( .A1(n2661), .A2(n2660), .ZN(n3494) );
  INV_X1 U2688 ( .A(n2828), .ZN(n2390) );
  INV_X1 U2689 ( .A(n2539), .ZN(n2095) );
  INV_X1 U2690 ( .A(n3315), .ZN(n3525) );
  INV_X1 U2691 ( .A(n2073), .ZN(n3053) );
  NAND2_X1 U2692 ( .A1(n2474), .A2(n2135), .ZN(n2134) );
  NAND2_X1 U2693 ( .A1(n2134), .A2(n2976), .ZN(n3383) );
  AOI21_X1 U2694 ( .B1(n3148), .B2(n3147), .A(n2175), .ZN(n3166) );
  INV_X1 U2695 ( .A(n3545), .ZN(n2080) );
  AOI21_X1 U2696 ( .B1(n3304), .B2(n3626), .A(n3303), .ZN(n3317) );
  OAI21_X1 U2697 ( .B1(n4450), .B2(n3204), .A(n3203), .ZN(n3258) );
  INV_X1 U2698 ( .A(n3477), .ZN(n2149) );
  INV_X1 U2699 ( .A(n2163), .ZN(n3328) );
  INV_X1 U2700 ( .A(IR_REG_10__SCAN_IN), .ZN(n2245) );
  NOR2_X1 U2701 ( .A1(n3328), .A2(n3797), .ZN(n2166) );
  INV_X1 U2702 ( .A(IR_REG_14__SCAN_IN), .ZN(n2157) );
  INV_X1 U2703 ( .A(IR_REG_15__SCAN_IN), .ZN(n2156) );
  NOR2_X1 U2704 ( .A1(n4365), .A2(n4364), .ZN(n2047) );
  AND2_X1 U2705 ( .A1(n2121), .A2(n2120), .ZN(n2048) );
  NAND2_X1 U2706 ( .A1(n4508), .A2(n2845), .ZN(n3018) );
  AND4_X1 U2707 ( .A1(n2894), .A2(n2893), .A3(n2892), .A4(n2891), .ZN(n2988)
         );
  INV_X1 U2708 ( .A(n2987), .ZN(n4502) );
  NAND2_X1 U2709 ( .A1(n2937), .A2(n2464), .ZN(n2946) );
  NAND2_X1 U2710 ( .A1(n2279), .A2(IR_REG_31__SCAN_IN), .ZN(n2308) );
  NAND2_X1 U2711 ( .A1(n2474), .A2(n2473), .ZN(n2974) );
  NAND2_X1 U2712 ( .A1(n2068), .A2(n2071), .ZN(n3104) );
  AND2_X1 U2713 ( .A1(n2964), .A2(n2968), .ZN(n2965) );
  INV_X1 U2714 ( .A(n2392), .ZN(n4508) );
  INV_X1 U2715 ( .A(IR_REG_0__SCAN_IN), .ZN(n2090) );
  INV_X1 U2716 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2113) );
  NAND2_X1 U2717 ( .A1(n2150), .A2(n2049), .ZN(n2152) );
  AND2_X2 U2718 ( .A1(n2053), .A2(n2046), .ZN(n3888) );
  OR2_X1 U2719 ( .A1(n3952), .A2(n3811), .ZN(n2055) );
  NAND2_X1 U2720 ( .A1(n2995), .A2(n2994), .ZN(n3132) );
  OR2_X1 U2721 ( .A1(n3137), .A2(n3708), .ZN(n2071) );
  OAI21_X2 U2722 ( .B1(n3819), .B2(n2072), .A(n3820), .ZN(n3838) );
  NAND3_X1 U2723 ( .A1(n4495), .A2(n2989), .A3(n2073), .ZN(n3052) );
  NAND2_X1 U2724 ( .A1(n2998), .A2(n4496), .ZN(n4495) );
  AOI21_X1 U2725 ( .B1(n3053), .B2(n2078), .A(n2077), .ZN(n2076) );
  AND2_X2 U2726 ( .A1(n4336), .A2(n2370), .ZN(n2692) );
  NAND2_X1 U2727 ( .A1(n3287), .A2(n3546), .ZN(n2081) );
  OAI21_X1 U2728 ( .B1(n3189), .B2(n3188), .A(n3581), .ZN(n3226) );
  NAND2_X1 U2729 ( .A1(n3189), .A2(n3581), .ZN(n2084) );
  NAND4_X1 U2730 ( .A1(n2034), .A2(n2159), .A3(n2086), .A4(n2162), .ZN(n2367)
         );
  NAND3_X1 U2731 ( .A1(n2103), .A2(n2106), .A3(n2100), .ZN(n4439) );
  NAND3_X1 U2732 ( .A1(n2103), .A2(n2101), .A3(n2100), .ZN(n2108) );
  NAND2_X1 U2733 ( .A1(n4425), .A2(n2262), .ZN(n2266) );
  NOR2_X1 U2734 ( .A1(n2107), .A2(n4541), .ZN(n2105) );
  NAND2_X1 U2735 ( .A1(n2107), .A2(n4541), .ZN(n2106) );
  INV_X1 U2736 ( .A(n2262), .ZN(n2107) );
  INV_X1 U2737 ( .A(n2108), .ZN(n4438) );
  INV_X1 U2738 ( .A(n2115), .ZN(n2920) );
  INV_X1 U2739 ( .A(n2231), .ZN(n2120) );
  NAND2_X1 U2740 ( .A1(n2231), .A2(n2118), .ZN(n2117) );
  INV_X1 U2741 ( .A(n2121), .ZN(n4384) );
  OAI211_X2 U2742 ( .C1(n2388), .C2(IR_REG_20__SCAN_IN), .A(n2124), .B(n2123), 
        .ZN(n2845) );
  NAND2_X1 U2743 ( .A1(n2463), .A2(n2464), .ZN(n2939) );
  NAND2_X1 U2744 ( .A1(n2447), .A2(n2446), .ZN(n2936) );
  NAND2_X1 U2745 ( .A1(n2125), .A2(n2447), .ZN(n2937) );
  AND3_X1 U2746 ( .A1(n2463), .A2(n2446), .A3(n2464), .ZN(n2125) );
  INV_X1 U2747 ( .A(n3384), .ZN(n2133) );
  INV_X1 U2748 ( .A(n2132), .ZN(n2129) );
  OAI22_X1 U2749 ( .A1(n3404), .A2(n3405), .B1(n2674), .B2(n2673), .ZN(n3475)
         );
  NAND2_X1 U2750 ( .A1(n2626), .A2(n2625), .ZN(n3519) );
  AOI21_X1 U2751 ( .B1(n2379), .B2(n2378), .A(n2365), .ZN(n2387) );
  NOR2_X1 U2752 ( .A1(n2252), .A2(n2251), .ZN(n2378) );
  MUX2_X1 U2753 ( .A(REG1_REG_29__SCAN_IN), .B(n2158), .S(n4621), .Z(U3547) );
  MUX2_X1 U2754 ( .A(REG0_REG_29__SCAN_IN), .B(n2158), .S(n4606), .Z(U3515) );
  NAND2_X1 U2755 ( .A1(n4075), .A2(n4076), .ZN(n2158) );
  INV_X1 U2756 ( .A(n2166), .ZN(n4052) );
  NAND2_X1 U2757 ( .A1(n2197), .A2(n2402), .ZN(n2198) );
  NAND2_X1 U2758 ( .A1(n4413), .A2(REG2_REG_14__SCAN_IN), .ZN(n4412) );
  OR2_X1 U2759 ( .A1(n2437), .A2(n2449), .ZN(n2450) );
  NAND2_X1 U2760 ( .A1(n2442), .A2(n2441), .ZN(n2444) );
  NAND2_X1 U2761 ( .A1(n3100), .A2(n3099), .ZN(n3159) );
  NOR2_X1 U2762 ( .A1(n4376), .A2(n4375), .ZN(n4374) );
  NAND2_X1 U2763 ( .A1(n4027), .A2(n4019), .ZN(n4018) );
  MUX2_X1 U2764 ( .A(n2188), .B(DATAI_2_), .S(n2454), .Z(n3055) );
  NOR2_X1 U2765 ( .A1(n4354), .A2(n4355), .ZN(n4353) );
  XNOR2_X1 U2766 ( .A(n2440), .B(n2793), .ZN(n2443) );
  AND2_X1 U2767 ( .A1(n2351), .A2(n2350), .ZN(n2170) );
  AND2_X1 U2768 ( .A1(n2170), .A2(n2360), .ZN(n2171) );
  OR2_X1 U2769 ( .A1(n4351), .A2(n3723), .ZN(n4431) );
  INV_X1 U2770 ( .A(n4431), .ZN(n2349) );
  AND2_X1 U2771 ( .A1(n2204), .A2(n2203), .ZN(n4338) );
  INV_X1 U2772 ( .A(n4338), .ZN(n2207) );
  OR2_X1 U2773 ( .A1(n2255), .A2(n2580), .ZN(n2172) );
  OR2_X1 U2774 ( .A1(n4544), .A2(n4131), .ZN(n2173) );
  AND4_X1 U2775 ( .A1(n2640), .A2(n2639), .A3(n2638), .A4(n2637), .ZN(n4036)
         );
  AND2_X1 U2776 ( .A1(n3821), .A2(n3841), .ZN(n2174) );
  NOR2_X1 U2777 ( .A1(n3146), .A2(n3621), .ZN(n2175) );
  OAI211_X1 U2778 ( .C1(n3862), .C2(n2023), .A(n2775), .B(n2774), .ZN(n3831)
         );
  AND4_X1 U2779 ( .A1(n2623), .A2(n2622), .A3(n2621), .A4(n2620), .ZN(n3528)
         );
  INV_X1 U2780 ( .A(n2603), .ZN(n2257) );
  INV_X1 U2781 ( .A(n3797), .ZN(n3329) );
  AND2_X1 U2782 ( .A1(n2826), .A2(n3523), .ZN(n2176) );
  INV_X1 U2783 ( .A(n3851), .ZN(n3860) );
  AND2_X1 U2784 ( .A1(n3852), .A2(n3871), .ZN(n2177) );
  AND2_X1 U2785 ( .A1(n3443), .A2(n2645), .ZN(n2178) );
  OR2_X1 U2786 ( .A1(n2319), .A2(n4556), .ZN(n2179) );
  INV_X1 U2787 ( .A(n4033), .ZN(n4029) );
  AND2_X1 U2788 ( .A1(n2557), .A2(REG2_REG_11__SCAN_IN), .ZN(n2180) );
  INV_X1 U2789 ( .A(n2557), .ZN(n4549) );
  INV_X1 U2790 ( .A(IR_REG_22__SCAN_IN), .ZN(n2276) );
  OAI22_X1 U2791 ( .A1(n2988), .A2(n2496), .B1(n2439), .B2(n4502), .ZN(n2440)
         );
  INV_X1 U2792 ( .A(n3396), .ZN(n2735) );
  NAND2_X1 U2793 ( .A1(n3710), .A2(n2427), .ZN(n2442) );
  AND2_X1 U2794 ( .A1(n2274), .A2(n2377), .ZN(n2275) );
  NAND2_X1 U2795 ( .A1(n3137), .A2(n2393), .ZN(n2417) );
  AND2_X1 U2796 ( .A1(n2590), .A2(n2591), .ZN(n3239) );
  INV_X1 U2797 ( .A(n2758), .ZN(n2757) );
  NAND2_X1 U2798 ( .A1(n2743), .A2(REG3_REG_25__SCAN_IN), .ZN(n2758) );
  INV_X1 U2799 ( .A(n2498), .ZN(n2781) );
  OR2_X1 U2800 ( .A1(n2437), .A2(n2395), .ZN(n2401) );
  NAND2_X1 U2801 ( .A1(n2317), .A2(n2402), .ZN(n2318) );
  NAND2_X1 U2802 ( .A1(n2757), .A2(REG3_REG_26__SCAN_IN), .ZN(n2772) );
  OR2_X1 U2803 ( .A1(n2729), .A2(n4187), .ZN(n2744) );
  INV_X1 U2804 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2549) );
  NAND2_X1 U2805 ( .A1(n2522), .A2(REG3_REG_9__SCAN_IN), .ZN(n2532) );
  MUX2_X1 U2806 ( .A(n2402), .B(DATAI_4_), .S(n2454), .Z(n3043) );
  INV_X1 U2807 ( .A(n2387), .ZN(n2381) );
  AND2_X1 U2808 ( .A1(n2693), .A2(REG3_REG_21__SCAN_IN), .ZN(n2707) );
  OR2_X1 U2809 ( .A1(n2663), .A2(n2662), .ZN(n2676) );
  INV_X1 U2810 ( .A(n3055), .ZN(n3062) );
  AND2_X1 U2811 ( .A1(n2847), .A2(n4057), .ZN(n3526) );
  OR2_X1 U2812 ( .A1(n3426), .A2(n2023), .ZN(n2750) );
  AND4_X1 U2813 ( .A1(n2401), .A2(n2400), .A3(n2399), .A4(n2398), .ZN(n2948)
         );
  NOR2_X1 U2814 ( .A1(n2914), .A2(n2915), .ZN(n2913) );
  NAND2_X1 U2815 ( .A1(n2244), .A2(n2223), .ZN(n2242) );
  INV_X1 U2816 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3529) );
  AND4_X1 U2817 ( .A1(n2700), .A2(n2699), .A3(n2698), .A4(n2697), .ZN(n3990)
         );
  NAND2_X1 U2818 ( .A1(n4036), .A2(n4055), .ZN(n3802) );
  OR2_X1 U2819 ( .A1(n2550), .A2(n2549), .ZN(n2566) );
  OAI21_X1 U2820 ( .B1(n3068), .B2(n2993), .A(n2992), .ZN(n3026) );
  OR2_X1 U2821 ( .A1(n2881), .A2(D_REG_0__SCAN_IN), .ZN(n2803) );
  NAND2_X1 U2822 ( .A1(n2384), .A2(n4535), .ZN(n2889) );
  NOR2_X1 U2823 ( .A1(n2251), .A2(IR_REG_5__SCAN_IN), .ZN(n2221) );
  OR2_X1 U2824 ( .A1(n2717), .A2(n3399), .ZN(n2729) );
  INV_X1 U2825 ( .A(n3527), .ZN(n3499) );
  INV_X1 U2826 ( .A(n3526), .ZN(n3500) );
  NAND2_X1 U2827 ( .A1(n2475), .A2(REG3_REG_6__SCAN_IN), .ZN(n2507) );
  AND2_X1 U2828 ( .A1(n2835), .A2(STATE_REG_SCAN_IN), .ZN(n3514) );
  AND4_X1 U2829 ( .A1(n2734), .A2(n2733), .A3(n2732), .A4(n2731), .ZN(n3814)
         );
  AND4_X1 U2830 ( .A1(n2653), .A2(n2652), .A3(n2651), .A4(n2650), .ZN(n4047)
         );
  AND4_X1 U2831 ( .A1(n2556), .A2(n2555), .A3(n2554), .A4(n2553), .ZN(n3228)
         );
  INV_X1 U2832 ( .A(n3369), .ZN(n3170) );
  OAI21_X1 U2833 ( .B1(n2341), .B2(n4442), .A(n2340), .ZN(n2342) );
  AND2_X1 U2834 ( .A1(n4508), .A2(n3690), .ZN(n4489) );
  OR2_X1 U2835 ( .A1(n2889), .A2(n3012), .ZN(n4057) );
  AND2_X1 U2836 ( .A1(n4621), .A2(n4596), .ZN(n4079) );
  AND2_X1 U2837 ( .A1(n2803), .A2(n2802), .ZN(n3020) );
  INV_X1 U2838 ( .A(n3813), .ZN(n3917) );
  INV_X1 U2839 ( .A(n3018), .ZN(n4596) );
  AND2_X1 U2840 ( .A1(n4510), .A2(n2828), .ZN(n4603) );
  INV_X1 U2841 ( .A(IR_REG_30__SCAN_IN), .ZN(n3346) );
  AND2_X1 U2842 ( .A1(n2234), .A2(n2235), .ZN(n2557) );
  INV_X1 U2843 ( .A(n2402), .ZN(n3751) );
  AND2_X1 U2844 ( .A1(n2339), .A2(n2338), .ZN(n4435) );
  NAND2_X1 U2845 ( .A1(n2849), .A2(n2820), .ZN(n3517) );
  INV_X1 U2846 ( .A(n3854), .ZN(n3821) );
  OAI211_X1 U2847 ( .C1(n2839), .C2(n3883), .A(n2763), .B(n2762), .ZN(n3852)
         );
  INV_X1 U2848 ( .A(n3528), .ZN(n4049) );
  OR2_X1 U2849 ( .A1(n2225), .A2(n2224), .ZN(n3122) );
  INV_X1 U2850 ( .A(n2342), .ZN(n2343) );
  INV_X1 U2851 ( .A(n3878), .ZN(n4063) );
  NAND2_X1 U2852 ( .A1(n3032), .A2(n4057), .ZN(n4519) );
  INV_X1 U2853 ( .A(n4079), .ZN(n4133) );
  INV_X1 U2854 ( .A(n4148), .ZN(n4331) );
  INV_X1 U2855 ( .A(n4606), .ZN(n4604) );
  INV_X1 U2856 ( .A(n4530), .ZN(n4534) );
  AND2_X1 U2857 ( .A1(n2301), .A2(STATE_REG_SCAN_IN), .ZN(n4535) );
  AND2_X1 U2858 ( .A1(n2254), .A2(n2253), .ZN(n4337) );
  INV_X1 U2859 ( .A(n3726), .ZN(U4043) );
  NAND2_X1 U2860 ( .A1(n2344), .A2(n2343), .ZN(U3257) );
  INV_X2 U2861 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U2862 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4376) );
  NAND2_X1 U2863 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2181)
         );
  INV_X1 U2864 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2183) );
  NAND2_X1 U2865 ( .A1(n4339), .A2(n2183), .ZN(n2185) );
  NAND2_X1 U2866 ( .A1(n2185), .A2(n2184), .ZN(n3717) );
  NAND2_X1 U2867 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3729) );
  INV_X1 U2868 ( .A(n3729), .ZN(n3716) );
  NAND2_X1 U2869 ( .A1(n3717), .A2(n3716), .ZN(n3715) );
  NAND2_X1 U2870 ( .A1(n4339), .A2(REG2_REG_1__SCAN_IN), .ZN(n2186) );
  NAND2_X1 U2871 ( .A1(n3715), .A2(n2186), .ZN(n3736) );
  INV_X1 U2872 ( .A(REG2_REG_2__SCAN_IN), .ZN(n4192) );
  MUX2_X1 U2873 ( .A(REG2_REG_2__SCAN_IN), .B(n4192), .S(n2188), .Z(n3737) );
  NAND2_X1 U2874 ( .A1(n3736), .A2(n3737), .ZN(n3735) );
  NAND2_X1 U2875 ( .A1(n2188), .A2(REG2_REG_2__SCAN_IN), .ZN(n2189) );
  NAND2_X1 U2876 ( .A1(n3735), .A2(n2189), .ZN(n2192) );
  NAND2_X1 U2877 ( .A1(n2191), .A2(IR_REG_31__SCAN_IN), .ZN(n2194) );
  INV_X1 U2878 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2915) );
  AND2_X1 U2879 ( .A1(n2192), .A2(n2858), .ZN(n2193) );
  NAND2_X1 U2880 ( .A1(n2194), .A2(n2200), .ZN(n2195) );
  NAND2_X1 U2881 ( .A1(n2195), .A2(IR_REG_31__SCAN_IN), .ZN(n2196) );
  XNOR2_X1 U2882 ( .A(n2196), .B(IR_REG_4__SCAN_IN), .ZN(n2402) );
  INV_X1 U2883 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2205) );
  NAND2_X1 U2884 ( .A1(n2251), .A2(IR_REG_31__SCAN_IN), .ZN(n2202) );
  MUX2_X1 U2885 ( .A(n2202), .B(IR_REG_31__SCAN_IN), .S(n2246), .Z(n2204) );
  INV_X1 U2886 ( .A(n2221), .ZN(n2203) );
  MUX2_X1 U2887 ( .A(REG2_REG_5__SCAN_IN), .B(n2205), .S(n4338), .Z(n2206) );
  INV_X1 U2888 ( .A(n2206), .ZN(n2921) );
  OR2_X1 U2889 ( .A1(n2221), .A2(n2365), .ZN(n2208) );
  XNOR2_X1 U2890 ( .A(n2208), .B(IR_REG_6__SCAN_IN), .ZN(n2480) );
  INV_X1 U2891 ( .A(n2480), .ZN(n4556) );
  NOR2_X1 U2892 ( .A1(n2026), .A2(n4556), .ZN(n2209) );
  XNOR2_X1 U2893 ( .A(n2026), .B(n4556), .ZN(n4354) );
  INV_X1 U2894 ( .A(REG2_REG_6__SCAN_IN), .ZN(n4355) );
  INV_X1 U2895 ( .A(IR_REG_6__SCAN_IN), .ZN(n2210) );
  NAND2_X1 U2896 ( .A1(n2221), .A2(n2210), .ZN(n2211) );
  NAND2_X1 U2897 ( .A1(n2211), .A2(IR_REG_31__SCAN_IN), .ZN(n2214) );
  XNOR2_X1 U2898 ( .A(n2214), .B(IR_REG_7__SCAN_IN), .ZN(n4368) );
  NAND2_X1 U2899 ( .A1(n4368), .A2(REG2_REG_7__SCAN_IN), .ZN(n2212) );
  OAI21_X1 U2900 ( .B1(n4368), .B2(REG2_REG_7__SCAN_IN), .A(n2212), .ZN(n4364)
         );
  INV_X1 U2901 ( .A(IR_REG_7__SCAN_IN), .ZN(n2213) );
  NAND2_X1 U2902 ( .A1(n2214), .A2(n2213), .ZN(n2215) );
  NAND2_X1 U2903 ( .A1(n2215), .A2(IR_REG_31__SCAN_IN), .ZN(n2216) );
  XNOR2_X1 U2904 ( .A(n2216), .B(IR_REG_8__SCAN_IN), .ZN(n2513) );
  INV_X1 U2905 ( .A(n2513), .ZN(n4552) );
  NOR2_X1 U2906 ( .A1(n2217), .A2(n4552), .ZN(n2218) );
  NOR2_X1 U2907 ( .A1(n4374), .A2(n2218), .ZN(n3118) );
  INV_X1 U2908 ( .A(IR_REG_8__SCAN_IN), .ZN(n2219) );
  AND2_X1 U2909 ( .A1(n2247), .A2(n2219), .ZN(n2220) );
  NOR2_X1 U2910 ( .A1(n2223), .A2(n2365), .ZN(n2222) );
  MUX2_X1 U2911 ( .A(n2365), .B(n2222), .S(IR_REG_9__SCAN_IN), .Z(n2225) );
  INV_X1 U2912 ( .A(n2242), .ZN(n2224) );
  NAND2_X1 U2913 ( .A1(n2528), .A2(REG2_REG_9__SCAN_IN), .ZN(n2227) );
  INV_X1 U2914 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3160) );
  NAND2_X1 U2915 ( .A1(n3122), .A2(n3160), .ZN(n2226) );
  NAND2_X1 U2916 ( .A1(n2227), .A2(n2226), .ZN(n3117) );
  NAND2_X1 U2917 ( .A1(n2242), .A2(IR_REG_31__SCAN_IN), .ZN(n2228) );
  XNOR2_X1 U2918 ( .A(n2228), .B(IR_REG_10__SCAN_IN), .ZN(n2539) );
  INV_X1 U2919 ( .A(REG2_REG_10__SCAN_IN), .ZN(n4386) );
  INV_X1 U2920 ( .A(n2229), .ZN(n2230) );
  NOR2_X1 U2921 ( .A1(n2230), .A2(n2095), .ZN(n2231) );
  NAND2_X1 U2922 ( .A1(n2232), .A2(IR_REG_31__SCAN_IN), .ZN(n2233) );
  OR2_X1 U2923 ( .A1(n2233), .A2(n2240), .ZN(n2234) );
  NAND2_X1 U2924 ( .A1(n2233), .A2(n2240), .ZN(n2235) );
  INV_X1 U2925 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4252) );
  AOI22_X1 U2926 ( .A1(n2557), .A2(n4252), .B1(REG2_REG_11__SCAN_IN), .B2(
        n4549), .ZN(n4394) );
  NAND2_X1 U2927 ( .A1(n2235), .A2(IR_REG_31__SCAN_IN), .ZN(n2236) );
  XNOR2_X1 U2928 ( .A(n2236), .B(IR_REG_12__SCAN_IN), .ZN(n2572) );
  INV_X1 U2929 ( .A(n2572), .ZN(n4547) );
  NOR2_X1 U2930 ( .A1(n2237), .A2(n4547), .ZN(n2238) );
  INV_X1 U2931 ( .A(REG2_REG_12__SCAN_IN), .ZN(n4405) );
  XNOR2_X1 U2932 ( .A(n4547), .B(n2237), .ZN(n4404) );
  INV_X1 U2933 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3268) );
  INV_X1 U2934 ( .A(IR_REG_12__SCAN_IN), .ZN(n2239) );
  NAND3_X1 U2935 ( .A1(n2240), .A2(n2245), .A3(n2239), .ZN(n2241) );
  OAI21_X1 U2936 ( .B1(n2242), .B2(n2241), .A(IR_REG_31__SCAN_IN), .ZN(n2243)
         );
  MUX2_X1 U2937 ( .A(IR_REG_31__SCAN_IN), .B(n2243), .S(IR_REG_13__SCAN_IN), 
        .Z(n2254) );
  INV_X1 U2938 ( .A(n2378), .ZN(n2253) );
  INV_X1 U2939 ( .A(n4337), .ZN(n2255) );
  OR2_X1 U2940 ( .A1(n2378), .A2(n2365), .ZN(n2256) );
  XNOR2_X1 U2941 ( .A(n2256), .B(IR_REG_14__SCAN_IN), .ZN(n2603) );
  NAND2_X1 U2942 ( .A1(n2603), .A2(n2258), .ZN(n2259) );
  NAND2_X1 U2943 ( .A1(n4412), .A2(n2259), .ZN(n4427) );
  NAND2_X1 U2944 ( .A1(n2378), .A2(n2157), .ZN(n2260) );
  NAND2_X1 U2945 ( .A1(n2260), .A2(IR_REG_31__SCAN_IN), .ZN(n2263) );
  XNOR2_X1 U2946 ( .A(n2263), .B(IR_REG_15__SCAN_IN), .ZN(n2614) );
  INV_X1 U2947 ( .A(n2614), .ZN(n4544) );
  INV_X1 U2948 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2261) );
  AOI22_X1 U2949 ( .A1(REG2_REG_15__SCAN_IN), .A2(n2614), .B1(n4544), .B2(
        n2261), .ZN(n4428) );
  NAND2_X1 U2950 ( .A1(n4427), .A2(n4428), .ZN(n4425) );
  NAND2_X1 U2951 ( .A1(REG2_REG_15__SCAN_IN), .A2(n2614), .ZN(n2262) );
  NAND2_X1 U2952 ( .A1(n2263), .A2(n2156), .ZN(n2264) );
  NAND2_X1 U2953 ( .A1(n2264), .A2(IR_REG_31__SCAN_IN), .ZN(n2265) );
  XNOR2_X1 U2954 ( .A(n2265), .B(IR_REG_16__SCAN_IN), .ZN(n4541) );
  NAND2_X1 U2955 ( .A1(n2378), .A2(n2273), .ZN(n2267) );
  NAND2_X1 U2956 ( .A1(n2267), .A2(IR_REG_31__SCAN_IN), .ZN(n2268) );
  XNOR2_X1 U2957 ( .A(n2268), .B(IR_REG_17__SCAN_IN), .ZN(n2641) );
  INV_X1 U2958 ( .A(n2641), .ZN(n4540) );
  INV_X1 U2959 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2352) );
  AOI22_X1 U2960 ( .A1(REG2_REG_17__SCAN_IN), .A2(n4540), .B1(n2641), .B2(
        n2352), .ZN(n2269) );
  AOI21_X1 U2961 ( .B1(n2270), .B2(n2269), .A(n2354), .ZN(n2309) );
  AND2_X1 U2962 ( .A1(n2304), .A2(n2303), .ZN(n2277) );
  NAND2_X1 U2963 ( .A1(n2305), .A2(n2278), .ZN(n2279) );
  NAND2_X1 U2964 ( .A1(n2363), .A2(IR_REG_27__SCAN_IN), .ZN(n2280) );
  OR2_X2 U2965 ( .A1(n2295), .A2(n2365), .ZN(n2284) );
  INV_X1 U2966 ( .A(IR_REG_23__SCAN_IN), .ZN(n2283) );
  NAND2_X1 U2967 ( .A1(n2284), .A2(n2283), .ZN(n2292) );
  OR2_X1 U2968 ( .A1(n2284), .A2(n2283), .ZN(n2285) );
  NAND2_X1 U2969 ( .A1(n2292), .A2(n2285), .ZN(n2301) );
  INV_X1 U2970 ( .A(n2305), .ZN(n2289) );
  NAND2_X1 U2971 ( .A1(n2289), .A2(IR_REG_31__SCAN_IN), .ZN(n2286) );
  NAND2_X1 U2972 ( .A1(n2378), .A2(n2364), .ZN(n2287) );
  NAND2_X1 U2973 ( .A1(n2287), .A2(IR_REG_31__SCAN_IN), .ZN(n2288) );
  AND2_X1 U2974 ( .A1(n2390), .A2(n3687), .ZN(n3008) );
  NAND2_X1 U2975 ( .A1(n2301), .A2(n3008), .ZN(n2291) );
  AND2_X1 U2976 ( .A1(n3349), .A2(n2291), .ZN(n2337) );
  NAND2_X1 U2977 ( .A1(n2292), .A2(IR_REG_31__SCAN_IN), .ZN(n2294) );
  INV_X1 U2978 ( .A(IR_REG_24__SCAN_IN), .ZN(n2293) );
  NAND2_X1 U2979 ( .A1(n2295), .A2(n2303), .ZN(n2298) );
  NAND2_X1 U2980 ( .A1(n2298), .A2(IR_REG_31__SCAN_IN), .ZN(n2297) );
  INV_X1 U2981 ( .A(IR_REG_25__SCAN_IN), .ZN(n2296) );
  NOR2_X1 U2982 ( .A1(n2799), .A2(n2884), .ZN(n2300) );
  NAND2_X1 U2983 ( .A1(n2300), .A2(n2798), .ZN(n2384) );
  INV_X1 U2984 ( .A(n2384), .ZN(n2428) );
  INV_X1 U2985 ( .A(n2301), .ZN(n2832) );
  NAND2_X1 U2986 ( .A1(n2832), .A2(STATE_REG_SCAN_IN), .ZN(n3697) );
  NAND2_X1 U2987 ( .A1(n2889), .A2(n3697), .ZN(n2338) );
  NAND2_X1 U2988 ( .A1(n2337), .A2(n2338), .ZN(n4351) );
  AND2_X1 U2989 ( .A1(n2305), .A2(n2362), .ZN(n2306) );
  OR2_X1 U2990 ( .A1(n2306), .A2(n2365), .ZN(n2307) );
  XNOR2_X1 U2991 ( .A(n2307), .B(n2363), .ZN(n4341) );
  XNOR2_X1 U2992 ( .A(n2308), .B(IR_REG_27__SCAN_IN), .ZN(n4348) );
  INV_X1 U2993 ( .A(n4348), .ZN(n3722) );
  OR2_X1 U2994 ( .A1(n4341), .A2(n3722), .ZN(n3730) );
  NOR2_X1 U2995 ( .A1(n4351), .A2(n3730), .ZN(n4426) );
  INV_X1 U2996 ( .A(n4341), .ZN(n3723) );
  OAI22_X1 U2997 ( .A1(n2309), .A2(n4440), .B1(n4540), .B2(n4431), .ZN(n2310)
         );
  NAND2_X1 U2998 ( .A1(n2528), .A2(REG1_REG_9__SCAN_IN), .ZN(n2323) );
  INV_X1 U2999 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2521) );
  MUX2_X1 U3000 ( .A(n2521), .B(REG1_REG_9__SCAN_IN), .S(n3122), .Z(n3113) );
  INV_X1 U3001 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4608) );
  AND2_X1 U3002 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3713)
         );
  NAND2_X1 U3003 ( .A1(n3714), .A2(n3713), .ZN(n3712) );
  NAND2_X1 U3004 ( .A1(n4339), .A2(REG1_REG_1__SCAN_IN), .ZN(n2314) );
  NAND2_X1 U3005 ( .A1(n3712), .A2(n2314), .ZN(n3739) );
  INV_X1 U3006 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4610) );
  NAND2_X1 U3007 ( .A1(n2188), .A2(REG1_REG_2__SCAN_IN), .ZN(n2315) );
  INV_X1 U3008 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4612) );
  INV_X1 U3009 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2412) );
  MUX2_X1 U3010 ( .A(n2412), .B(REG1_REG_5__SCAN_IN), .S(n4338), .Z(n2926) );
  NOR2_X1 U3011 ( .A1(n2925), .A2(n2926), .ZN(n2924) );
  AOI21_X1 U3012 ( .B1(n4338), .B2(REG1_REG_5__SCAN_IN), .A(n2924), .ZN(n2319)
         );
  XNOR2_X1 U3013 ( .A(n2319), .B(n4556), .ZN(n4359) );
  INV_X1 U3014 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4360) );
  INV_X1 U3015 ( .A(n4358), .ZN(n2320) );
  INV_X1 U3016 ( .A(n4368), .ZN(n4554) );
  NAND2_X1 U3017 ( .A1(n2513), .A2(n2321), .ZN(n2322) );
  NAND2_X1 U3018 ( .A1(REG1_REG_8__SCAN_IN), .A2(n4381), .ZN(n4380) );
  NAND2_X1 U3019 ( .A1(n2322), .A2(n4380), .ZN(n3114) );
  NAND2_X1 U3020 ( .A1(n3113), .A2(n3114), .ZN(n3112) );
  NAND2_X1 U3021 ( .A1(n2323), .A2(n3112), .ZN(n2324) );
  NAND2_X1 U3022 ( .A1(n2539), .A2(n2324), .ZN(n2325) );
  INV_X1 U3023 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4619) );
  AOI22_X1 U3024 ( .A1(n2557), .A2(REG1_REG_11__SCAN_IN), .B1(n4619), .B2(
        n4549), .ZN(n4400) );
  NAND2_X1 U3025 ( .A1(n2572), .A2(n2327), .ZN(n2328) );
  XNOR2_X1 U3026 ( .A(n4337), .B(REG1_REG_13__SCAN_IN), .ZN(n3335) );
  INV_X1 U3027 ( .A(REG1_REG_13__SCAN_IN), .ZN(n2580) );
  NAND2_X1 U3028 ( .A1(n2603), .A2(n2331), .ZN(n2332) );
  INV_X1 U3029 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U3030 ( .A1(REG1_REG_15__SCAN_IN), .A2(n2614), .B1(n4544), .B2(
        n4131), .ZN(n4424) );
  XNOR2_X1 U3031 ( .A(n2333), .B(n4541), .ZN(n4437) );
  NOR2_X1 U3032 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4437), .ZN(n4436) );
  NOR2_X1 U3033 ( .A1(n4541), .A2(n2333), .ZN(n2334) );
  INV_X1 U3034 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4123) );
  AOI22_X1 U3035 ( .A1(REG1_REG_17__SCAN_IN), .A2(n4540), .B1(n2641), .B2(
        n4123), .ZN(n2335) );
  AOI21_X1 U3036 ( .B1(n2336), .B2(n2335), .A(n2035), .ZN(n2341) );
  OR2_X1 U3037 ( .A1(n4351), .A2(n4348), .ZN(n4442) );
  INV_X1 U3038 ( .A(n2337), .ZN(n2339) );
  AND2_X1 U3039 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n3446) );
  NAND2_X1 U3040 ( .A1(n2378), .A2(n2376), .ZN(n2345) );
  NAND2_X1 U3041 ( .A1(n2345), .A2(IR_REG_31__SCAN_IN), .ZN(n2346) );
  XNOR2_X1 U3042 ( .A(n2346), .B(IR_REG_18__SCAN_IN), .ZN(n2654) );
  INV_X1 U3043 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3762) );
  INV_X1 U3044 ( .A(n2654), .ZN(n4538) );
  AOI22_X1 U3045 ( .A1(n2654), .A2(REG1_REG_18__SCAN_IN), .B1(n3762), .B2(
        n4538), .ZN(n2347) );
  OAI211_X1 U3046 ( .C1(n2348), .C2(n2347), .A(n3761), .B(n4422), .ZN(n2351)
         );
  NAND2_X1 U3047 ( .A1(n2349), .A2(n2654), .ZN(n2350) );
  NOR2_X1 U3048 ( .A1(n2354), .A2(n2353), .ZN(n2355) );
  INV_X1 U3049 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4263) );
  AOI22_X1 U3050 ( .A1(n2654), .A2(REG2_REG_18__SCAN_IN), .B1(n4263), .B2(
        n4538), .ZN(n2356) );
  NAND2_X1 U3051 ( .A1(n2355), .A2(n2356), .ZN(n3758) );
  INV_X1 U3052 ( .A(n2355), .ZN(n2358) );
  INV_X1 U3053 ( .A(n2356), .ZN(n2357) );
  NAND2_X1 U3054 ( .A1(n2358), .A2(n2357), .ZN(n2359) );
  NAND3_X1 U3055 ( .A1(n3758), .A2(n2359), .A3(n4426), .ZN(n2360) );
  INV_X1 U3056 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4261) );
  NOR2_X1 U3057 ( .A1(STATE_REG_SCAN_IN), .A2(n4261), .ZN(n3497) );
  AOI21_X1 U3058 ( .B1(n4435), .B2(ADDR_REG_18__SCAN_IN), .A(n3497), .ZN(n2361) );
  NAND2_X1 U3059 ( .A1(n2171), .A2(n2361), .ZN(U3258) );
  NAND2_X1 U3060 ( .A1(n2367), .A2(IR_REG_31__SCAN_IN), .ZN(n2368) );
  NAND2_X1 U3061 ( .A1(n2692), .A2(REG1_REG_3__SCAN_IN), .ZN(n2375) );
  OR2_X1 U3062 ( .A1(n2023), .A2(REG3_REG_3__SCAN_IN), .ZN(n2374) );
  OR2_X1 U3063 ( .A1(n2746), .A2(n2915), .ZN(n2373) );
  INV_X1 U3064 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2371) );
  OR2_X1 U3065 ( .A1(n2437), .A2(n2371), .ZN(n2372) );
  AND2_X1 U3066 ( .A1(n2377), .A2(n2376), .ZN(n2379) );
  INV_X1 U3067 ( .A(IR_REG_19__SCAN_IN), .ZN(n2380) );
  INV_X1 U3068 ( .A(IR_REG_20__SCAN_IN), .ZN(n2382) );
  NAND2_X1 U3069 ( .A1(n2384), .A2(n2383), .ZN(n2496) );
  NAND2_X1 U3070 ( .A1(n3056), .A2(n2456), .ZN(n2386) );
  MUX2_X1 U3071 ( .A(n2858), .B(DATAI_3_), .S(n2454), .Z(n3558) );
  NAND2_X1 U3072 ( .A1(n3558), .A2(n2393), .ZN(n2385) );
  NAND2_X1 U3073 ( .A1(n2386), .A2(n2385), .ZN(n2391) );
  NAND2_X1 U3074 ( .A1(n2387), .A2(IR_REG_19__SCAN_IN), .ZN(n2389) );
  NAND2_X1 U3075 ( .A1(n2390), .A2(n3768), .ZN(n2840) );
  XNOR2_X1 U3076 ( .A(n2391), .B(n2778), .ZN(n2466) );
  INV_X1 U3077 ( .A(n2466), .ZN(n2394) );
  INV_X1 U3078 ( .A(n3687), .ZN(n2829) );
  NAND2_X1 U3079 ( .A1(n2829), .A2(n2828), .ZN(n2392) );
  INV_X1 U3080 ( .A(n2498), .ZN(n2427) );
  AOI22_X1 U3081 ( .A1(n3056), .A2(n2427), .B1(n2456), .B2(n3558), .ZN(n2465)
         );
  NAND2_X1 U3082 ( .A1(n2394), .A2(n2465), .ZN(n2964) );
  INV_X1 U3083 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2395) );
  INV_X1 U3084 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2396) );
  OR2_X1 U3085 ( .A1(n2397), .A2(n2396), .ZN(n2400) );
  XNOR2_X1 U3086 ( .A(REG3_REG_4__SCAN_IN), .B(REG3_REG_3__SCAN_IN), .ZN(n3045) );
  OR2_X1 U3087 ( .A1(n2023), .A2(n3045), .ZN(n2399) );
  OR2_X1 U3088 ( .A1(n2746), .A2(n2113), .ZN(n2398) );
  INV_X1 U3089 ( .A(n3043), .ZN(n2970) );
  XNOR2_X1 U3090 ( .A(n2403), .B(n2793), .ZN(n2406) );
  OR2_X1 U3091 ( .A1(n2948), .A2(n2498), .ZN(n2405) );
  NAND2_X1 U3092 ( .A1(n3043), .A2(n2456), .ZN(n2404) );
  NAND2_X1 U3093 ( .A1(n2405), .A2(n2404), .ZN(n2407) );
  XNOR2_X1 U3094 ( .A(n2406), .B(n2407), .ZN(n2968) );
  INV_X1 U3095 ( .A(n2406), .ZN(n2408) );
  NAND2_X1 U3096 ( .A1(n2408), .A2(n2407), .ZN(n2467) );
  INV_X1 U3097 ( .A(n2467), .ZN(n2409) );
  OR2_X1 U3098 ( .A1(n2965), .A2(n2409), .ZN(n2954) );
  AOI21_X1 U3099 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        REG3_REG_5__SCAN_IN), .ZN(n2410) );
  NOR2_X1 U3100 ( .A1(n2410), .A2(n2475), .ZN(n3141) );
  NAND2_X1 U3101 ( .A1(n2025), .A2(n3141), .ZN(n2416) );
  INV_X1 U3102 ( .A(REG0_REG_5__SCAN_IN), .ZN(n2411) );
  OR2_X1 U3103 ( .A1(n2437), .A2(n2411), .ZN(n2415) );
  OR2_X1 U3104 ( .A1(n2397), .A2(n2412), .ZN(n2414) );
  OR2_X1 U3105 ( .A1(n2746), .A2(n2205), .ZN(n2413) );
  NAND2_X1 U3106 ( .A1(n3708), .A2(n2456), .ZN(n2418) );
  MUX2_X1 U3107 ( .A(n4338), .B(DATAI_5_), .S(n3349), .Z(n3137) );
  NAND2_X1 U3108 ( .A1(n2418), .A2(n2417), .ZN(n2419) );
  AOI22_X1 U3109 ( .A1(n3708), .A2(n2781), .B1(n2456), .B2(n3137), .ZN(n2470)
         );
  XNOR2_X1 U3110 ( .A(n2472), .B(n2470), .ZN(n2956) );
  AND2_X1 U3111 ( .A1(n2954), .A2(n2956), .ZN(n2469) );
  NAND2_X1 U3112 ( .A1(n2692), .A2(REG1_REG_0__SCAN_IN), .ZN(n2426) );
  INV_X1 U3113 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2420) );
  OR2_X1 U3114 ( .A1(n2023), .A2(n2420), .ZN(n2425) );
  INV_X1 U3115 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2421) );
  OR2_X1 U3116 ( .A1(n2746), .A2(n2421), .ZN(n2424) );
  INV_X1 U3117 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2422) );
  OR2_X1 U3118 ( .A1(n2437), .A2(n2422), .ZN(n2423) );
  NAND2_X1 U3119 ( .A1(n3711), .A2(n2427), .ZN(n2430) );
  MUX2_X1 U3120 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2454), .Z(n2999) );
  AOI22_X1 U3121 ( .A1(n2999), .A2(n2456), .B1(n2428), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2429) );
  NAND2_X1 U3122 ( .A1(n2430), .A2(n2429), .ZN(n2887) );
  INV_X1 U3123 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2432) );
  NAND2_X1 U3124 ( .A1(n3711), .A2(n2456), .ZN(n2431) );
  NAND2_X1 U3125 ( .A1(n2999), .A2(n2393), .ZN(n2433) );
  NAND2_X1 U3126 ( .A1(n2887), .A2(n2886), .ZN(n2435) );
  NAND2_X1 U3127 ( .A1(n2433), .A2(n2793), .ZN(n2434) );
  NAND2_X1 U3128 ( .A1(n2435), .A2(n2434), .ZN(n2931) );
  INV_X1 U3129 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2436) );
  OR2_X1 U3130 ( .A1(n2437), .A2(n2436), .ZN(n2894) );
  OR2_X1 U3131 ( .A1(n2746), .A2(n2183), .ZN(n2892) );
  INV_X1 U3132 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2438) );
  OR2_X1 U3133 ( .A1(n2023), .A2(n2438), .ZN(n2891) );
  MUX2_X1 U3134 ( .A(n4339), .B(DATAI_1_), .S(n2454), .Z(n2987) );
  NAND2_X1 U3135 ( .A1(n2987), .A2(n2456), .ZN(n2441) );
  XNOR2_X1 U3136 ( .A(n2443), .B(n2444), .ZN(n2930) );
  NAND2_X1 U3137 ( .A1(n2931), .A2(n2930), .ZN(n2447) );
  INV_X1 U3138 ( .A(n2443), .ZN(n2445) );
  NAND2_X1 U3139 ( .A1(n2445), .A2(n2444), .ZN(n2446) );
  NAND2_X1 U3140 ( .A1(n2692), .A2(REG1_REG_2__SCAN_IN), .ZN(n2453) );
  INV_X1 U3141 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2448) );
  OR2_X1 U3142 ( .A1(n2023), .A2(n2448), .ZN(n2452) );
  OR2_X1 U3143 ( .A1(n2746), .A2(n4192), .ZN(n2451) );
  INV_X1 U3144 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2449) );
  OAI22_X1 U3145 ( .A1(n2990), .A2(n2496), .B1(n2439), .B2(n3062), .ZN(n2455)
         );
  XNOR2_X1 U3146 ( .A(n2455), .B(n2793), .ZN(n2462) );
  INV_X1 U3147 ( .A(n2462), .ZN(n2460) );
  OR2_X1 U31480 ( .A1(n2990), .A2(n2498), .ZN(n2458) );
  NAND2_X1 U31490 ( .A1(n3055), .A2(n2456), .ZN(n2457) );
  AND2_X1 U3150 ( .A1(n2458), .A2(n2457), .ZN(n2461) );
  INV_X1 U3151 ( .A(n2461), .ZN(n2459) );
  NAND2_X1 U3152 ( .A1(n2462), .A2(n2461), .ZN(n2464) );
  XNOR2_X1 U3153 ( .A(n2466), .B(n2465), .ZN(n2945) );
  AND2_X1 U3154 ( .A1(n2945), .A2(n2467), .ZN(n2468) );
  NAND2_X1 U3155 ( .A1(n2946), .A2(n2468), .ZN(n2953) );
  NAND2_X1 U3156 ( .A1(n2469), .A2(n2953), .ZN(n2474) );
  INV_X1 U3157 ( .A(n2470), .ZN(n2471) );
  NAND2_X1 U3158 ( .A1(n2472), .A2(n2471), .ZN(n2473) );
  NAND2_X1 U3159 ( .A1(n3609), .A2(REG0_REG_6__SCAN_IN), .ZN(n2479) );
  OR2_X1 U3160 ( .A1(n2397), .A2(n4360), .ZN(n2478) );
  OAI21_X1 U3161 ( .B1(n2475), .B2(REG3_REG_6__SCAN_IN), .A(n2507), .ZN(n3125)
         );
  OR2_X1 U3162 ( .A1(n2024), .A2(n3125), .ZN(n2477) );
  OR2_X1 U3163 ( .A1(n2746), .A2(n4355), .ZN(n2476) );
  NAND4_X1 U3164 ( .A1(n2479), .A2(n2478), .A3(n2477), .A4(n2476), .ZN(n3707)
         );
  NAND2_X1 U3165 ( .A1(n3707), .A2(n2456), .ZN(n2482) );
  MUX2_X1 U3166 ( .A(n2480), .B(DATAI_6_), .S(n3349), .Z(n3105) );
  NAND2_X1 U3167 ( .A1(n3105), .A2(n2393), .ZN(n2481) );
  NAND2_X1 U3168 ( .A1(n2482), .A2(n2481), .ZN(n2483) );
  XNOR2_X1 U3169 ( .A(n2483), .B(n2778), .ZN(n2486) );
  NAND2_X1 U3170 ( .A1(n3707), .A2(n2781), .ZN(n2485) );
  NAND2_X1 U3171 ( .A1(n3105), .A2(n2456), .ZN(n2484) );
  NAND2_X1 U3172 ( .A1(n2485), .A2(n2484), .ZN(n2487) );
  AND2_X1 U3173 ( .A1(n2486), .A2(n2487), .ZN(n2975) );
  INV_X1 U3174 ( .A(n2486), .ZN(n2489) );
  INV_X1 U3175 ( .A(n2487), .ZN(n2488) );
  NAND2_X1 U3176 ( .A1(n2489), .A2(n2488), .ZN(n2976) );
  NAND2_X1 U3177 ( .A1(n3609), .A2(REG0_REG_7__SCAN_IN), .ZN(n2495) );
  INV_X1 U3178 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2490) );
  OR2_X1 U3179 ( .A1(n2397), .A2(n2490), .ZN(n2494) );
  INV_X1 U3180 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2491) );
  XNOR2_X1 U3181 ( .A(n2507), .B(n2491), .ZN(n3388) );
  OR2_X1 U3182 ( .A1(n2024), .A2(n3388), .ZN(n2493) );
  INV_X1 U3183 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3102) );
  OR2_X1 U3184 ( .A1(n2839), .A2(n3102), .ZN(n2492) );
  MUX2_X1 U3185 ( .A(n4368), .B(DATAI_7_), .S(n3349), .Z(n3387) );
  OAI22_X1 U3186 ( .A1(n3369), .A2(n2843), .B1(n2792), .B2(n3099), .ZN(n2497)
         );
  XNOR2_X1 U3187 ( .A(n2497), .B(n2778), .ZN(n2502) );
  OR2_X1 U3188 ( .A1(n3369), .A2(n2795), .ZN(n2500) );
  NAND2_X1 U3189 ( .A1(n3387), .A2(n2456), .ZN(n2499) );
  NAND2_X1 U3190 ( .A1(n2500), .A2(n2499), .ZN(n2501) );
  XNOR2_X1 U3191 ( .A(n2502), .B(n2501), .ZN(n3384) );
  NAND2_X1 U3192 ( .A1(n2502), .A2(n2501), .ZN(n2503) );
  NAND2_X1 U3193 ( .A1(n3609), .A2(REG0_REG_8__SCAN_IN), .ZN(n2512) );
  INV_X1 U3194 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2504) );
  OR2_X1 U3195 ( .A1(n2397), .A2(n2504), .ZN(n2511) );
  INV_X1 U3196 ( .A(n2507), .ZN(n2505) );
  AOI21_X1 U3197 ( .B1(n2505), .B2(REG3_REG_7__SCAN_IN), .A(
        REG3_REG_8__SCAN_IN), .ZN(n2508) );
  NAND2_X1 U3198 ( .A1(REG3_REG_7__SCAN_IN), .A2(REG3_REG_8__SCAN_IN), .ZN(
        n2506) );
  OR2_X1 U3199 ( .A1(n2508), .A2(n2522), .ZN(n3366) );
  OR2_X1 U3200 ( .A1(n2024), .A2(n3366), .ZN(n2510) );
  OR2_X1 U3201 ( .A1(n2839), .A2(n4376), .ZN(n2509) );
  NAND4_X1 U3202 ( .A1(n2512), .A2(n2511), .A3(n2510), .A4(n2509), .ZN(n3706)
         );
  NAND2_X1 U3203 ( .A1(n3706), .A2(n2781), .ZN(n2515) );
  MUX2_X1 U3204 ( .A(n2513), .B(DATAI_8_), .S(n3349), .Z(n3367) );
  NAND2_X1 U3205 ( .A1(n3367), .A2(n2456), .ZN(n2514) );
  NAND2_X1 U3206 ( .A1(n2515), .A2(n2514), .ZN(n3363) );
  NAND2_X1 U3207 ( .A1(n3706), .A2(n2456), .ZN(n2517) );
  NAND2_X1 U3208 ( .A1(n3367), .A2(n2393), .ZN(n2516) );
  NAND2_X1 U3209 ( .A1(n2517), .A2(n2516), .ZN(n2518) );
  XNOR2_X1 U32100 ( .A(n2518), .B(n2778), .ZN(n3362) );
  NAND2_X1 U32110 ( .A1(n3365), .A2(n3363), .ZN(n2519) );
  NAND2_X1 U32120 ( .A1(n2520), .A2(n2519), .ZN(n3462) );
  NAND2_X1 U32130 ( .A1(n3609), .A2(REG0_REG_9__SCAN_IN), .ZN(n2527) );
  OR2_X1 U32140 ( .A1(n2397), .A2(n2521), .ZN(n2526) );
  OR2_X1 U32150 ( .A1(n2522), .A2(REG3_REG_9__SCAN_IN), .ZN(n2523) );
  NAND2_X1 U32160 ( .A1(n2532), .A2(n2523), .ZN(n3468) );
  OR2_X1 U32170 ( .A1(n2024), .A2(n3468), .ZN(n2525) );
  OR2_X1 U32180 ( .A1(n2839), .A2(n3160), .ZN(n2524) );
  NAND4_X1 U32190 ( .A1(n2527), .A2(n2526), .A3(n2525), .A4(n2524), .ZN(n3705)
         );
  NAND2_X1 U32200 ( .A1(n3705), .A2(n2456), .ZN(n2530) );
  MUX2_X1 U32210 ( .A(n2528), .B(DATAI_9_), .S(n3349), .Z(n3467) );
  NAND2_X1 U32220 ( .A1(n3467), .A2(n2393), .ZN(n2529) );
  NAND2_X1 U32230 ( .A1(n2530), .A2(n2529), .ZN(n2531) );
  XNOR2_X1 U32240 ( .A(n2531), .B(n2793), .ZN(n2544) );
  AOI22_X1 U32250 ( .A1(n3705), .A2(n2781), .B1(n2456), .B2(n3467), .ZN(n2543)
         );
  XNOR2_X1 U32260 ( .A(n2544), .B(n2543), .ZN(n3464) );
  NAND2_X1 U32270 ( .A1(n3609), .A2(REG0_REG_10__SCAN_IN), .ZN(n2538) );
  NAND2_X1 U32280 ( .A1(n2532), .A2(n3089), .ZN(n2533) );
  AND2_X1 U32290 ( .A1(n2550), .A2(n2533), .ZN(n4472) );
  INV_X1 U32300 ( .A(n4472), .ZN(n3093) );
  OR2_X1 U32310 ( .A1(n2024), .A2(n3093), .ZN(n2537) );
  INV_X1 U32320 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2534) );
  OR2_X1 U32330 ( .A1(n2397), .A2(n2534), .ZN(n2536) );
  OR2_X1 U32340 ( .A1(n2839), .A2(n4386), .ZN(n2535) );
  NAND4_X1 U32350 ( .A1(n2538), .A2(n2537), .A3(n2536), .A4(n2535), .ZN(n4459)
         );
  NAND2_X1 U32360 ( .A1(n4459), .A2(n2456), .ZN(n2541) );
  MUX2_X1 U32370 ( .A(n2539), .B(DATAI_10_), .S(n3349), .Z(n3205) );
  NAND2_X1 U32380 ( .A1(n3205), .A2(n2393), .ZN(n2540) );
  NAND2_X1 U32390 ( .A1(n2541), .A2(n2540), .ZN(n2542) );
  XNOR2_X1 U32400 ( .A(n2542), .B(n2778), .ZN(n2548) );
  AOI22_X1 U32410 ( .A1(n4459), .A2(n2781), .B1(n2456), .B2(n3205), .ZN(n2546)
         );
  XNOR2_X1 U32420 ( .A(n2548), .B(n2546), .ZN(n3087) );
  NAND2_X1 U32430 ( .A1(n2544), .A2(n2543), .ZN(n3085) );
  AND2_X1 U32440 ( .A1(n3087), .A2(n3085), .ZN(n2545) );
  INV_X1 U32450 ( .A(n2546), .ZN(n2547) );
  NAND2_X1 U32460 ( .A1(n3609), .A2(REG0_REG_11__SCAN_IN), .ZN(n2556) );
  OR2_X1 U32470 ( .A1(n2397), .A2(n4619), .ZN(n2555) );
  NAND2_X1 U32480 ( .A1(n2550), .A2(n2549), .ZN(n2551) );
  AND2_X1 U32490 ( .A1(n2566), .A2(n2551), .ZN(n4465) );
  INV_X1 U32500 ( .A(n4465), .ZN(n2552) );
  OR2_X1 U32510 ( .A1(n2024), .A2(n2552), .ZN(n2554) );
  OR2_X1 U32520 ( .A1(n2839), .A2(n4252), .ZN(n2553) );
  MUX2_X1 U32530 ( .A(n2557), .B(DATAI_11_), .S(n3349), .Z(n3212) );
  OAI22_X1 U32540 ( .A1(n3228), .A2(n2843), .B1(n2792), .B2(n4467), .ZN(n2558)
         );
  XNOR2_X1 U32550 ( .A(n2558), .B(n2793), .ZN(n2561) );
  OR2_X1 U32560 ( .A1(n3228), .A2(n2795), .ZN(n2560) );
  NAND2_X1 U32570 ( .A1(n3212), .A2(n2456), .ZN(n2559) );
  NAND2_X1 U32580 ( .A1(n2561), .A2(n2562), .ZN(n3217) );
  NAND2_X1 U32590 ( .A1(n3216), .A2(n3217), .ZN(n3215) );
  INV_X1 U32600 ( .A(n2561), .ZN(n2564) );
  INV_X1 U32610 ( .A(n2562), .ZN(n2563) );
  NAND2_X1 U32620 ( .A1(n2564), .A2(n2563), .ZN(n3219) );
  NAND2_X1 U32630 ( .A1(n3609), .A2(REG0_REG_12__SCAN_IN), .ZN(n2571) );
  INV_X1 U32640 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4271) );
  OR2_X1 U32650 ( .A1(n2397), .A2(n4271), .ZN(n2570) );
  INV_X1 U32660 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4202) );
  NAND2_X1 U32670 ( .A1(n2566), .A2(n4202), .ZN(n2567) );
  NAND2_X1 U32680 ( .A1(n2597), .A2(n2567), .ZN(n3208) );
  OR2_X1 U32690 ( .A1(n2024), .A2(n3208), .ZN(n2569) );
  OR2_X1 U32700 ( .A1(n2839), .A2(n4405), .ZN(n2568) );
  NAND2_X1 U32710 ( .A1(n3703), .A2(n2456), .ZN(n2574) );
  MUX2_X1 U32720 ( .A(n2572), .B(DATAI_12_), .S(n3349), .Z(n3257) );
  NAND2_X1 U32730 ( .A1(n3257), .A2(n2393), .ZN(n2573) );
  NAND2_X1 U32740 ( .A1(n2574), .A2(n2573), .ZN(n2575) );
  XNOR2_X1 U32750 ( .A(n2575), .B(n2778), .ZN(n3180) );
  NAND2_X1 U32760 ( .A1(n3703), .A2(n2781), .ZN(n2577) );
  NAND2_X1 U32770 ( .A1(n3257), .A2(n2456), .ZN(n2576) );
  NAND2_X1 U32780 ( .A1(n2577), .A2(n2576), .ZN(n3179) );
  OAI21_X1 U32790 ( .B1(n3182), .B2(n3180), .A(n3179), .ZN(n2579) );
  NAND2_X1 U32800 ( .A1(n3182), .A2(n3180), .ZN(n2578) );
  NAND2_X1 U32810 ( .A1(n2579), .A2(n2578), .ZN(n3238) );
  NAND2_X1 U32820 ( .A1(n3609), .A2(REG0_REG_13__SCAN_IN), .ZN(n2584) );
  OR2_X1 U32830 ( .A1(n2397), .A2(n2580), .ZN(n2583) );
  XNOR2_X1 U32840 ( .A(n2597), .B(n2595), .ZN(n3267) );
  OR2_X1 U32850 ( .A1(n2024), .A2(n3267), .ZN(n2582) );
  OR2_X1 U32860 ( .A1(n2839), .A2(n3268), .ZN(n2581) );
  NAND4_X1 U32870 ( .A1(n2584), .A2(n2583), .A3(n2582), .A4(n2581), .ZN(n3702)
         );
  NAND2_X1 U32880 ( .A1(n3702), .A2(n2456), .ZN(n2586) );
  MUX2_X1 U32890 ( .A(n4337), .B(DATAI_13_), .S(n3349), .Z(n3281) );
  NAND2_X1 U32900 ( .A1(n3281), .A2(n2393), .ZN(n2585) );
  NAND2_X1 U32910 ( .A1(n2586), .A2(n2585), .ZN(n2587) );
  XNOR2_X1 U32920 ( .A(n2587), .B(n2778), .ZN(n2590) );
  NAND2_X1 U32930 ( .A1(n3702), .A2(n2781), .ZN(n2589) );
  NAND2_X1 U32940 ( .A1(n3281), .A2(n2456), .ZN(n2588) );
  NAND2_X1 U32950 ( .A1(n2589), .A2(n2588), .ZN(n2591) );
  INV_X1 U32960 ( .A(n2590), .ZN(n2593) );
  INV_X1 U32970 ( .A(n2591), .ZN(n2592) );
  NAND2_X1 U32980 ( .A1(n2593), .A2(n2592), .ZN(n3240) );
  NAND2_X1 U32990 ( .A1(n3609), .A2(REG0_REG_14__SCAN_IN), .ZN(n2602) );
  INV_X1 U33000 ( .A(REG1_REG_14__SCAN_IN), .ZN(n2594) );
  OR2_X1 U33010 ( .A1(n2397), .A2(n2594), .ZN(n2601) );
  OAI21_X1 U33020 ( .B1(n2597), .B2(n2595), .A(n2596), .ZN(n2598) );
  NAND2_X1 U33030 ( .A1(n2598), .A2(n2608), .ZN(n3297) );
  OR2_X1 U33040 ( .A1(n2024), .A2(n3297), .ZN(n2600) );
  INV_X1 U33050 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3298) );
  OR2_X1 U33060 ( .A1(n2839), .A2(n3298), .ZN(n2599) );
  MUX2_X1 U33070 ( .A(n2603), .B(DATAI_14_), .S(n3349), .Z(n3295) );
  OAI22_X1 U33080 ( .A1(n3532), .A2(n2843), .B1(n2792), .B2(n3302), .ZN(n2604)
         );
  OR2_X1 U33090 ( .A1(n3532), .A2(n2795), .ZN(n2606) );
  NAND2_X1 U33100 ( .A1(n3295), .A2(n2456), .ZN(n2605) );
  NAND2_X1 U33110 ( .A1(n2606), .A2(n2605), .ZN(n3274) );
  INV_X1 U33120 ( .A(n3273), .ZN(n2607) );
  NAND2_X1 U33130 ( .A1(n3609), .A2(REG0_REG_15__SCAN_IN), .ZN(n2613) );
  OR2_X1 U33140 ( .A1(n2397), .A2(n4131), .ZN(n2612) );
  INV_X1 U33150 ( .A(n2635), .ZN(n2633) );
  NAND2_X1 U33160 ( .A1(n2608), .A2(n3529), .ZN(n2609) );
  NAND2_X1 U33170 ( .A1(n2633), .A2(n2609), .ZN(n3537) );
  OR2_X1 U33180 ( .A1(n2024), .A2(n3537), .ZN(n2611) );
  OR2_X1 U33190 ( .A1(n2839), .A2(n2261), .ZN(n2610) );
  NAND4_X1 U33200 ( .A1(n2613), .A2(n2612), .A3(n2611), .A4(n2610), .ZN(n3325)
         );
  NAND2_X1 U33210 ( .A1(n3325), .A2(n2456), .ZN(n2616) );
  MUX2_X1 U33220 ( .A(n2614), .B(DATAI_15_), .S(n3349), .Z(n3315) );
  NAND2_X1 U33230 ( .A1(n3315), .A2(n2393), .ZN(n2615) );
  NAND2_X1 U33240 ( .A1(n2616), .A2(n2615), .ZN(n2617) );
  XNOR2_X1 U33250 ( .A(n2617), .B(n2778), .ZN(n2625) );
  NOR2_X1 U33260 ( .A1(n2626), .A2(n2625), .ZN(n3432) );
  AND2_X1 U33270 ( .A1(n3315), .A2(n2456), .ZN(n2618) );
  AOI21_X1 U33280 ( .B1(n3325), .B2(n2781), .A(n2618), .ZN(n3521) );
  NAND2_X1 U33290 ( .A1(n3609), .A2(REG0_REG_16__SCAN_IN), .ZN(n2623) );
  INV_X1 U33300 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2632) );
  XNOR2_X1 U33310 ( .A(n2633), .B(n2632), .ZN(n3330) );
  OR2_X1 U33320 ( .A1(n2024), .A2(n3330), .ZN(n2622) );
  INV_X1 U33330 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4127) );
  OR2_X1 U33340 ( .A1(n2397), .A2(n4127), .ZN(n2621) );
  INV_X1 U33350 ( .A(REG2_REG_16__SCAN_IN), .ZN(n2619) );
  OR2_X1 U33360 ( .A1(n2839), .A2(n2619), .ZN(n2620) );
  MUX2_X1 U33370 ( .A(n4541), .B(DATAI_16_), .S(n3349), .Z(n3797) );
  OAI22_X1 U33380 ( .A1(n3528), .A2(n2795), .B1(n2843), .B2(n3329), .ZN(n2627)
         );
  OAI22_X1 U33390 ( .A1(n3528), .A2(n2843), .B1(n2792), .B2(n3329), .ZN(n2624)
         );
  XNOR2_X1 U33400 ( .A(n2624), .B(n2778), .ZN(n2628) );
  XOR2_X1 U33410 ( .A(n2627), .B(n2628), .Z(n3433) );
  OAI211_X1 U33420 ( .C1(n3432), .C2(n3521), .A(n3433), .B(n3519), .ZN(n2630)
         );
  NAND2_X1 U33430 ( .A1(n2630), .A2(n2629), .ZN(n3441) );
  NAND2_X1 U33440 ( .A1(n3609), .A2(REG0_REG_17__SCAN_IN), .ZN(n2640) );
  OR2_X1 U33450 ( .A1(n2397), .A2(n4123), .ZN(n2639) );
  INV_X1 U33460 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2631) );
  OAI21_X1 U33470 ( .B1(n2633), .B2(n2632), .A(n2631), .ZN(n2636) );
  AND2_X1 U33480 ( .A1(REG3_REG_16__SCAN_IN), .A2(REG3_REG_17__SCAN_IN), .ZN(
        n2634) );
  INV_X1 U33490 ( .A(n2647), .ZN(n2648) );
  NAND2_X1 U33500 ( .A1(n2636), .A2(n2648), .ZN(n4058) );
  OR2_X1 U33510 ( .A1(n2024), .A2(n4058), .ZN(n2638) );
  OR2_X1 U33520 ( .A1(n2839), .A2(n2352), .ZN(n2637) );
  MUX2_X1 U3353 ( .A(n2641), .B(DATAI_17_), .S(n3349), .Z(n3801) );
  INV_X1 U33540 ( .A(n3801), .ZN(n4055) );
  OAI22_X1 U3355 ( .A1(n4036), .A2(n2843), .B1(n2792), .B2(n4055), .ZN(n2642)
         );
  XNOR2_X1 U3356 ( .A(n2642), .B(n2793), .ZN(n3443) );
  OR2_X1 U3357 ( .A1(n4036), .A2(n2795), .ZN(n2644) );
  NAND2_X1 U3358 ( .A1(n3801), .A2(n2456), .ZN(n2643) );
  INV_X1 U3359 ( .A(n3443), .ZN(n2646) );
  INV_X1 U3360 ( .A(n2645), .ZN(n3442) );
  NAND2_X1 U3361 ( .A1(n3609), .A2(REG0_REG_18__SCAN_IN), .ZN(n2653) );
  OR2_X1 U3362 ( .A1(n2397), .A2(n3762), .ZN(n2652) );
  NAND2_X1 U3363 ( .A1(n2648), .A2(n4261), .ZN(n2649) );
  NAND2_X1 U3364 ( .A1(n2663), .A2(n2649), .ZN(n4030) );
  OR2_X1 U3365 ( .A1(n2024), .A2(n4030), .ZN(n2651) );
  OR2_X1 U3366 ( .A1(n2839), .A2(n4263), .ZN(n2650) );
  MUX2_X1 U3367 ( .A(n2654), .B(DATAI_18_), .S(n3349), .Z(n4033) );
  OAI22_X1 U3368 ( .A1(n4047), .A2(n2843), .B1(n2792), .B2(n4029), .ZN(n2655)
         );
  XNOR2_X1 U3369 ( .A(n2655), .B(n2793), .ZN(n2661) );
  INV_X1 U3370 ( .A(n2661), .ZN(n2659) );
  OR2_X1 U3371 ( .A1(n4047), .A2(n2795), .ZN(n2657) );
  NAND2_X1 U3372 ( .A1(n4033), .A2(n2456), .ZN(n2656) );
  AND2_X1 U3373 ( .A1(n2657), .A2(n2656), .ZN(n2660) );
  INV_X1 U3374 ( .A(n2660), .ZN(n2658) );
  NAND2_X1 U3375 ( .A1(n2659), .A2(n2658), .ZN(n3493) );
  INV_X1 U3376 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4316) );
  OR2_X1 U3377 ( .A1(n2437), .A2(n4316), .ZN(n2668) );
  INV_X1 U3378 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4210) );
  OR2_X1 U3379 ( .A1(n2397), .A2(n4210), .ZN(n2667) );
  INV_X1 U3380 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2662) );
  NAND2_X1 U3381 ( .A1(n2663), .A2(n2662), .ZN(n2664) );
  NAND2_X1 U3382 ( .A1(n2676), .A2(n2664), .ZN(n4020) );
  OR2_X1 U3383 ( .A1(n2024), .A2(n4020), .ZN(n2666) );
  INV_X1 U3384 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4021) );
  OR2_X1 U3385 ( .A1(n2839), .A2(n4021), .ZN(n2665) );
  NAND4_X1 U3386 ( .A1(n2668), .A2(n2667), .A3(n2666), .A4(n2665), .ZN(n4034)
         );
  NAND2_X1 U3387 ( .A1(n4034), .A2(n2456), .ZN(n2671) );
  INV_X1 U3388 ( .A(DATAI_19_), .ZN(n2669) );
  MUX2_X1 U3389 ( .A(n3768), .B(n2669), .S(n3349), .Z(n4019) );
  NAND2_X1 U3390 ( .A1(n4014), .A2(n2393), .ZN(n2670) );
  NAND2_X1 U3391 ( .A1(n2671), .A2(n2670), .ZN(n2672) );
  XNOR2_X1 U3392 ( .A(n2672), .B(n2778), .ZN(n2674) );
  INV_X1 U3393 ( .A(n4034), .ZN(n3804) );
  OAI22_X1 U3394 ( .A1(n3804), .A2(n2795), .B1(n2843), .B2(n4019), .ZN(n2673)
         );
  XNOR2_X1 U3395 ( .A(n2674), .B(n2673), .ZN(n3405) );
  NAND2_X1 U3396 ( .A1(n3609), .A2(REG0_REG_20__SCAN_IN), .ZN(n2681) );
  INV_X1 U3397 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4113) );
  OR2_X1 U3398 ( .A1(n2397), .A2(n4113), .ZN(n2680) );
  INV_X1 U3399 ( .A(REG3_REG_20__SCAN_IN), .ZN(n2675) );
  INV_X1 U3400 ( .A(n2693), .ZN(n2695) );
  NAND2_X1 U3401 ( .A1(n2676), .A2(n2675), .ZN(n2677) );
  NAND2_X1 U3402 ( .A1(n2695), .A2(n2677), .ZN(n3997) );
  OR2_X1 U3403 ( .A1(n2024), .A2(n3997), .ZN(n2679) );
  INV_X1 U3404 ( .A(REG2_REG_20__SCAN_IN), .ZN(n3998) );
  OR2_X1 U3405 ( .A1(n2839), .A2(n3998), .ZN(n2678) );
  NAND2_X1 U3406 ( .A1(n4015), .A2(n2456), .ZN(n2684) );
  NAND2_X1 U3407 ( .A1(n3349), .A2(DATAI_20_), .ZN(n3995) );
  NAND2_X1 U3408 ( .A1(n3632), .A2(n2393), .ZN(n2683) );
  NAND2_X1 U3409 ( .A1(n2684), .A2(n2683), .ZN(n2685) );
  XNOR2_X1 U3410 ( .A(n2685), .B(n2778), .ZN(n2688) );
  NAND2_X1 U3411 ( .A1(n4015), .A2(n2781), .ZN(n2687) );
  NAND2_X1 U3412 ( .A1(n3632), .A2(n2456), .ZN(n2686) );
  NAND2_X1 U3413 ( .A1(n2687), .A2(n2686), .ZN(n2689) );
  NAND2_X1 U3414 ( .A1(n2688), .A2(n2689), .ZN(n3476) );
  NAND2_X1 U3415 ( .A1(n3475), .A2(n3476), .ZN(n3474) );
  INV_X1 U3416 ( .A(n2688), .ZN(n2691) );
  INV_X1 U3417 ( .A(n2689), .ZN(n2690) );
  NAND2_X1 U3418 ( .A1(n2691), .A2(n2690), .ZN(n3477) );
  NAND2_X1 U3419 ( .A1(n2692), .A2(REG1_REG_21__SCAN_IN), .ZN(n2700) );
  INV_X1 U3420 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4308) );
  OR2_X1 U3421 ( .A1(n2437), .A2(n4308), .ZN(n2699) );
  INV_X1 U3422 ( .A(n2707), .ZN(n2708) );
  INV_X1 U3423 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2694) );
  NAND2_X1 U3424 ( .A1(n2695), .A2(n2694), .ZN(n2696) );
  NAND2_X1 U3425 ( .A1(n2708), .A2(n2696), .ZN(n3978) );
  OR2_X1 U3426 ( .A1(n2024), .A2(n3978), .ZN(n2698) );
  INV_X1 U3427 ( .A(REG2_REG_21__SCAN_IN), .ZN(n3979) );
  OR2_X1 U3428 ( .A1(n2839), .A2(n3979), .ZN(n2697) );
  AND2_X1 U3429 ( .A1(n3349), .A2(DATAI_21_), .ZN(n3598) );
  INV_X1 U3430 ( .A(n3598), .ZN(n3977) );
  OAI22_X1 U3431 ( .A1(n3990), .A2(n2843), .B1(n2792), .B2(n3977), .ZN(n2701)
         );
  XNOR2_X1 U3432 ( .A(n2701), .B(n2778), .ZN(n3412) );
  OR2_X1 U3433 ( .A1(n3990), .A2(n2795), .ZN(n2703) );
  NAND2_X1 U3434 ( .A1(n3598), .A2(n2456), .ZN(n2702) );
  NAND2_X1 U3435 ( .A1(n2703), .A2(n2702), .ZN(n2704) );
  NOR2_X1 U3436 ( .A1(n3412), .A2(n2704), .ZN(n2705) );
  INV_X1 U3437 ( .A(n2704), .ZN(n3411) );
  NAND2_X1 U3438 ( .A1(n3609), .A2(REG0_REG_22__SCAN_IN), .ZN(n2713) );
  INV_X1 U3439 ( .A(REG1_REG_22__SCAN_IN), .ZN(n2706) );
  OR2_X1 U3440 ( .A1(n2397), .A2(n2706), .ZN(n2712) );
  INV_X1 U3441 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3487) );
  NAND2_X1 U3442 ( .A1(n2708), .A2(n3487), .ZN(n2709) );
  NAND2_X1 U3443 ( .A1(n2717), .A2(n2709), .ZN(n3964) );
  OR2_X1 U3444 ( .A1(n2024), .A2(n3964), .ZN(n2711) );
  INV_X1 U3445 ( .A(REG2_REG_22__SCAN_IN), .ZN(n3965) );
  OR2_X1 U3446 ( .A1(n2839), .A2(n3965), .ZN(n2710) );
  AND2_X1 U3447 ( .A1(n3349), .A2(DATAI_22_), .ZN(n3963) );
  INV_X1 U3448 ( .A(n3963), .ZN(n3601) );
  OAI22_X1 U3449 ( .A1(n3972), .A2(n2843), .B1(n2792), .B2(n3601), .ZN(n2714)
         );
  XNOR2_X1 U3450 ( .A(n2714), .B(n2778), .ZN(n2716) );
  OAI22_X1 U3451 ( .A1(n3972), .A2(n2795), .B1(n2843), .B2(n3601), .ZN(n2715)
         );
  XNOR2_X1 U3452 ( .A(n2716), .B(n2715), .ZN(n3486) );
  NOR2_X1 U3453 ( .A1(n2716), .A2(n2715), .ZN(n3396) );
  NAND2_X1 U3454 ( .A1(n2692), .A2(REG1_REG_23__SCAN_IN), .ZN(n2722) );
  INV_X1 U3455 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4303) );
  OR2_X1 U3456 ( .A1(n2437), .A2(n4303), .ZN(n2721) );
  INV_X1 U3457 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3399) );
  NAND2_X1 U34580 ( .A1(n2717), .A2(n3399), .ZN(n2718) );
  NAND2_X1 U34590 ( .A1(n2729), .A2(n2718), .ZN(n3944) );
  OR2_X1 U3460 ( .A1(n2024), .A2(n3944), .ZN(n2720) );
  INV_X1 U3461 ( .A(REG2_REG_23__SCAN_IN), .ZN(n3945) );
  OR2_X1 U3462 ( .A1(n2839), .A2(n3945), .ZN(n2719) );
  NAND4_X1 U3463 ( .A1(n2722), .A2(n2721), .A3(n2720), .A4(n2719), .ZN(n3953)
         );
  NAND2_X1 U3464 ( .A1(n3953), .A2(n2456), .ZN(n2724) );
  AND2_X1 U3465 ( .A1(n3349), .A2(DATAI_23_), .ZN(n3808) );
  NAND2_X1 U3466 ( .A1(n3808), .A2(n2393), .ZN(n2723) );
  NAND2_X1 U34670 ( .A1(n2724), .A2(n2723), .ZN(n2725) );
  XNOR2_X1 U3468 ( .A(n2725), .B(n2793), .ZN(n2728) );
  AND2_X1 U34690 ( .A1(n3808), .A2(n2456), .ZN(n2726) );
  AOI21_X1 U3470 ( .B1(n3953), .B2(n2781), .A(n2726), .ZN(n2727) );
  XNOR2_X1 U34710 ( .A(n2728), .B(n2727), .ZN(n3395) );
  NOR2_X1 U3472 ( .A1(n2728), .A2(n2727), .ZN(n2738) );
  NAND2_X1 U34730 ( .A1(n3609), .A2(REG0_REG_24__SCAN_IN), .ZN(n2734) );
  INV_X1 U3474 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4187) );
  NAND2_X1 U34750 ( .A1(n2729), .A2(n4187), .ZN(n2730) );
  NAND2_X1 U3476 ( .A1(n2744), .A2(n2730), .ZN(n3919) );
  OR2_X1 U34770 ( .A1(n3919), .A2(n2024), .ZN(n2733) );
  INV_X1 U3478 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4096) );
  OR2_X1 U34790 ( .A1(n2397), .A2(n4096), .ZN(n2732) );
  INV_X1 U3480 ( .A(REG2_REG_24__SCAN_IN), .ZN(n3920) );
  OR2_X1 U34810 ( .A1(n2839), .A2(n3920), .ZN(n2731) );
  AND2_X1 U3482 ( .A1(n3349), .A2(DATAI_24_), .ZN(n3813) );
  OAI22_X1 U34830 ( .A1(n3814), .A2(n2795), .B1(n2843), .B2(n3917), .ZN(n2737)
         );
  OAI21_X1 U3484 ( .B1(n3394), .B2(n2738), .A(n2737), .ZN(n3453) );
  OAI22_X1 U34850 ( .A1(n3814), .A2(n2843), .B1(n2792), .B2(n3917), .ZN(n2741)
         );
  XNOR2_X1 U3486 ( .A(n2741), .B(n2778), .ZN(n3454) );
  NAND2_X1 U34870 ( .A1(n3452), .A2(n3454), .ZN(n2742) );
  NAND2_X1 U3488 ( .A1(n3453), .A2(n2742), .ZN(n3421) );
  INV_X1 U34890 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3427) );
  NAND2_X1 U3490 ( .A1(n2744), .A2(n3427), .ZN(n2745) );
  NAND2_X1 U34910 ( .A1(n2758), .A2(n2745), .ZN(n3426) );
  NAND2_X1 U3492 ( .A1(n2692), .A2(REG1_REG_25__SCAN_IN), .ZN(n2749) );
  NAND2_X1 U34930 ( .A1(n2786), .A2(REG2_REG_25__SCAN_IN), .ZN(n2748) );
  INV_X1 U3494 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4295) );
  OR2_X1 U34950 ( .A1(n2437), .A2(n4295), .ZN(n2747) );
  NAND2_X1 U3496 ( .A1(n3913), .A2(n2456), .ZN(n2752) );
  AND2_X1 U34970 ( .A1(n3349), .A2(DATAI_25_), .ZN(n3899) );
  NAND2_X1 U3498 ( .A1(n3899), .A2(n2393), .ZN(n2751) );
  NAND2_X1 U34990 ( .A1(n2752), .A2(n2751), .ZN(n2753) );
  XNOR2_X1 U3500 ( .A(n2753), .B(n2793), .ZN(n2756) );
  AND2_X1 U35010 ( .A1(n3899), .A2(n2456), .ZN(n2754) );
  AOI21_X1 U3502 ( .B1(n3913), .B2(n2781), .A(n2754), .ZN(n2755) );
  NAND2_X1 U35030 ( .A1(n2756), .A2(n2755), .ZN(n3422) );
  NOR2_X1 U3504 ( .A1(n2756), .A2(n2755), .ZN(n3424) );
  INV_X1 U35050 ( .A(REG2_REG_26__SCAN_IN), .ZN(n3883) );
  INV_X1 U35060 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3511) );
  NAND2_X1 U35070 ( .A1(n2758), .A2(n3511), .ZN(n2759) );
  NAND2_X1 U35080 ( .A1(n2772), .A2(n2759), .ZN(n3882) );
  NAND2_X1 U35090 ( .A1(n3609), .A2(REG0_REG_26__SCAN_IN), .ZN(n2761) );
  NAND2_X1 U35100 ( .A1(n2692), .A2(REG1_REG_26__SCAN_IN), .ZN(n2760) );
  AND2_X1 U35110 ( .A1(n2761), .A2(n2760), .ZN(n2762) );
  NAND2_X1 U35120 ( .A1(n3852), .A2(n2456), .ZN(n2765) );
  AND2_X1 U35130 ( .A1(n3349), .A2(DATAI_26_), .ZN(n3871) );
  NAND2_X1 U35140 ( .A1(n3871), .A2(n2393), .ZN(n2764) );
  NAND2_X1 U35150 ( .A1(n2765), .A2(n2764), .ZN(n2766) );
  XNOR2_X1 U35160 ( .A(n2766), .B(n2793), .ZN(n2771) );
  INV_X1 U35170 ( .A(n2771), .ZN(n2769) );
  AND2_X1 U35180 ( .A1(n3871), .A2(n2456), .ZN(n2767) );
  AOI21_X1 U35190 ( .B1(n3852), .B2(n2781), .A(n2767), .ZN(n2770) );
  INV_X1 U35200 ( .A(n2770), .ZN(n2768) );
  NAND2_X1 U35210 ( .A1(n2769), .A2(n2768), .ZN(n3507) );
  AND2_X1 U35220 ( .A1(n2771), .A2(n2770), .ZN(n3506) );
  INV_X1 U35230 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3377) );
  NAND2_X1 U35240 ( .A1(n2772), .A2(n3377), .ZN(n2773) );
  NAND2_X1 U35250 ( .A1(n2784), .A2(n2773), .ZN(n3862) );
  AOI22_X1 U35260 ( .A1(n3609), .A2(REG0_REG_27__SCAN_IN), .B1(n2692), .B2(
        REG1_REG_27__SCAN_IN), .ZN(n2775) );
  NAND2_X1 U35270 ( .A1(n2786), .A2(REG2_REG_27__SCAN_IN), .ZN(n2774) );
  NAND2_X1 U35280 ( .A1(n3831), .A2(n2456), .ZN(n2777) );
  AND2_X1 U35290 ( .A1(n3349), .A2(DATAI_27_), .ZN(n3851) );
  NAND2_X1 U35300 ( .A1(n3851), .A2(n2393), .ZN(n2776) );
  NAND2_X1 U35310 ( .A1(n2777), .A2(n2776), .ZN(n2779) );
  XNOR2_X1 U35320 ( .A(n2779), .B(n2778), .ZN(n2824) );
  AND2_X1 U35330 ( .A1(n3851), .A2(n2456), .ZN(n2780) );
  AOI21_X1 U35340 ( .B1(n3831), .B2(n2781), .A(n2780), .ZN(n2822) );
  XNOR2_X1 U35350 ( .A(n2824), .B(n2822), .ZN(n3375) );
  NAND2_X1 U35360 ( .A1(n3376), .A2(n3375), .ZN(n2857) );
  INV_X1 U35370 ( .A(n2784), .ZN(n2782) );
  NAND2_X1 U35380 ( .A1(n2782), .A2(REG3_REG_28__SCAN_IN), .ZN(n3773) );
  INV_X1 U35390 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2783) );
  NAND2_X1 U35400 ( .A1(n2784), .A2(n2783), .ZN(n2785) );
  NAND2_X1 U35410 ( .A1(n3773), .A2(n2785), .ZN(n3843) );
  INV_X1 U35420 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4254) );
  NAND2_X1 U35430 ( .A1(n3609), .A2(REG0_REG_28__SCAN_IN), .ZN(n2788) );
  NAND2_X1 U35440 ( .A1(n2786), .A2(REG2_REG_28__SCAN_IN), .ZN(n2787) );
  OAI211_X1 U35450 ( .C1(n2397), .C2(n4254), .A(n2788), .B(n2787), .ZN(n2789)
         );
  INV_X1 U35460 ( .A(n2789), .ZN(n2790) );
  AND2_X1 U35470 ( .A1(n3349), .A2(DATAI_28_), .ZN(n3841) );
  INV_X1 U35480 ( .A(n3841), .ZN(n3604) );
  OAI22_X1 U35490 ( .A1(n3854), .A2(n2843), .B1(n2792), .B2(n3604), .ZN(n2794)
         );
  XNOR2_X1 U35500 ( .A(n2794), .B(n2793), .ZN(n2797) );
  OAI22_X1 U35510 ( .A1(n3854), .A2(n2795), .B1(n2843), .B2(n3604), .ZN(n2796)
         );
  XNOR2_X1 U35520 ( .A(n2797), .B(n2796), .ZN(n2827) );
  INV_X1 U35530 ( .A(n2827), .ZN(n2821) );
  NAND2_X1 U35540 ( .A1(n2799), .A2(n2884), .ZN(n2800) );
  MUX2_X1 U35550 ( .A(n2799), .B(n2800), .S(B_REG_SCAN_IN), .Z(n2801) );
  INV_X1 U35560 ( .A(n2798), .ZN(n2814) );
  NAND2_X1 U35570 ( .A1(n2814), .A2(n2799), .ZN(n2802) );
  NOR4_X1 U35580 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_29__SCAN_IN), .ZN(n2812) );
  NOR4_X1 U35590 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2811) );
  INV_X1 U35600 ( .A(D_REG_20__SCAN_IN), .ZN(n4525) );
  INV_X1 U35610 ( .A(D_REG_4__SCAN_IN), .ZN(n4531) );
  INV_X1 U35620 ( .A(D_REG_13__SCAN_IN), .ZN(n4528) );
  INV_X1 U35630 ( .A(D_REG_22__SCAN_IN), .ZN(n4524) );
  NAND4_X1 U35640 ( .A1(n4525), .A2(n4531), .A3(n4528), .A4(n4524), .ZN(n2809)
         );
  NOR4_X1 U35650 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2807) );
  NOR4_X1 U35660 ( .A1(D_REG_8__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_7__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2806) );
  NOR4_X1 U35670 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2805) );
  NOR4_X1 U35680 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2804) );
  NAND4_X1 U35690 ( .A1(n2807), .A2(n2806), .A3(n2805), .A4(n2804), .ZN(n2808)
         );
  NOR4_X1 U35700 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(n2809), 
        .A4(n2808), .ZN(n2810) );
  AND3_X1 U35710 ( .A1(n2812), .A2(n2811), .A3(n2810), .ZN(n2813) );
  NOR2_X1 U35720 ( .A1(n2881), .A2(n2813), .ZN(n3027) );
  OR2_X1 U35730 ( .A1(n2881), .A2(D_REG_1__SCAN_IN), .ZN(n2816) );
  NAND2_X1 U35740 ( .A1(n2814), .A2(n2884), .ZN(n2815) );
  NAND2_X1 U35750 ( .A1(n2816), .A2(n2815), .ZN(n3014) );
  NOR2_X1 U35760 ( .A1(n3027), .A2(n3014), .ZN(n2817) );
  INV_X1 U35770 ( .A(n3008), .ZN(n3007) );
  NAND2_X1 U35780 ( .A1(n2845), .A2(n3768), .ZN(n2831) );
  NAND2_X1 U35790 ( .A1(n4508), .A2(n2831), .ZN(n2818) );
  NAND2_X1 U35800 ( .A1(n3007), .A2(n2818), .ZN(n2819) );
  NOR2_X1 U35810 ( .A1(n2889), .A2(n2819), .ZN(n2820) );
  NAND2_X1 U3582 ( .A1(n2821), .A2(n3523), .ZN(n2856) );
  INV_X1 U3583 ( .A(n2822), .ZN(n2823) );
  NAND2_X1 U3584 ( .A1(n2824), .A2(n2823), .ZN(n2826) );
  NAND2_X1 U3585 ( .A1(n2857), .A2(n2825), .ZN(n2855) );
  NOR3_X1 U3586 ( .A1(n2827), .A2(n3517), .A3(n2826), .ZN(n2853) );
  INV_X1 U3587 ( .A(n2849), .ZN(n2830) );
  AND2_X1 U3588 ( .A1(n2845), .A2(n3763), .ZN(n4510) );
  NAND2_X1 U3589 ( .A1(n4603), .A2(n2829), .ZN(n3012) );
  NAND2_X1 U3590 ( .A1(n2830), .A2(n3012), .ZN(n2890) );
  AND2_X1 U3591 ( .A1(n3008), .A2(n2831), .ZN(n2888) );
  NOR2_X1 U3592 ( .A1(n2888), .A2(n2832), .ZN(n2833) );
  AND2_X1 U3593 ( .A1(n2384), .A2(n2833), .ZN(n2834) );
  NAND2_X1 U3594 ( .A1(n2890), .A2(n2834), .ZN(n2835) );
  INV_X1 U3595 ( .A(REG2_REG_29__SCAN_IN), .ZN(n2838) );
  OR2_X1 U3596 ( .A1(n3773), .A2(n2024), .ZN(n2837) );
  AOI22_X1 U3597 ( .A1(n3609), .A2(REG0_REG_29__SCAN_IN), .B1(n2692), .B2(
        REG1_REG_29__SCAN_IN), .ZN(n2836) );
  OAI211_X1 U3598 ( .C1(n2839), .C2(n2838), .A(n2837), .B(n2836), .ZN(n3832)
         );
  INV_X1 U3599 ( .A(n2840), .ZN(n2841) );
  NAND2_X1 U3600 ( .A1(n4535), .A2(n2841), .ZN(n2842) );
  OR2_X1 U3601 ( .A1(n2843), .A2(n2842), .ZN(n3694) );
  NOR2_X1 U3602 ( .A1(n3723), .A2(n3694), .ZN(n2844) );
  NAND2_X1 U3603 ( .A1(n2849), .A2(n2844), .ZN(n3527) );
  INV_X1 U3604 ( .A(n2845), .ZN(n3690) );
  NOR2_X1 U3605 ( .A1(n2889), .A2(n4456), .ZN(n2846) );
  NAND2_X1 U3606 ( .A1(n2849), .A2(n2846), .ZN(n2847) );
  AOI22_X1 U3607 ( .A1(n3832), .A2(n3499), .B1(n3841), .B2(n3500), .ZN(n2851)
         );
  NOR2_X1 U3608 ( .A1(n3694), .A2(n4341), .ZN(n2848) );
  NAND2_X1 U3609 ( .A1(n2849), .A2(n2848), .ZN(n3531) );
  AOI22_X1 U3610 ( .A1(n3831), .A2(n3498), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n2850) );
  OAI211_X1 U3611 ( .C1(n3538), .C2(n3843), .A(n2851), .B(n2850), .ZN(n2852)
         );
  NOR2_X1 U3612 ( .A1(n2853), .A2(n2852), .ZN(n2854) );
  OAI211_X1 U3613 ( .C1(n2857), .C2(n2856), .A(n2855), .B(n2854), .ZN(U3217)
         );
  INV_X1 U3614 ( .A(n4535), .ZN(n2883) );
  INV_X1 U3615 ( .A(DATAI_3_), .ZN(n2859) );
  INV_X1 U3616 ( .A(n2858), .ZN(n2912) );
  MUX2_X1 U3617 ( .A(n2859), .B(n2912), .S(STATE_REG_SCAN_IN), .Z(n2860) );
  INV_X1 U3618 ( .A(n2860), .ZN(U3349) );
  INV_X1 U3619 ( .A(DATAI_4_), .ZN(n2861) );
  MUX2_X1 U3620 ( .A(n2861), .B(n3751), .S(STATE_REG_SCAN_IN), .Z(n2862) );
  INV_X1 U3621 ( .A(n2862), .ZN(U3348) );
  INV_X1 U3622 ( .A(DATAI_21_), .ZN(n2864) );
  NAND2_X1 U3623 ( .A1(n3687), .A2(STATE_REG_SCAN_IN), .ZN(n2863) );
  OAI21_X1 U3624 ( .B1(STATE_REG_SCAN_IN), .B2(n2864), .A(n2863), .ZN(U3331)
         );
  INV_X1 U3625 ( .A(DATAI_22_), .ZN(n2866) );
  NAND2_X1 U3626 ( .A1(n2390), .A2(STATE_REG_SCAN_IN), .ZN(n2865) );
  OAI21_X1 U3627 ( .B1(STATE_REG_SCAN_IN), .B2(n2866), .A(n2865), .ZN(U3330)
         );
  MUX2_X1 U3628 ( .A(n3768), .B(n2669), .S(U3149), .Z(n2867) );
  INV_X1 U3629 ( .A(n2867), .ZN(U3333) );
  INV_X1 U3630 ( .A(DATAI_27_), .ZN(n2869) );
  NAND2_X1 U3631 ( .A1(n4348), .A2(STATE_REG_SCAN_IN), .ZN(n2868) );
  OAI21_X1 U3632 ( .B1(STATE_REG_SCAN_IN), .B2(n2869), .A(n2868), .ZN(U3325)
         );
  INV_X1 U3633 ( .A(DATAI_20_), .ZN(n2871) );
  NAND2_X1 U3634 ( .A1(n3690), .A2(STATE_REG_SCAN_IN), .ZN(n2870) );
  OAI21_X1 U3635 ( .B1(STATE_REG_SCAN_IN), .B2(n2871), .A(n2870), .ZN(U3332)
         );
  INV_X1 U3636 ( .A(DATAI_9_), .ZN(n2872) );
  MUX2_X1 U3637 ( .A(n3122), .B(n2872), .S(U3149), .Z(n2873) );
  INV_X1 U3638 ( .A(n2873), .ZN(U3343) );
  INV_X1 U3639 ( .A(DATAI_25_), .ZN(n2876) );
  INV_X1 U3640 ( .A(n2884), .ZN(n2874) );
  NAND2_X1 U3641 ( .A1(n2874), .A2(STATE_REG_SCAN_IN), .ZN(n2875) );
  OAI21_X1 U3642 ( .B1(STATE_REG_SCAN_IN), .B2(n2876), .A(n2875), .ZN(U3327)
         );
  INV_X1 U3643 ( .A(DATAI_24_), .ZN(n2877) );
  MUX2_X1 U3644 ( .A(n2877), .B(n2799), .S(STATE_REG_SCAN_IN), .Z(n2878) );
  INV_X1 U3645 ( .A(n2878), .ZN(U3328) );
  INV_X1 U3646 ( .A(DATAI_26_), .ZN(n2880) );
  NAND2_X1 U3647 ( .A1(n2798), .A2(STATE_REG_SCAN_IN), .ZN(n2879) );
  OAI21_X1 U3648 ( .B1(STATE_REG_SCAN_IN), .B2(n2880), .A(n2879), .ZN(U3326)
         );
  INV_X1 U3649 ( .A(n2889), .ZN(n2882) );
  INV_X1 U3650 ( .A(D_REG_1__SCAN_IN), .ZN(n2885) );
  NOR2_X1 U3651 ( .A1(n2883), .A2(n2798), .ZN(n3373) );
  AOI22_X1 U3652 ( .A1(n4530), .A2(n2885), .B1(n3373), .B2(n2884), .ZN(U3459)
         );
  NOR2_X1 U3653 ( .A1(n4435), .A2(U4043), .ZN(U3148) );
  XNOR2_X1 U3654 ( .A(n2887), .B(n2886), .ZN(n3724) );
  NOR2_X1 U3655 ( .A1(n2889), .A2(n2888), .ZN(n3028) );
  NAND2_X1 U3656 ( .A1(n2890), .A2(n3028), .ZN(n2942) );
  NAND4_X1 U3657 ( .A1(n2894), .A2(n2893), .A3(n2892), .A4(n2891), .ZN(n3710)
         );
  OAI22_X1 U3658 ( .A1(n2988), .A2(n3527), .B1(n3526), .B2(n4509), .ZN(n2895)
         );
  AOI21_X1 U3659 ( .B1(REG3_REG_0__SCAN_IN), .B2(n2942), .A(n2895), .ZN(n2896)
         );
  OAI21_X1 U3660 ( .B1(n3724), .B2(n3517), .A(n2896), .ZN(U3229) );
  INV_X1 U3661 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n2898) );
  NAND2_X1 U3662 ( .A1(n3170), .A2(U4043), .ZN(n2897) );
  OAI21_X1 U3663 ( .B1(U4043), .B2(n2898), .A(n2897), .ZN(U3557) );
  INV_X1 U3664 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n2900) );
  INV_X1 U3665 ( .A(n4036), .ZN(n3800) );
  NAND2_X1 U3666 ( .A1(n3800), .A2(U4043), .ZN(n2899) );
  OAI21_X1 U3667 ( .B1(U4043), .B2(n2900), .A(n2899), .ZN(U3567) );
  INV_X1 U3668 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n2903) );
  INV_X1 U3669 ( .A(n3990), .ZN(n2901) );
  NAND2_X1 U3670 ( .A1(n2901), .A2(U4043), .ZN(n2902) );
  OAI21_X1 U3671 ( .B1(U4043), .B2(n2903), .A(n2902), .ZN(U3571) );
  INV_X1 U3672 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n4233) );
  NAND2_X1 U3673 ( .A1(n3325), .A2(U4043), .ZN(n2904) );
  OAI21_X1 U3674 ( .B1(U4043), .B2(n4233), .A(n2904), .ZN(U3565) );
  INV_X1 U3675 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n2906) );
  NAND2_X1 U3676 ( .A1(n3056), .A2(U4043), .ZN(n2905) );
  OAI21_X1 U3677 ( .B1(U4043), .B2(n2906), .A(n2905), .ZN(U3553) );
  INV_X1 U3678 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n2908) );
  INV_X1 U3679 ( .A(n3972), .ZN(n3810) );
  NAND2_X1 U3680 ( .A1(n3810), .A2(U4043), .ZN(n2907) );
  OAI21_X1 U3681 ( .B1(U4043), .B2(n2908), .A(n2907), .ZN(U3572) );
  AOI21_X1 U3682 ( .B1(n4612), .B2(n2910), .A(n2909), .ZN(n2918) );
  INV_X1 U3683 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3078) );
  NOR2_X1 U3684 ( .A1(STATE_REG_SCAN_IN), .A2(n3078), .ZN(n2950) );
  AOI21_X1 U3685 ( .B1(n4435), .B2(ADDR_REG_3__SCAN_IN), .A(n2950), .ZN(n2911)
         );
  OAI21_X1 U3686 ( .B1(n2912), .B2(n4431), .A(n2911), .ZN(n2917) );
  AOI211_X1 U3687 ( .C1(n2915), .C2(n2914), .A(n2913), .B(n4440), .ZN(n2916)
         );
  AOI211_X1 U3688 ( .C1(n4422), .C2(n2918), .A(n2917), .B(n2916), .ZN(n2919)
         );
  INV_X1 U3689 ( .A(n2919), .ZN(U3243) );
  AND2_X1 U3690 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n2958) );
  AOI211_X1 U3691 ( .C1(n2922), .C2(n2921), .A(n2920), .B(n4440), .ZN(n2923)
         );
  AOI211_X1 U3692 ( .C1(n4435), .C2(ADDR_REG_5__SCAN_IN), .A(n2958), .B(n2923), 
        .ZN(n2929) );
  AOI21_X1 U3693 ( .B1(n2926), .B2(n2925), .A(n2924), .ZN(n2927) );
  NAND2_X1 U3694 ( .A1(n4422), .A2(n2927), .ZN(n2928) );
  OAI211_X1 U3695 ( .C1(n4431), .C2(n2207), .A(n2929), .B(n2928), .ZN(U3245)
         );
  XNOR2_X1 U3696 ( .A(n2931), .B(n2930), .ZN(n2935) );
  AOI22_X1 U3697 ( .A1(n4491), .A2(n3499), .B1(n3498), .B2(n3711), .ZN(n2932)
         );
  OAI21_X1 U3698 ( .B1(n3526), .B2(n4502), .A(n2932), .ZN(n2933) );
  AOI21_X1 U3699 ( .B1(REG3_REG_1__SCAN_IN), .B2(n2942), .A(n2933), .ZN(n2934)
         );
  OAI21_X1 U3700 ( .B1(n2935), .B2(n3517), .A(n2934), .ZN(U3219) );
  INV_X1 U3701 ( .A(n2937), .ZN(n2938) );
  AOI21_X1 U3702 ( .B1(n2936), .B2(n2939), .A(n2938), .ZN(n2944) );
  AOI22_X1 U3703 ( .A1(n3710), .A2(n3498), .B1(n3499), .B2(n3056), .ZN(n2940)
         );
  OAI21_X1 U3704 ( .B1(n3526), .B2(n3062), .A(n2940), .ZN(n2941) );
  AOI21_X1 U3705 ( .B1(REG3_REG_2__SCAN_IN), .B2(n2942), .A(n2941), .ZN(n2943)
         );
  OAI21_X1 U3706 ( .B1(n2944), .B2(n3517), .A(n2943), .ZN(U3234) );
  NAND2_X1 U3707 ( .A1(n2946), .A2(n2945), .ZN(n2966) );
  OAI21_X1 U3708 ( .B1(n2945), .B2(n2946), .A(n2966), .ZN(n2947) );
  NAND2_X1 U3709 ( .A1(n2947), .A2(n3523), .ZN(n2952) );
  OAI22_X1 U3710 ( .A1(n2948), .A2(n3527), .B1(n3526), .B2(n3077), .ZN(n2949)
         );
  AOI211_X1 U3711 ( .C1(n3498), .C2(n4491), .A(n2950), .B(n2949), .ZN(n2951)
         );
  OAI211_X1 U3712 ( .C1(REG3_REG_3__SCAN_IN), .C2(n3538), .A(n2952), .B(n2951), 
        .ZN(U3215) );
  AND2_X1 U3713 ( .A1(n2954), .A2(n2953), .ZN(n2955) );
  XNOR2_X1 U3714 ( .A(n2956), .B(n2955), .ZN(n2961) );
  INV_X1 U3715 ( .A(n2948), .ZN(n3709) );
  INV_X1 U3716 ( .A(n3707), .ZN(n2997) );
  INV_X1 U3717 ( .A(n3137), .ZN(n3003) );
  OAI22_X1 U3718 ( .A1(n2997), .A2(n3527), .B1(n3526), .B2(n3003), .ZN(n2957)
         );
  AOI211_X1 U3719 ( .C1(n3498), .C2(n3709), .A(n2958), .B(n2957), .ZN(n2960)
         );
  NAND2_X1 U3720 ( .A1(n3514), .A2(n3141), .ZN(n2959) );
  OAI211_X1 U3721 ( .C1(n2961), .C2(n3517), .A(n2960), .B(n2959), .ZN(U3224)
         );
  INV_X1 U3722 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n2963) );
  NAND2_X1 U3723 ( .A1(n3913), .A2(U4043), .ZN(n2962) );
  OAI21_X1 U3724 ( .B1(U4043), .B2(n2963), .A(n2962), .ZN(U3575) );
  AND2_X1 U3725 ( .A1(n2964), .A2(n2966), .ZN(n2969) );
  NAND2_X1 U3726 ( .A1(n2966), .A2(n2965), .ZN(n2967) );
  OAI211_X1 U3727 ( .C1(n2969), .C2(n2968), .A(n3523), .B(n2967), .ZN(n2973)
         );
  AND2_X1 U3728 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3748) );
  INV_X1 U3729 ( .A(n3708), .ZN(n3004) );
  OAI22_X1 U3730 ( .A1(n3004), .A2(n3527), .B1(n3526), .B2(n2970), .ZN(n2971)
         );
  AOI211_X1 U3731 ( .C1(n3498), .C2(n3056), .A(n3748), .B(n2971), .ZN(n2972)
         );
  OAI211_X1 U3732 ( .C1(n3538), .C2(n3045), .A(n2973), .B(n2972), .ZN(U3227)
         );
  INV_X1 U3733 ( .A(n2975), .ZN(n2977) );
  NAND2_X1 U3734 ( .A1(n2977), .A2(n2976), .ZN(n2978) );
  XNOR2_X1 U3735 ( .A(n2974), .B(n2978), .ZN(n2979) );
  NAND2_X1 U3736 ( .A1(n2979), .A2(n3523), .ZN(n2985) );
  NAND2_X1 U3737 ( .A1(n3500), .A2(n3105), .ZN(n2982) );
  INV_X1 U3738 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2980) );
  NOR2_X1 U3739 ( .A1(STATE_REG_SCAN_IN), .A2(n2980), .ZN(n4356) );
  AOI21_X1 U3740 ( .B1(n3498), .B2(n3708), .A(n4356), .ZN(n2981) );
  OAI211_X1 U3741 ( .C1(n3369), .C2(n3527), .A(n2982), .B(n2981), .ZN(n2983)
         );
  INV_X1 U3742 ( .A(n2983), .ZN(n2984) );
  OAI211_X1 U3743 ( .C1(n3538), .C2(n3125), .A(n2985), .B(n2984), .ZN(U3236)
         );
  XNOR2_X1 U3744 ( .A(n3033), .B(n2390), .ZN(n2986) );
  NAND2_X1 U3745 ( .A1(n2986), .A2(n3768), .ZN(n4497) );
  INV_X1 U3746 ( .A(n4603), .ZN(n4572) );
  NAND2_X1 U3747 ( .A1(n4497), .A2(n4572), .ZN(n4588) );
  NAND2_X1 U3748 ( .A1(n2988), .A2(n2987), .ZN(n3000) );
  NAND2_X1 U3749 ( .A1(n3710), .A2(n4502), .ZN(n3552) );
  NAND2_X1 U3750 ( .A1(n3000), .A2(n3552), .ZN(n2998) );
  AND2_X1 U3751 ( .A1(n3711), .A2(n2999), .ZN(n4496) );
  NAND2_X1 U3752 ( .A1(n3710), .A2(n2987), .ZN(n2989) );
  NAND2_X1 U3753 ( .A1(n2990), .A2(n3055), .ZN(n3553) );
  NAND2_X1 U3754 ( .A1(n2990), .A2(n3062), .ZN(n2991) );
  NOR2_X1 U3755 ( .A1(n3056), .A2(n3558), .ZN(n2993) );
  NAND2_X1 U3756 ( .A1(n3056), .A2(n3558), .ZN(n2992) );
  NAND2_X1 U3757 ( .A1(n2948), .A2(n3043), .ZN(n3560) );
  NAND2_X1 U3758 ( .A1(n3709), .A2(n2970), .ZN(n3563) );
  NAND2_X1 U3759 ( .A1(n3560), .A2(n3563), .ZN(n3624) );
  NAND2_X1 U3760 ( .A1(n3026), .A2(n3624), .ZN(n2995) );
  NAND2_X1 U3761 ( .A1(n3709), .A2(n3043), .ZN(n2994) );
  AND2_X1 U3762 ( .A1(n3708), .A2(n3137), .ZN(n2996) );
  NAND2_X1 U3763 ( .A1(n2997), .A2(n3105), .ZN(n3565) );
  NAND2_X1 U3764 ( .A1(n3707), .A2(n3016), .ZN(n3568) );
  NAND2_X1 U3765 ( .A1(n3565), .A2(n3568), .ZN(n3623) );
  XNOR2_X1 U3766 ( .A(n3104), .B(n3623), .ZN(n3123) );
  INV_X1 U3767 ( .A(n3711), .ZN(n4494) );
  NAND2_X1 U3768 ( .A1(n4494), .A2(n2999), .ZN(n3647) );
  XNOR2_X1 U3769 ( .A(n3056), .B(n3558), .ZN(n3652) );
  NAND2_X1 U3770 ( .A1(n3001), .A2(n3652), .ZN(n3072) );
  INV_X1 U3771 ( .A(n3056), .ZN(n3557) );
  NAND2_X1 U3772 ( .A1(n3557), .A2(n3558), .ZN(n3559) );
  INV_X1 U3773 ( .A(n3560), .ZN(n3002) );
  AND2_X1 U3774 ( .A1(n3708), .A2(n3003), .ZN(n3131) );
  NAND2_X1 U3775 ( .A1(n3004), .A2(n3137), .ZN(n3569) );
  XNOR2_X1 U3776 ( .A(n3094), .B(n3623), .ZN(n3011) );
  NAND2_X1 U3777 ( .A1(n2390), .A2(n3763), .ZN(n3006) );
  NAND2_X1 U3778 ( .A1(n3687), .A2(n3690), .ZN(n3005) );
  NAND2_X1 U3779 ( .A1(n4341), .A2(n3008), .ZN(n4514) );
  OAI22_X1 U3780 ( .A1(n3369), .A2(n4514), .B1(n4456), .B2(n3016), .ZN(n3009)
         );
  AOI21_X1 U3781 ( .B1(n4460), .B2(n3708), .A(n3009), .ZN(n3010) );
  OAI21_X1 U3782 ( .B1(n3011), .B2(n4462), .A(n3010), .ZN(n3124) );
  AOI21_X1 U3783 ( .B1(n4588), .B2(n3123), .A(n3124), .ZN(n3025) );
  NAND2_X1 U3784 ( .A1(n3028), .A2(n3012), .ZN(n3013) );
  INV_X1 U3785 ( .A(n3140), .ZN(n3017) );
  AOI21_X1 U3786 ( .B1(n3105), .B2(n3017), .A(n3100), .ZN(n3127) );
  AOI22_X1 U3787 ( .A1(n3127), .A2(n4079), .B1(n4618), .B2(REG1_REG_6__SCAN_IN), .ZN(n3019) );
  OAI21_X1 U3788 ( .B1(n3025), .B2(n4618), .A(n3019), .ZN(U3524) );
  INV_X1 U3789 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3022) );
  NOR2_X1 U3790 ( .A1(n4606), .A2(n3022), .ZN(n3023) );
  AOI21_X1 U3791 ( .B1(n3127), .B2(n4148), .A(n3023), .ZN(n3024) );
  OAI21_X1 U3792 ( .B1(n3025), .B2(n4604), .A(n3024), .ZN(U3479) );
  INV_X1 U3793 ( .A(n3624), .ZN(n3035) );
  XNOR2_X1 U3794 ( .A(n3026), .B(n3035), .ZN(n4576) );
  INV_X1 U3795 ( .A(n4576), .ZN(n3049) );
  INV_X1 U3796 ( .A(n3027), .ZN(n3030) );
  NAND4_X1 U3797 ( .A1(n3031), .A2(n3030), .A3(n3029), .A4(n3028), .ZN(n3032)
         );
  INV_X2 U3798 ( .A(n4519), .ZN(n4521) );
  NOR2_X1 U3799 ( .A1(n3033), .A2(n3768), .ZN(n3034) );
  NAND2_X1 U3800 ( .A1(n4061), .A2(n3034), .ZN(n3108) );
  NAND2_X1 U3801 ( .A1(n4576), .A2(n4512), .ZN(n3042) );
  XNOR2_X1 U3802 ( .A(n3036), .B(n3035), .ZN(n3040) );
  NAND2_X1 U3803 ( .A1(n3056), .A2(n4460), .ZN(n3038) );
  INV_X1 U3804 ( .A(n4514), .ZN(n4490) );
  NAND2_X1 U3805 ( .A1(n3708), .A2(n4490), .ZN(n3037) );
  OAI211_X1 U3806 ( .C1(n4456), .C2(n2970), .A(n3038), .B(n3037), .ZN(n3039)
         );
  AOI21_X1 U3807 ( .B1(n3040), .B2(n4511), .A(n3039), .ZN(n3041) );
  NAND2_X1 U3808 ( .A1(n3042), .A2(n3041), .ZN(n4580) );
  AOI21_X1 U3809 ( .B1(n3076), .B2(n3043), .A(n3018), .ZN(n3044) );
  NAND2_X1 U3810 ( .A1(n3044), .A2(n3138), .ZN(n4577) );
  OAI22_X1 U3811 ( .A1(n4577), .A2(n3763), .B1(n4057), .B2(n3045), .ZN(n3046)
         );
  OAI21_X1 U3812 ( .B1(n4580), .B2(n3046), .A(n4061), .ZN(n3048) );
  NAND2_X1 U3813 ( .A1(n4521), .A2(REG2_REG_4__SCAN_IN), .ZN(n3047) );
  OAI211_X1 U3814 ( .C1(n3049), .C2(n3108), .A(n3048), .B(n3047), .ZN(U3286)
         );
  NAND2_X1 U3815 ( .A1(n3050), .A2(n3053), .ZN(n3051) );
  NAND2_X1 U3816 ( .A1(n3052), .A2(n3051), .ZN(n4570) );
  INV_X1 U3817 ( .A(n4570), .ZN(n3067) );
  NAND3_X1 U3818 ( .A1(n2073), .A2(n3000), .A3(n4486), .ZN(n3054) );
  NAND2_X1 U3819 ( .A1(n3070), .A2(n3054), .ZN(n3059) );
  AOI22_X1 U3820 ( .A1(n3056), .A2(n4490), .B1(n3055), .B2(n4489), .ZN(n3057)
         );
  OAI21_X1 U3821 ( .B1(n2988), .B2(n4493), .A(n3057), .ZN(n3058) );
  AOI21_X1 U3822 ( .B1(n3059), .B2(n4511), .A(n3058), .ZN(n3061) );
  NAND2_X1 U3823 ( .A1(n4570), .A2(n4512), .ZN(n3060) );
  AND2_X1 U3824 ( .A1(n3061), .A2(n3060), .ZN(n4567) );
  MUX2_X1 U3825 ( .A(n4567), .B(n4192), .S(n4521), .Z(n3066) );
  INV_X1 U3826 ( .A(n4057), .ZN(n4516) );
  AND2_X1 U3827 ( .A1(n4519), .A2(n3768), .ZN(n4041) );
  INV_X1 U3828 ( .A(n4501), .ZN(n3063) );
  NOR2_X1 U3829 ( .A1(n3063), .A2(n3062), .ZN(n4566) );
  NOR3_X1 U3830 ( .A1(n4056), .A2(n4565), .A3(n4566), .ZN(n3064) );
  AOI21_X1 U3831 ( .B1(n4516), .B2(REG3_REG_2__SCAN_IN), .A(n3064), .ZN(n3065)
         );
  OAI211_X1 U3832 ( .C1(n3067), .C2(n3108), .A(n3066), .B(n3065), .ZN(U3288)
         );
  XNOR2_X1 U3833 ( .A(n3068), .B(n3652), .ZN(n4573) );
  OAI22_X1 U3834 ( .A1(n2948), .A2(n4514), .B1(n4456), .B2(n3077), .ZN(n3074)
         );
  INV_X1 U3835 ( .A(n3652), .ZN(n3069) );
  NAND3_X1 U3836 ( .A1(n3070), .A2(n3553), .A3(n3069), .ZN(n3071) );
  AOI21_X1 U3837 ( .B1(n3072), .B2(n3071), .A(n4462), .ZN(n3073) );
  AOI211_X1 U3838 ( .C1(n4460), .C2(n4491), .A(n3074), .B(n3073), .ZN(n3075)
         );
  OAI21_X1 U3839 ( .B1(n4573), .B2(n4497), .A(n3075), .ZN(n4575) );
  INV_X1 U3840 ( .A(n4575), .ZN(n3083) );
  INV_X1 U3841 ( .A(n4573), .ZN(n3081) );
  INV_X1 U3842 ( .A(n3108), .ZN(n4517) );
  OAI21_X1 U3843 ( .B1(n4565), .B2(n3077), .A(n3076), .ZN(n4571) );
  AOI22_X1 U3844 ( .A1(n4521), .A2(REG2_REG_3__SCAN_IN), .B1(n4516), .B2(n3078), .ZN(n3079) );
  OAI21_X1 U3845 ( .B1(n4056), .B2(n4571), .A(n3079), .ZN(n3080) );
  AOI21_X1 U3846 ( .B1(n3081), .B2(n4517), .A(n3080), .ZN(n3082) );
  OAI21_X1 U3847 ( .B1(n3083), .B2(n4521), .A(n3082), .ZN(U3287) );
  AND2_X1 U3848 ( .A1(n3084), .A2(n3085), .ZN(n3088) );
  OAI211_X1 U3849 ( .C1(n3088), .C2(n3087), .A(n3523), .B(n3086), .ZN(n3092)
         );
  NOR2_X1 U3850 ( .A1(STATE_REG_SCAN_IN), .A2(n3089), .ZN(n4387) );
  INV_X1 U3851 ( .A(n3205), .ZN(n3227) );
  OAI22_X1 U3852 ( .A1(n3228), .A2(n3527), .B1(n3526), .B2(n3227), .ZN(n3090)
         );
  AOI211_X1 U3853 ( .C1(n3498), .C2(n3705), .A(n4387), .B(n3090), .ZN(n3091)
         );
  OAI211_X1 U3854 ( .C1(n3538), .C2(n3093), .A(n3092), .B(n3091), .ZN(U3214)
         );
  NAND2_X1 U3855 ( .A1(n3094), .A2(n3568), .ZN(n3095) );
  NAND2_X1 U3856 ( .A1(n3369), .A2(n3387), .ZN(n3151) );
  NAND2_X1 U3857 ( .A1(n3170), .A2(n3099), .ZN(n3574) );
  NAND2_X1 U3858 ( .A1(n3151), .A2(n3574), .ZN(n3621) );
  XNOR2_X1 U3859 ( .A(n3153), .B(n3621), .ZN(n3098) );
  INV_X1 U3860 ( .A(n3706), .ZN(n3154) );
  OAI22_X1 U3861 ( .A1(n3154), .A2(n4514), .B1(n4456), .B2(n3099), .ZN(n3096)
         );
  AOI21_X1 U3862 ( .B1(n4460), .B2(n3707), .A(n3096), .ZN(n3097) );
  OAI21_X1 U3863 ( .B1(n3098), .B2(n4462), .A(n3097), .ZN(n4586) );
  INV_X1 U3864 ( .A(n4586), .ZN(n3111) );
  INV_X1 U3865 ( .A(n3100), .ZN(n3101) );
  INV_X1 U3866 ( .A(n3159), .ZN(n3165) );
  AOI211_X1 U3867 ( .C1(n3387), .C2(n3101), .A(n3018), .B(n3165), .ZN(n4587)
         );
  OAI22_X1 U3868 ( .A1(n4061), .A2(n3102), .B1(n3388), .B2(n4057), .ZN(n3103)
         );
  AOI21_X1 U3869 ( .B1(n4587), .B2(n4041), .A(n3103), .ZN(n3110) );
  NAND2_X1 U3870 ( .A1(n3707), .A2(n3105), .ZN(n3144) );
  NAND2_X1 U3871 ( .A1(n3148), .A2(n3144), .ZN(n3106) );
  XOR2_X1 U3872 ( .A(n3621), .B(n3106), .Z(n4589) );
  NAND2_X1 U3873 ( .A1(n4061), .A2(n4512), .ZN(n3107) );
  NAND2_X1 U3874 ( .A1(n3108), .A2(n3107), .ZN(n3878) );
  NAND2_X1 U3875 ( .A1(n4589), .A2(n3878), .ZN(n3109) );
  OAI211_X1 U3876 ( .C1(n3111), .C2(n4521), .A(n3110), .B(n3109), .ZN(U3283)
         );
  OAI211_X1 U3877 ( .C1(n3114), .C2(n3113), .A(n4422), .B(n3112), .ZN(n3121)
         );
  INV_X1 U3878 ( .A(REG3_REG_9__SCAN_IN), .ZN(n4212) );
  NOR2_X1 U3879 ( .A1(STATE_REG_SCAN_IN), .A2(n4212), .ZN(n3466) );
  INV_X1 U3880 ( .A(n3115), .ZN(n3116) );
  AOI211_X1 U3881 ( .C1(n3118), .C2(n3117), .A(n3116), .B(n4440), .ZN(n3119)
         );
  AOI211_X1 U3882 ( .C1(n4435), .C2(ADDR_REG_9__SCAN_IN), .A(n3466), .B(n3119), 
        .ZN(n3120) );
  OAI211_X1 U3883 ( .C1(n4431), .C2(n3122), .A(n3121), .B(n3120), .ZN(U3249)
         );
  INV_X1 U3884 ( .A(n3123), .ZN(n3130) );
  NAND2_X1 U3885 ( .A1(n3124), .A2(n4519), .ZN(n3129) );
  OAI22_X1 U3886 ( .A1(n4061), .A2(n4355), .B1(n3125), .B2(n4057), .ZN(n3126)
         );
  AOI21_X1 U3887 ( .B1(n3127), .B2(n4504), .A(n3126), .ZN(n3128) );
  OAI211_X1 U3888 ( .C1(n4063), .C2(n3130), .A(n3129), .B(n3128), .ZN(U3284)
         );
  INV_X1 U3889 ( .A(n3131), .ZN(n3562) );
  NAND2_X1 U3890 ( .A1(n3562), .A2(n3569), .ZN(n3618) );
  XNOR2_X1 U3891 ( .A(n3132), .B(n3618), .ZN(n4581) );
  XNOR2_X1 U3892 ( .A(n3133), .B(n3618), .ZN(n3136) );
  AOI22_X1 U3893 ( .A1(n3707), .A2(n4490), .B1(n4489), .B2(n3137), .ZN(n3134)
         );
  OAI21_X1 U3894 ( .B1(n2948), .B2(n4493), .A(n3134), .ZN(n3135) );
  AOI21_X1 U3895 ( .B1(n3136), .B2(n4511), .A(n3135), .ZN(n4582) );
  MUX2_X1 U3896 ( .A(n4582), .B(n2205), .S(n4521), .Z(n3143) );
  AND2_X1 U3897 ( .A1(n3138), .A2(n3137), .ZN(n3139) );
  NOR2_X1 U3898 ( .A1(n3140), .A2(n3139), .ZN(n4585) );
  AOI22_X1 U3899 ( .A1(n4585), .A2(n4504), .B1(n3141), .B2(n4516), .ZN(n3142)
         );
  OAI211_X1 U3900 ( .C1(n4063), .C2(n4581), .A(n3143), .B(n3142), .ZN(U3285)
         );
  INV_X1 U3901 ( .A(n3467), .ZN(n3195) );
  AND2_X1 U3902 ( .A1(n3705), .A2(n3195), .ZN(n3188) );
  INV_X1 U3903 ( .A(n3188), .ZN(n3582) );
  INV_X1 U3904 ( .A(n3705), .ZN(n3196) );
  NAND2_X1 U3905 ( .A1(n3196), .A2(n3467), .ZN(n3581) );
  NAND2_X1 U3906 ( .A1(n3582), .A2(n3581), .ZN(n3619) );
  NAND2_X1 U3907 ( .A1(n3170), .A2(n3387), .ZN(n3145) );
  AND2_X1 U3908 ( .A1(n3144), .A2(n3145), .ZN(n3147) );
  INV_X1 U3909 ( .A(n3145), .ZN(n3146) );
  AND2_X1 U3910 ( .A1(n3706), .A2(n3367), .ZN(n3150) );
  INV_X1 U3911 ( .A(n3367), .ZN(n3168) );
  NAND2_X1 U3912 ( .A1(n3154), .A2(n3168), .ZN(n3149) );
  OAI21_X1 U3913 ( .B1(n3166), .B2(n3150), .A(n3149), .ZN(n3198) );
  XOR2_X1 U3914 ( .A(n3619), .B(n3198), .Z(n4592) );
  INV_X1 U3915 ( .A(n3151), .ZN(n3152) );
  NAND2_X1 U3916 ( .A1(n3154), .A2(n3367), .ZN(n3580) );
  NAND2_X1 U3917 ( .A1(n3706), .A2(n3168), .ZN(n3575) );
  NAND2_X1 U3918 ( .A1(n3155), .A2(n3575), .ZN(n3189) );
  XOR2_X1 U3919 ( .A(n3619), .B(n3189), .Z(n3158) );
  INV_X1 U3920 ( .A(n4459), .ZN(n3214) );
  OAI22_X1 U3921 ( .A1(n3214), .A2(n4514), .B1(n4456), .B2(n3195), .ZN(n3156)
         );
  AOI21_X1 U3922 ( .B1(n4460), .B2(n3706), .A(n3156), .ZN(n3157) );
  OAI21_X1 U3923 ( .B1(n3158), .B2(n4462), .A(n3157), .ZN(n4594) );
  NAND2_X1 U3924 ( .A1(n4594), .A2(n4519), .ZN(n3163) );
  INV_X1 U3925 ( .A(n3206), .ZN(n3225) );
  AOI21_X1 U3926 ( .B1(n3467), .B2(n3164), .A(n3225), .ZN(n4595) );
  OAI22_X1 U3927 ( .A1(n4061), .A2(n3160), .B1(n3468), .B2(n4057), .ZN(n3161)
         );
  AOI21_X1 U3928 ( .B1(n4595), .B2(n4504), .A(n3161), .ZN(n3162) );
  OAI211_X1 U3929 ( .C1(n4063), .C2(n4592), .A(n3163), .B(n3162), .ZN(U3281)
         );
  OAI21_X1 U3930 ( .B1(n3165), .B2(n3168), .A(n3164), .ZN(n4480) );
  INV_X1 U3931 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3175) );
  NAND2_X1 U3932 ( .A1(n3580), .A2(n3575), .ZN(n3639) );
  XOR2_X1 U3933 ( .A(n3639), .B(n3166), .Z(n4482) );
  XOR2_X1 U3934 ( .A(n3639), .B(n3167), .Z(n3172) );
  OAI22_X1 U3935 ( .A1(n3196), .A2(n4514), .B1(n4456), .B2(n3168), .ZN(n3169)
         );
  AOI21_X1 U3936 ( .B1(n4460), .B2(n3170), .A(n3169), .ZN(n3171) );
  OAI21_X1 U3937 ( .B1(n3172), .B2(n4462), .A(n3171), .ZN(n3173) );
  AOI21_X1 U3938 ( .B1(n4512), .B2(n4482), .A(n3173), .ZN(n4485) );
  INV_X1 U3939 ( .A(n4485), .ZN(n3174) );
  AOI21_X1 U3940 ( .B1(n4603), .B2(n4482), .A(n3174), .ZN(n3177) );
  MUX2_X1 U3941 ( .A(n3175), .B(n3177), .S(n4606), .Z(n3176) );
  OAI21_X1 U3942 ( .B1(n4480), .B2(n4331), .A(n3176), .ZN(U3483) );
  MUX2_X1 U3943 ( .A(n2504), .B(n3177), .S(n4621), .Z(n3178) );
  OAI21_X1 U3944 ( .B1(n4480), .B2(n4133), .A(n3178), .ZN(U3526) );
  XNOR2_X1 U3945 ( .A(n3180), .B(n3179), .ZN(n3181) );
  XNOR2_X1 U3946 ( .A(n3182), .B(n3181), .ZN(n3186) );
  INV_X1 U3947 ( .A(n3228), .ZN(n3704) );
  NOR2_X1 U3948 ( .A1(STATE_REG_SCAN_IN), .A2(n4202), .ZN(n4406) );
  AOI21_X1 U3949 ( .B1(n3704), .B2(n3498), .A(n4406), .ZN(n3184) );
  AOI22_X1 U3950 ( .A1(n3500), .A2(n3257), .B1(n3499), .B2(n3702), .ZN(n3183)
         );
  OAI211_X1 U3951 ( .C1(n3208), .C2(n3538), .A(n3184), .B(n3183), .ZN(n3185)
         );
  AOI21_X1 U3952 ( .B1(n3186), .B2(n3523), .A(n3185), .ZN(n3187) );
  INV_X1 U3953 ( .A(n3187), .ZN(U3221) );
  NAND2_X1 U3954 ( .A1(n4459), .A2(n3227), .ZN(n3542) );
  NAND2_X1 U3955 ( .A1(n3214), .A2(n3205), .ZN(n3541) );
  NAND2_X1 U3956 ( .A1(n3704), .A2(n4467), .ZN(n3543) );
  NAND2_X1 U3957 ( .A1(n4455), .A2(n3543), .ZN(n3190) );
  NAND2_X1 U3958 ( .A1(n3228), .A2(n3212), .ZN(n3545) );
  INV_X1 U3959 ( .A(n3257), .ZN(n3260) );
  XNOR2_X1 U3960 ( .A(n3703), .B(n3260), .ZN(n3654) );
  INV_X1 U3961 ( .A(n3654), .ZN(n3191) );
  XNOR2_X1 U3962 ( .A(n3259), .B(n3191), .ZN(n3194) );
  AOI22_X1 U3963 ( .A1(n3702), .A2(n4490), .B1(n4489), .B2(n3257), .ZN(n3192)
         );
  OAI21_X1 U3964 ( .B1(n3228), .B2(n4493), .A(n3192), .ZN(n3193) );
  AOI21_X1 U3965 ( .B1(n3194), .B2(n4511), .A(n3193), .ZN(n3250) );
  NOR2_X1 U3966 ( .A1(n3705), .A2(n3467), .ZN(n3197) );
  OAI22_X2 U3967 ( .A1(n3198), .A2(n3197), .B1(n3196), .B2(n3195), .ZN(n4450)
         );
  AND2_X1 U3968 ( .A1(n4459), .A2(n3205), .ZN(n4449) );
  NAND2_X1 U3969 ( .A1(n3228), .A2(n4467), .ZN(n3200) );
  INV_X1 U3970 ( .A(n3200), .ZN(n3199) );
  NAND2_X1 U3971 ( .A1(n3545), .A2(n3543), .ZN(n4454) );
  NOR2_X1 U3972 ( .A1(n3199), .A2(n4454), .ZN(n3202) );
  OR2_X1 U3973 ( .A1(n4449), .A2(n3202), .ZN(n3204) );
  NAND2_X1 U3974 ( .A1(n3214), .A2(n3227), .ZN(n4451) );
  AND2_X1 U3975 ( .A1(n4451), .A2(n3200), .ZN(n3201) );
  OR2_X1 U3976 ( .A1(n3202), .A2(n3201), .ZN(n3203) );
  XNOR2_X1 U3977 ( .A(n3258), .B(n3654), .ZN(n3249) );
  NAND2_X1 U3978 ( .A1(n4466), .A2(n3257), .ZN(n3207) );
  NAND2_X1 U3979 ( .A1(n3265), .A2(n3207), .ZN(n3256) );
  NOR2_X1 U3980 ( .A1(n3256), .A2(n4056), .ZN(n3210) );
  OAI22_X1 U3981 ( .A1(n4061), .A2(n4405), .B1(n3208), .B2(n4057), .ZN(n3209)
         );
  AOI211_X1 U3982 ( .C1(n3249), .C2(n3878), .A(n3210), .B(n3209), .ZN(n3211)
         );
  OAI21_X1 U3983 ( .B1(n4521), .B2(n3250), .A(n3211), .ZN(U3278) );
  AOI22_X1 U3984 ( .A1(n3500), .A2(n3212), .B1(n3499), .B2(n3703), .ZN(n3213)
         );
  NAND2_X1 U3985 ( .A1(REG3_REG_11__SCAN_IN), .A2(U3149), .ZN(n4395) );
  OAI211_X1 U3986 ( .C1(n3214), .C2(n3531), .A(n3213), .B(n4395), .ZN(n3222)
         );
  INV_X1 U3987 ( .A(n3215), .ZN(n3220) );
  AOI21_X1 U3988 ( .B1(n3219), .B2(n3217), .A(n3216), .ZN(n3218) );
  AOI211_X1 U3989 ( .C1(n3220), .C2(n3219), .A(n3517), .B(n3218), .ZN(n3221)
         );
  AOI211_X1 U3990 ( .C1(n3514), .C2(n4465), .A(n3222), .B(n3221), .ZN(n3223)
         );
  INV_X1 U3991 ( .A(n3223), .ZN(U3233) );
  INV_X1 U3992 ( .A(n4468), .ZN(n3224) );
  OAI21_X1 U3993 ( .B1(n3225), .B2(n3227), .A(n3224), .ZN(n4473) );
  INV_X1 U3994 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3234) );
  NAND2_X1 U3995 ( .A1(n3541), .A2(n3542), .ZN(n3620) );
  XOR2_X1 U3996 ( .A(n3620), .B(n4450), .Z(n4475) );
  XNOR2_X1 U3997 ( .A(n3226), .B(n3620), .ZN(n3231) );
  OAI22_X1 U3998 ( .A1(n3228), .A2(n4514), .B1(n4456), .B2(n3227), .ZN(n3229)
         );
  AOI21_X1 U3999 ( .B1(n4460), .B2(n3705), .A(n3229), .ZN(n3230) );
  OAI21_X1 U4000 ( .B1(n3231), .B2(n4462), .A(n3230), .ZN(n3232) );
  AOI21_X1 U4001 ( .B1(n4475), .B2(n4512), .A(n3232), .ZN(n4478) );
  INV_X1 U4002 ( .A(n4478), .ZN(n3233) );
  AOI21_X1 U4003 ( .B1(n4603), .B2(n4475), .A(n3233), .ZN(n3236) );
  MUX2_X1 U4004 ( .A(n3234), .B(n3236), .S(n4606), .Z(n3235) );
  OAI21_X1 U4005 ( .B1(n4473), .B2(n4331), .A(n3235), .ZN(U3487) );
  MUX2_X1 U4006 ( .A(n2534), .B(n3236), .S(n4621), .Z(n3237) );
  OAI21_X1 U4007 ( .B1(n4473), .B2(n4133), .A(n3237), .ZN(U3528) );
  INV_X1 U4008 ( .A(n3239), .ZN(n3241) );
  NAND2_X1 U4009 ( .A1(n3241), .A2(n3240), .ZN(n3242) );
  XNOR2_X1 U4010 ( .A(n3238), .B(n3242), .ZN(n3243) );
  NAND2_X1 U4011 ( .A1(n3243), .A2(n3523), .ZN(n3248) );
  NAND2_X1 U4012 ( .A1(n3500), .A2(n3281), .ZN(n3245) );
  AND2_X1 U4013 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n3337) );
  AOI21_X1 U4014 ( .B1(n3498), .B2(n3703), .A(n3337), .ZN(n3244) );
  OAI211_X1 U4015 ( .C1(n3532), .C2(n3527), .A(n3245), .B(n3244), .ZN(n3246)
         );
  INV_X1 U4016 ( .A(n3246), .ZN(n3247) );
  OAI211_X1 U4017 ( .C1(n3538), .C2(n3267), .A(n3248), .B(n3247), .ZN(U3231)
         );
  NAND2_X1 U4018 ( .A1(n3249), .A2(n4588), .ZN(n3251) );
  AND2_X1 U4019 ( .A1(n3251), .A2(n3250), .ZN(n3253) );
  MUX2_X1 U4020 ( .A(n4271), .B(n3253), .S(n4621), .Z(n3252) );
  OAI21_X1 U4021 ( .B1(n4133), .B2(n3256), .A(n3252), .ZN(U3530) );
  INV_X1 U4022 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3254) );
  MUX2_X1 U4023 ( .A(n3254), .B(n3253), .S(n4606), .Z(n3255) );
  OAI21_X1 U4024 ( .B1(n3256), .B2(n4331), .A(n3255), .ZN(U3491) );
  INV_X1 U4025 ( .A(n3703), .ZN(n4457) );
  INV_X1 U4026 ( .A(n3702), .ZN(n3292) );
  NAND2_X1 U4027 ( .A1(n3292), .A2(n3281), .ZN(n3548) );
  NAND2_X1 U4028 ( .A1(n3702), .A2(n2165), .ZN(n3286) );
  NAND2_X1 U4029 ( .A1(n3548), .A2(n3286), .ZN(n3638) );
  XNOR2_X1 U4030 ( .A(n3284), .B(n3638), .ZN(n4143) );
  NOR2_X1 U4031 ( .A1(n3703), .A2(n3260), .ZN(n3547) );
  NAND2_X1 U4032 ( .A1(n3703), .A2(n3260), .ZN(n3285) );
  NAND2_X1 U4033 ( .A1(n3287), .A2(n3285), .ZN(n3261) );
  XOR2_X1 U4034 ( .A(n3638), .B(n3261), .Z(n3264) );
  OAI22_X1 U4035 ( .A1(n3532), .A2(n4514), .B1(n4456), .B2(n2165), .ZN(n3262)
         );
  AOI21_X1 U4036 ( .B1(n4460), .B2(n3703), .A(n3262), .ZN(n3263) );
  OAI21_X1 U4037 ( .B1(n3264), .B2(n4462), .A(n3263), .ZN(n4140) );
  NAND2_X1 U4038 ( .A1(n4140), .A2(n4519), .ZN(n3271) );
  AND2_X1 U4039 ( .A1(n3265), .A2(n3281), .ZN(n3266) );
  NOR2_X1 U4040 ( .A1(n3294), .A2(n3266), .ZN(n4141) );
  OAI22_X1 U4041 ( .A1(n4061), .A2(n3268), .B1(n3267), .B2(n4057), .ZN(n3269)
         );
  AOI21_X1 U4042 ( .B1(n4141), .B2(n4504), .A(n3269), .ZN(n3270) );
  OAI211_X1 U40430 ( .C1(n4063), .C2(n4143), .A(n3271), .B(n3270), .ZN(U3277)
         );
  XOR2_X1 U4044 ( .A(n3274), .B(n3273), .Z(n3275) );
  XNOR2_X1 U4045 ( .A(n3272), .B(n3275), .ZN(n3280) );
  INV_X1 U4046 ( .A(n3297), .ZN(n3278) );
  AOI22_X1 U4047 ( .A1(n3500), .A2(n3295), .B1(n3499), .B2(n3325), .ZN(n3276)
         );
  NAND2_X1 U4048 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4415) );
  OAI211_X1 U4049 ( .C1(n3292), .C2(n3531), .A(n3276), .B(n4415), .ZN(n3277)
         );
  AOI21_X1 U4050 ( .B1(n3278), .B2(n3514), .A(n3277), .ZN(n3279) );
  OAI21_X1 U4051 ( .B1(n3280), .B2(n3517), .A(n3279), .ZN(U3212) );
  AND2_X1 U4052 ( .A1(n3702), .A2(n3281), .ZN(n3283) );
  NAND2_X1 U4053 ( .A1(n3292), .A2(n2165), .ZN(n3282) );
  NAND2_X1 U4054 ( .A1(n3532), .A2(n3295), .ZN(n3657) );
  INV_X1 U4055 ( .A(n3532), .ZN(n3701) );
  NAND2_X1 U4056 ( .A1(n3701), .A2(n3302), .ZN(n3539) );
  NAND2_X1 U4057 ( .A1(n3657), .A2(n3539), .ZN(n3626) );
  XNOR2_X1 U4058 ( .A(n3304), .B(n3626), .ZN(n4134) );
  INV_X1 U4059 ( .A(n3626), .ZN(n3288) );
  AND2_X1 U4060 ( .A1(n3286), .A2(n3285), .ZN(n3546) );
  OAI21_X1 U4061 ( .B1(n3288), .B2(n3660), .A(n3322), .ZN(n3289) );
  NAND2_X1 U4062 ( .A1(n3289), .A2(n4511), .ZN(n3291) );
  AOI22_X1 U4063 ( .A1(n3325), .A2(n4490), .B1(n4489), .B2(n3295), .ZN(n3290)
         );
  OAI211_X1 U4064 ( .C1(n3292), .C2(n4493), .A(n3291), .B(n3290), .ZN(n3293)
         );
  AOI21_X1 U4065 ( .B1(n4134), .B2(n4512), .A(n3293), .ZN(n4138) );
  INV_X1 U4066 ( .A(n3309), .ZN(n4136) );
  INV_X1 U4067 ( .A(n3294), .ZN(n3296) );
  NAND2_X1 U4068 ( .A1(n3296), .A2(n3295), .ZN(n4135) );
  AND3_X1 U4069 ( .A1(n4136), .A2(n4504), .A3(n4135), .ZN(n3300) );
  OAI22_X1 U4070 ( .A1(n4061), .A2(n3298), .B1(n3297), .B2(n4057), .ZN(n3299)
         );
  AOI211_X1 U4071 ( .C1(n4134), .C2(n4517), .A(n3300), .B(n3299), .ZN(n3301)
         );
  OAI21_X1 U4072 ( .B1(n4138), .B2(n4521), .A(n3301), .ZN(U3276) );
  INV_X1 U4073 ( .A(n3325), .ZN(n3436) );
  NAND2_X1 U4074 ( .A1(n3436), .A2(n3315), .ZN(n3656) );
  NAND2_X1 U4075 ( .A1(n3325), .A2(n3525), .ZN(n3540) );
  NAND2_X1 U4076 ( .A1(n3656), .A2(n3540), .ZN(n3625) );
  XOR2_X1 U4077 ( .A(n3317), .B(n3625), .Z(n4130) );
  INV_X1 U4078 ( .A(n4130), .ZN(n3314) );
  NAND2_X1 U4079 ( .A1(n3322), .A2(n3657), .ZN(n3305) );
  XNOR2_X1 U4080 ( .A(n3305), .B(n3625), .ZN(n3308) );
  OAI22_X1 U4081 ( .A1(n3528), .A2(n4514), .B1(n4456), .B2(n3525), .ZN(n3306)
         );
  AOI21_X1 U4082 ( .B1(n4460), .B2(n3701), .A(n3306), .ZN(n3307) );
  OAI21_X1 U4083 ( .B1(n3308), .B2(n4462), .A(n3307), .ZN(n4129) );
  OR2_X1 U4084 ( .A1(n3309), .A2(n3525), .ZN(n3310) );
  NAND2_X1 U4085 ( .A1(n3328), .A2(n3310), .ZN(n4332) );
  NOR2_X1 U4086 ( .A1(n4332), .A2(n4056), .ZN(n3312) );
  OAI22_X1 U4087 ( .A1(n4061), .A2(n2261), .B1(n3537), .B2(n4057), .ZN(n3311)
         );
  AOI211_X1 U4088 ( .C1(n4129), .C2(n4061), .A(n3312), .B(n3311), .ZN(n3313)
         );
  OAI21_X1 U4089 ( .B1(n3314), .B2(n4063), .A(n3313), .ZN(U3275) );
  NAND2_X1 U4090 ( .A1(n3317), .A2(n3316), .ZN(n3319) );
  NAND2_X1 U4091 ( .A1(n3319), .A2(n3318), .ZN(n3799) );
  NAND2_X1 U4092 ( .A1(n3528), .A2(n3797), .ZN(n3662) );
  NAND2_X1 U4093 ( .A1(n4049), .A2(n3329), .ZN(n3776) );
  NAND2_X1 U4094 ( .A1(n3662), .A2(n3776), .ZN(n3798) );
  INV_X1 U4095 ( .A(n3798), .ZN(n3774) );
  XNOR2_X1 U4096 ( .A(n3799), .B(n3774), .ZN(n4126) );
  INV_X1 U4097 ( .A(n4126), .ZN(n3334) );
  INV_X1 U4098 ( .A(n3657), .ZN(n3320) );
  NOR2_X1 U4099 ( .A1(n3625), .A2(n3320), .ZN(n3321) );
  NAND2_X1 U4100 ( .A1(n3322), .A2(n3321), .ZN(n3323) );
  NAND2_X1 U4101 ( .A1(n3323), .A2(n3540), .ZN(n3775) );
  XNOR2_X1 U4102 ( .A(n3775), .B(n3774), .ZN(n3327) );
  OAI22_X1 U4103 ( .A1(n4036), .A2(n4514), .B1(n4456), .B2(n3329), .ZN(n3324)
         );
  AOI21_X1 U4104 ( .B1(n4460), .B2(n3325), .A(n3324), .ZN(n3326) );
  OAI21_X1 U4105 ( .B1(n3327), .B2(n4462), .A(n3326), .ZN(n4125) );
  OAI21_X1 U4106 ( .B1(n2163), .B2(n3329), .A(n4052), .ZN(n4327) );
  INV_X1 U4107 ( .A(n3330), .ZN(n3438) );
  AOI22_X1 U4108 ( .A1(n4521), .A2(REG2_REG_16__SCAN_IN), .B1(n3438), .B2(
        n4516), .ZN(n3331) );
  OAI21_X1 U4109 ( .B1(n4327), .B2(n4056), .A(n3331), .ZN(n3332) );
  AOI21_X1 U4110 ( .B1(n4125), .B2(n4519), .A(n3332), .ZN(n3333) );
  OAI21_X1 U4111 ( .B1(n3334), .B2(n4063), .A(n3333), .ZN(U3274) );
  XNOR2_X1 U4112 ( .A(n3336), .B(n3335), .ZN(n3344) );
  AOI21_X1 U4113 ( .B1(n4435), .B2(ADDR_REG_13__SCAN_IN), .A(n3337), .ZN(n3338) );
  OAI21_X1 U4114 ( .B1(n2255), .B2(n4431), .A(n3338), .ZN(n3343) );
  XNOR2_X1 U4115 ( .A(n4337), .B(REG2_REG_13__SCAN_IN), .ZN(n3340) );
  OAI21_X1 U4116 ( .B1(n3341), .B2(n3340), .A(n4426), .ZN(n3339) );
  AOI21_X1 U4117 ( .B1(n3341), .B2(n3340), .A(n3339), .ZN(n3342) );
  AOI211_X1 U4118 ( .C1(n4422), .C2(n3344), .A(n3343), .B(n3342), .ZN(n3345)
         );
  INV_X1 U4119 ( .A(n3345), .ZN(U3253) );
  NAND3_X1 U4120 ( .A1(n3346), .A2(STATE_REG_SCAN_IN), .A3(IR_REG_31__SCAN_IN), 
        .ZN(n3348) );
  INV_X1 U4121 ( .A(DATAI_31_), .ZN(n3347) );
  OAI22_X1 U4122 ( .A1(n2152), .A2(n3348), .B1(STATE_REG_SCAN_IN), .B2(n3347), 
        .ZN(U3321) );
  NAND2_X1 U4123 ( .A1(n3349), .A2(DATAI_31_), .ZN(n3683) );
  NAND2_X1 U4124 ( .A1(n3349), .A2(DATAI_29_), .ZN(n3631) );
  INV_X1 U4125 ( .A(n3631), .ZN(n3824) );
  NAND2_X1 U4126 ( .A1(n3349), .A2(DATAI_30_), .ZN(n4066) );
  NAND2_X1 U4127 ( .A1(n4067), .A2(n4066), .ZN(n4065) );
  XOR2_X1 U4128 ( .A(n3683), .B(n4065), .Z(n3361) );
  INV_X1 U4129 ( .A(REG1_REG_31__SCAN_IN), .ZN(n3355) );
  INV_X1 U4130 ( .A(REG2_REG_31__SCAN_IN), .ZN(n3350) );
  OR2_X1 U4131 ( .A1(n2839), .A2(n3350), .ZN(n3352) );
  NAND2_X1 U4132 ( .A1(n3609), .A2(REG0_REG_31__SCAN_IN), .ZN(n3351) );
  OAI211_X1 U4133 ( .C1(n2397), .C2(n3355), .A(n3352), .B(n3351), .ZN(n3699)
         );
  AOI21_X1 U4134 ( .B1(n4348), .B2(B_REG_SCAN_IN), .A(n4514), .ZN(n3791) );
  NAND2_X1 U4135 ( .A1(n3699), .A2(n3791), .ZN(n4068) );
  OAI21_X1 U4136 ( .B1(n3683), .B2(n4456), .A(n4068), .ZN(n3359) );
  NAND2_X1 U4137 ( .A1(n3359), .A2(n4606), .ZN(n3354) );
  NAND2_X1 U4138 ( .A1(n4604), .A2(REG0_REG_31__SCAN_IN), .ZN(n3353) );
  OAI211_X1 U4139 ( .C1(n3361), .C2(n4331), .A(n3354), .B(n3353), .ZN(U3517)
         );
  NOR2_X1 U4140 ( .A1(n4621), .A2(n3355), .ZN(n3356) );
  AOI21_X1 U4141 ( .B1(n4621), .B2(n3359), .A(n3356), .ZN(n3357) );
  OAI21_X1 U4142 ( .B1(n3361), .B2(n4133), .A(n3357), .ZN(U3549) );
  NOR2_X1 U4143 ( .A1(n4061), .A2(n3350), .ZN(n3358) );
  AOI21_X1 U4144 ( .B1(n3359), .B2(n4519), .A(n3358), .ZN(n3360) );
  OAI21_X1 U4145 ( .B1(n3361), .B2(n4056), .A(n3360), .ZN(U3260) );
  XOR2_X1 U4146 ( .A(n3363), .B(n3362), .Z(n3364) );
  XNOR2_X1 U4147 ( .A(n3365), .B(n3364), .ZN(n3372) );
  INV_X1 U4148 ( .A(n3366), .ZN(n4479) );
  AOI22_X1 U4149 ( .A1(n3500), .A2(n3367), .B1(n3499), .B2(n3705), .ZN(n3368)
         );
  NAND2_X1 U4150 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n4377) );
  OAI211_X1 U4151 ( .C1(n3369), .C2(n3531), .A(n3368), .B(n4377), .ZN(n3370)
         );
  AOI21_X1 U4152 ( .B1(n4479), .B2(n3514), .A(n3370), .ZN(n3371) );
  OAI21_X1 U4153 ( .B1(n3372), .B2(n3517), .A(n3371), .ZN(U3218) );
  INV_X1 U4154 ( .A(D_REG_0__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4155 ( .A1(n4530), .A2(n3374), .B1(n3373), .B2(n2799), .ZN(U3458)
         );
  XNOR2_X1 U4156 ( .A(n3376), .B(n3375), .ZN(n3382) );
  INV_X1 U4157 ( .A(n3862), .ZN(n3380) );
  OAI22_X1 U4158 ( .A1(n3895), .A2(n3531), .B1(STATE_REG_SCAN_IN), .B2(n3377), 
        .ZN(n3379) );
  OAI22_X1 U4159 ( .A1(n3854), .A2(n3527), .B1(n3526), .B2(n3860), .ZN(n3378)
         );
  AOI211_X1 U4160 ( .C1(n3380), .C2(n3514), .A(n3379), .B(n3378), .ZN(n3381)
         );
  OAI21_X1 U4161 ( .B1(n3382), .B2(n3517), .A(n3381), .ZN(U3211) );
  AOI21_X1 U4162 ( .B1(n3383), .B2(n3384), .A(n3517), .ZN(n3386) );
  OR2_X1 U4163 ( .A1(n3383), .A2(n3384), .ZN(n3385) );
  NAND2_X1 U4164 ( .A1(n3386), .A2(n3385), .ZN(n3393) );
  NOR2_X1 U4165 ( .A1(STATE_REG_SCAN_IN), .A2(n2491), .ZN(n4366) );
  AOI21_X1 U4166 ( .B1(n3498), .B2(n3707), .A(n4366), .ZN(n3392) );
  AOI22_X1 U4167 ( .A1(n3500), .A2(n3387), .B1(n3499), .B2(n3706), .ZN(n3391)
         );
  INV_X1 U4168 ( .A(n3388), .ZN(n3389) );
  NAND2_X1 U4169 ( .A1(n3514), .A2(n3389), .ZN(n3390) );
  NAND4_X1 U4170 ( .A1(n3393), .A2(n3392), .A3(n3391), .A4(n3390), .ZN(U3210)
         );
  INV_X1 U4171 ( .A(n3394), .ZN(n3398) );
  OAI21_X1 U4172 ( .B1(n2022), .B2(n3396), .A(n3395), .ZN(n3397) );
  NAND3_X1 U4173 ( .A1(n3398), .A2(n3523), .A3(n3397), .ZN(n3403) );
  OAI22_X1 U4174 ( .A1(n3814), .A2(n3527), .B1(n3526), .B2(n3941), .ZN(n3401)
         );
  OAI22_X1 U4175 ( .A1(n3972), .A2(n3531), .B1(STATE_REG_SCAN_IN), .B2(n3399), 
        .ZN(n3400) );
  NOR2_X1 U4176 ( .A1(n3401), .A2(n3400), .ZN(n3402) );
  OAI211_X1 U4177 ( .C1(n3538), .C2(n3944), .A(n3403), .B(n3402), .ZN(U3213)
         );
  XOR2_X1 U4178 ( .A(n3405), .B(n3404), .Z(n3410) );
  INV_X1 U4179 ( .A(n4020), .ZN(n3408) );
  AOI22_X1 U4180 ( .A1(n3500), .A2(n4014), .B1(n3499), .B2(n4015), .ZN(n3406)
         );
  NAND2_X1 U4181 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3766) );
  OAI211_X1 U4182 ( .C1(n4047), .C2(n3531), .A(n3406), .B(n3766), .ZN(n3407)
         );
  AOI21_X1 U4183 ( .B1(n3408), .B2(n3514), .A(n3407), .ZN(n3409) );
  OAI21_X1 U4184 ( .B1(n3410), .B2(n3517), .A(n3409), .ZN(U3216) );
  XNOR2_X1 U4185 ( .A(n3412), .B(n3411), .ZN(n3413) );
  XNOR2_X1 U4186 ( .A(n3414), .B(n3413), .ZN(n3415) );
  NAND2_X1 U4187 ( .A1(n3415), .A2(n3523), .ZN(n3420) );
  AOI22_X1 U4188 ( .A1(n3498), .A2(n4015), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3417) );
  NAND2_X1 U4189 ( .A1(n3500), .A2(n3598), .ZN(n3416) );
  OAI211_X1 U4190 ( .C1(n3972), .C2(n3527), .A(n3417), .B(n3416), .ZN(n3418)
         );
  INV_X1 U4191 ( .A(n3418), .ZN(n3419) );
  OAI211_X1 U4192 ( .C1(n3538), .C2(n3978), .A(n3420), .B(n3419), .ZN(U3220)
         );
  INV_X1 U4193 ( .A(n3422), .ZN(n3423) );
  NOR2_X1 U4194 ( .A1(n3424), .A2(n3423), .ZN(n3425) );
  XNOR2_X1 U4195 ( .A(n3421), .B(n3425), .ZN(n3431) );
  INV_X1 U4196 ( .A(n3426), .ZN(n3902) );
  INV_X1 U4197 ( .A(n3899), .ZN(n3894) );
  OAI22_X1 U4198 ( .A1(n3814), .A2(n3531), .B1(n3526), .B2(n3894), .ZN(n3429)
         );
  OAI22_X1 U4199 ( .A1(n3895), .A2(n3527), .B1(STATE_REG_SCAN_IN), .B2(n3427), 
        .ZN(n3428) );
  AOI211_X1 U4200 ( .C1(n3902), .C2(n3514), .A(n3429), .B(n3428), .ZN(n3430)
         );
  OAI21_X1 U4201 ( .B1(n3431), .B2(n3517), .A(n3430), .ZN(U3222) );
  AOI21_X1 U4202 ( .B1(n3521), .B2(n3519), .A(n3432), .ZN(n3434) );
  XNOR2_X1 U4203 ( .A(n3434), .B(n3433), .ZN(n3440) );
  AOI22_X1 U4204 ( .A1(n3800), .A2(n3499), .B1(n3500), .B2(n3797), .ZN(n3435)
         );
  NAND2_X1 U4205 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4445) );
  OAI211_X1 U4206 ( .C1(n3436), .C2(n3531), .A(n3435), .B(n4445), .ZN(n3437)
         );
  AOI21_X1 U4207 ( .B1(n3438), .B2(n3514), .A(n3437), .ZN(n3439) );
  OAI21_X1 U4208 ( .B1(n3440), .B2(n3517), .A(n3439), .ZN(U3223) );
  XNOR2_X1 U4209 ( .A(n3443), .B(n3442), .ZN(n3444) );
  XNOR2_X1 U4210 ( .A(n3441), .B(n3444), .ZN(n3445) );
  NAND2_X1 U4211 ( .A1(n3445), .A2(n3523), .ZN(n3451) );
  OAI22_X1 U4212 ( .A1(n4047), .A2(n3527), .B1(n3526), .B2(n4055), .ZN(n3449)
         );
  INV_X1 U4213 ( .A(n3446), .ZN(n3447) );
  OAI21_X1 U4214 ( .B1(n3528), .B2(n3531), .A(n3447), .ZN(n3448) );
  NOR2_X1 U4215 ( .A1(n3449), .A2(n3448), .ZN(n3450) );
  OAI211_X1 U4216 ( .C1(n3538), .C2(n4058), .A(n3451), .B(n3450), .ZN(U3225)
         );
  NAND2_X1 U4217 ( .A1(n3453), .A2(n3452), .ZN(n3455) );
  XNOR2_X1 U4218 ( .A(n3455), .B(n3454), .ZN(n3456) );
  NAND2_X1 U4219 ( .A1(n3456), .A2(n3523), .ZN(n3461) );
  AOI22_X1 U4220 ( .A1(n3498), .A2(n3953), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3460) );
  AOI22_X1 U4221 ( .A1(n3500), .A2(n3813), .B1(n3499), .B2(n3913), .ZN(n3459)
         );
  INV_X1 U4222 ( .A(n3919), .ZN(n3457) );
  NAND2_X1 U4223 ( .A1(n3514), .A2(n3457), .ZN(n3458) );
  NAND4_X1 U4224 ( .A1(n3461), .A2(n3460), .A3(n3459), .A4(n3458), .ZN(U3226)
         );
  INV_X1 U4225 ( .A(n3084), .ZN(n3463) );
  AOI21_X1 U4226 ( .B1(n3464), .B2(n3462), .A(n3463), .ZN(n3465) );
  OR2_X1 U4227 ( .A1(n3465), .A2(n3517), .ZN(n3473) );
  AOI21_X1 U4228 ( .B1(n3498), .B2(n3706), .A(n3466), .ZN(n3472) );
  AOI22_X1 U4229 ( .A1(n3500), .A2(n3467), .B1(n3499), .B2(n4459), .ZN(n3471)
         );
  INV_X1 U4230 ( .A(n3468), .ZN(n3469) );
  NAND2_X1 U4231 ( .A1(n3514), .A2(n3469), .ZN(n3470) );
  NAND4_X1 U4232 ( .A1(n3473), .A2(n3472), .A3(n3471), .A4(n3470), .ZN(U3228)
         );
  NOR2_X1 U4233 ( .A1(n3474), .A2(n2149), .ZN(n3479) );
  AOI21_X1 U4234 ( .B1(n3477), .B2(n3476), .A(n3475), .ZN(n3478) );
  OAI21_X1 U4235 ( .B1(n3479), .B2(n3478), .A(n3523), .ZN(n3484) );
  AOI22_X1 U4236 ( .A1(n3498), .A2(n4034), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n3481) );
  NAND2_X1 U4237 ( .A1(n3500), .A2(n3632), .ZN(n3480) );
  OAI211_X1 U4238 ( .C1(n3990), .C2(n3527), .A(n3481), .B(n3480), .ZN(n3482)
         );
  INV_X1 U4239 ( .A(n3482), .ZN(n3483) );
  OAI211_X1 U4240 ( .C1(n3538), .C2(n3997), .A(n3484), .B(n3483), .ZN(U3230)
         );
  AOI21_X1 U4241 ( .B1(n3486), .B2(n3485), .A(n2022), .ZN(n3492) );
  INV_X1 U4242 ( .A(n3964), .ZN(n3490) );
  OAI22_X1 U4243 ( .A1(n3990), .A2(n3531), .B1(STATE_REG_SCAN_IN), .B2(n3487), 
        .ZN(n3489) );
  INV_X1 U4244 ( .A(n3953), .ZN(n3911) );
  OAI22_X1 U4245 ( .A1(n3911), .A2(n3527), .B1(n3526), .B2(n3601), .ZN(n3488)
         );
  AOI211_X1 U4246 ( .C1(n3490), .C2(n3514), .A(n3489), .B(n3488), .ZN(n3491)
         );
  OAI21_X1 U4247 ( .B1(n3492), .B2(n3517), .A(n3491), .ZN(U3232) );
  INV_X1 U4248 ( .A(n3493), .ZN(n3495) );
  NOR2_X1 U4249 ( .A1(n3495), .A2(n3494), .ZN(n3496) );
  XNOR2_X1 U4250 ( .A(n2045), .B(n3496), .ZN(n3504) );
  AOI21_X1 U4251 ( .B1(n3800), .B2(n3498), .A(n3497), .ZN(n3502) );
  AOI22_X1 U4252 ( .A1(n3500), .A2(n4033), .B1(n3499), .B2(n4034), .ZN(n3501)
         );
  OAI211_X1 U4253 ( .C1(n4030), .C2(n3538), .A(n3502), .B(n3501), .ZN(n3503)
         );
  AOI21_X1 U4254 ( .B1(n3504), .B2(n3523), .A(n3503), .ZN(n3505) );
  INV_X1 U4255 ( .A(n3505), .ZN(U3235) );
  INV_X1 U4256 ( .A(n3506), .ZN(n3508) );
  NAND2_X1 U4257 ( .A1(n3508), .A2(n3507), .ZN(n3509) );
  XNOR2_X1 U4258 ( .A(n3510), .B(n3509), .ZN(n3518) );
  INV_X1 U4259 ( .A(n3882), .ZN(n3515) );
  OAI22_X1 U4260 ( .A1(n3817), .A2(n3531), .B1(n3526), .B2(n3881), .ZN(n3513)
         );
  INV_X1 U4261 ( .A(n3831), .ZN(n3873) );
  OAI22_X1 U4262 ( .A1(n3873), .A2(n3527), .B1(STATE_REG_SCAN_IN), .B2(n3511), 
        .ZN(n3512) );
  AOI211_X1 U4263 ( .C1(n3515), .C2(n3514), .A(n3513), .B(n3512), .ZN(n3516)
         );
  OAI21_X1 U4264 ( .B1(n3518), .B2(n3517), .A(n3516), .ZN(U3237) );
  INV_X1 U4265 ( .A(n3519), .ZN(n3520) );
  NOR2_X1 U4266 ( .A1(n3432), .A2(n3520), .ZN(n3522) );
  XNOR2_X1 U4267 ( .A(n3522), .B(n3521), .ZN(n3524) );
  NAND2_X1 U4268 ( .A1(n3524), .A2(n3523), .ZN(n3536) );
  OAI22_X1 U4269 ( .A1(n3528), .A2(n3527), .B1(n3526), .B2(n3525), .ZN(n3534)
         );
  NOR2_X1 U4270 ( .A1(STATE_REG_SCAN_IN), .A2(n3529), .ZN(n4433) );
  INV_X1 U4271 ( .A(n4433), .ZN(n3530) );
  OAI21_X1 U4272 ( .B1(n3532), .B2(n3531), .A(n3530), .ZN(n3533) );
  NOR2_X1 U4273 ( .A1(n3534), .A2(n3533), .ZN(n3535) );
  OAI211_X1 U4274 ( .C1(n3538), .C2(n3537), .A(n3536), .B(n3535), .ZN(U3238)
         );
  NOR2_X1 U4275 ( .A1(n3990), .A2(n3598), .ZN(n3930) );
  NAND2_X1 U4276 ( .A1(n3540), .A2(n3539), .ZN(n3579) );
  NAND2_X1 U4277 ( .A1(n3579), .A2(n3656), .ZN(n3658) );
  INV_X1 U4278 ( .A(n3658), .ZN(n3588) );
  INV_X1 U4279 ( .A(n3541), .ZN(n3551) );
  AND2_X1 U4280 ( .A1(n3543), .A2(n3542), .ZN(n3544) );
  AND2_X1 U4281 ( .A1(n3546), .A2(n3544), .ZN(n3583) );
  OAI21_X1 U4282 ( .B1(n2080), .B2(n3547), .A(n3546), .ZN(n3549) );
  NAND4_X1 U4283 ( .A1(n3549), .A2(n3657), .A3(n3548), .A4(n3656), .ZN(n3550)
         );
  AOI21_X1 U4284 ( .B1(n3551), .B2(n3583), .A(n3550), .ZN(n3587) );
  INV_X1 U4285 ( .A(n3647), .ZN(n4487) );
  NAND2_X1 U4286 ( .A1(n3711), .A2(n4509), .ZN(n3646) );
  OAI211_X1 U4287 ( .C1(n4487), .C2(n3687), .A(n3646), .B(n3552), .ZN(n3554)
         );
  NAND3_X1 U4288 ( .A1(n3554), .A2(n3553), .A3(n3000), .ZN(n3556) );
  OAI211_X1 U4289 ( .C1(n3558), .C2(n3557), .A(n3556), .B(n3555), .ZN(n3561)
         );
  NAND3_X1 U4290 ( .A1(n3561), .A2(n3560), .A3(n3559), .ZN(n3564) );
  NAND4_X1 U4291 ( .A1(n3564), .A2(n3563), .A3(n3562), .A4(n3568), .ZN(n3567)
         );
  INV_X1 U4292 ( .A(n3621), .ZN(n3566) );
  NAND3_X1 U4293 ( .A1(n3567), .A2(n3566), .A3(n3565), .ZN(n3573) );
  INV_X1 U4294 ( .A(n3579), .ZN(n3572) );
  INV_X1 U4295 ( .A(n3568), .ZN(n3570) );
  NOR2_X1 U4296 ( .A1(n3570), .A2(n3569), .ZN(n3571) );
  AOI22_X1 U4297 ( .A1(n3573), .A2(n3572), .B1(n3571), .B2(n3658), .ZN(n3578)
         );
  INV_X1 U4298 ( .A(n3574), .ZN(n3577) );
  INV_X1 U4299 ( .A(n3575), .ZN(n3576) );
  NOR3_X1 U4300 ( .A1(n3578), .A2(n3577), .A3(n3576), .ZN(n3585) );
  AOI21_X1 U4301 ( .B1(n3581), .B2(n3580), .A(n3579), .ZN(n3584) );
  OAI211_X1 U4302 ( .C1(n3585), .C2(n3584), .A(n3583), .B(n3582), .ZN(n3586)
         );
  OAI21_X1 U4303 ( .B1(n3588), .B2(n3587), .A(n3586), .ZN(n3589) );
  NAND2_X1 U4304 ( .A1(n3589), .A2(n3776), .ZN(n3591) );
  NAND2_X1 U4305 ( .A1(n4015), .A2(n3995), .ZN(n3664) );
  INV_X1 U4306 ( .A(n3664), .ZN(n3779) );
  INV_X1 U4307 ( .A(n4047), .ZN(n3700) );
  NAND2_X1 U4308 ( .A1(n3700), .A2(n4029), .ZN(n4009) );
  NAND2_X1 U4309 ( .A1(n4034), .A2(n4019), .ZN(n3590) );
  AND2_X1 U4310 ( .A1(n4009), .A2(n3590), .ZN(n3592) );
  OR2_X1 U4311 ( .A1(n4036), .A2(n3801), .ZN(n4005) );
  NAND2_X1 U4312 ( .A1(n3592), .A2(n4005), .ZN(n3778) );
  AOI211_X1 U4313 ( .C1(n3591), .C2(n3662), .A(n3779), .B(n3778), .ZN(n3597)
         );
  NAND2_X1 U4314 ( .A1(n4047), .A2(n4033), .ZN(n4008) );
  NAND2_X1 U4315 ( .A1(n4036), .A2(n3801), .ZN(n4006) );
  NAND2_X1 U4316 ( .A1(n4008), .A2(n4006), .ZN(n3593) );
  NAND2_X1 U4317 ( .A1(n3593), .A2(n3592), .ZN(n3595) );
  NAND2_X1 U4318 ( .A1(n3804), .A2(n4014), .ZN(n3594) );
  NAND2_X1 U4319 ( .A1(n3595), .A2(n3594), .ZN(n3985) );
  NOR2_X1 U4320 ( .A1(n4015), .A2(n3995), .ZN(n3596) );
  OR2_X1 U4321 ( .A1(n3985), .A2(n3596), .ZN(n3665) );
  AND2_X1 U4322 ( .A1(n3665), .A2(n3664), .ZN(n3780) );
  NOR2_X1 U4323 ( .A1(n3597), .A2(n3780), .ZN(n3599) );
  NAND2_X1 U4324 ( .A1(n3972), .A2(n3963), .ZN(n3934) );
  NAND2_X1 U4325 ( .A1(n3990), .A2(n3598), .ZN(n3932) );
  AND2_X1 U4326 ( .A1(n3934), .A2(n3932), .ZN(n3782) );
  OAI21_X1 U4327 ( .B1(n3930), .B2(n3599), .A(n3782), .ZN(n3600) );
  INV_X1 U4328 ( .A(n3600), .ZN(n3602) );
  NAND2_X1 U4329 ( .A1(n3810), .A2(n3601), .ZN(n3622) );
  NAND2_X1 U4330 ( .A1(n3953), .A2(n3941), .ZN(n3637) );
  NAND2_X1 U4331 ( .A1(n3622), .A2(n3637), .ZN(n3667) );
  NAND2_X1 U4332 ( .A1(n3895), .A2(n3871), .ZN(n3634) );
  NAND2_X1 U4333 ( .A1(n3817), .A2(n3899), .ZN(n3868) );
  NAND2_X1 U4334 ( .A1(n3634), .A2(n3868), .ZN(n3603) );
  INV_X1 U4335 ( .A(n3603), .ZN(n3787) );
  NAND2_X1 U4336 ( .A1(n3911), .A2(n3808), .ZN(n3907) );
  NAND2_X1 U4337 ( .A1(n3814), .A2(n3813), .ZN(n3636) );
  OAI211_X1 U4338 ( .C1(n3602), .C2(n3667), .A(n3787), .B(n3785), .ZN(n3607)
         );
  NAND2_X1 U4339 ( .A1(n3913), .A2(n3894), .ZN(n3635) );
  NAND2_X1 U4340 ( .A1(n3938), .A2(n3917), .ZN(n3889) );
  AND2_X1 U4341 ( .A1(n3635), .A2(n3889), .ZN(n3867) );
  NAND2_X1 U4342 ( .A1(n3852), .A2(n3881), .ZN(n3676) );
  OAI21_X1 U4343 ( .B1(n3603), .B2(n3867), .A(n3676), .ZN(n3786) );
  INV_X1 U4344 ( .A(n3786), .ZN(n3606) );
  NAND2_X1 U4345 ( .A1(n3821), .A2(n3604), .ZN(n3788) );
  INV_X1 U4346 ( .A(n3788), .ZN(n3605) );
  AOI21_X1 U4347 ( .B1(n3832), .B2(n3631), .A(n3605), .ZN(n3675) );
  NAND2_X1 U4348 ( .A1(n3831), .A2(n3860), .ZN(n3644) );
  NAND4_X1 U4349 ( .A1(n3607), .A2(n3606), .A3(n3675), .A4(n3644), .ZN(n3616)
         );
  NAND2_X1 U4350 ( .A1(n3854), .A2(n3841), .ZN(n3617) );
  OR2_X1 U4351 ( .A1(n3831), .A2(n3860), .ZN(n3828) );
  NAND2_X1 U4352 ( .A1(n3617), .A2(n3828), .ZN(n3789) );
  INV_X1 U4353 ( .A(n3832), .ZN(n3613) );
  INV_X1 U4354 ( .A(REG1_REG_30__SCAN_IN), .ZN(n3612) );
  INV_X1 U4355 ( .A(REG2_REG_30__SCAN_IN), .ZN(n3608) );
  OR2_X1 U4356 ( .A1(n2839), .A2(n3608), .ZN(n3611) );
  NAND2_X1 U4357 ( .A1(n3609), .A2(REG0_REG_30__SCAN_IN), .ZN(n3610) );
  OAI211_X1 U4358 ( .C1(n2397), .C2(n3612), .A(n3611), .B(n3610), .ZN(n3792)
         );
  NAND2_X1 U4359 ( .A1(n3699), .A2(n3683), .ZN(n3615) );
  OAI21_X1 U4360 ( .B1(n3792), .B2(n4066), .A(n3615), .ZN(n3649) );
  AOI21_X1 U4361 ( .B1(n3613), .B2(n3824), .A(n3649), .ZN(n3672) );
  INV_X1 U4362 ( .A(n3672), .ZN(n3614) );
  AOI21_X1 U4363 ( .B1(n3675), .B2(n3789), .A(n3614), .ZN(n3677) );
  NAND2_X1 U4364 ( .A1(n3792), .A2(n4066), .ZN(n3684) );
  OAI21_X1 U4365 ( .B1(n3699), .B2(n3683), .A(n3684), .ZN(n3648) );
  AOI22_X1 U4366 ( .A1(n3616), .A2(n3677), .B1(n3615), .B2(n3648), .ZN(n3692)
         );
  NAND2_X1 U4367 ( .A1(n3617), .A2(n3788), .ZN(n3836) );
  NOR3_X1 U4368 ( .A1(n3836), .A2(n3619), .A3(n3618), .ZN(n3630) );
  NAND2_X1 U4369 ( .A1(n4008), .A2(n4009), .ZN(n4032) );
  NOR4_X1 U4370 ( .A1(n4032), .A2(n4454), .A3(n3621), .A4(n3620), .ZN(n3629)
         );
  INV_X1 U4371 ( .A(n3952), .ZN(n3960) );
  NOR4_X1 U4372 ( .A1(n3960), .A2(n3798), .A3(n3624), .A4(n3623), .ZN(n3628)
         );
  NOR4_X1 U4373 ( .A1(n2073), .A2(n3626), .A3(n2998), .A4(n3625), .ZN(n3627)
         );
  AND4_X1 U4374 ( .A1(n3630), .A2(n3629), .A3(n3628), .A4(n3627), .ZN(n3643)
         );
  XNOR2_X1 U4375 ( .A(n3832), .B(n3631), .ZN(n3822) );
  INV_X1 U4376 ( .A(n3822), .ZN(n3642) );
  NOR2_X1 U4377 ( .A1(n4015), .A2(n3632), .ZN(n3806) );
  NAND2_X1 U4378 ( .A1(n4015), .A2(n3632), .ZN(n3807) );
  INV_X1 U4379 ( .A(n3807), .ZN(n3633) );
  NOR2_X1 U4380 ( .A1(n3806), .A2(n3633), .ZN(n3988) );
  NAND2_X1 U4381 ( .A1(n3634), .A2(n3676), .ZN(n3877) );
  NAND2_X1 U4382 ( .A1(n3868), .A2(n3635), .ZN(n3892) );
  NAND2_X1 U4383 ( .A1(n3889), .A2(n3636), .ZN(n3909) );
  NOR4_X1 U4384 ( .A1(n3988), .A2(n3877), .A3(n3892), .A4(n3909), .ZN(n3641)
         );
  NAND2_X1 U4385 ( .A1(n3907), .A2(n3637), .ZN(n3935) );
  NAND2_X1 U4386 ( .A1(n4005), .A2(n4006), .ZN(n4046) );
  NOR4_X1 U4387 ( .A1(n3935), .A2(n4046), .A3(n3639), .A4(n3638), .ZN(n3640)
         );
  NAND4_X1 U4388 ( .A1(n3643), .A2(n3642), .A3(n3641), .A4(n3640), .ZN(n3655)
         );
  XNOR2_X1 U4389 ( .A(n4034), .B(n4014), .ZN(n4003) );
  INV_X1 U4390 ( .A(n4003), .ZN(n4011) );
  INV_X1 U4391 ( .A(n3932), .ZN(n3645) );
  OR2_X1 U4392 ( .A1(n3930), .A2(n3645), .ZN(n3970) );
  NAND2_X1 U4393 ( .A1(n3647), .A2(n3646), .ZN(n4559) );
  NOR2_X1 U4394 ( .A1(n3970), .A2(n4559), .ZN(n3651) );
  NOR2_X1 U4395 ( .A1(n3649), .A2(n3648), .ZN(n3650) );
  NAND4_X1 U4396 ( .A1(n3857), .A2(n3652), .A3(n3651), .A4(n3650), .ZN(n3653)
         );
  NOR4_X1 U4397 ( .A1(n3655), .A2(n3654), .A3(n4011), .A4(n3653), .ZN(n3689)
         );
  NAND2_X1 U4398 ( .A1(n3657), .A2(n3656), .ZN(n3659) );
  OAI21_X1 U4399 ( .B1(n3660), .B2(n3659), .A(n3658), .ZN(n3663) );
  INV_X1 U4400 ( .A(n3776), .ZN(n3661) );
  AOI211_X1 U4401 ( .C1(n3663), .C2(n3662), .A(n3661), .B(n3778), .ZN(n3666)
         );
  OAI21_X1 U4402 ( .B1(n3666), .B2(n3665), .A(n3664), .ZN(n3669) );
  AOI21_X1 U4403 ( .B1(n3930), .B2(n3934), .A(n3667), .ZN(n3783) );
  INV_X1 U4404 ( .A(n3783), .ZN(n3668) );
  AOI21_X1 U4405 ( .B1(n3669), .B2(n3782), .A(n3668), .ZN(n3671) );
  INV_X1 U4406 ( .A(n3785), .ZN(n3670) );
  OAI21_X1 U4407 ( .B1(n3671), .B2(n3670), .A(n3867), .ZN(n3674) );
  INV_X1 U4408 ( .A(n3789), .ZN(n3673) );
  NAND4_X1 U4409 ( .A1(n3674), .A2(n3673), .A3(n3787), .A4(n3672), .ZN(n3682)
         );
  INV_X1 U4410 ( .A(n3675), .ZN(n3679) );
  NAND2_X1 U4411 ( .A1(n3857), .A2(n3676), .ZN(n3678) );
  OAI21_X1 U4412 ( .B1(n3679), .B2(n3678), .A(n3677), .ZN(n3681) );
  INV_X1 U4413 ( .A(n4066), .ZN(n4070) );
  INV_X1 U4414 ( .A(n3699), .ZN(n3680) );
  AOI22_X1 U4415 ( .A1(n3682), .A2(n3681), .B1(n4070), .B2(n3680), .ZN(n3686)
         );
  AOI21_X1 U4416 ( .B1(n3684), .B2(n3699), .A(n3683), .ZN(n3685) );
  NOR2_X1 U4417 ( .A1(n3686), .A2(n3685), .ZN(n3688) );
  MUX2_X1 U4418 ( .A(n3689), .B(n3688), .S(n3687), .Z(n3691) );
  MUX2_X1 U4419 ( .A(n3692), .B(n3691), .S(n3690), .Z(n3693) );
  XNOR2_X1 U4420 ( .A(n3693), .B(n3763), .ZN(n3698) );
  NOR2_X1 U4421 ( .A1(n3730), .A2(n3694), .ZN(n3696) );
  OAI21_X1 U4422 ( .B1(n3697), .B2(n2390), .A(B_REG_SCAN_IN), .ZN(n3695) );
  OAI22_X1 U4423 ( .A1(n3698), .A2(n3697), .B1(n3696), .B2(n3695), .ZN(U3239)
         );
  MUX2_X1 U4424 ( .A(n3699), .B(DATAO_REG_31__SCAN_IN), .S(n3726), .Z(U3581)
         );
  MUX2_X1 U4425 ( .A(n3792), .B(DATAO_REG_30__SCAN_IN), .S(n3726), .Z(U3580)
         );
  MUX2_X1 U4426 ( .A(n3832), .B(DATAO_REG_29__SCAN_IN), .S(n3726), .Z(U3579)
         );
  MUX2_X1 U4427 ( .A(n3821), .B(DATAO_REG_28__SCAN_IN), .S(n3726), .Z(U3578)
         );
  MUX2_X1 U4428 ( .A(n3831), .B(DATAO_REG_27__SCAN_IN), .S(n3726), .Z(U3577)
         );
  MUX2_X1 U4429 ( .A(n3852), .B(DATAO_REG_26__SCAN_IN), .S(n3726), .Z(U3576)
         );
  MUX2_X1 U4430 ( .A(n3938), .B(DATAO_REG_24__SCAN_IN), .S(n3726), .Z(U3574)
         );
  MUX2_X1 U4431 ( .A(n3953), .B(DATAO_REG_23__SCAN_IN), .S(n3726), .Z(U3573)
         );
  MUX2_X1 U4432 ( .A(n4015), .B(DATAO_REG_20__SCAN_IN), .S(n3726), .Z(U3570)
         );
  MUX2_X1 U4433 ( .A(n4034), .B(DATAO_REG_19__SCAN_IN), .S(n3726), .Z(U3569)
         );
  MUX2_X1 U4434 ( .A(DATAO_REG_18__SCAN_IN), .B(n3700), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4435 ( .A(DATAO_REG_16__SCAN_IN), .B(n4049), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4436 ( .A(DATAO_REG_14__SCAN_IN), .B(n3701), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4437 ( .A(n3702), .B(DATAO_REG_13__SCAN_IN), .S(n3726), .Z(U3563)
         );
  MUX2_X1 U4438 ( .A(n3703), .B(DATAO_REG_12__SCAN_IN), .S(n3726), .Z(U3562)
         );
  MUX2_X1 U4439 ( .A(DATAO_REG_11__SCAN_IN), .B(n3704), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4440 ( .A(n4459), .B(DATAO_REG_10__SCAN_IN), .S(n3726), .Z(U3560)
         );
  MUX2_X1 U4441 ( .A(n3705), .B(DATAO_REG_9__SCAN_IN), .S(n3726), .Z(U3559) );
  MUX2_X1 U4442 ( .A(n3706), .B(DATAO_REG_8__SCAN_IN), .S(n3726), .Z(U3558) );
  MUX2_X1 U4443 ( .A(n3707), .B(DATAO_REG_6__SCAN_IN), .S(n3726), .Z(U3556) );
  MUX2_X1 U4444 ( .A(n3708), .B(DATAO_REG_5__SCAN_IN), .S(n3726), .Z(U3555) );
  MUX2_X1 U4445 ( .A(DATAO_REG_4__SCAN_IN), .B(n3709), .S(U4043), .Z(U3554) );
  MUX2_X1 U4446 ( .A(DATAO_REG_2__SCAN_IN), .B(n4491), .S(U4043), .Z(U3552) );
  MUX2_X1 U4447 ( .A(DATAO_REG_1__SCAN_IN), .B(n3710), .S(U4043), .Z(U3551) );
  MUX2_X1 U4448 ( .A(n3711), .B(DATAO_REG_0__SCAN_IN), .S(n3726), .Z(U3550) );
  OAI211_X1 U4449 ( .C1(n3714), .C2(n3713), .A(n4422), .B(n3712), .ZN(n3721)
         );
  OAI211_X1 U4450 ( .C1(n3717), .C2(n3716), .A(n4426), .B(n3715), .ZN(n3720)
         );
  AOI22_X1 U4451 ( .A1(n4435), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3719) );
  NAND2_X1 U4452 ( .A1(n2349), .A2(n4339), .ZN(n3718) );
  NAND4_X1 U4453 ( .A1(n3721), .A2(n3720), .A3(n3719), .A4(n3718), .ZN(U3241)
         );
  NAND3_X1 U4454 ( .A1(n3724), .A2(n3723), .A3(n3722), .ZN(n3728) );
  AND2_X1 U4455 ( .A1(n4348), .A2(n2421), .ZN(n3725) );
  OR2_X1 U4456 ( .A1(n4341), .A2(n3725), .ZN(n4346) );
  AOI21_X1 U4457 ( .B1(n4346), .B2(n2090), .A(n3726), .ZN(n3727) );
  OAI211_X1 U4458 ( .C1(n3730), .C2(n3729), .A(n3728), .B(n3727), .ZN(n3757)
         );
  INV_X1 U4459 ( .A(n2188), .ZN(n3733) );
  NAND2_X1 U4460 ( .A1(n4435), .A2(ADDR_REG_2__SCAN_IN), .ZN(n3732) );
  NAND2_X1 U4461 ( .A1(U3149), .A2(REG3_REG_2__SCAN_IN), .ZN(n3731) );
  OAI211_X1 U4462 ( .C1(n4431), .C2(n3733), .A(n3732), .B(n3731), .ZN(n3734)
         );
  INV_X1 U4463 ( .A(n3734), .ZN(n3743) );
  OAI211_X1 U4464 ( .C1(n3737), .C2(n3736), .A(n4426), .B(n3735), .ZN(n3742)
         );
  OAI211_X1 U4465 ( .C1(n3740), .C2(n3739), .A(n4422), .B(n3738), .ZN(n3741)
         );
  NAND4_X1 U4466 ( .A1(n3757), .A2(n3743), .A3(n3742), .A4(n3741), .ZN(U3242)
         );
  INV_X1 U4467 ( .A(n3744), .ZN(n3745) );
  NAND2_X1 U4468 ( .A1(n3745), .A2(n2113), .ZN(n3746) );
  NAND3_X1 U4469 ( .A1(n4426), .A2(n3747), .A3(n3746), .ZN(n3750) );
  AOI21_X1 U4470 ( .B1(n4435), .B2(ADDR_REG_4__SCAN_IN), .A(n3748), .ZN(n3749)
         );
  OAI211_X1 U4471 ( .C1(n4431), .C2(n3751), .A(n3750), .B(n3749), .ZN(n3752)
         );
  INV_X1 U4472 ( .A(n3752), .ZN(n3756) );
  OAI211_X1 U4473 ( .C1(REG1_REG_4__SCAN_IN), .C2(n3754), .A(n4422), .B(n3753), 
        .ZN(n3755) );
  NAND3_X1 U4474 ( .A1(n3757), .A2(n3756), .A3(n3755), .ZN(U3244) );
  OAI21_X1 U4475 ( .B1(n4263), .B2(n4538), .A(n3758), .ZN(n3760) );
  MUX2_X1 U4476 ( .A(n4021), .B(REG2_REG_19__SCAN_IN), .S(n3768), .Z(n3759) );
  XNOR2_X1 U4477 ( .A(n3760), .B(n3759), .ZN(n3772) );
  OAI21_X1 U4478 ( .B1(n3762), .B2(n4538), .A(n3761), .ZN(n3765) );
  XNOR2_X1 U4479 ( .A(n3763), .B(REG1_REG_19__SCAN_IN), .ZN(n3764) );
  XNOR2_X1 U4480 ( .A(n3765), .B(n3764), .ZN(n3770) );
  NAND2_X1 U4481 ( .A1(n4435), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3767) );
  OAI211_X1 U4482 ( .C1(n4431), .C2(n3768), .A(n3767), .B(n3766), .ZN(n3769)
         );
  AOI21_X1 U4483 ( .B1(n3770), .B2(n4422), .A(n3769), .ZN(n3771) );
  OAI21_X1 U4484 ( .B1(n3772), .B2(n4440), .A(n3771), .ZN(U3259) );
  INV_X1 U4485 ( .A(n3773), .ZN(n3796) );
  NAND2_X1 U4486 ( .A1(n3775), .A2(n3774), .ZN(n3777) );
  INV_X1 U4487 ( .A(n3780), .ZN(n3781) );
  INV_X1 U4488 ( .A(n3782), .ZN(n3784) );
  OAI21_X1 U4489 ( .B1(n3971), .B2(n3784), .A(n3783), .ZN(n3908) );
  OAI21_X1 U4490 ( .B1(n3850), .B2(n3789), .A(n3788), .ZN(n3790) );
  XOR2_X1 U4491 ( .A(n3822), .B(n3790), .Z(n3795) );
  AOI22_X1 U4492 ( .A1(n3792), .A2(n3791), .B1(n4489), .B2(n3824), .ZN(n3794)
         );
  NAND2_X1 U4493 ( .A1(n3821), .A2(n4460), .ZN(n3793) );
  OAI211_X1 U4494 ( .C1(n3795), .C2(n4462), .A(n3794), .B(n3793), .ZN(n4073)
         );
  AOI21_X1 U4495 ( .B1(n4516), .B2(n3796), .A(n4073), .ZN(n3827) );
  NAND2_X1 U4496 ( .A1(n3804), .A2(n4019), .ZN(n3805) );
  NAND2_X1 U4497 ( .A1(n3990), .A2(n3977), .ZN(n3926) );
  NOR2_X1 U4498 ( .A1(n3990), .A2(n3977), .ZN(n3927) );
  AOI21_X1 U4499 ( .B1(n3925), .B2(n3926), .A(n3927), .ZN(n3809) );
  NOR2_X1 U4500 ( .A1(n3953), .A2(n3808), .ZN(n3811) );
  NAND2_X1 U4501 ( .A1(n3810), .A2(n3963), .ZN(n3928) );
  OAI22_X1 U4502 ( .A1(n3811), .A2(n3928), .B1(n3911), .B2(n3941), .ZN(n3812)
         );
  NAND2_X1 U4503 ( .A1(n3938), .A2(n3813), .ZN(n3815) );
  OAI21_X1 U4504 ( .B1(n3817), .B2(n3894), .A(n3816), .ZN(n3876) );
  OAI21_X1 U4505 ( .B1(n3876), .B2(n2177), .A(n3818), .ZN(n3819) );
  XNOR2_X1 U4506 ( .A(n3823), .B(n3822), .ZN(n4072) );
  NAND2_X1 U4507 ( .A1(n4072), .A2(n3878), .ZN(n3826) );
  AOI21_X1 U4508 ( .B1(n3824), .B2(n3839), .A(n4067), .ZN(n4074) );
  AOI22_X1 U4509 ( .A1(n4074), .A2(n4504), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4521), .ZN(n3825) );
  OAI211_X1 U4510 ( .C1(n4521), .C2(n3827), .A(n3826), .B(n3825), .ZN(U3354)
         );
  INV_X1 U4511 ( .A(n3850), .ZN(n3829) );
  NAND2_X1 U4512 ( .A1(n3829), .A2(n3828), .ZN(n3830) );
  XNOR2_X1 U4513 ( .A(n3830), .B(n3836), .ZN(n3835) );
  AOI22_X1 U4514 ( .A1(n3831), .A2(n4460), .B1(n3841), .B2(n4489), .ZN(n3834)
         );
  NAND2_X1 U4515 ( .A1(n3832), .A2(n4490), .ZN(n3833) );
  OAI211_X1 U4516 ( .C1(n3835), .C2(n4462), .A(n3834), .B(n3833), .ZN(n4077)
         );
  INV_X1 U4517 ( .A(n4077), .ZN(n3847) );
  INV_X1 U4518 ( .A(n3836), .ZN(n3837) );
  XNOR2_X1 U4519 ( .A(n3838), .B(n3837), .ZN(n4078) );
  NAND2_X1 U4520 ( .A1(n4078), .A2(n3878), .ZN(n3846) );
  INV_X1 U4521 ( .A(n3839), .ZN(n3840) );
  AOI21_X1 U4522 ( .B1(n3841), .B2(n3859), .A(n3840), .ZN(n4149) );
  INV_X1 U4523 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3842) );
  OAI22_X1 U4524 ( .A1(n3843), .A2(n4057), .B1(n3842), .B2(n4061), .ZN(n3844)
         );
  AOI21_X1 U4525 ( .B1(n4149), .B2(n4504), .A(n3844), .ZN(n3845) );
  OAI211_X1 U4526 ( .C1(n3847), .C2(n4521), .A(n3846), .B(n3845), .ZN(U3262)
         );
  NOR2_X1 U4527 ( .A1(n3848), .A2(n3857), .ZN(n3849) );
  OR2_X1 U4528 ( .A1(n3850), .A2(n3849), .ZN(n3856) );
  AOI22_X1 U4529 ( .A1(n3852), .A2(n4460), .B1(n3851), .B2(n4489), .ZN(n3853)
         );
  OAI21_X1 U4530 ( .B1(n3854), .B2(n4514), .A(n3853), .ZN(n3855) );
  AOI21_X1 U4531 ( .B1(n3856), .B2(n4511), .A(n3855), .ZN(n4083) );
  XNOR2_X1 U4532 ( .A(n3858), .B(n3857), .ZN(n4082) );
  NAND2_X1 U4533 ( .A1(n4082), .A2(n3878), .ZN(n3866) );
  OAI21_X1 U4534 ( .B1(n3879), .B2(n3860), .A(n3859), .ZN(n4085) );
  INV_X1 U4535 ( .A(n4085), .ZN(n3864) );
  INV_X1 U4536 ( .A(REG2_REG_27__SCAN_IN), .ZN(n3861) );
  OAI22_X1 U4537 ( .A1(n3862), .A2(n4057), .B1(n4519), .B2(n3861), .ZN(n3863)
         );
  AOI21_X1 U4538 ( .B1(n3864), .B2(n4504), .A(n3863), .ZN(n3865) );
  OAI211_X1 U4539 ( .C1(n4083), .C2(n4521), .A(n3866), .B(n3865), .ZN(U3263)
         );
  INV_X1 U4540 ( .A(n3867), .ZN(n3869) );
  OAI21_X1 U4541 ( .B1(n3891), .B2(n3869), .A(n3868), .ZN(n3870) );
  XOR2_X1 U4542 ( .A(n3877), .B(n3870), .Z(n3875) );
  AOI22_X1 U4543 ( .A1(n3913), .A2(n4460), .B1(n3871), .B2(n4489), .ZN(n3872)
         );
  OAI21_X1 U4544 ( .B1(n3873), .B2(n4514), .A(n3872), .ZN(n3874) );
  AOI21_X1 U4545 ( .B1(n3875), .B2(n4511), .A(n3874), .ZN(n4087) );
  XOR2_X1 U4546 ( .A(n3877), .B(n3876), .Z(n4086) );
  NAND2_X1 U4547 ( .A1(n4086), .A2(n3878), .ZN(n3887) );
  INV_X1 U4548 ( .A(n3879), .ZN(n3880) );
  OAI21_X1 U4549 ( .B1(n3900), .B2(n3881), .A(n3880), .ZN(n4089) );
  INV_X1 U4550 ( .A(n4089), .ZN(n3885) );
  OAI22_X1 U4551 ( .A1(n4519), .A2(n3883), .B1(n3882), .B2(n4057), .ZN(n3884)
         );
  AOI21_X1 U4552 ( .B1(n3885), .B2(n4504), .A(n3884), .ZN(n3886) );
  OAI211_X1 U4553 ( .C1(n4521), .C2(n4087), .A(n3887), .B(n3886), .ZN(U3264)
         );
  XOR2_X1 U4554 ( .A(n3892), .B(n3888), .Z(n4091) );
  INV_X1 U4555 ( .A(n4091), .ZN(n3906) );
  INV_X1 U4556 ( .A(n3889), .ZN(n3890) );
  NOR2_X1 U4557 ( .A1(n3891), .A2(n3890), .ZN(n3893) );
  XNOR2_X1 U4558 ( .A(n3893), .B(n3892), .ZN(n3898) );
  OAI22_X1 U4559 ( .A1(n3895), .A2(n4514), .B1(n4456), .B2(n3894), .ZN(n3896)
         );
  AOI21_X1 U4560 ( .B1(n4460), .B2(n3938), .A(n3896), .ZN(n3897) );
  OAI21_X1 U4561 ( .B1(n3898), .B2(n4462), .A(n3897), .ZN(n4090) );
  AND2_X1 U4562 ( .A1(n3916), .A2(n3899), .ZN(n3901) );
  OR2_X1 U4563 ( .A1(n3901), .A2(n3900), .ZN(n4297) );
  AOI22_X1 U4564 ( .A1(n4521), .A2(REG2_REG_25__SCAN_IN), .B1(n3902), .B2(
        n4516), .ZN(n3903) );
  OAI21_X1 U4565 ( .B1(n4297), .B2(n4056), .A(n3903), .ZN(n3904) );
  AOI21_X1 U4566 ( .B1(n4090), .B2(n4519), .A(n3904), .ZN(n3905) );
  OAI21_X1 U4567 ( .B1(n3906), .B2(n4063), .A(n3905), .ZN(U3265) );
  XNOR2_X1 U4568 ( .A(n2032), .B(n3909), .ZN(n4095) );
  INV_X1 U4569 ( .A(n4095), .ZN(n3924) );
  NAND2_X1 U4570 ( .A1(n3908), .A2(n3907), .ZN(n3910) );
  XNOR2_X1 U4571 ( .A(n3910), .B(n3909), .ZN(n3915) );
  OAI22_X1 U4572 ( .A1(n3911), .A2(n4493), .B1(n4456), .B2(n3917), .ZN(n3912)
         );
  AOI21_X1 U4573 ( .B1(n4490), .B2(n3913), .A(n3912), .ZN(n3914) );
  OAI21_X1 U4574 ( .B1(n3915), .B2(n4462), .A(n3914), .ZN(n4094) );
  INV_X1 U4575 ( .A(n3943), .ZN(n3918) );
  OAI21_X1 U4576 ( .B1(n3918), .B2(n3917), .A(n3916), .ZN(n4301) );
  NOR2_X1 U4577 ( .A1(n4301), .A2(n4056), .ZN(n3922) );
  OAI22_X1 U4578 ( .A1(n4519), .A2(n3920), .B1(n3919), .B2(n4057), .ZN(n3921)
         );
  AOI211_X1 U4579 ( .C1(n4094), .C2(n4519), .A(n3922), .B(n3921), .ZN(n3923)
         );
  OAI21_X1 U4580 ( .B1(n3924), .B2(n4063), .A(n3923), .ZN(U3266) );
  OAI21_X1 U4581 ( .B1(n3925), .B2(n3927), .A(n3926), .ZN(n3958) );
  OR2_X1 U4582 ( .A1(n3958), .A2(n3952), .ZN(n3959) );
  NAND2_X1 U4583 ( .A1(n3959), .A2(n3928), .ZN(n3929) );
  XOR2_X1 U4584 ( .A(n3935), .B(n3929), .Z(n4099) );
  INV_X1 U4585 ( .A(n4099), .ZN(n3949) );
  INV_X1 U4586 ( .A(n3930), .ZN(n3931) );
  NAND2_X1 U4587 ( .A1(n3971), .A2(n3931), .ZN(n3933) );
  NAND2_X1 U4588 ( .A1(n3933), .A2(n3932), .ZN(n3951) );
  NAND2_X1 U4589 ( .A1(n3951), .A2(n3952), .ZN(n3950) );
  NAND2_X1 U4590 ( .A1(n3950), .A2(n3934), .ZN(n3936) );
  XNOR2_X1 U4591 ( .A(n3936), .B(n3935), .ZN(n3940) );
  OAI22_X1 U4592 ( .A1(n3972), .A2(n4493), .B1(n4456), .B2(n3941), .ZN(n3937)
         );
  AOI21_X1 U4593 ( .B1(n4490), .B2(n3938), .A(n3937), .ZN(n3939) );
  OAI21_X1 U4594 ( .B1(n3940), .B2(n4462), .A(n3939), .ZN(n4098) );
  OR2_X1 U4595 ( .A1(n3962), .A2(n3941), .ZN(n3942) );
  NAND2_X1 U4596 ( .A1(n3943), .A2(n3942), .ZN(n4305) );
  NOR2_X1 U4597 ( .A1(n4305), .A2(n4056), .ZN(n3947) );
  OAI22_X1 U4598 ( .A1(n4519), .A2(n3945), .B1(n3944), .B2(n4057), .ZN(n3946)
         );
  AOI211_X1 U4599 ( .C1(n4098), .C2(n4519), .A(n3947), .B(n3946), .ZN(n3948)
         );
  OAI21_X1 U4600 ( .B1(n3949), .B2(n4063), .A(n3948), .ZN(U3267) );
  OAI21_X1 U4601 ( .B1(n3952), .B2(n3951), .A(n3950), .ZN(n3957) );
  NAND2_X1 U4602 ( .A1(n3963), .A2(n4489), .ZN(n3955) );
  NAND2_X1 U4603 ( .A1(n3953), .A2(n4490), .ZN(n3954) );
  OAI211_X1 U4604 ( .C1(n3990), .C2(n4493), .A(n3955), .B(n3954), .ZN(n3956)
         );
  AOI21_X1 U4605 ( .B1(n3957), .B2(n4511), .A(n3956), .ZN(n4105) );
  INV_X1 U4606 ( .A(n3958), .ZN(n3961) );
  OAI21_X1 U4607 ( .B1(n3961), .B2(n3960), .A(n3959), .ZN(n4106) );
  OR2_X1 U4608 ( .A1(n4106), .A2(n4063), .ZN(n3969) );
  INV_X1 U4609 ( .A(n3962), .ZN(n4103) );
  NAND2_X1 U4610 ( .A1(n3976), .A2(n3963), .ZN(n4102) );
  AND2_X1 U4611 ( .A1(n4102), .A2(n4504), .ZN(n3967) );
  OAI22_X1 U4612 ( .A1(n4519), .A2(n3965), .B1(n3964), .B2(n4057), .ZN(n3966)
         );
  AOI21_X1 U4613 ( .B1(n4103), .B2(n3967), .A(n3966), .ZN(n3968) );
  OAI211_X1 U4614 ( .C1(n4521), .C2(n4105), .A(n3969), .B(n3968), .ZN(U3268)
         );
  XOR2_X1 U4615 ( .A(n3970), .B(n3925), .Z(n4108) );
  INV_X1 U4616 ( .A(n4108), .ZN(n3983) );
  XNOR2_X1 U4617 ( .A(n3971), .B(n3970), .ZN(n3975) );
  OAI22_X1 U4618 ( .A1(n3972), .A2(n4514), .B1(n4456), .B2(n3977), .ZN(n3973)
         );
  AOI21_X1 U4619 ( .B1(n4460), .B2(n4015), .A(n3973), .ZN(n3974) );
  OAI21_X1 U4620 ( .B1(n3975), .B2(n4462), .A(n3974), .ZN(n4107) );
  OAI21_X1 U4621 ( .B1(n2169), .B2(n3977), .A(n3976), .ZN(n4310) );
  NOR2_X1 U4622 ( .A1(n4310), .A2(n4056), .ZN(n3981) );
  OAI22_X1 U4623 ( .A1(n4061), .A2(n3979), .B1(n3978), .B2(n4057), .ZN(n3980)
         );
  AOI211_X1 U4624 ( .C1(n4107), .C2(n4061), .A(n3981), .B(n3980), .ZN(n3982)
         );
  OAI21_X1 U4625 ( .B1(n3983), .B2(n4063), .A(n3982), .ZN(U3269) );
  XNOR2_X1 U4626 ( .A(n3984), .B(n3988), .ZN(n4112) );
  INV_X1 U4627 ( .A(n4112), .ZN(n4002) );
  INV_X1 U4628 ( .A(n3985), .ZN(n3986) );
  NAND2_X1 U4629 ( .A1(n3987), .A2(n3986), .ZN(n3989) );
  XNOR2_X1 U4630 ( .A(n3989), .B(n3988), .ZN(n3993) );
  OAI22_X1 U4631 ( .A1(n3990), .A2(n4514), .B1(n4456), .B2(n3995), .ZN(n3991)
         );
  AOI21_X1 U4632 ( .B1(n4460), .B2(n4034), .A(n3991), .ZN(n3992) );
  OAI21_X1 U4633 ( .B1(n3993), .B2(n4462), .A(n3992), .ZN(n4111) );
  INV_X1 U4634 ( .A(n4018), .ZN(n3996) );
  OAI21_X1 U4635 ( .B1(n3996), .B2(n3995), .A(n3994), .ZN(n4314) );
  NOR2_X1 U4636 ( .A1(n4314), .A2(n4056), .ZN(n4000) );
  OAI22_X1 U4637 ( .A1(n4519), .A2(n3998), .B1(n3997), .B2(n4057), .ZN(n3999)
         );
  AOI211_X1 U4638 ( .C1(n4111), .C2(n4061), .A(n4000), .B(n3999), .ZN(n4001)
         );
  OAI21_X1 U4639 ( .B1(n4002), .B2(n4063), .A(n4001), .ZN(U3270) );
  XNOR2_X1 U4640 ( .A(n4004), .B(n4003), .ZN(n4116) );
  INV_X1 U4641 ( .A(n4116), .ZN(n4025) );
  INV_X1 U4642 ( .A(n4005), .ZN(n4007) );
  OAI21_X1 U4643 ( .B1(n4045), .B2(n4007), .A(n4006), .ZN(n4031) );
  INV_X1 U4644 ( .A(n4008), .ZN(n4010) );
  OAI21_X1 U4645 ( .B1(n4031), .B2(n4010), .A(n4009), .ZN(n4012) );
  XNOR2_X1 U4646 ( .A(n4012), .B(n4011), .ZN(n4013) );
  NAND2_X1 U4647 ( .A1(n4013), .A2(n4511), .ZN(n4017) );
  AOI22_X1 U4648 ( .A1(n4015), .A2(n4490), .B1(n4489), .B2(n4014), .ZN(n4016)
         );
  OAI211_X1 U4649 ( .C1(n4047), .C2(n4493), .A(n4017), .B(n4016), .ZN(n4115)
         );
  OAI21_X1 U4650 ( .B1(n4027), .B2(n4019), .A(n4018), .ZN(n4318) );
  NOR2_X1 U4651 ( .A1(n4318), .A2(n4056), .ZN(n4023) );
  OAI22_X1 U4652 ( .A1(n4061), .A2(n4021), .B1(n4020), .B2(n4057), .ZN(n4022)
         );
  AOI211_X1 U4653 ( .C1(n4115), .C2(n4061), .A(n4023), .B(n4022), .ZN(n4024)
         );
  OAI21_X1 U4654 ( .B1(n4025), .B2(n4063), .A(n4024), .ZN(U3271) );
  XOR2_X1 U4655 ( .A(n4032), .B(n4026), .Z(n4120) );
  INV_X1 U4656 ( .A(n4027), .ZN(n4028) );
  OAI211_X1 U4657 ( .C1(n4053), .C2(n4029), .A(n4028), .B(n4596), .ZN(n4118)
         );
  INV_X1 U4658 ( .A(n4118), .ZN(n4042) );
  OAI22_X1 U4659 ( .A1(n4061), .A2(n4263), .B1(n4030), .B2(n4057), .ZN(n4040)
         );
  XOR2_X1 U4660 ( .A(n4032), .B(n4031), .Z(n4038) );
  AOI22_X1 U4661 ( .A1(n4034), .A2(n4490), .B1(n4033), .B2(n4489), .ZN(n4035)
         );
  OAI21_X1 U4662 ( .B1(n4036), .B2(n4493), .A(n4035), .ZN(n4037) );
  AOI21_X1 U4663 ( .B1(n4038), .B2(n4511), .A(n4037), .ZN(n4119) );
  NOR2_X1 U4664 ( .A1(n4119), .A2(n4521), .ZN(n4039) );
  AOI211_X1 U4665 ( .C1(n4042), .C2(n4041), .A(n4040), .B(n4039), .ZN(n4043)
         );
  OAI21_X1 U4666 ( .B1(n4063), .B2(n4120), .A(n4043), .ZN(U3272) );
  XNOR2_X1 U4667 ( .A(n4044), .B(n4046), .ZN(n4122) );
  INV_X1 U4668 ( .A(n4122), .ZN(n4064) );
  XOR2_X1 U4669 ( .A(n4046), .B(n4045), .Z(n4051) );
  OAI22_X1 U4670 ( .A1(n4047), .A2(n4514), .B1(n4456), .B2(n4055), .ZN(n4048)
         );
  AOI21_X1 U4671 ( .B1(n4460), .B2(n4049), .A(n4048), .ZN(n4050) );
  OAI21_X1 U4672 ( .B1(n4051), .B2(n4462), .A(n4050), .ZN(n4121) );
  INV_X1 U4673 ( .A(n4053), .ZN(n4054) );
  OAI21_X1 U4674 ( .B1(n2166), .B2(n4055), .A(n4054), .ZN(n4323) );
  NOR2_X1 U4675 ( .A1(n4323), .A2(n4056), .ZN(n4060) );
  OAI22_X1 U4676 ( .A1(n4061), .A2(n2352), .B1(n4058), .B2(n4057), .ZN(n4059)
         );
  AOI211_X1 U4677 ( .C1(n4121), .C2(n4061), .A(n4060), .B(n4059), .ZN(n4062)
         );
  OAI21_X1 U4678 ( .B1(n4064), .B2(n4063), .A(n4062), .ZN(U3273) );
  OAI21_X1 U4679 ( .B1(n4067), .B2(n4066), .A(n4065), .ZN(n4342) );
  INV_X1 U4680 ( .A(n4068), .ZN(n4069) );
  AOI21_X1 U4681 ( .B1(n4070), .B2(n4489), .A(n4069), .ZN(n4345) );
  MUX2_X1 U4682 ( .A(n3612), .B(n4345), .S(n4621), .Z(n4071) );
  OAI21_X1 U4683 ( .B1(n4342), .B2(n4133), .A(n4071), .ZN(U3548) );
  NAND2_X1 U4684 ( .A1(n4072), .A2(n4588), .ZN(n4076) );
  AOI21_X1 U4685 ( .B1(n4078), .B2(n4588), .A(n4077), .ZN(n4146) );
  MUX2_X1 U4686 ( .A(n4254), .B(n4146), .S(n4621), .Z(n4081) );
  NAND2_X1 U4687 ( .A1(n4149), .A2(n4079), .ZN(n4080) );
  NAND2_X1 U4688 ( .A1(n4081), .A2(n4080), .ZN(U3546) );
  NAND2_X1 U4689 ( .A1(n4082), .A2(n4588), .ZN(n4084) );
  OAI211_X1 U4690 ( .C1(n3018), .C2(n4085), .A(n4084), .B(n4083), .ZN(n4152)
         );
  MUX2_X1 U4691 ( .A(REG1_REG_27__SCAN_IN), .B(n4152), .S(n4621), .Z(U3545) );
  NAND2_X1 U4692 ( .A1(n4086), .A2(n4588), .ZN(n4088) );
  OAI211_X1 U4693 ( .C1(n3018), .C2(n4089), .A(n4088), .B(n4087), .ZN(n4153)
         );
  MUX2_X1 U4694 ( .A(REG1_REG_26__SCAN_IN), .B(n4153), .S(n4621), .Z(U3544) );
  INV_X1 U4695 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4092) );
  AOI21_X1 U4696 ( .B1(n4091), .B2(n4588), .A(n4090), .ZN(n4294) );
  MUX2_X1 U4697 ( .A(n4092), .B(n4294), .S(n4621), .Z(n4093) );
  OAI21_X1 U4698 ( .B1(n4133), .B2(n4297), .A(n4093), .ZN(U3543) );
  AOI21_X1 U4699 ( .B1(n4095), .B2(n4588), .A(n4094), .ZN(n4298) );
  MUX2_X1 U4700 ( .A(n4096), .B(n4298), .S(n4621), .Z(n4097) );
  OAI21_X1 U4701 ( .B1(n4133), .B2(n4301), .A(n4097), .ZN(U3542) );
  INV_X1 U4702 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4100) );
  AOI21_X1 U4703 ( .B1(n4099), .B2(n4588), .A(n4098), .ZN(n4302) );
  MUX2_X1 U4704 ( .A(n4100), .B(n4302), .S(n4621), .Z(n4101) );
  OAI21_X1 U4705 ( .B1(n4133), .B2(n4305), .A(n4101), .ZN(U3541) );
  INV_X1 U4706 ( .A(n4588), .ZN(n4591) );
  NAND3_X1 U4707 ( .A1(n4103), .A2(n4596), .A3(n4102), .ZN(n4104) );
  OAI211_X1 U4708 ( .C1(n4106), .C2(n4591), .A(n4105), .B(n4104), .ZN(n4306)
         );
  MUX2_X1 U4709 ( .A(REG1_REG_22__SCAN_IN), .B(n4306), .S(n4621), .Z(U3540) );
  INV_X1 U4710 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4109) );
  AOI21_X1 U4711 ( .B1(n4108), .B2(n4588), .A(n4107), .ZN(n4307) );
  MUX2_X1 U4712 ( .A(n4109), .B(n4307), .S(n4621), .Z(n4110) );
  OAI21_X1 U4713 ( .B1(n4133), .B2(n4310), .A(n4110), .ZN(U3539) );
  AOI21_X1 U4714 ( .B1(n4112), .B2(n4588), .A(n4111), .ZN(n4311) );
  MUX2_X1 U4715 ( .A(n4113), .B(n4311), .S(n4621), .Z(n4114) );
  OAI21_X1 U4716 ( .B1(n4133), .B2(n4314), .A(n4114), .ZN(U3538) );
  AOI21_X1 U4717 ( .B1(n4116), .B2(n4588), .A(n4115), .ZN(n4315) );
  MUX2_X1 U4718 ( .A(n4210), .B(n4315), .S(n4621), .Z(n4117) );
  OAI21_X1 U4719 ( .B1(n4133), .B2(n4318), .A(n4117), .ZN(U3537) );
  OAI211_X1 U4720 ( .C1(n4120), .C2(n4591), .A(n4119), .B(n4118), .ZN(n4319)
         );
  MUX2_X1 U4721 ( .A(REG1_REG_18__SCAN_IN), .B(n4319), .S(n4621), .Z(U3536) );
  AOI21_X1 U4722 ( .B1(n4122), .B2(n4588), .A(n4121), .ZN(n4320) );
  MUX2_X1 U4723 ( .A(n4123), .B(n4320), .S(n4621), .Z(n4124) );
  OAI21_X1 U4724 ( .B1(n4133), .B2(n4323), .A(n4124), .ZN(U3535) );
  AOI21_X1 U4725 ( .B1(n4126), .B2(n4588), .A(n4125), .ZN(n4324) );
  MUX2_X1 U4726 ( .A(n4127), .B(n4324), .S(n4621), .Z(n4128) );
  OAI21_X1 U4727 ( .B1(n4133), .B2(n4327), .A(n4128), .ZN(U3534) );
  AOI21_X1 U4728 ( .B1(n4130), .B2(n4588), .A(n4129), .ZN(n4328) );
  MUX2_X1 U4729 ( .A(n4131), .B(n4328), .S(n4621), .Z(n4132) );
  OAI21_X1 U4730 ( .B1(n4133), .B2(n4332), .A(n4132), .ZN(U3533) );
  INV_X1 U4731 ( .A(n4134), .ZN(n4139) );
  NAND3_X1 U4732 ( .A1(n4136), .A2(n4596), .A3(n4135), .ZN(n4137) );
  OAI211_X1 U4733 ( .C1(n4139), .C2(n4572), .A(n4138), .B(n4137), .ZN(n4333)
         );
  MUX2_X1 U4734 ( .A(REG1_REG_14__SCAN_IN), .B(n4333), .S(n4621), .Z(U3532) );
  AOI21_X1 U4735 ( .B1(n4596), .B2(n4141), .A(n4140), .ZN(n4142) );
  OAI21_X1 U4736 ( .B1(n4591), .B2(n4143), .A(n4142), .ZN(n4334) );
  MUX2_X1 U4737 ( .A(REG1_REG_13__SCAN_IN), .B(n4334), .S(n4621), .Z(U3531) );
  INV_X1 U4738 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4144) );
  MUX2_X1 U4739 ( .A(n4144), .B(n4345), .S(n4606), .Z(n4145) );
  OAI21_X1 U4740 ( .B1(n4342), .B2(n4331), .A(n4145), .ZN(U3516) );
  INV_X1 U4741 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4147) );
  MUX2_X1 U4742 ( .A(n4147), .B(n4146), .S(n4606), .Z(n4151) );
  NAND2_X1 U4743 ( .A1(n4149), .A2(n4148), .ZN(n4150) );
  NAND2_X1 U4744 ( .A1(n4151), .A2(n4150), .ZN(U3514) );
  MUX2_X1 U4745 ( .A(REG0_REG_27__SCAN_IN), .B(n4152), .S(n4606), .Z(U3513) );
  MUX2_X1 U4746 ( .A(REG0_REG_26__SCAN_IN), .B(n4153), .S(n4606), .Z(n4293) );
  INV_X1 U4747 ( .A(keyinput62), .ZN(n4160) );
  NOR2_X1 U4748 ( .A1(keyinput10), .A2(keyinput3), .ZN(n4158) );
  NAND2_X1 U4749 ( .A1(keyinput6), .A2(keyinput26), .ZN(n4156) );
  INV_X1 U4750 ( .A(keyinput31), .ZN(n4154) );
  NAND4_X1 U4751 ( .A1(keyinput18), .A2(keyinput19), .A3(keyinput30), .A4(
        n4154), .ZN(n4155) );
  NOR4_X1 U4752 ( .A1(keyinput15), .A2(keyinput23), .A3(n4156), .A4(n4155), 
        .ZN(n4157) );
  NAND4_X1 U4753 ( .A1(keyinput2), .A2(keyinput11), .A3(n4158), .A4(n4157), 
        .ZN(n4159) );
  NOR4_X1 U4754 ( .A1(keyinput14), .A2(keyinput7), .A3(n4160), .A4(n4159), 
        .ZN(n4175) );
  NAND3_X1 U4755 ( .A1(keyinput1), .A2(keyinput5), .A3(keyinput21), .ZN(n4162)
         );
  NAND3_X1 U4756 ( .A1(keyinput41), .A2(keyinput53), .A3(keyinput49), .ZN(
        n4161) );
  NOR4_X1 U4757 ( .A1(keyinput17), .A2(keyinput45), .A3(n4162), .A4(n4161), 
        .ZN(n4174) );
  NAND2_X1 U4758 ( .A1(keyinput22), .A2(keyinput9), .ZN(n4164) );
  NAND4_X1 U4759 ( .A1(keyinput25), .A2(keyinput29), .A3(keyinput33), .A4(
        keyinput37), .ZN(n4163) );
  NOR4_X1 U4760 ( .A1(keyinput27), .A2(keyinput13), .A3(n4164), .A4(n4163), 
        .ZN(n4173) );
  NAND2_X1 U4761 ( .A1(keyinput32), .A2(keyinput0), .ZN(n4171) );
  NOR2_X1 U4762 ( .A1(keyinput54), .A2(keyinput35), .ZN(n4169) );
  NAND2_X1 U4763 ( .A1(keyinput46), .A2(keyinput59), .ZN(n4167) );
  INV_X1 U4764 ( .A(keyinput58), .ZN(n4165) );
  NAND4_X1 U4765 ( .A1(keyinput34), .A2(keyinput42), .A3(keyinput51), .A4(
        n4165), .ZN(n4166) );
  NOR4_X1 U4766 ( .A1(keyinput50), .A2(keyinput63), .A3(n4167), .A4(n4166), 
        .ZN(n4168) );
  NAND4_X1 U4767 ( .A1(keyinput47), .A2(keyinput38), .A3(n4169), .A4(n4168), 
        .ZN(n4170) );
  NOR4_X1 U4768 ( .A1(keyinput55), .A2(keyinput39), .A3(n4171), .A4(n4170), 
        .ZN(n4172) );
  NAND4_X1 U4769 ( .A1(n4175), .A2(n4174), .A3(n4173), .A4(n4172), .ZN(n4183)
         );
  NAND3_X1 U4770 ( .A1(keyinput12), .A2(keyinput61), .A3(keyinput57), .ZN(
        n4176) );
  NOR2_X1 U4771 ( .A1(keyinput4), .A2(n4176), .ZN(n4181) );
  NOR3_X1 U4772 ( .A1(keyinput20), .A2(keyinput28), .A3(keyinput24), .ZN(n4180) );
  NAND3_X1 U4773 ( .A1(keyinput36), .A2(keyinput16), .A3(keyinput40), .ZN(
        n4178) );
  NAND3_X1 U4774 ( .A1(keyinput52), .A2(keyinput60), .A3(keyinput48), .ZN(
        n4177) );
  NOR4_X1 U4775 ( .A1(keyinput44), .A2(keyinput56), .A3(n4178), .A4(n4177), 
        .ZN(n4179) );
  NAND4_X1 U4776 ( .A1(n4181), .A2(keyinput8), .A3(n4180), .A4(n4179), .ZN(
        n4182) );
  OAI21_X1 U4777 ( .B1(n4183), .B2(n4182), .A(keyinput43), .ZN(n4184) );
  NAND2_X1 U4778 ( .A1(n4184), .A2(REG2_REG_31__SCAN_IN), .ZN(n4291) );
  INV_X1 U4779 ( .A(keyinput39), .ZN(n4186) );
  AOI22_X1 U4780 ( .A1(n4187), .A2(keyinput54), .B1(DATAO_REG_7__SCAN_IN), 
        .B2(n4186), .ZN(n4185) );
  OAI221_X1 U4781 ( .B1(n4187), .B2(keyinput54), .C1(n4186), .C2(
        DATAO_REG_7__SCAN_IN), .A(n4185), .ZN(n4196) );
  INV_X1 U4782 ( .A(IR_REG_26__SCAN_IN), .ZN(n4189) );
  AOI22_X1 U4783 ( .A1(n4189), .A2(keyinput0), .B1(keyinput55), .B2(n3842), 
        .ZN(n4188) );
  OAI221_X1 U4784 ( .B1(n4189), .B2(keyinput0), .C1(n3842), .C2(keyinput55), 
        .A(n4188), .ZN(n4195) );
  AOI22_X1 U4785 ( .A1(n4308), .A2(keyinput38), .B1(n4316), .B2(keyinput46), 
        .ZN(n4190) );
  OAI221_X1 U4786 ( .B1(n4308), .B2(keyinput38), .C1(n4316), .C2(keyinput46), 
        .A(n4190), .ZN(n4194) );
  AOI22_X1 U4787 ( .A1(n2396), .A2(keyinput47), .B1(keyinput35), .B2(n4192), 
        .ZN(n4191) );
  OAI221_X1 U4788 ( .B1(n2396), .B2(keyinput47), .C1(n4192), .C2(keyinput35), 
        .A(n4191), .ZN(n4193) );
  NOR4_X1 U4789 ( .A1(n4196), .A2(n4195), .A3(n4194), .A4(n4193), .ZN(n4290)
         );
  INV_X1 U4790 ( .A(D_REG_23__SCAN_IN), .ZN(n4523) );
  INV_X1 U4791 ( .A(keyinput4), .ZN(n4198) );
  AOI22_X1 U4792 ( .A1(n4523), .A2(keyinput20), .B1(DATAO_REG_29__SCAN_IN), 
        .B2(n4198), .ZN(n4197) );
  OAI221_X1 U4793 ( .B1(n4523), .B2(keyinput20), .C1(n4198), .C2(
        DATAO_REG_29__SCAN_IN), .A(n4197), .ZN(n4208) );
  INV_X1 U4794 ( .A(D_REG_10__SCAN_IN), .ZN(n4529) );
  INV_X1 U4795 ( .A(keyinput12), .ZN(n4200) );
  AOI22_X1 U4796 ( .A1(n4529), .A2(keyinput57), .B1(DATAO_REG_25__SCAN_IN), 
        .B2(n4200), .ZN(n4199) );
  OAI221_X1 U4797 ( .B1(n4529), .B2(keyinput57), .C1(n4200), .C2(
        DATAO_REG_25__SCAN_IN), .A(n4199), .ZN(n4207) );
  AOI22_X1 U4798 ( .A1(n2491), .A2(keyinput24), .B1(n4202), .B2(keyinput36), 
        .ZN(n4201) );
  OAI221_X1 U4799 ( .B1(n2491), .B2(keyinput24), .C1(n4202), .C2(keyinput36), 
        .A(n4201), .ZN(n4206) );
  INV_X1 U4800 ( .A(DATAI_2_), .ZN(n4204) );
  AOI22_X1 U4801 ( .A1(n4204), .A2(keyinput8), .B1(keyinput28), .B2(n4610), 
        .ZN(n4203) );
  OAI221_X1 U4802 ( .B1(n4204), .B2(keyinput8), .C1(n4610), .C2(keyinput28), 
        .A(n4203), .ZN(n4205) );
  NOR4_X1 U4803 ( .A1(n4208), .A2(n4207), .A3(n4206), .A4(n4205), .ZN(n4289)
         );
  AOI22_X1 U4804 ( .A1(n4524), .A2(keyinput27), .B1(keyinput9), .B2(n4210), 
        .ZN(n4209) );
  OAI221_X1 U4805 ( .B1(n4524), .B2(keyinput27), .C1(n4210), .C2(keyinput9), 
        .A(n4209), .ZN(n4218) );
  AOI22_X1 U4806 ( .A1(n4212), .A2(keyinput13), .B1(keyinput1), .B2(n2619), 
        .ZN(n4211) );
  OAI221_X1 U4807 ( .B1(n4212), .B2(keyinput13), .C1(n2619), .C2(keyinput1), 
        .A(n4211), .ZN(n4217) );
  AOI22_X1 U4808 ( .A1(n3883), .A2(keyinput5), .B1(keyinput17), .B2(n3945), 
        .ZN(n4213) );
  OAI221_X1 U4809 ( .B1(n3883), .B2(keyinput5), .C1(n3945), .C2(keyinput17), 
        .A(n4213), .ZN(n4216) );
  INV_X1 U4810 ( .A(D_REG_18__SCAN_IN), .ZN(n4526) );
  INV_X1 U4811 ( .A(DATAI_12_), .ZN(n4546) );
  AOI22_X1 U4812 ( .A1(n4526), .A2(keyinput21), .B1(keyinput25), .B2(n4546), 
        .ZN(n4214) );
  OAI221_X1 U4813 ( .B1(n4526), .B2(keyinput21), .C1(n4546), .C2(keyinput25), 
        .A(n4214), .ZN(n4215) );
  NOR4_X1 U4814 ( .A1(n4218), .A2(n4217), .A3(n4216), .A4(n4215), .ZN(n4231)
         );
  AOI22_X1 U4815 ( .A1(n4531), .A2(keyinput6), .B1(keyinput26), .B2(n4386), 
        .ZN(n4219) );
  OAI221_X1 U4816 ( .B1(n4531), .B2(keyinput6), .C1(n4386), .C2(keyinput26), 
        .A(n4219), .ZN(n4229) );
  INV_X1 U4817 ( .A(keyinput19), .ZN(n4221) );
  AOI22_X1 U4818 ( .A1(n2412), .A2(keyinput23), .B1(DATAO_REG_17__SCAN_IN), 
        .B2(n4221), .ZN(n4220) );
  OAI221_X1 U4819 ( .B1(n2412), .B2(keyinput23), .C1(n4221), .C2(
        DATAO_REG_17__SCAN_IN), .A(n4220), .ZN(n4228) );
  INV_X1 U4820 ( .A(keyinput18), .ZN(n4223) );
  AOI22_X1 U4821 ( .A1(n3612), .A2(keyinput31), .B1(DATAO_REG_21__SCAN_IN), 
        .B2(n4223), .ZN(n4222) );
  OAI221_X1 U4822 ( .B1(n3612), .B2(keyinput31), .C1(n4223), .C2(
        DATAO_REG_21__SCAN_IN), .A(n4222), .ZN(n4227) );
  INV_X1 U4823 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4225) );
  AOI22_X1 U4824 ( .A1(n4225), .A2(keyinput30), .B1(n4528), .B2(keyinput22), 
        .ZN(n4224) );
  OAI221_X1 U4825 ( .B1(n4225), .B2(keyinput30), .C1(n4528), .C2(keyinput22), 
        .A(n4224), .ZN(n4226) );
  NOR4_X1 U4826 ( .A1(n4229), .A2(n4228), .A3(n4227), .A4(n4226), .ZN(n4230)
         );
  NAND2_X1 U4827 ( .A1(n4231), .A2(n4230), .ZN(n4287) );
  AOI22_X1 U4828 ( .A1(keyinput43), .A2(n3350), .B1(keyinput14), .B2(n4233), 
        .ZN(n4232) );
  OAI21_X1 U4829 ( .B1(keyinput14), .B2(n4233), .A(n4232), .ZN(n4244) );
  INV_X1 U4830 ( .A(keyinput7), .ZN(n4236) );
  INV_X1 U4831 ( .A(keyinput2), .ZN(n4235) );
  AOI22_X1 U4832 ( .A1(n4236), .A2(ADDR_REG_1__SCAN_IN), .B1(
        ADDR_REG_4__SCAN_IN), .B2(n4235), .ZN(n4234) );
  OAI221_X1 U4833 ( .B1(n4236), .B2(ADDR_REG_1__SCAN_IN), .C1(n4235), .C2(
        ADDR_REG_4__SCAN_IN), .A(n4234), .ZN(n4243) );
  INV_X1 U4834 ( .A(keyinput10), .ZN(n4238) );
  AOI22_X1 U4835 ( .A1(n4376), .A2(keyinput11), .B1(ADDR_REG_16__SCAN_IN), 
        .B2(n4238), .ZN(n4237) );
  OAI221_X1 U4836 ( .B1(n4376), .B2(keyinput11), .C1(n4238), .C2(
        ADDR_REG_16__SCAN_IN), .A(n4237), .ZN(n4242) );
  INV_X1 U4837 ( .A(REG0_REG_29__SCAN_IN), .ZN(n4240) );
  AOI22_X1 U4838 ( .A1(n4240), .A2(keyinput3), .B1(n4525), .B2(keyinput15), 
        .ZN(n4239) );
  OAI221_X1 U4839 ( .B1(n4240), .B2(keyinput3), .C1(n4525), .C2(keyinput15), 
        .A(n4239), .ZN(n4241) );
  NOR4_X1 U4840 ( .A1(n4244), .A2(n4243), .A3(n4242), .A4(n4241), .ZN(n4285)
         );
  INV_X1 U4841 ( .A(D_REG_29__SCAN_IN), .ZN(n4522) );
  INV_X1 U4842 ( .A(keyinput44), .ZN(n4246) );
  AOI22_X1 U4843 ( .A1(n4522), .A2(keyinput16), .B1(DATAO_REG_22__SCAN_IN), 
        .B2(n4246), .ZN(n4245) );
  OAI221_X1 U4844 ( .B1(n4522), .B2(keyinput16), .C1(n4246), .C2(
        DATAO_REG_22__SCAN_IN), .A(n4245), .ZN(n4250) );
  INV_X1 U4845 ( .A(keyinput37), .ZN(n4248) );
  AOI22_X1 U4846 ( .A1(n2422), .A2(keyinput41), .B1(DATAO_REG_3__SCAN_IN), 
        .B2(n4248), .ZN(n4247) );
  OAI221_X1 U4847 ( .B1(n2422), .B2(keyinput41), .C1(n4248), .C2(
        DATAO_REG_3__SCAN_IN), .A(n4247), .ZN(n4249) );
  NOR2_X1 U4848 ( .A1(n4250), .A2(n4249), .ZN(n4284) );
  INV_X1 U4849 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4590) );
  AOI22_X1 U4850 ( .A1(n4590), .A2(keyinput49), .B1(n4252), .B2(keyinput61), 
        .ZN(n4251) );
  OAI221_X1 U4851 ( .B1(n4590), .B2(keyinput49), .C1(n4252), .C2(keyinput61), 
        .A(n4251), .ZN(n4259) );
  AOI22_X1 U4852 ( .A1(n4303), .A2(keyinput40), .B1(n4254), .B2(keyinput52), 
        .ZN(n4253) );
  OAI221_X1 U4853 ( .B1(n4303), .B2(keyinput40), .C1(n4254), .C2(keyinput52), 
        .A(n4253), .ZN(n4258) );
  XNOR2_X1 U4854 ( .A(keyinput56), .B(REG1_REG_6__SCAN_IN), .ZN(n4256) );
  XNOR2_X1 U4855 ( .A(keyinput53), .B(REG1_REG_7__SCAN_IN), .ZN(n4255) );
  NAND2_X1 U4856 ( .A1(n4256), .A2(n4255), .ZN(n4257) );
  NOR3_X1 U4857 ( .A1(n4259), .A2(n4258), .A3(n4257), .ZN(n4283) );
  INV_X1 U4858 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4597) );
  AOI22_X1 U4859 ( .A1(n4261), .A2(keyinput50), .B1(keyinput63), .B2(n4597), 
        .ZN(n4260) );
  OAI221_X1 U4860 ( .B1(n4261), .B2(keyinput50), .C1(n4597), .C2(keyinput63), 
        .A(n4260), .ZN(n4265) );
  AOI22_X1 U4861 ( .A1(n2411), .A2(keyinput29), .B1(n4263), .B2(keyinput33), 
        .ZN(n4262) );
  OAI221_X1 U4862 ( .B1(n2411), .B2(keyinput29), .C1(n4263), .C2(keyinput33), 
        .A(n4262), .ZN(n4264) );
  NOR2_X1 U4863 ( .A1(n4265), .A2(n4264), .ZN(n4281) );
  INV_X1 U4864 ( .A(D_REG_17__SCAN_IN), .ZN(n4527) );
  AOI22_X1 U4865 ( .A1(n4295), .A2(keyinput58), .B1(n4527), .B2(keyinput42), 
        .ZN(n4266) );
  OAI221_X1 U4866 ( .B1(n4295), .B2(keyinput58), .C1(n4527), .C2(keyinput42), 
        .A(n4266), .ZN(n4269) );
  INV_X1 U4867 ( .A(D_REG_2__SCAN_IN), .ZN(n4533) );
  INV_X1 U4868 ( .A(D_REG_3__SCAN_IN), .ZN(n4532) );
  AOI22_X1 U4869 ( .A1(n4533), .A2(keyinput62), .B1(n4532), .B2(keyinput51), 
        .ZN(n4267) );
  OAI221_X1 U4870 ( .B1(n4533), .B2(keyinput62), .C1(n4532), .C2(keyinput51), 
        .A(n4267), .ZN(n4268) );
  NOR2_X1 U4871 ( .A1(n4269), .A2(n4268), .ZN(n4280) );
  INV_X1 U4872 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4272) );
  AOI22_X1 U4873 ( .A1(n4272), .A2(keyinput48), .B1(keyinput32), .B2(n4271), 
        .ZN(n4270) );
  OAI221_X1 U4874 ( .B1(n4272), .B2(keyinput48), .C1(n4271), .C2(keyinput32), 
        .A(n4270), .ZN(n4278) );
  XNOR2_X1 U4875 ( .A(IR_REG_25__SCAN_IN), .B(keyinput45), .ZN(n4276) );
  XNOR2_X1 U4876 ( .A(IR_REG_1__SCAN_IN), .B(keyinput59), .ZN(n4275) );
  XNOR2_X1 U4877 ( .A(DATAI_23_), .B(keyinput34), .ZN(n4274) );
  XNOR2_X1 U4878 ( .A(IR_REG_17__SCAN_IN), .B(keyinput60), .ZN(n4273) );
  NAND4_X1 U4879 ( .A1(n4276), .A2(n4275), .A3(n4274), .A4(n4273), .ZN(n4277)
         );
  NOR2_X1 U4880 ( .A1(n4278), .A2(n4277), .ZN(n4279) );
  AND3_X1 U4881 ( .A1(n4281), .A2(n4280), .A3(n4279), .ZN(n4282) );
  NAND4_X1 U4882 ( .A1(n4285), .A2(n4284), .A3(n4283), .A4(n4282), .ZN(n4286)
         );
  NOR2_X1 U4883 ( .A1(n4287), .A2(n4286), .ZN(n4288) );
  NAND4_X1 U4884 ( .A1(n4291), .A2(n4290), .A3(n4289), .A4(n4288), .ZN(n4292)
         );
  XNOR2_X1 U4885 ( .A(n4293), .B(n4292), .ZN(U3512) );
  MUX2_X1 U4886 ( .A(n4295), .B(n4294), .S(n4606), .Z(n4296) );
  OAI21_X1 U4887 ( .B1(n4297), .B2(n4331), .A(n4296), .ZN(U3511) );
  INV_X1 U4888 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4299) );
  MUX2_X1 U4889 ( .A(n4299), .B(n4298), .S(n4606), .Z(n4300) );
  OAI21_X1 U4890 ( .B1(n4301), .B2(n4331), .A(n4300), .ZN(U3510) );
  MUX2_X1 U4891 ( .A(n4303), .B(n4302), .S(n4606), .Z(n4304) );
  OAI21_X1 U4892 ( .B1(n4305), .B2(n4331), .A(n4304), .ZN(U3509) );
  MUX2_X1 U4893 ( .A(REG0_REG_22__SCAN_IN), .B(n4306), .S(n4606), .Z(U3508) );
  MUX2_X1 U4894 ( .A(n4308), .B(n4307), .S(n4606), .Z(n4309) );
  OAI21_X1 U4895 ( .B1(n4310), .B2(n4331), .A(n4309), .ZN(U3507) );
  INV_X1 U4896 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4312) );
  MUX2_X1 U4897 ( .A(n4312), .B(n4311), .S(n4606), .Z(n4313) );
  OAI21_X1 U4898 ( .B1(n4314), .B2(n4331), .A(n4313), .ZN(U3506) );
  MUX2_X1 U4899 ( .A(n4316), .B(n4315), .S(n4606), .Z(n4317) );
  OAI21_X1 U4900 ( .B1(n4318), .B2(n4331), .A(n4317), .ZN(U3505) );
  MUX2_X1 U4901 ( .A(REG0_REG_18__SCAN_IN), .B(n4319), .S(n4606), .Z(U3503) );
  INV_X1 U4902 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4321) );
  MUX2_X1 U4903 ( .A(n4321), .B(n4320), .S(n4606), .Z(n4322) );
  OAI21_X1 U4904 ( .B1(n4323), .B2(n4331), .A(n4322), .ZN(U3501) );
  INV_X1 U4905 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4325) );
  MUX2_X1 U4906 ( .A(n4325), .B(n4324), .S(n4606), .Z(n4326) );
  OAI21_X1 U4907 ( .B1(n4327), .B2(n4331), .A(n4326), .ZN(U3499) );
  INV_X1 U4908 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4329) );
  MUX2_X1 U4909 ( .A(n4329), .B(n4328), .S(n4606), .Z(n4330) );
  OAI21_X1 U4910 ( .B1(n4332), .B2(n4331), .A(n4330), .ZN(U3497) );
  MUX2_X1 U4911 ( .A(REG0_REG_14__SCAN_IN), .B(n4333), .S(n4606), .Z(U3495) );
  MUX2_X1 U4912 ( .A(REG0_REG_13__SCAN_IN), .B(n4334), .S(n4606), .Z(U3493) );
  MUX2_X1 U4913 ( .A(DATAI_30_), .B(n4335), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4914 ( .A(DATAI_29_), .B(n4336), .S(STATE_REG_SCAN_IN), .Z(U3323)
         );
  MUX2_X1 U4915 ( .A(n4337), .B(DATAI_13_), .S(U3149), .Z(U3339) );
  MUX2_X1 U4916 ( .A(n4338), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U4917 ( .A(n2188), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4918 ( .A(n4339), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U4919 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(STATE_REG_SCAN_IN), 
        .Z(U3352) );
  INV_X1 U4920 ( .A(DATAI_28_), .ZN(n4340) );
  AOI22_X1 U4921 ( .A1(STATE_REG_SCAN_IN), .A2(n4341), .B1(n4340), .B2(U3149), 
        .ZN(U3324) );
  INV_X1 U4922 ( .A(n4342), .ZN(n4343) );
  OAI21_X1 U4923 ( .B1(n4521), .B2(n4345), .A(n4344), .ZN(U3261) );
  INV_X1 U4924 ( .A(n4346), .ZN(n4347) );
  OAI21_X1 U4925 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4348), .A(n4347), .ZN(n4349)
         );
  XOR2_X1 U4926 ( .A(n4349), .B(IR_REG_0__SCAN_IN), .Z(n4352) );
  AOI22_X1 U4927 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4435), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4350) );
  OAI21_X1 U4928 ( .B1(n4352), .B2(n4351), .A(n4350), .ZN(U3240) );
  AOI211_X1 U4929 ( .C1(n4355), .C2(n4354), .A(n4353), .B(n4440), .ZN(n4357)
         );
  AOI211_X1 U4930 ( .C1(n4435), .C2(ADDR_REG_6__SCAN_IN), .A(n4357), .B(n4356), 
        .ZN(n4363) );
  AOI21_X1 U4931 ( .B1(n4360), .B2(n4359), .A(n4358), .ZN(n4361) );
  NAND2_X1 U4932 ( .A1(n4422), .A2(n4361), .ZN(n4362) );
  OAI211_X1 U4933 ( .C1(n4431), .C2(n4556), .A(n4363), .B(n4362), .ZN(U3246)
         );
  AOI211_X1 U4934 ( .C1(n4365), .C2(n4364), .A(n2047), .B(n4440), .ZN(n4367)
         );
  AOI211_X1 U4935 ( .C1(n4435), .C2(ADDR_REG_7__SCAN_IN), .A(n4367), .B(n4366), 
        .ZN(n4373) );
  AOI22_X1 U4936 ( .A1(n4368), .A2(n2490), .B1(REG1_REG_7__SCAN_IN), .B2(n4554), .ZN(n4370) );
  AOI21_X1 U4937 ( .B1(n4371), .B2(n4370), .A(n4442), .ZN(n4369) );
  OAI21_X1 U4938 ( .B1(n4371), .B2(n4370), .A(n4369), .ZN(n4372) );
  OAI211_X1 U4939 ( .C1(n4431), .C2(n4554), .A(n4373), .B(n4372), .ZN(U3247)
         );
  AOI211_X1 U4940 ( .C1(n4376), .C2(n4375), .A(n4374), .B(n4440), .ZN(n4379)
         );
  INV_X1 U4941 ( .A(n4377), .ZN(n4378) );
  AOI211_X1 U4942 ( .C1(n4435), .C2(ADDR_REG_8__SCAN_IN), .A(n4379), .B(n4378), 
        .ZN(n4383) );
  OAI211_X1 U4943 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4381), .A(n4422), .B(n4380), 
        .ZN(n4382) );
  OAI211_X1 U4944 ( .C1(n4431), .C2(n4552), .A(n4383), .B(n4382), .ZN(U3248)
         );
  AOI211_X1 U4945 ( .C1(n4386), .C2(n4385), .A(n4384), .B(n4440), .ZN(n4388)
         );
  AOI211_X1 U4946 ( .C1(n4435), .C2(ADDR_REG_10__SCAN_IN), .A(n4388), .B(n4387), .ZN(n4392) );
  OAI211_X1 U4947 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4390), .A(n4422), .B(n4389), .ZN(n4391) );
  OAI211_X1 U4948 ( .C1(n4431), .C2(n2095), .A(n4392), .B(n4391), .ZN(U3250)
         );
  AOI211_X1 U4949 ( .C1(n2048), .C2(n4394), .A(n4393), .B(n4440), .ZN(n4397)
         );
  INV_X1 U4950 ( .A(n4395), .ZN(n4396) );
  AOI211_X1 U4951 ( .C1(n4435), .C2(ADDR_REG_11__SCAN_IN), .A(n4397), .B(n4396), .ZN(n4402) );
  OAI211_X1 U4952 ( .C1(n4400), .C2(n4399), .A(n4422), .B(n4398), .ZN(n4401)
         );
  OAI211_X1 U4953 ( .C1(n4431), .C2(n4549), .A(n4402), .B(n4401), .ZN(U3251)
         );
  AOI211_X1 U4954 ( .C1(n4405), .C2(n4404), .A(n4403), .B(n4440), .ZN(n4407)
         );
  AOI211_X1 U4955 ( .C1(n4435), .C2(ADDR_REG_12__SCAN_IN), .A(n4407), .B(n4406), .ZN(n4411) );
  OAI211_X1 U4956 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4409), .A(n4422), .B(n4408), .ZN(n4410) );
  OAI211_X1 U4957 ( .C1(n4431), .C2(n4547), .A(n4411), .B(n4410), .ZN(U3252)
         );
  OAI211_X1 U4958 ( .C1(REG2_REG_14__SCAN_IN), .C2(n4413), .A(n4426), .B(n4412), .ZN(n4414) );
  NAND2_X1 U4959 ( .A1(n4415), .A2(n4414), .ZN(n4416) );
  AOI21_X1 U4960 ( .B1(n4435), .B2(ADDR_REG_14__SCAN_IN), .A(n4416), .ZN(n4420) );
  OAI211_X1 U4961 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4418), .A(n4422), .B(n4417), .ZN(n4419) );
  OAI211_X1 U4962 ( .C1(n4431), .C2(n2257), .A(n4420), .B(n4419), .ZN(U3254)
         );
  OAI211_X1 U4963 ( .C1(n4424), .C2(n4423), .A(n4422), .B(n4421), .ZN(n4430)
         );
  OAI211_X1 U4964 ( .C1(n4428), .C2(n4427), .A(n4426), .B(n4425), .ZN(n4429)
         );
  OAI211_X1 U4965 ( .C1(n4431), .C2(n4544), .A(n4430), .B(n4429), .ZN(n4432)
         );
  AOI211_X1 U4966 ( .C1(n4435), .C2(ADDR_REG_15__SCAN_IN), .A(n4433), .B(n4432), .ZN(n4434) );
  INV_X1 U4967 ( .A(n4434), .ZN(U3255) );
  INV_X1 U4968 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n4448) );
  INV_X1 U4969 ( .A(n4435), .ZN(n4447) );
  AOI21_X1 U4970 ( .B1(REG1_REG_16__SCAN_IN), .B2(n4437), .A(n4436), .ZN(n4443) );
  AOI21_X1 U4971 ( .B1(REG2_REG_16__SCAN_IN), .B2(n4439), .A(n4438), .ZN(n4441) );
  OAI22_X1 U4972 ( .A1(n4443), .A2(n4442), .B1(n4441), .B2(n4440), .ZN(n4444)
         );
  AOI21_X1 U4973 ( .B1(n4541), .B2(n2349), .A(n4444), .ZN(n4446) );
  OAI211_X1 U4974 ( .C1(n4448), .C2(n4447), .A(n4446), .B(n4445), .ZN(U3256)
         );
  OR2_X1 U4975 ( .A1(n4450), .A2(n4449), .ZN(n4452) );
  NAND2_X1 U4976 ( .A1(n4452), .A2(n4451), .ZN(n4453) );
  XNOR2_X1 U4977 ( .A(n4453), .B(n4454), .ZN(n4602) );
  XNOR2_X1 U4978 ( .A(n4455), .B(n4454), .ZN(n4463) );
  OAI22_X1 U4979 ( .A1(n4457), .A2(n4514), .B1(n4456), .B2(n4467), .ZN(n4458)
         );
  AOI21_X1 U4980 ( .B1(n4460), .B2(n4459), .A(n4458), .ZN(n4461) );
  OAI21_X1 U4981 ( .B1(n4463), .B2(n4462), .A(n4461), .ZN(n4464) );
  AOI21_X1 U4982 ( .B1(n4512), .B2(n4602), .A(n4464), .ZN(n4599) );
  AOI22_X1 U4983 ( .A1(n4465), .A2(n4516), .B1(REG2_REG_11__SCAN_IN), .B2(
        n4521), .ZN(n4471) );
  OAI21_X1 U4984 ( .B1(n4468), .B2(n4467), .A(n4466), .ZN(n4598) );
  INV_X1 U4985 ( .A(n4598), .ZN(n4469) );
  AOI22_X1 U4986 ( .A1(n4602), .A2(n4517), .B1(n4504), .B2(n4469), .ZN(n4470)
         );
  OAI211_X1 U4987 ( .C1(n4521), .C2(n4599), .A(n4471), .B(n4470), .ZN(U3279)
         );
  AOI22_X1 U4988 ( .A1(n4472), .A2(n4516), .B1(REG2_REG_10__SCAN_IN), .B2(
        n4521), .ZN(n4477) );
  INV_X1 U4989 ( .A(n4473), .ZN(n4474) );
  AOI22_X1 U4990 ( .A1(n4475), .A2(n4517), .B1(n4504), .B2(n4474), .ZN(n4476)
         );
  OAI211_X1 U4991 ( .C1(n4521), .C2(n4478), .A(n4477), .B(n4476), .ZN(U3280)
         );
  AOI22_X1 U4992 ( .A1(n4479), .A2(n4516), .B1(REG2_REG_8__SCAN_IN), .B2(n4521), .ZN(n4484) );
  INV_X1 U4993 ( .A(n4480), .ZN(n4481) );
  AOI22_X1 U4994 ( .A1(n4482), .A2(n4517), .B1(n4504), .B2(n4481), .ZN(n4483)
         );
  OAI211_X1 U4995 ( .C1(n4521), .C2(n4485), .A(n4484), .B(n4483), .ZN(U3282)
         );
  INV_X1 U4996 ( .A(n2998), .ZN(n4488) );
  OAI21_X1 U4997 ( .B1(n4488), .B2(n4487), .A(n4486), .ZN(n4500) );
  AOI22_X1 U4998 ( .A1(n4491), .A2(n4490), .B1(n4489), .B2(n2987), .ZN(n4492)
         );
  OAI21_X1 U4999 ( .B1(n4494), .B2(n4493), .A(n4492), .ZN(n4499) );
  OAI21_X1 U5000 ( .B1(n2998), .B2(n4496), .A(n4495), .ZN(n4562) );
  NOR2_X1 U5001 ( .A1(n4562), .A2(n4497), .ZN(n4498) );
  AOI211_X1 U5002 ( .C1(n4511), .C2(n4500), .A(n4499), .B(n4498), .ZN(n4560)
         );
  AOI22_X1 U5003 ( .A1(REG3_REG_1__SCAN_IN), .A2(n4516), .B1(
        REG2_REG_1__SCAN_IN), .B2(n4521), .ZN(n4507) );
  INV_X1 U5004 ( .A(n4562), .ZN(n4505) );
  OAI21_X1 U5005 ( .B1(n4502), .B2(n4509), .A(n4501), .ZN(n4561) );
  INV_X1 U5006 ( .A(n4561), .ZN(n4503) );
  AOI22_X1 U5007 ( .A1(n4505), .A2(n4517), .B1(n4504), .B2(n4503), .ZN(n4506)
         );
  OAI211_X1 U5008 ( .C1(n4521), .C2(n4560), .A(n4507), .B(n4506), .ZN(U3289)
         );
  NOR2_X1 U5009 ( .A1(n4509), .A2(n2392), .ZN(n4558) );
  INV_X1 U5010 ( .A(n4510), .ZN(n4515) );
  OAI21_X1 U5011 ( .B1(n4512), .B2(n4511), .A(n4559), .ZN(n4513) );
  OAI21_X1 U5012 ( .B1(n2988), .B2(n4514), .A(n4513), .ZN(n4557) );
  AOI21_X1 U5013 ( .B1(n4558), .B2(n4515), .A(n4557), .ZN(n4520) );
  AOI22_X1 U5014 ( .A1(n4559), .A2(n4517), .B1(REG3_REG_0__SCAN_IN), .B2(n4516), .ZN(n4518) );
  OAI221_X1 U5015 ( .B1(n4521), .B2(n4520), .C1(n4519), .C2(n2421), .A(n4518), 
        .ZN(U3290) );
  AND2_X1 U5016 ( .A1(D_REG_31__SCAN_IN), .A2(n4530), .ZN(U3291) );
  AND2_X1 U5017 ( .A1(D_REG_30__SCAN_IN), .A2(n4530), .ZN(U3292) );
  NOR2_X1 U5018 ( .A1(n4534), .A2(n4522), .ZN(U3293) );
  AND2_X1 U5019 ( .A1(D_REG_28__SCAN_IN), .A2(n4530), .ZN(U3294) );
  AND2_X1 U5020 ( .A1(D_REG_27__SCAN_IN), .A2(n4530), .ZN(U3295) );
  AND2_X1 U5021 ( .A1(D_REG_26__SCAN_IN), .A2(n4530), .ZN(U3296) );
  AND2_X1 U5022 ( .A1(D_REG_25__SCAN_IN), .A2(n4530), .ZN(U3297) );
  AND2_X1 U5023 ( .A1(D_REG_24__SCAN_IN), .A2(n4530), .ZN(U3298) );
  NOR2_X1 U5024 ( .A1(n4534), .A2(n4523), .ZN(U3299) );
  NOR2_X1 U5025 ( .A1(n4534), .A2(n4524), .ZN(U3300) );
  AND2_X1 U5026 ( .A1(D_REG_21__SCAN_IN), .A2(n4530), .ZN(U3301) );
  NOR2_X1 U5027 ( .A1(n4534), .A2(n4525), .ZN(U3302) );
  AND2_X1 U5028 ( .A1(D_REG_19__SCAN_IN), .A2(n4530), .ZN(U3303) );
  NOR2_X1 U5029 ( .A1(n4534), .A2(n4526), .ZN(U3304) );
  NOR2_X1 U5030 ( .A1(n4534), .A2(n4527), .ZN(U3305) );
  AND2_X1 U5031 ( .A1(D_REG_16__SCAN_IN), .A2(n4530), .ZN(U3306) );
  AND2_X1 U5032 ( .A1(D_REG_15__SCAN_IN), .A2(n4530), .ZN(U3307) );
  AND2_X1 U5033 ( .A1(D_REG_14__SCAN_IN), .A2(n4530), .ZN(U3308) );
  NOR2_X1 U5034 ( .A1(n4534), .A2(n4528), .ZN(U3309) );
  AND2_X1 U5035 ( .A1(D_REG_12__SCAN_IN), .A2(n4530), .ZN(U3310) );
  AND2_X1 U5036 ( .A1(D_REG_11__SCAN_IN), .A2(n4530), .ZN(U3311) );
  NOR2_X1 U5037 ( .A1(n4534), .A2(n4529), .ZN(U3312) );
  AND2_X1 U5038 ( .A1(D_REG_9__SCAN_IN), .A2(n4530), .ZN(U3313) );
  AND2_X1 U5039 ( .A1(D_REG_8__SCAN_IN), .A2(n4530), .ZN(U3314) );
  AND2_X1 U5040 ( .A1(D_REG_7__SCAN_IN), .A2(n4530), .ZN(U3315) );
  AND2_X1 U5041 ( .A1(D_REG_6__SCAN_IN), .A2(n4530), .ZN(U3316) );
  AND2_X1 U5042 ( .A1(D_REG_5__SCAN_IN), .A2(n4530), .ZN(U3317) );
  NOR2_X1 U5043 ( .A1(n4534), .A2(n4531), .ZN(U3318) );
  NOR2_X1 U5044 ( .A1(n4534), .A2(n4532), .ZN(U3319) );
  NOR2_X1 U5045 ( .A1(n4534), .A2(n4533), .ZN(U3320) );
  INV_X1 U5046 ( .A(DATAI_23_), .ZN(n4536) );
  AOI21_X1 U5047 ( .B1(U3149), .B2(n4536), .A(n4535), .ZN(U3329) );
  INV_X1 U5048 ( .A(DATAI_18_), .ZN(n4537) );
  AOI22_X1 U5049 ( .A1(STATE_REG_SCAN_IN), .A2(n4538), .B1(n4537), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U5050 ( .A(DATAI_17_), .ZN(n4539) );
  AOI22_X1 U5051 ( .A1(STATE_REG_SCAN_IN), .A2(n4540), .B1(n4539), .B2(U3149), 
        .ZN(U3335) );
  OAI22_X1 U5052 ( .A1(U3149), .A2(n4541), .B1(DATAI_16_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4542) );
  INV_X1 U5053 ( .A(n4542), .ZN(U3336) );
  INV_X1 U5054 ( .A(DATAI_15_), .ZN(n4543) );
  AOI22_X1 U5055 ( .A1(STATE_REG_SCAN_IN), .A2(n4544), .B1(n4543), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5056 ( .A(DATAI_14_), .ZN(n4545) );
  AOI22_X1 U5057 ( .A1(STATE_REG_SCAN_IN), .A2(n2257), .B1(n4545), .B2(U3149), 
        .ZN(U3338) );
  AOI22_X1 U5058 ( .A1(STATE_REG_SCAN_IN), .A2(n4547), .B1(n4546), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5059 ( .A(DATAI_11_), .ZN(n4548) );
  AOI22_X1 U5060 ( .A1(STATE_REG_SCAN_IN), .A2(n4549), .B1(n4548), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5061 ( .A(DATAI_10_), .ZN(n4550) );
  AOI22_X1 U5062 ( .A1(STATE_REG_SCAN_IN), .A2(n2095), .B1(n4550), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5063 ( .A(DATAI_8_), .ZN(n4551) );
  AOI22_X1 U5064 ( .A1(STATE_REG_SCAN_IN), .A2(n4552), .B1(n4551), .B2(U3149), 
        .ZN(U3344) );
  INV_X1 U5065 ( .A(DATAI_7_), .ZN(n4553) );
  AOI22_X1 U5066 ( .A1(STATE_REG_SCAN_IN), .A2(n4554), .B1(n4553), .B2(U3149), 
        .ZN(U3345) );
  INV_X1 U5067 ( .A(DATAI_6_), .ZN(n4555) );
  AOI22_X1 U5068 ( .A1(STATE_REG_SCAN_IN), .A2(n4556), .B1(n4555), .B2(U3149), 
        .ZN(U3346) );
  AOI211_X1 U5069 ( .C1(n4603), .C2(n4559), .A(n4558), .B(n4557), .ZN(n4607)
         );
  AOI22_X1 U5070 ( .A1(n4606), .A2(n4607), .B1(n2422), .B2(n4604), .ZN(U3467)
         );
  INV_X1 U5071 ( .A(n4560), .ZN(n4564) );
  OAI22_X1 U5072 ( .A1(n4562), .A2(n4572), .B1(n3018), .B2(n4561), .ZN(n4563)
         );
  NOR2_X1 U5073 ( .A1(n4564), .A2(n4563), .ZN(n4609) );
  AOI22_X1 U5074 ( .A1(n4606), .A2(n4609), .B1(n2436), .B2(n4604), .ZN(U3469)
         );
  NOR3_X1 U5075 ( .A1(n4566), .A2(n4565), .A3(n3018), .ZN(n4569) );
  INV_X1 U5076 ( .A(n4567), .ZN(n4568) );
  AOI211_X1 U5077 ( .C1(n4603), .C2(n4570), .A(n4569), .B(n4568), .ZN(n4611)
         );
  AOI22_X1 U5078 ( .A1(n4606), .A2(n4611), .B1(n2449), .B2(n4604), .ZN(U3471)
         );
  OAI22_X1 U5079 ( .A1(n4573), .A2(n4572), .B1(n3018), .B2(n4571), .ZN(n4574)
         );
  NOR2_X1 U5080 ( .A1(n4575), .A2(n4574), .ZN(n4613) );
  AOI22_X1 U5081 ( .A1(n4606), .A2(n4613), .B1(n2371), .B2(n4604), .ZN(U3473)
         );
  NAND2_X1 U5082 ( .A1(n4576), .A2(n4603), .ZN(n4578) );
  NAND2_X1 U5083 ( .A1(n4578), .A2(n4577), .ZN(n4579) );
  NOR2_X1 U5084 ( .A1(n4580), .A2(n4579), .ZN(n4614) );
  AOI22_X1 U5085 ( .A1(n4606), .A2(n4614), .B1(n2395), .B2(n4604), .ZN(U3475)
         );
  NOR2_X1 U5086 ( .A1(n4581), .A2(n4591), .ZN(n4584) );
  INV_X1 U5087 ( .A(n4582), .ZN(n4583) );
  AOI211_X1 U5088 ( .C1(n4596), .C2(n4585), .A(n4584), .B(n4583), .ZN(n4615)
         );
  AOI22_X1 U5089 ( .A1(n4606), .A2(n4615), .B1(n2411), .B2(n4604), .ZN(U3477)
         );
  AOI211_X1 U5090 ( .C1(n4589), .C2(n4588), .A(n4587), .B(n4586), .ZN(n4616)
         );
  AOI22_X1 U5091 ( .A1(n4606), .A2(n4616), .B1(n4590), .B2(n4604), .ZN(U3481)
         );
  NOR2_X1 U5092 ( .A1(n4592), .A2(n4591), .ZN(n4593) );
  AOI211_X1 U5093 ( .C1(n4596), .C2(n4595), .A(n4594), .B(n4593), .ZN(n4617)
         );
  AOI22_X1 U5094 ( .A1(n4606), .A2(n4617), .B1(n4597), .B2(n4604), .ZN(U3485)
         );
  NOR2_X1 U5095 ( .A1(n4598), .A2(n3018), .ZN(n4601) );
  INV_X1 U5096 ( .A(n4599), .ZN(n4600) );
  AOI211_X1 U5097 ( .C1(n4603), .C2(n4602), .A(n4601), .B(n4600), .ZN(n4620)
         );
  INV_X1 U5098 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4605) );
  AOI22_X1 U5099 ( .A1(n4606), .A2(n4620), .B1(n4605), .B2(n4604), .ZN(U3489)
         );
  AOI22_X1 U5100 ( .A1(n4621), .A2(n4607), .B1(n2432), .B2(n4618), .ZN(U3518)
         );
  AOI22_X1 U5101 ( .A1(n4621), .A2(n4609), .B1(n4608), .B2(n4618), .ZN(U3519)
         );
  AOI22_X1 U5102 ( .A1(n4621), .A2(n4611), .B1(n4610), .B2(n4618), .ZN(U3520)
         );
  AOI22_X1 U5103 ( .A1(n4621), .A2(n4613), .B1(n4612), .B2(n4618), .ZN(U3521)
         );
  AOI22_X1 U5104 ( .A1(n4621), .A2(n4614), .B1(n2396), .B2(n4618), .ZN(U3522)
         );
  AOI22_X1 U5105 ( .A1(n4621), .A2(n4615), .B1(n2412), .B2(n4618), .ZN(U3523)
         );
  AOI22_X1 U5106 ( .A1(n4621), .A2(n4616), .B1(n2490), .B2(n4618), .ZN(U3525)
         );
  AOI22_X1 U5107 ( .A1(n4621), .A2(n4617), .B1(n2521), .B2(n4618), .ZN(U3527)
         );
  AOI22_X1 U5108 ( .A1(n4621), .A2(n4620), .B1(n4619), .B2(n4618), .ZN(U3529)
         );
  INV_X2 U2267 ( .A(n2793), .ZN(n2778) );
  CLKBUF_X1 U2273 ( .A(n2498), .Z(n2795) );
  CLKBUF_X1 U2278 ( .A(n2496), .Z(n2843) );
  CLKBUF_X1 U2292 ( .A(n2746), .Z(n2839) );
endmodule

