

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6441, n6442, n6443, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15883, n15884;

  NAND2_X1 U7188 ( .A1(n14781), .A2(n14769), .ZN(n14763) );
  NAND2_X1 U7189 ( .A1(n12794), .A2(n9270), .ZN(n9271) );
  NAND2_X1 U7190 ( .A1(n14815), .A2(n14683), .ZN(n14791) );
  INV_X1 U7191 ( .A(n13720), .ZN(n13966) );
  NAND2_X1 U7192 ( .A1(n8495), .A2(n8029), .ZN(n15168) );
  INV_X2 U7193 ( .A(n12267), .ZN(n12269) );
  INV_X1 U7194 ( .A(n8131), .ZN(n8531) );
  INV_X1 U7195 ( .A(n15591), .ZN(n15620) );
  INV_X1 U7196 ( .A(n9425), .ZN(n9924) );
  AND4_X1 U7197 ( .A1(n8843), .A2(n8842), .A3(n8841), .A4(n8840), .ZN(n15608)
         );
  OAI21_X1 U7198 ( .B1(n10318), .B2(n9907), .A(n9477), .ZN(n11104) );
  INV_X1 U7199 ( .A(n10847), .ZN(n15592) );
  INV_X1 U7200 ( .A(n10254), .ZN(n8113) );
  NAND2_X1 U7201 ( .A1(n8610), .A2(n8558), .ZN(n13742) );
  INV_X2 U7202 ( .A(n9955), .ZN(n10085) );
  INV_X2 U7203 ( .A(n10002), .ZN(n9955) );
  INV_X2 U7204 ( .A(n13744), .ZN(n8610) );
  XNOR2_X1 U7205 ( .A(n10756), .B(n10386), .ZN(n10755) );
  NAND2_X1 U7206 ( .A1(n14817), .A2(n15176), .ZN(n10974) );
  NOR2_X2 U7207 ( .A1(n9352), .A2(n9351), .ZN(n9458) );
  NAND2_X2 U7208 ( .A1(n7140), .A2(n7137), .ZN(n15167) );
  NOR2_X1 U7209 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n9299) );
  NOR2_X1 U7210 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n9298) );
  NOR2_X1 U7211 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n9297) );
  NOR2_X1 U7213 ( .A1(n8344), .A2(n7598), .ZN(n7597) );
  NOR2_X1 U7214 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n9322) );
  OR2_X1 U7215 ( .A1(n12772), .A2(n12796), .ZN(n12783) );
  INV_X1 U7217 ( .A(n9745), .ZN(n12427) );
  AND2_X1 U7218 ( .A1(n14853), .A2(n14833), .ZN(n14835) );
  AND2_X1 U7219 ( .A1(n7767), .A2(n7766), .ZN(n15014) );
  AND4_X1 U7220 ( .A1(n9302), .A2(n9301), .A3(n9371), .A4(n9612), .ZN(n9304)
         );
  CLKBUF_X2 U7221 ( .A(n8897), .Z(n6448) );
  AND2_X1 U7222 ( .A1(n12158), .A2(n12783), .ZN(n12536) );
  OR2_X1 U7223 ( .A1(n9145), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9166) );
  AND4_X1 U7224 ( .A1(n8885), .A2(n8884), .A3(n8883), .A4(n8882), .ZN(n15623)
         );
  NAND2_X1 U7225 ( .A1(n10853), .A2(n12165), .ZN(n13018) );
  INV_X1 U7226 ( .A(n13811), .ZN(n13985) );
  INV_X1 U7227 ( .A(n14026), .ZN(n13986) );
  CLKBUF_X3 U7228 ( .A(n8113), .Z(n8532) );
  INV_X2 U7229 ( .A(n14181), .ZN(n15561) );
  AND2_X1 U7230 ( .A1(n7566), .A2(n7567), .ZN(n13535) );
  NAND2_X1 U7231 ( .A1(n14469), .A2(n14470), .ZN(n7908) );
  NOR4_X1 U7232 ( .A1(n9954), .A2(n9953), .A3(n9952), .A4(n9951), .ZN(n9979)
         );
  BUF_X1 U7233 ( .A(n9443), .Z(n6445) );
  AND2_X1 U7234 ( .A1(n9352), .A2(n9351), .ZN(n9443) );
  NAND2_X1 U7235 ( .A1(n6616), .A2(n14745), .ZN(n15021) );
  NAND2_X1 U7236 ( .A1(n7754), .A2(n15040), .ZN(n14796) );
  AND2_X1 U7237 ( .A1(n14912), .A2(n14899), .ZN(n14894) );
  INV_X1 U7238 ( .A(n10657), .ZN(n9891) );
  NAND2_X1 U7239 ( .A1(n7024), .A2(n7023), .ZN(n9473) );
  AND2_X1 U7240 ( .A1(n9188), .A2(n9187), .ZN(n13051) );
  AND2_X1 U7241 ( .A1(n9108), .A2(n9107), .ZN(n13070) );
  NAND2_X1 U7242 ( .A1(n8373), .A2(n8372), .ZN(n14127) );
  NAND2_X2 U7243 ( .A1(n9872), .A2(n9871), .ZN(n15027) );
  AND4_X1 U7244 ( .A1(n9448), .A2(n9447), .A3(n9446), .A4(n9445), .ZN(n9892)
         );
  XNOR2_X1 U7245 ( .A(n8889), .B(n8888), .ZN(n10436) );
  NAND2_X1 U7246 ( .A1(n8522), .A2(n8521), .ZN(n13809) );
  INV_X1 U7247 ( .A(n15496), .ZN(n13828) );
  INV_X1 U7248 ( .A(n15580), .ZN(n15578) );
  NAND2_X1 U7249 ( .A1(n14650), .A2(n15328), .ZN(n15003) );
  XOR2_X1 U7250 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10367), .Z(n15847) );
  CLKBUF_X3 U7251 ( .A(n8897), .Z(n6449) );
  INV_X2 U7252 ( .A(n15831), .ZN(n14180) );
  AOI21_X2 U7253 ( .B1(n12814), .B2(n9268), .A(n6605), .ZN(n12795) );
  NAND2_X2 U7254 ( .A1(n11955), .A2(n12326), .ZN(n8948) );
  OAI21_X2 U7255 ( .B1(n8711), .B2(P3_D_REG_0__SCAN_IN), .A(n8710), .ZN(n10848) );
  INV_X2 U7256 ( .A(n8111), .ZN(n8535) );
  OR2_X4 U7257 ( .A1(n9363), .A2(n9745), .ZN(n9800) );
  NAND2_X2 U7258 ( .A1(n8991), .A2(n12208), .ZN(n12982) );
  NAND2_X2 U7259 ( .A1(n12995), .A2(n12997), .ZN(n8991) );
  CLKBUF_X1 U7261 ( .A(n7698), .Z(n6441) );
  INV_X1 U7262 ( .A(n7699), .ZN(n7698) );
  XNOR2_X2 U7263 ( .A(n10760), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(n15179) );
  NAND2_X2 U7264 ( .A1(n7164), .A2(n7458), .ZN(n10760) );
  NOR2_X2 U7265 ( .A1(n9271), .A2(n12536), .ZN(n12768) );
  AOI21_X2 U7266 ( .B1(n7708), .B2(n6489), .A(n6727), .ZN(n14688) );
  BUF_X4 U7267 ( .A(n7966), .Z(n6442) );
  BUF_X4 U7268 ( .A(n7966), .Z(n6443) );
  NAND2_X2 U7269 ( .A1(n7604), .A2(n7603), .ZN(n7966) );
  XNOR2_X2 U7270 ( .A(n10383), .B(n10364), .ZN(n10382) );
  NAND2_X2 U7271 ( .A1(n10363), .A2(n10362), .ZN(n10383) );
  OAI21_X2 U7272 ( .B1(n12927), .B2(n9111), .A(n9110), .ZN(n9112) );
  NAND2_X2 U7273 ( .A1(n9062), .A2(n12228), .ZN(n12927) );
  AOI21_X2 U7274 ( .B1(n7597), .B2(n7595), .A(n7594), .ZN(n7593) );
  NAND2_X2 U7275 ( .A1(n10385), .A2(n10384), .ZN(n10756) );
  OAI22_X2 U7276 ( .A1(n14112), .A2(n8594), .B1(n14262), .B2(n13815), .ZN(
        n14098) );
  XNOR2_X2 U7277 ( .A(n11282), .B(n11283), .ZN(n15183) );
  XNOR2_X2 U7278 ( .A(n8838), .B(P3_IR_REG_1__SCAN_IN), .ZN(n10440) );
  XNOR2_X1 U7279 ( .A(n13828), .B(n13535), .ZN(n13763) );
  AND2_X1 U7280 ( .A1(n7868), .A2(n7867), .ZN(n7866) );
  XNOR2_X1 U7281 ( .A(n9223), .B(n9222), .ZN(n12453) );
  AND2_X1 U7282 ( .A1(n7233), .A2(n12792), .ZN(n12800) );
  INV_X1 U7283 ( .A(n13810), .ZN(n13719) );
  AND2_X1 U7284 ( .A1(n9221), .A2(n9220), .ZN(n12796) );
  NAND2_X1 U7285 ( .A1(n9213), .A2(n9212), .ZN(n13036) );
  NAND2_X1 U7287 ( .A1(n8073), .A2(n8072), .ZN(n14008) );
  NAND2_X1 U7288 ( .A1(n14881), .A2(n14679), .ZN(n14866) );
  INV_X1 U7289 ( .A(n14004), .ZN(n8606) );
  OR2_X1 U7290 ( .A1(n8028), .A2(n8027), .ZN(n8495) );
  AND2_X1 U7291 ( .A1(n12175), .A2(n12176), .ZN(n12327) );
  NAND2_X2 U7292 ( .A1(n12180), .A2(n12181), .ZN(n12320) );
  INV_X1 U7293 ( .A(n15623), .ZN(n15639) );
  AND3_X1 U7294 ( .A1(n8864), .A2(n8863), .A3(n8862), .ZN(n15615) );
  CLKBUF_X1 U7295 ( .A(n10847), .Z(n12646) );
  OR2_X1 U7296 ( .A1(n10389), .A2(n10388), .ZN(n7458) );
  INV_X1 U7297 ( .A(n13762), .ZN(n15545) );
  INV_X1 U7298 ( .A(n13379), .ZN(n13314) );
  INV_X2 U7299 ( .A(n9800), .ZN(n9434) );
  INV_X1 U7300 ( .A(n10980), .ZN(n14510) );
  NAND4_X2 U7301 ( .A1(n9472), .A2(n9471), .A3(n9470), .A4(n9469), .ZN(n14509)
         );
  INV_X2 U7302 ( .A(n13515), .ZN(n15533) );
  INV_X1 U7303 ( .A(n13829), .ZN(n11298) );
  AND2_X1 U7305 ( .A1(n8093), .A2(n6602), .ZN(n15496) );
  AND3_X1 U7306 ( .A1(n9460), .A2(n7734), .A3(n7733), .ZN(n10980) );
  NAND2_X2 U7307 ( .A1(n13243), .A2(n13246), .ZN(n8938) );
  INV_X1 U7308 ( .A(n8823), .ZN(n13238) );
  NAND2_X2 U7309 ( .A1(n9942), .A2(n11710), .ZN(n15344) );
  CLKBUF_X2 U7310 ( .A(n8126), .Z(n8530) );
  NAND2_X1 U7311 ( .A1(n9810), .A2(n9339), .ZN(n10296) );
  AOI21_X2 U7312 ( .B1(n8805), .B2(n6495), .A(n7392), .ZN(n7391) );
  INV_X1 U7313 ( .A(n9352), .ZN(n15158) );
  NAND2_X2 U7314 ( .A1(n10339), .A2(P1_U3086), .ZN(n15169) );
  AND2_X1 U7315 ( .A1(n8683), .A2(n7396), .ZN(n7184) );
  AND2_X1 U7316 ( .A1(n8046), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8180) );
  INV_X1 U7317 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7438) );
  OR2_X1 U7319 ( .A1(n7731), .A2(n6572), .ZN(n7039) );
  OAI211_X1 U7320 ( .C1(n6736), .C2(n6735), .A(n8623), .B(n8624), .ZN(n8667)
         );
  AOI21_X1 U7321 ( .B1(n7866), .B2(n7863), .A(n6650), .ZN(n7862) );
  AND2_X1 U7322 ( .A1(n7422), .A2(n12779), .ZN(n13136) );
  OAI211_X1 U7323 ( .C1(n10267), .C2(n7940), .A(n7513), .B(n6550), .ZN(n13954)
         );
  NAND2_X1 U7324 ( .A1(n9280), .A2(n9281), .ZN(n7868) );
  INV_X1 U7325 ( .A(n6916), .ZN(n6915) );
  NAND2_X1 U7326 ( .A1(n10267), .A2(n6536), .ZN(n7513) );
  OAI21_X1 U7327 ( .B1(n12453), .B2(n13138), .A(n15676), .ZN(n7790) );
  INV_X1 U7328 ( .A(n6481), .ZN(n6446) );
  AND2_X1 U7329 ( .A1(n14771), .A2(n14772), .ZN(n7358) );
  NOR2_X1 U7330 ( .A1(n15014), .A2(n15013), .ZN(n15015) );
  NAND2_X1 U7331 ( .A1(n12790), .A2(n12791), .ZN(n12792) );
  INV_X1 U7332 ( .A(n7766), .ZN(n14725) );
  NAND2_X1 U7333 ( .A1(n14459), .A2(n9751), .ZN(n14389) );
  NAND2_X1 U7334 ( .A1(n6994), .A2(n6992), .ZN(n14444) );
  AND2_X1 U7335 ( .A1(n7265), .A2(n6977), .ZN(n12726) );
  XNOR2_X1 U7336 ( .A(n12492), .B(n12490), .ZN(n12599) );
  NAND2_X1 U7337 ( .A1(n15207), .A2(n15206), .ZN(n15212) );
  NAND2_X1 U7338 ( .A1(n15199), .A2(n7145), .ZN(n15207) );
  NAND2_X1 U7339 ( .A1(n12383), .A2(n12382), .ZN(n12381) );
  AOI21_X1 U7340 ( .B1(n12454), .B2(n10248), .A(n6669), .ZN(n14314) );
  NAND2_X1 U7341 ( .A1(n7773), .A2(n9263), .ZN(n12846) );
  OR2_X1 U7342 ( .A1(n12914), .A2(n12885), .ZN(n12903) );
  NAND2_X2 U7343 ( .A1(n8498), .A2(n8497), .ZN(n13974) );
  XNOR2_X1 U7344 ( .A(n14638), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n7334) );
  NAND2_X1 U7345 ( .A1(n7069), .A2(n6539), .ZN(n13305) );
  NOR2_X1 U7346 ( .A1(n12915), .A2(n6867), .ZN(n12914) );
  XNOR2_X1 U7347 ( .A(n8508), .B(n8496), .ZN(n12448) );
  NAND2_X1 U7348 ( .A1(n6922), .A2(n6919), .ZN(n14893) );
  OR2_X1 U7349 ( .A1(n13382), .A2(n8530), .ZN(n8538) );
  NAND2_X1 U7350 ( .A1(n15185), .A2(n15184), .ZN(n7464) );
  OR2_X1 U7351 ( .A1(n9214), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n12761) );
  NAND2_X1 U7352 ( .A1(n9790), .A2(n9789), .ZN(n14795) );
  NAND2_X1 U7353 ( .A1(n8482), .A2(n8481), .ZN(n14217) );
  NOR2_X1 U7354 ( .A1(n14849), .A2(n7722), .ZN(n7721) );
  NAND2_X2 U7355 ( .A1(n12241), .A2(n12242), .ZN(n12887) );
  OR2_X1 U7356 ( .A1(n13484), .A2(n13485), .ZN(n13489) );
  AND2_X1 U7357 ( .A1(n9173), .A2(n9172), .ZN(n13050) );
  NAND2_X1 U7358 ( .A1(n8449), .A2(n8448), .ZN(n14059) );
  NAND2_X1 U7359 ( .A1(n7085), .A2(n7084), .ZN(n7083) );
  INV_X1 U7360 ( .A(n14854), .ZN(n15058) );
  OAI21_X1 U7361 ( .B1(n11991), .B2(n6800), .A(n7800), .ZN(n12508) );
  NAND2_X1 U7362 ( .A1(n8420), .A2(n8419), .ZN(n14092) );
  AND2_X1 U7363 ( .A1(n15177), .A2(n7215), .ZN(n14854) );
  NAND2_X1 U7364 ( .A1(n8405), .A2(n8404), .ZN(n14105) );
  NAND2_X1 U7365 ( .A1(n9125), .A2(n9124), .ZN(n12908) );
  OR2_X1 U7366 ( .A1(n7448), .A2(n7450), .ZN(n7447) );
  XNOR2_X1 U7367 ( .A(n14597), .B(n7339), .ZN(n14600) );
  OAI21_X1 U7368 ( .B1(n11840), .B2(n11841), .A(n7425), .ZN(n11844) );
  NAND2_X1 U7369 ( .A1(n8430), .A2(n8418), .ZN(n12447) );
  NAND2_X1 U7370 ( .A1(n9671), .A2(n9670), .ZN(n15083) );
  AND2_X1 U7371 ( .A1(n14668), .A2(n7705), .ZN(n7704) );
  NAND2_X1 U7372 ( .A1(n11275), .A2(n11274), .ZN(n11282) );
  INV_X1 U7373 ( .A(n14671), .ZN(n14943) );
  NAND2_X1 U7374 ( .A1(n11831), .A2(n11830), .ZN(n15290) );
  AOI21_X1 U7375 ( .B1(n7401), .B2(n7783), .A(n6515), .ZN(n7399) );
  NAND2_X1 U7376 ( .A1(n7166), .A2(n7206), .ZN(n11275) );
  NOR2_X2 U7377 ( .A1(n14194), .A2(n14296), .ZN(n14193) );
  AND2_X1 U7378 ( .A1(n6781), .A2(n6779), .ZN(n11640) );
  AND2_X1 U7379 ( .A1(n7165), .A2(n11274), .ZN(n7166) );
  NAND2_X1 U7380 ( .A1(n7315), .A2(n7317), .ZN(n7105) );
  NAND2_X1 U7381 ( .A1(n9632), .A2(n9631), .ZN(n15103) );
  NAND2_X1 U7382 ( .A1(n11523), .A2(n12327), .ZN(n8875) );
  NAND2_X1 U7383 ( .A1(n7419), .A2(n6457), .ZN(n7418) );
  NAND2_X1 U7384 ( .A1(n7461), .A2(n7459), .ZN(n11274) );
  OR2_X1 U7385 ( .A1(n9091), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9102) );
  AND2_X1 U7386 ( .A1(n7427), .A2(n11466), .ZN(n10150) );
  NAND2_X1 U7387 ( .A1(n8273), .A2(n8272), .ZN(n13585) );
  XNOR2_X1 U7388 ( .A(n8316), .B(n8318), .ZN(n10554) );
  NAND2_X1 U7389 ( .A1(n9581), .A2(n9580), .ZN(n15116) );
  NOR2_X1 U7390 ( .A1(n12322), .A2(n7781), .ZN(n7780) );
  NAND2_X1 U7391 ( .A1(n11280), .A2(n11279), .ZN(n11286) );
  NAND2_X1 U7392 ( .A1(n8955), .A2(n8954), .ZN(n12057) );
  NAND2_X1 U7393 ( .A1(n15630), .A2(n8928), .ZN(n12182) );
  NAND2_X1 U7394 ( .A1(n10775), .A2(n10774), .ZN(n11277) );
  NAND4_X1 U7395 ( .A1(n8978), .A2(n8977), .A3(n8976), .A4(n8975), .ZN(n12998)
         );
  NAND2_X1 U7397 ( .A1(n8911), .A2(n6684), .ZN(n15636) );
  AND3_X1 U7398 ( .A1(n8895), .A2(n8894), .A3(n8893), .ZN(n11541) );
  NOR2_X2 U7399 ( .A1(n6493), .A2(n7424), .ZN(n15619) );
  INV_X1 U7400 ( .A(n11310), .ZN(n15356) );
  INV_X1 U7401 ( .A(n15608), .ZN(n13012) );
  AND3_X1 U7402 ( .A1(n8849), .A2(n8848), .A3(n8847), .ZN(n15585) );
  AOI21_X1 U7403 ( .B1(n10768), .B2(n10767), .A(n10766), .ZN(n10773) );
  NOR2_X1 U7404 ( .A1(n9844), .A2(n11046), .ZN(n14491) );
  OAI211_X1 U7405 ( .C1(n9038), .C2(n10421), .A(n8830), .B(n8829), .ZN(n11397)
         );
  OAI211_X1 U7406 ( .C1(n8837), .C2(n9038), .A(n7405), .B(n6809), .ZN(n13014)
         );
  NAND3_X1 U7407 ( .A1(n7775), .A2(n8833), .A3(n7774), .ZN(n10847) );
  NAND4_X1 U7408 ( .A1(n8963), .A2(n8962), .A3(n8961), .A4(n8960), .ZN(n12643)
         );
  AND4_X1 U7409 ( .A1(n8856), .A2(n8855), .A3(n8854), .A4(n8853), .ZN(n15591)
         );
  NAND2_X1 U7410 ( .A1(n6703), .A2(n6702), .ZN(n8985) );
  AND2_X1 U7411 ( .A1(n8835), .A2(n8834), .ZN(n7774) );
  BUF_X2 U7412 ( .A(n8851), .Z(n9058) );
  NAND4_X1 U7413 ( .A1(n8235), .A2(n8234), .A3(n8233), .A4(n8232), .ZN(n13823)
         );
  INV_X4 U7414 ( .A(n12300), .ZN(n7776) );
  NAND4_X1 U7415 ( .A1(n8117), .A2(n8116), .A3(n8115), .A4(n8114), .ZN(n13508)
         );
  NAND4_X1 U7416 ( .A1(n8085), .A2(n8084), .A3(n8083), .A4(n8082), .ZN(n13829)
         );
  NAND2_X2 U7417 ( .A1(n12461), .A2(n13238), .ZN(n8880) );
  AOI21_X1 U7418 ( .B1(n7571), .B2(n8261), .A(n7569), .ZN(n7568) );
  NAND2_X1 U7419 ( .A1(n9424), .A2(n9423), .ZN(n14512) );
  NAND2_X2 U7421 ( .A1(n10296), .A2(n10973), .ZN(n9745) );
  NAND2_X1 U7422 ( .A1(n8818), .A2(n8804), .ZN(n13243) );
  AND2_X2 U7423 ( .A1(n12456), .A2(n14363), .ZN(n8111) );
  AND2_X1 U7424 ( .A1(n8820), .A2(n13232), .ZN(n8823) );
  NAND2_X1 U7425 ( .A1(n7202), .A2(n7201), .ZN(n8804) );
  INV_X2 U7426 ( .A(n8123), .ZN(n10248) );
  NAND2_X1 U7427 ( .A1(n9362), .A2(n9361), .ZN(n11050) );
  NAND2_X1 U7428 ( .A1(n7195), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8275) );
  XNOR2_X1 U7429 ( .A(n8686), .B(P3_IR_REG_20__SCAN_IN), .ZN(n9286) );
  NAND2_X1 U7430 ( .A1(n8699), .A2(n8698), .ZN(n11818) );
  NAND2_X1 U7431 ( .A1(n8546), .A2(n8545), .ZN(n13744) );
  NAND2_X1 U7432 ( .A1(n7818), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8676) );
  NAND2_X1 U7433 ( .A1(n9338), .A2(n9337), .ZN(n15171) );
  AND2_X1 U7434 ( .A1(n9342), .A2(n9358), .ZN(n10987) );
  INV_X1 U7435 ( .A(n7249), .ZN(n15173) );
  NAND2_X1 U7436 ( .A1(n6937), .A2(n6940), .ZN(n15162) );
  XNOR2_X1 U7437 ( .A(n9348), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9352) );
  OR2_X1 U7438 ( .A1(n9311), .A2(n9310), .ZN(n7140) );
  OAI21_X1 U7439 ( .B1(n9824), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9327) );
  XNOR2_X1 U7440 ( .A(n8149), .B(n8151), .ZN(n13861) );
  AND2_X1 U7441 ( .A1(n9343), .A2(n9374), .ZN(n9940) );
  XNOR2_X1 U7442 ( .A(n6734), .B(n8058), .ZN(n8615) );
  NAND2_X1 U7443 ( .A1(n9347), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9348) );
  OAI21_X1 U7444 ( .B1(n6499), .B2(n9368), .A(n9372), .ZN(n9374) );
  AND2_X1 U7445 ( .A1(n8332), .A2(n6609), .ZN(n8401) );
  CLKBUF_X1 U7446 ( .A(n8332), .Z(n8626) );
  NOR2_X1 U7447 ( .A1(n8540), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n7514) );
  NAND2_X1 U7448 ( .A1(n10358), .A2(n10357), .ZN(n10371) );
  OAI211_X2 U7449 ( .C1(n10139), .C2(n7645), .A(n7646), .B(n7642), .ZN(n10947)
         );
  NAND2_X1 U7450 ( .A1(n8180), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8229) );
  AND3_X1 U7451 ( .A1(n8036), .A2(n8348), .A3(n8285), .ZN(n8041) );
  AND2_X1 U7452 ( .A1(n10359), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n7157) );
  INV_X1 U7453 ( .A(n7814), .ZN(n7813) );
  AND3_X1 U7454 ( .A1(n8682), .A2(n7395), .A3(n7394), .ZN(n7396) );
  AND3_X1 U7455 ( .A1(n13832), .A2(n8035), .A3(n8086), .ZN(n8036) );
  AND3_X1 U7456 ( .A1(n8034), .A2(n8302), .A3(n8033), .ZN(n8348) );
  NOR2_X1 U7457 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n8285) );
  INV_X1 U7458 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9335) );
  INV_X1 U7459 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9377) );
  INV_X4 U7460 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7461 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n8216) );
  INV_X1 U7462 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9612) );
  INV_X1 U7463 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8891) );
  NOR2_X1 U7464 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n8670) );
  NOR2_X1 U7465 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n8671) );
  NOR2_X1 U7466 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n8669) );
  NOR2_X1 U7467 ( .A1(P3_IR_REG_24__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n7395) );
  INV_X1 U7468 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n15774) );
  INV_X4 U7469 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7470 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9371) );
  NOR2_X1 U7471 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n9302) );
  NOR2_X1 U7472 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n9301) );
  NOR2_X1 U7473 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n7811) );
  NOR2_X1 U7474 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n8674) );
  INV_X1 U7475 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8673) );
  INV_X1 U7476 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7439) );
  INV_X1 U7477 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9022) );
  NOR2_X1 U7478 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), .ZN(
        n8679) );
  INV_X4 U7479 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7480 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8097) );
  INV_X1 U7481 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8098) );
  NAND3_X1 U7482 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n8182) );
  NOR2_X1 U7483 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .ZN(
        n8682) );
  OR2_X2 U7484 ( .A1(n9450), .A2(n15153), .ZN(n9451) );
  NOR2_X2 U7485 ( .A1(n8308), .A2(n8307), .ZN(n7196) );
  NAND2_X1 U7486 ( .A1(n8048), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8308) );
  AOI21_X1 U7487 ( .B1(n7500), .B2(n7499), .A(n8608), .ZN(n7498) );
  AND2_X2 U7488 ( .A1(n10518), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n10365) );
  OAI21_X2 U7490 ( .B1(n8948), .B2(n7872), .A(n7869), .ZN(n12995) );
  AND4_X2 U7491 ( .A1(n8870), .A2(n8869), .A3(n8868), .A4(n8867), .ZN(n15628)
         );
  INV_X1 U7492 ( .A(n8880), .ZN(n6447) );
  AND2_X1 U7493 ( .A1(n8821), .A2(n8823), .ZN(n8897) );
  NAND2_X1 U7494 ( .A1(n12231), .A2(n12896), .ZN(n7611) );
  OR2_X1 U7495 ( .A1(n13139), .A2(n12539), .ZN(n12345) );
  OR2_X1 U7496 ( .A1(n13002), .A2(n12642), .ZN(n12208) );
  INV_X1 U7497 ( .A(n8459), .ZN(n7561) );
  INV_X1 U7498 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8302) );
  AND2_X1 U7499 ( .A1(n12398), .A2(n12392), .ZN(n12395) );
  NOR2_X1 U7500 ( .A1(n7765), .A2(n14726), .ZN(n7764) );
  NAND2_X1 U7501 ( .A1(n15020), .A2(n14769), .ZN(n7765) );
  AND3_X1 U7502 ( .A1(n6909), .A2(n6908), .A3(n6907), .ZN(n9328) );
  NOR2_X1 U7503 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n6909) );
  NOR2_X1 U7504 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n6908) );
  INV_X1 U7505 ( .A(n11769), .ZN(n7521) );
  INV_X1 U7506 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n13832) );
  INV_X1 U7507 ( .A(n13785), .ZN(n10283) );
  NAND2_X1 U7508 ( .A1(n13996), .A2(n6543), .ZN(n7301) );
  AOI21_X1 U7509 ( .B1(n7552), .B2(n7549), .A(n6549), .ZN(n7548) );
  INV_X1 U7510 ( .A(n6484), .ZN(n7549) );
  XNOR2_X1 U7511 ( .A(n15033), .B(n14800), .ZN(n14779) );
  AOI21_X1 U7512 ( .B1(n14772), .B2(n7710), .A(n6575), .ZN(n7709) );
  INV_X1 U7513 ( .A(n14685), .ZN(n7710) );
  OAI211_X1 U7514 ( .C1(n13838), .C2(n6966), .A(n10582), .B(n6965), .ZN(n13834) );
  NAND2_X1 U7515 ( .A1(n13838), .A2(n6966), .ZN(n6965) );
  AND2_X1 U7516 ( .A1(n7026), .A2(n7025), .ZN(n7744) );
  NAND2_X1 U7517 ( .A1(n10002), .A2(n11104), .ZN(n7025) );
  NAND2_X1 U7518 ( .A1(n9955), .A2(n14509), .ZN(n7026) );
  NAND2_X1 U7519 ( .A1(n13517), .A2(n13516), .ZN(n13525) );
  INV_X1 U7520 ( .A(n7031), .ZN(n7030) );
  INV_X1 U7521 ( .A(n12173), .ZN(n7619) );
  INV_X1 U7522 ( .A(n13582), .ZN(n6715) );
  AOI21_X1 U7523 ( .B1(n6864), .B2(n6865), .A(n12240), .ZN(n6863) );
  INV_X1 U7524 ( .A(n7611), .ZN(n6865) );
  AOI21_X1 U7525 ( .B1(n8011), .B2(n7582), .A(n7585), .ZN(n7584) );
  NAND2_X1 U7526 ( .A1(n7099), .A2(n7102), .ZN(n7587) );
  INV_X1 U7527 ( .A(n8462), .ZN(n7585) );
  NOR2_X1 U7528 ( .A1(n7606), .A2(n12847), .ZN(n7605) );
  AND2_X1 U7529 ( .A1(n12263), .A2(n12269), .ZN(n6847) );
  NOR2_X1 U7530 ( .A1(n13473), .A2(n7173), .ZN(n13322) );
  INV_X1 U7531 ( .A(n13466), .ZN(n7173) );
  OR2_X1 U7532 ( .A1(n15107), .A2(n14981), .ZN(n14666) );
  NAND2_X1 U7533 ( .A1(n7761), .A2(n11242), .ZN(n7760) );
  NOR2_X1 U7534 ( .A1(n7102), .A2(n7588), .ZN(n7101) );
  INV_X1 U7535 ( .A(n8317), .ZN(n7993) );
  NAND2_X1 U7536 ( .A1(n7995), .A2(n10503), .ZN(n7998) );
  OAI21_X1 U7537 ( .B1(n6442), .B2(n10346), .A(n7238), .ZN(n7965) );
  NAND2_X1 U7538 ( .A1(n6442), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7238) );
  NOR2_X1 U7539 ( .A1(n9166), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n7170) );
  OR2_X1 U7540 ( .A1(n10143), .A2(n10423), .ZN(n10144) );
  NAND2_X1 U7541 ( .A1(n10811), .A2(n10810), .ZN(n7632) );
  NAND2_X1 U7542 ( .A1(n7632), .A2(n7631), .ZN(n7630) );
  NAND2_X1 U7543 ( .A1(n10436), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7631) );
  OR2_X1 U7544 ( .A1(n10230), .A2(n13112), .ZN(n7629) );
  NAND2_X1 U7545 ( .A1(n7367), .A2(n7365), .ZN(n7363) );
  OR2_X1 U7546 ( .A1(n9193), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9207) );
  NAND2_X1 U7547 ( .A1(n15619), .A2(n15628), .ZN(n12176) );
  AND2_X1 U7548 ( .A1(n12345), .A2(n12349), .ZN(n12771) );
  XNOR2_X1 U7549 ( .A(n12801), .B(n13036), .ZN(n12791) );
  OR2_X1 U7550 ( .A1(n13168), .A2(n12860), .ZN(n12243) );
  NAND2_X1 U7551 ( .A1(n9099), .A2(n10440), .ZN(n6809) );
  OR2_X1 U7552 ( .A1(n7404), .A2(n10441), .ZN(n7405) );
  NOR2_X1 U7553 ( .A1(n9141), .A2(n7669), .ZN(n7668) );
  INV_X1 U7554 ( .A(n8788), .ZN(n7669) );
  NAND2_X1 U7555 ( .A1(n10346), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8754) );
  AND2_X1 U7556 ( .A1(n13735), .A2(n13734), .ZN(n7478) );
  AND2_X1 U7557 ( .A1(n7581), .A2(n7580), .ZN(n13732) );
  AND2_X1 U7558 ( .A1(n13966), .A2(n7914), .ZN(n7915) );
  NOR2_X1 U7559 ( .A1(n13983), .A2(n7254), .ZN(n7253) );
  NAND2_X1 U7560 ( .A1(n8055), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8500) );
  OR2_X1 U7561 ( .A1(n8485), .A2(n8074), .ZN(n8076) );
  NAND2_X1 U7562 ( .A1(n8054), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8485) );
  INV_X1 U7563 ( .A(n8483), .ZN(n8054) );
  NOR2_X1 U7564 ( .A1(n7554), .A2(n8315), .ZN(n7552) );
  OR2_X1 U7565 ( .A1(n11700), .A2(n6777), .ZN(n6774) );
  INV_X1 U7566 ( .A(n8573), .ZN(n6777) );
  AND2_X1 U7567 ( .A1(n7294), .A2(n8174), .ZN(n7543) );
  AND2_X1 U7568 ( .A1(n8141), .A2(n8139), .ZN(n7293) );
  INV_X1 U7569 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8039) );
  INV_X1 U7570 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n8038) );
  NOR3_X1 U7571 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .A3(
        P2_IR_REG_22__SCAN_IN), .ZN(n8031) );
  AND2_X1 U7572 ( .A1(n8549), .A2(n8030), .ZN(n8539) );
  NOR2_X1 U7573 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n8030) );
  NOR3_X1 U7574 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n8032) );
  INV_X1 U7575 ( .A(n14445), .ZN(n7223) );
  NOR2_X1 U7576 ( .A1(n11720), .A2(n7019), .ZN(n11722) );
  AND2_X1 U7577 ( .A1(n11721), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7019) );
  AOI21_X1 U7578 ( .B1(n7704), .B2(n7707), .A(n7703), .ZN(n7702) );
  INV_X1 U7579 ( .A(n14670), .ZN(n7703) );
  INV_X1 U7580 ( .A(n12028), .ZN(n7353) );
  NOR2_X1 U7581 ( .A1(n11237), .A2(n7120), .ZN(n7119) );
  INV_X1 U7582 ( .A(n11108), .ZN(n7120) );
  AND2_X1 U7583 ( .A1(n11250), .A2(n7762), .ZN(n7761) );
  NAND2_X1 U7584 ( .A1(n6570), .A2(n11106), .ZN(n7118) );
  NAND2_X1 U7585 ( .A1(n9852), .A2(n9851), .ZN(n9912) );
  OAI21_X1 U7586 ( .B1(n8524), .B2(n8523), .A(n8513), .ZN(n9852) );
  INV_X1 U7587 ( .A(n7998), .ZN(n7594) );
  INV_X1 U7588 ( .A(n7599), .ZN(n7595) );
  NAND2_X1 U7589 ( .A1(n7093), .A2(n7091), .ZN(n8299) );
  AOI21_X1 U7590 ( .B1(n7095), .B2(n7941), .A(n7094), .ZN(n7093) );
  AND2_X1 U7591 ( .A1(n7941), .A2(n7975), .ZN(n7092) );
  XNOR2_X1 U7592 ( .A(n7965), .B(SI_7_), .ZN(n8200) );
  XNOR2_X1 U7593 ( .A(n7961), .B(SI_5_), .ZN(n8158) );
  AOI21_X1 U7594 ( .B1(n11498), .B2(n7451), .A(n7455), .ZN(n7450) );
  NAND2_X1 U7595 ( .A1(n7796), .A2(n7795), .ZN(n7794) );
  NAND2_X1 U7596 ( .A1(n12343), .A2(n10849), .ZN(n10850) );
  NAND2_X1 U7597 ( .A1(n6796), .A2(n6797), .ZN(n12546) );
  AND2_X1 U7598 ( .A1(n6604), .A2(n6798), .ZN(n6797) );
  NAND2_X1 U7599 ( .A1(n7821), .A2(n12608), .ZN(n6798) );
  NOR2_X1 U7600 ( .A1(n12562), .A2(n7799), .ZN(n7798) );
  INV_X1 U7601 ( .A(n12473), .ZN(n7799) );
  NAND2_X1 U7602 ( .A1(n15804), .A2(n15680), .ZN(n8878) );
  AOI21_X1 U7603 ( .B1(n11654), .B2(n11746), .A(n6552), .ZN(n7809) );
  NAND2_X1 U7604 ( .A1(n11423), .A2(n6780), .ZN(n6779) );
  INV_X1 U7605 ( .A(n11420), .ZN(n6780) );
  NAND2_X1 U7606 ( .A1(n12499), .A2(n12498), .ZN(n7840) );
  NOR2_X1 U7607 ( .A1(n7627), .A2(n12275), .ZN(n7624) );
  XNOR2_X1 U7608 ( .A(n7630), .B(n6979), .ZN(n11124) );
  INV_X1 U7609 ( .A(n10808), .ZN(n7387) );
  NAND2_X1 U7610 ( .A1(n11782), .A2(n11781), .ZN(n11849) );
  AND2_X1 U7611 ( .A1(n11847), .A2(n10233), .ZN(n6836) );
  NAND2_X1 U7612 ( .A1(n11788), .A2(n10188), .ZN(n11846) );
  INV_X1 U7613 ( .A(n6838), .ZN(n6837) );
  OAI21_X1 U7614 ( .B1(n11847), .B2(n6635), .A(n6839), .ZN(n6838) );
  NAND2_X1 U7615 ( .A1(n6840), .A2(n10233), .ZN(n6839) );
  INV_X1 U7616 ( .A(n7629), .ZN(n6840) );
  NAND2_X1 U7617 ( .A1(n12690), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n12689) );
  NOR2_X1 U7618 ( .A1(n12697), .A2(n12696), .ZN(n12695) );
  AOI21_X1 U7619 ( .B1(n6459), .B2(n7368), .A(n6660), .ZN(n7367) );
  OAI21_X1 U7620 ( .B1(n12728), .B2(n13089), .A(n7256), .ZN(n12747) );
  NAND2_X1 U7621 ( .A1(n12704), .A2(n7638), .ZN(n7257) );
  INV_X1 U7622 ( .A(n9264), .ZN(n7415) );
  NAND2_X1 U7623 ( .A1(n12846), .A2(n12847), .ZN(n9265) );
  INV_X1 U7624 ( .A(n9058), .ZN(n9276) );
  INV_X2 U7625 ( .A(n8880), .ZN(n9273) );
  NAND2_X1 U7626 ( .A1(n9233), .A2(n9232), .ZN(n11956) );
  INV_X1 U7627 ( .A(n7778), .ZN(n7777) );
  OAI21_X1 U7628 ( .B1(n7780), .B2(n7779), .A(n11636), .ZN(n7778) );
  INV_X1 U7630 ( .A(n12771), .ZN(n12785) );
  AOI21_X1 U7631 ( .B1(n7881), .B2(n7880), .A(n7879), .ZN(n7878) );
  INV_X1 U7632 ( .A(n12241), .ZN(n7880) );
  INV_X1 U7633 ( .A(n12247), .ZN(n7879) );
  OR2_X1 U7634 ( .A1(n13073), .A2(n12528), .ZN(n12241) );
  AND2_X1 U7635 ( .A1(n7854), .A2(n12220), .ZN(n7853) );
  NAND2_X1 U7636 ( .A1(n7786), .A2(n9236), .ZN(n7784) );
  INV_X1 U7637 ( .A(n8711), .ZN(n12155) );
  AND2_X1 U7638 ( .A1(n7792), .A2(n8802), .ZN(n7791) );
  NAND2_X1 U7639 ( .A1(n9127), .A2(n9126), .ZN(n9129) );
  NAND3_X1 U7640 ( .A1(n6899), .A2(n7230), .A3(n8786), .ZN(n9115) );
  AOI21_X1 U7641 ( .B1(n6881), .B2(n6883), .A(n6878), .ZN(n6877) );
  INV_X1 U7642 ( .A(n8780), .ZN(n6878) );
  NAND2_X1 U7643 ( .A1(n9050), .A2(n8777), .ZN(n6880) );
  INV_X1 U7644 ( .A(n6897), .ZN(n6896) );
  NAND2_X1 U7645 ( .A1(n8922), .A2(n8754), .ZN(n8943) );
  NAND2_X1 U7646 ( .A1(n8943), .A2(n8942), .ZN(n8945) );
  NAND2_X1 U7647 ( .A1(n6888), .A2(n6886), .ZN(n8906) );
  INV_X1 U7648 ( .A(n6887), .ZN(n6886) );
  NAND2_X1 U7649 ( .A1(n10139), .A2(n8846), .ZN(n8859) );
  NAND2_X1 U7650 ( .A1(n7647), .A2(n8846), .ZN(n7646) );
  NAND2_X1 U7651 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7645) );
  AND2_X1 U7652 ( .A1(n11619), .A2(n11618), .ZN(n7244) );
  XNOR2_X1 U7653 ( .A(n13379), .B(n15524), .ZN(n10875) );
  XNOR2_X1 U7654 ( .A(n13974), .B(n13985), .ZN(n13785) );
  NAND2_X1 U7655 ( .A1(n8062), .A2(n8063), .ZN(n8126) );
  INV_X1 U7656 ( .A(n14363), .ZN(n8062) );
  NAND2_X1 U7657 ( .A1(n13901), .A2(n13902), .ZN(n13910) );
  INV_X1 U7658 ( .A(n13786), .ZN(n10274) );
  NAND2_X1 U7659 ( .A1(n7917), .A2(n7916), .ZN(n10271) );
  NOR2_X1 U7660 ( .A1(n13720), .A2(n13974), .ZN(n7916) );
  OR2_X1 U7661 ( .A1(n14008), .A2(n14026), .ZN(n8492) );
  AND3_X1 U7662 ( .A1(n6742), .A2(n6741), .A3(n6613), .ZN(n13996) );
  OR2_X1 U7663 ( .A1(n7558), .A2(n6743), .ZN(n6742) );
  NAND2_X1 U7664 ( .A1(n14065), .A2(n13755), .ZN(n6744) );
  OAI21_X1 U7665 ( .B1(n14065), .B2(n13757), .A(n13755), .ZN(n14053) );
  NOR2_X1 U7666 ( .A1(n7545), .A2(n7285), .ZN(n7284) );
  INV_X1 U7667 ( .A(n8366), .ZN(n7285) );
  NAND2_X1 U7668 ( .A1(n7548), .A2(n6807), .ZN(n7547) );
  AND2_X1 U7669 ( .A1(n11813), .A2(n6512), .ZN(n6807) );
  OR2_X1 U7670 ( .A1(n13590), .A2(n14189), .ZN(n7556) );
  NAND2_X1 U7671 ( .A1(n7300), .A2(n8210), .ZN(n7299) );
  INV_X1 U7672 ( .A(n8252), .ZN(n7300) );
  NAND2_X1 U7673 ( .A1(n11352), .A2(n11354), .ZN(n6770) );
  INV_X1 U7674 ( .A(n13826), .ZN(n15494) );
  CLKBUF_X1 U7675 ( .A(n10737), .Z(n15501) );
  INV_X1 U7677 ( .A(n10250), .ZN(n8403) );
  INV_X1 U7678 ( .A(n8202), .ZN(n10576) );
  NAND2_X1 U7679 ( .A1(n13744), .A2(n8559), .ZN(n15518) );
  INV_X1 U7680 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8035) );
  INV_X1 U7681 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8033) );
  AOI21_X1 U7682 ( .B1(n7889), .B2(n7890), .A(n6500), .ZN(n7888) );
  NAND2_X1 U7683 ( .A1(n11591), .A2(n11590), .ZN(n11589) );
  NAND2_X1 U7684 ( .A1(n12381), .A2(n7898), .ZN(n14404) );
  NOR2_X1 U7685 ( .A1(n14407), .A2(n7899), .ZN(n7898) );
  INV_X1 U7686 ( .A(n9718), .ZN(n7899) );
  OAI21_X1 U7687 ( .B1(n12447), .B2(n9907), .A(n9706), .ZN(n14702) );
  NAND2_X1 U7688 ( .A1(n7910), .A2(n7909), .ZN(n11930) );
  NOR2_X1 U7689 ( .A1(n11933), .A2(n9569), .ZN(n7909) );
  NOR2_X1 U7690 ( .A1(n9649), .A2(n7904), .ZN(n7903) );
  INV_X1 U7691 ( .A(n9610), .ZN(n7904) );
  AND2_X1 U7692 ( .A1(n9780), .A2(n9779), .ZN(n14798) );
  INV_X1 U7693 ( .A(n9458), .ZN(n9353) );
  NAND2_X1 U7694 ( .A1(n7125), .A2(n7123), .ZN(n14757) );
  AND2_X1 U7695 ( .A1(n7124), .A2(n14685), .ZN(n7123) );
  NAND2_X1 U7696 ( .A1(n14777), .A2(n6942), .ZN(n14716) );
  AND2_X1 U7697 ( .A1(n9874), .A2(n9836), .ZN(n14782) );
  AND2_X1 U7698 ( .A1(n7128), .A2(n14779), .ZN(n7127) );
  AOI21_X1 U7699 ( .B1(n7721), .B2(n7719), .A(n7718), .ZN(n7717) );
  INV_X1 U7700 ( .A(n7721), .ZN(n7720) );
  INV_X1 U7701 ( .A(n14681), .ZN(n7718) );
  AOI21_X1 U7702 ( .B1(n14893), .B2(n14697), .A(n6556), .ZN(n14880) );
  NAND2_X1 U7703 ( .A1(n14918), .A2(n14919), .ZN(n7143) );
  AOI21_X1 U7704 ( .B1(n6464), .B2(n7696), .A(n6555), .ZN(n7692) );
  NOR2_X1 U7705 ( .A1(n11829), .A2(n7725), .ZN(n7724) );
  INV_X1 U7706 ( .A(n14721), .ZN(n14717) );
  OAI22_X1 U7707 ( .A1(n14763), .A2(n7763), .B1(n15344), .B2(n14726), .ZN(
        n7767) );
  OR2_X1 U7708 ( .A1(n14748), .A2(n15344), .ZN(n7763) );
  AND2_X1 U7709 ( .A1(n9328), .A2(n6523), .ZN(n6453) );
  INV_X1 U7710 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9308) );
  INV_X1 U7711 ( .A(n9347), .ZN(n6939) );
  NAND2_X1 U7712 ( .A1(n9358), .A2(n7260), .ZN(n9362) );
  NOR2_X1 U7713 ( .A1(n9360), .A2(n9359), .ZN(n9361) );
  NOR2_X1 U7714 ( .A1(n9326), .A2(n15153), .ZN(n7260) );
  OAI21_X1 U7715 ( .B1(n9520), .B2(P1_IR_REG_8__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9533) );
  NAND2_X1 U7716 ( .A1(n10763), .A2(n10762), .ZN(n10770) );
  NAND2_X1 U7717 ( .A1(n15224), .A2(n15223), .ZN(n7162) );
  NAND2_X1 U7718 ( .A1(n8809), .A2(n8808), .ZN(n12772) );
  OR2_X1 U7719 ( .A1(n11164), .A2(n15628), .ZN(n7797) );
  OAI21_X1 U7720 ( .B1(n10951), .B2(n10932), .A(n10933), .ZN(n10935) );
  NAND2_X1 U7721 ( .A1(n10802), .A2(n10211), .ZN(n7388) );
  AND2_X1 U7722 ( .A1(n12772), .A2(n12991), .ZN(n6707) );
  NAND2_X1 U7723 ( .A1(n10583), .A2(n13834), .ZN(n13846) );
  NAND2_X1 U7724 ( .A1(n10287), .A2(n10286), .ZN(n10288) );
  NAND2_X1 U7725 ( .A1(n12448), .A2(n9461), .ZN(n9872) );
  NAND2_X1 U7726 ( .A1(n9889), .A2(n9888), .ZN(n14758) );
  OAI21_X1 U7727 ( .B1(n14766), .B2(n9876), .A(n9881), .ZN(n14741) );
  OAI211_X1 U7728 ( .C1(n13507), .C2(n13506), .A(n13505), .B(n13504), .ZN(
        n13518) );
  NAND2_X1 U7729 ( .A1(n7738), .A2(n7737), .ZN(n10006) );
  NAND2_X1 U7730 ( .A1(n7739), .A2(n7743), .ZN(n7737) );
  INV_X1 U7731 ( .A(n7744), .ZN(n7743) );
  NOR2_X1 U7732 ( .A1(n12031), .A2(n10027), .ZN(n10055) );
  OR2_X1 U7733 ( .A1(n10015), .A2(n10014), .ZN(n10016) );
  INV_X1 U7734 ( .A(n7028), .ZN(n7027) );
  OAI21_X1 U7735 ( .B1(n7030), .B2(n7029), .A(n10023), .ZN(n7028) );
  AND2_X1 U7736 ( .A1(n7750), .A2(n7032), .ZN(n7029) );
  NAND2_X1 U7737 ( .A1(n13544), .A2(n13546), .ZN(n7466) );
  AND2_X1 U7738 ( .A1(n6597), .A2(n6718), .ZN(n6716) );
  NAND2_X1 U7739 ( .A1(n6565), .A2(n13550), .ZN(n6718) );
  AND2_X1 U7740 ( .A1(n12327), .A2(n7616), .ZN(n7615) );
  NAND2_X1 U7741 ( .A1(n7217), .A2(n7216), .ZN(n10065) );
  INV_X1 U7742 ( .A(n10062), .ZN(n7216) );
  AND2_X1 U7743 ( .A1(n10069), .A2(n14919), .ZN(n10070) );
  OR2_X1 U7744 ( .A1(n12206), .A2(n12994), .ZN(n6816) );
  OR2_X1 U7745 ( .A1(n13572), .A2(n13571), .ZN(n13578) );
  NOR2_X1 U7746 ( .A1(n13577), .A2(n6506), .ZN(n6713) );
  NOR2_X1 U7747 ( .A1(n6490), .A2(n6715), .ZN(n6714) );
  OR3_X1 U7748 ( .A1(n13623), .A2(n13622), .A3(n13621), .ZN(n13645) );
  INV_X1 U7749 ( .A(n10095), .ZN(n7250) );
  NAND2_X1 U7750 ( .A1(n10091), .A2(n7045), .ZN(n7044) );
  AND2_X1 U7751 ( .A1(n10093), .A2(n7047), .ZN(n7046) );
  INV_X1 U7752 ( .A(n10091), .ZN(n7047) );
  AND2_X1 U7753 ( .A1(n7472), .A2(n13656), .ZN(n7469) );
  INV_X1 U7754 ( .A(n7473), .ZN(n7472) );
  AOI21_X1 U7755 ( .B1(n7473), .B2(n6470), .A(n6558), .ZN(n7471) );
  OR2_X1 U7756 ( .A1(n12226), .A2(n7613), .ZN(n7612) );
  NAND2_X1 U7757 ( .A1(n7614), .A2(n12228), .ZN(n7613) );
  NAND2_X1 U7758 ( .A1(n12227), .A2(n12269), .ZN(n7614) );
  AOI21_X1 U7759 ( .B1(n6863), .B2(n6861), .A(n6579), .ZN(n6860) );
  INV_X1 U7760 ( .A(n6864), .ZN(n6861) );
  INV_X1 U7761 ( .A(n12239), .ZN(n6866) );
  INV_X1 U7762 ( .A(n6863), .ZN(n6862) );
  NAND2_X1 U7763 ( .A1(n6723), .A2(n6724), .ZN(n13664) );
  NAND2_X1 U7764 ( .A1(n13660), .A2(n13661), .ZN(n6724) );
  NAND2_X1 U7765 ( .A1(n10104), .A2(n10106), .ZN(n7746) );
  INV_X1 U7766 ( .A(n10110), .ZN(n7753) );
  NOR2_X1 U7767 ( .A1(n7051), .A2(n10107), .ZN(n7052) );
  NAND2_X1 U7768 ( .A1(n10107), .A2(n7051), .ZN(n7050) );
  AND2_X1 U7769 ( .A1(n13132), .A2(n12760), .ZN(n12315) );
  NOR2_X1 U7770 ( .A1(n6849), .A2(n12269), .ZN(n6848) );
  INV_X1 U7771 ( .A(n12260), .ZN(n6849) );
  INV_X1 U7772 ( .A(n6843), .ZN(n6842) );
  OAI21_X1 U7773 ( .B1(n6573), .B2(n6845), .A(n12791), .ZN(n6843) );
  INV_X1 U7774 ( .A(n6847), .ZN(n6845) );
  INV_X1 U7775 ( .A(n11084), .ZN(n7435) );
  OAI21_X1 U7776 ( .B1(n10147), .B2(n7435), .A(n10149), .ZN(n7434) );
  NOR2_X1 U7777 ( .A1(n10186), .A2(n6830), .ZN(n6829) );
  INV_X1 U7778 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n6830) );
  INV_X1 U7779 ( .A(n9162), .ZN(n7663) );
  OR2_X1 U7780 ( .A1(n14314), .A2(n13736), .ZN(n7581) );
  NAND2_X1 U7781 ( .A1(n13714), .A2(n13808), .ZN(n7580) );
  NAND2_X1 U7782 ( .A1(n14210), .A2(n8606), .ZN(n8607) );
  AND2_X1 U7783 ( .A1(n8463), .A2(n8444), .ZN(n7277) );
  INV_X1 U7784 ( .A(n7568), .ZN(n7095) );
  OAI21_X1 U7785 ( .B1(n6442), .B2(P2_DATAO_REG_11__SCAN_IN), .A(n7261), .ZN(
        n7980) );
  OR2_X1 U7786 ( .A1(n10339), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7261) );
  OAI21_X1 U7787 ( .B1(n6443), .B2(n10401), .A(n7279), .ZN(n7978) );
  NAND2_X1 U7788 ( .A1(n6443), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7279) );
  NAND2_X1 U7789 ( .A1(n10377), .A2(n14546), .ZN(n10363) );
  INV_X1 U7790 ( .A(n10848), .ZN(n7796) );
  INV_X1 U7791 ( .A(n12361), .ZN(n7795) );
  NOR2_X1 U7792 ( .A1(n12465), .A2(n7806), .ZN(n7805) );
  INV_X1 U7793 ( .A(n11999), .ZN(n7806) );
  AND2_X1 U7794 ( .A1(n11420), .A2(n11162), .ZN(n6782) );
  NAND2_X1 U7795 ( .A1(n6693), .A2(n6692), .ZN(n6691) );
  NOR2_X1 U7796 ( .A1(n12900), .A2(n12884), .ZN(n6692) );
  INV_X1 U7797 ( .A(n12835), .ZN(n7259) );
  AOI21_X1 U7798 ( .B1(n12341), .B2(n12349), .A(n12357), .ZN(n12311) );
  NAND2_X1 U7799 ( .A1(n12342), .A2(n12312), .ZN(n12313) );
  INV_X1 U7800 ( .A(n12315), .ZN(n12348) );
  NOR2_X1 U7801 ( .A1(n11088), .A2(n10214), .ZN(n6853) );
  NOR2_X1 U7802 ( .A1(n11088), .A2(n6979), .ZN(n6852) );
  OR2_X1 U7803 ( .A1(n11194), .A2(n7428), .ZN(n7427) );
  AND2_X1 U7804 ( .A1(n10428), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7428) );
  AND2_X1 U7805 ( .A1(n11459), .A2(n6503), .ZN(n7379) );
  NOR2_X1 U7806 ( .A1(n11844), .A2(n6975), .ZN(n10154) );
  NOR2_X1 U7807 ( .A1(n10230), .A2(n10153), .ZN(n6975) );
  INV_X1 U7808 ( .A(n12705), .ZN(n7635) );
  INV_X1 U7809 ( .A(n6494), .ZN(n7411) );
  NAND2_X1 U7810 ( .A1(n9181), .A2(n9180), .ZN(n9193) );
  INV_X1 U7811 ( .A(n9182), .ZN(n9181) );
  OR2_X1 U7812 ( .A1(n13046), .A2(n13051), .ZN(n12261) );
  INV_X1 U7813 ( .A(n9229), .ZN(n7781) );
  OR2_X1 U7814 ( .A1(n13162), .A2(n12848), .ZN(n12250) );
  OR2_X1 U7815 ( .A1(n13094), .A2(n13097), .ZN(n12222) );
  NOR2_X1 U7816 ( .A1(n9017), .A2(n7860), .ZN(n7859) );
  INV_X1 U7817 ( .A(n12213), .ZN(n7860) );
  OR2_X1 U7818 ( .A1(n13206), .A2(n12985), .ZN(n12216) );
  XNOR2_X1 U7819 ( .A(n12057), .B(n12643), .ZN(n11920) );
  NAND2_X1 U7820 ( .A1(n11956), .A2(n7785), .ZN(n11919) );
  INV_X1 U7821 ( .A(n7786), .ZN(n7785) );
  OR2_X1 U7822 ( .A1(n9038), .A2(SI_4_), .ZN(n8874) );
  AND2_X1 U7823 ( .A1(n8702), .A2(n7793), .ZN(n7792) );
  INV_X1 U7824 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7793) );
  NOR2_X1 U7825 ( .A1(n8693), .A2(n8695), .ZN(n8691) );
  NOR2_X1 U7826 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n7817) );
  NAND2_X1 U7827 ( .A1(n7678), .A2(n7676), .ZN(n8785) );
  AOI21_X1 U7828 ( .B1(n7679), .B2(n7681), .A(n7677), .ZN(n7676) );
  INV_X1 U7829 ( .A(n8784), .ZN(n7677) );
  NAND2_X1 U7830 ( .A1(n10315), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8741) );
  AND2_X1 U7831 ( .A1(n13300), .A2(n13827), .ZN(n11472) );
  AOI21_X1 U7832 ( .B1(n13458), .B2(n7073), .A(n7072), .ZN(n7071) );
  INV_X1 U7833 ( .A(n13292), .ZN(n7072) );
  NOR2_X1 U7834 ( .A1(n13388), .A2(n13295), .ZN(n7528) );
  INV_X1 U7835 ( .A(n13442), .ZN(n7526) );
  INV_X1 U7836 ( .A(n7528), .ZN(n7527) );
  INV_X1 U7837 ( .A(n7071), .ZN(n7070) );
  OR2_X1 U7838 ( .A1(n7527), .A2(n7067), .ZN(n7066) );
  NAND2_X1 U7839 ( .A1(n7071), .A2(n7068), .ZN(n7067) );
  INV_X1 U7840 ( .A(n7073), .ZN(n7068) );
  NAND2_X2 U7841 ( .A1(n10737), .A2(n13742), .ZN(n13379) );
  INV_X1 U7842 ( .A(n13432), .ZN(n7535) );
  INV_X1 U7843 ( .A(n13322), .ZN(n7532) );
  NOR2_X1 U7844 ( .A1(n6974), .A2(n11378), .ZN(n6973) );
  INV_X1 U7845 ( .A(n11376), .ZN(n6974) );
  OR2_X1 U7846 ( .A1(n8500), .A2(n8499), .ZN(n8528) );
  NAND2_X1 U7847 ( .A1(n7496), .A2(n7495), .ZN(n7501) );
  NOR2_X1 U7848 ( .A1(n8603), .A2(n7499), .ZN(n7495) );
  NAND2_X1 U7849 ( .A1(n6767), .A2(n6765), .ZN(n13998) );
  NAND2_X1 U7850 ( .A1(n7504), .A2(n8598), .ZN(n6767) );
  NAND2_X1 U7851 ( .A1(n8053), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8483) );
  INV_X1 U7852 ( .A(n8468), .ZN(n8053) );
  NOR2_X1 U7853 ( .A1(n14100), .A2(n14092), .ZN(n7919) );
  AND2_X1 U7854 ( .A1(n6516), .A2(n12099), .ZN(n6958) );
  AOI21_X1 U7855 ( .B1(n8573), .B2(n6776), .A(n6524), .ZN(n6775) );
  INV_X1 U7856 ( .A(n8572), .ZN(n6776) );
  NOR2_X1 U7857 ( .A1(n13829), .A2(n15533), .ZN(n8566) );
  INV_X1 U7858 ( .A(n6762), .ZN(n6760) );
  OAI22_X1 U7859 ( .A1(n10283), .A2(n7557), .B1(n13985), .B2(n14318), .ZN(
        n6757) );
  AND2_X1 U7860 ( .A1(n14058), .A2(n6954), .ZN(n14011) );
  NOR2_X1 U7861 ( .A1(n6955), .A2(n14008), .ZN(n6954) );
  INV_X1 U7862 ( .A(n6956), .ZN(n6955) );
  NOR2_X1 U7863 ( .A1(n9773), .A2(n9772), .ZN(n6720) );
  NAND2_X1 U7864 ( .A1(n9919), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7735) );
  NAND2_X1 U7865 ( .A1(n14361), .A2(n9461), .ZN(n7110) );
  OR2_X1 U7866 ( .A1(n14748), .A2(n14758), .ZN(n14714) );
  NAND2_X1 U7867 ( .A1(n14748), .A2(n14758), .ZN(n14719) );
  NOR2_X1 U7868 ( .A1(n9694), .A2(n15744), .ZN(n6733) );
  NAND2_X1 U7869 ( .A1(n6925), .A2(n6928), .ZN(n6921) );
  NOR2_X1 U7870 ( .A1(n6492), .A2(n6924), .ZN(n6923) );
  INV_X1 U7871 ( .A(n6925), .ZN(n6924) );
  NOR2_X1 U7872 ( .A1(n14694), .A2(n6930), .ZN(n6929) );
  INV_X1 U7873 ( .A(n14693), .ZN(n6930) );
  AND2_X1 U7874 ( .A1(n14966), .A2(n14690), .ZN(n14671) );
  AND2_X1 U7875 ( .A1(n15103), .A2(n12018), .ZN(n14669) );
  NAND2_X1 U7876 ( .A1(n14663), .A2(n7706), .ZN(n7705) );
  INV_X1 U7877 ( .A(n7945), .ZN(n7714) );
  NOR2_X1 U7878 ( .A1(n7716), .A2(n7945), .ZN(n7715) );
  NOR2_X1 U7879 ( .A1(n15126), .A2(n15417), .ZN(n7771) );
  OAI21_X1 U7880 ( .B1(n11254), .B2(n7348), .A(n11829), .ZN(n7347) );
  INV_X1 U7881 ( .A(n11255), .ZN(n7348) );
  NOR2_X1 U7882 ( .A1(n7118), .A2(n6454), .ZN(n7117) );
  NAND2_X1 U7883 ( .A1(n10987), .A2(n11513), .ZN(n10973) );
  NOR2_X1 U7884 ( .A1(n7760), .A2(n11987), .ZN(n7757) );
  XNOR2_X1 U7885 ( .A(n14509), .B(n11104), .ZN(n11102) );
  NAND2_X1 U7886 ( .A1(n7090), .A2(n7600), .ZN(n8524) );
  AOI21_X1 U7887 ( .B1(n7602), .B2(n7601), .A(n6645), .ZN(n7600) );
  NAND2_X1 U7888 ( .A1(n8026), .A2(SI_26_), .ZN(n8494) );
  NAND2_X1 U7889 ( .A1(n8024), .A2(SI_24_), .ZN(n7576) );
  NAND2_X1 U7890 ( .A1(n7097), .A2(n7100), .ZN(n8016) );
  NAND2_X1 U7891 ( .A1(n7104), .A2(n7102), .ZN(n7100) );
  NOR2_X1 U7892 ( .A1(n7318), .A2(n7101), .ZN(n7098) );
  INV_X1 U7893 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9326) );
  NAND2_X1 U7894 ( .A1(n8012), .A2(n12379), .ZN(n8432) );
  AND4_X1 U7895 ( .A1(n7111), .A2(n7024), .A3(n9304), .A4(n9306), .ZN(n9313)
         );
  NOR2_X1 U7896 ( .A1(n9366), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n7111) );
  NAND2_X1 U7897 ( .A1(n7315), .A2(n7314), .ZN(n8429) );
  NOR2_X1 U7898 ( .A1(n7318), .A2(n10964), .ZN(n7314) );
  INV_X1 U7899 ( .A(n8380), .ZN(n7322) );
  AOI21_X1 U7900 ( .B1(n7593), .B2(n7596), .A(n7590), .ZN(n7589) );
  INV_X1 U7901 ( .A(n7942), .ZN(n7590) );
  INV_X1 U7902 ( .A(n7597), .ZN(n7596) );
  AND2_X1 U7903 ( .A1(n7991), .A2(n6599), .ZN(n7599) );
  NAND2_X1 U7904 ( .A1(n7998), .A2(n7997), .ZN(n8344) );
  NAND2_X1 U7905 ( .A1(n7988), .A2(n10510), .ZN(n7991) );
  NAND2_X1 U7906 ( .A1(n8299), .A2(n7937), .ZN(n7992) );
  NAND2_X1 U7907 ( .A1(n7976), .A2(n7975), .ZN(n8260) );
  NAND2_X1 U7908 ( .A1(n6586), .A2(n7200), .ZN(n7967) );
  INV_X1 U7909 ( .A(n8200), .ZN(n7200) );
  OAI21_X1 U7910 ( .B1(n7966), .B2(n10319), .A(n7252), .ZN(n8089) );
  NAND2_X1 U7911 ( .A1(n6443), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7252) );
  NAND2_X1 U7912 ( .A1(n7564), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n7604) );
  NAND3_X1 U7913 ( .A1(n7948), .A2(n14648), .A3(n7565), .ZN(n7564) );
  INV_X1 U7914 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7565) );
  INV_X1 U7915 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7563) );
  AND2_X1 U7916 ( .A1(n10360), .A2(n10370), .ZN(n7151) );
  AND2_X1 U7917 ( .A1(n11735), .A2(n11734), .ZN(n11739) );
  AND2_X1 U7918 ( .A1(n7835), .A2(n6623), .ZN(n7834) );
  NAND2_X1 U7919 ( .A1(n7837), .A2(n7836), .ZN(n7835) );
  INV_X1 U7920 ( .A(n7805), .ZN(n7804) );
  AOI21_X1 U7921 ( .B1(n7805), .B2(n11992), .A(n7803), .ZN(n7802) );
  INV_X1 U7922 ( .A(n12464), .ZN(n7803) );
  INV_X1 U7923 ( .A(n12534), .ZN(n7831) );
  OR2_X1 U7924 ( .A1(n7834), .A2(n7831), .ZN(n7830) );
  INV_X1 U7925 ( .A(n13014), .ZN(n10845) );
  AND2_X1 U7926 ( .A1(n10891), .A2(n10852), .ZN(n10857) );
  AOI21_X1 U7927 ( .B1(n7821), .B2(n7824), .A(n6567), .ZN(n7819) );
  AOI21_X1 U7928 ( .B1(n7798), .B2(n12625), .A(n6571), .ZN(n6786) );
  INV_X1 U7929 ( .A(n7798), .ZN(n6787) );
  INV_X1 U7930 ( .A(n9074), .ZN(n9089) );
  AND2_X1 U7931 ( .A1(n6482), .A2(n12481), .ZN(n7827) );
  NAND2_X1 U7932 ( .A1(n7826), .A2(n6482), .ZN(n7825) );
  INV_X1 U7933 ( .A(n12524), .ZN(n7826) );
  INV_X1 U7934 ( .A(n11991), .ZN(n11994) );
  NAND2_X1 U7935 ( .A1(n12546), .A2(n12488), .ZN(n12492) );
  AND2_X1 U7936 ( .A1(n10862), .A2(n12365), .ZN(n10844) );
  NAND2_X1 U7937 ( .A1(n12471), .A2(n12470), .ZN(n12622) );
  INV_X1 U7938 ( .A(n11291), .ZN(n12368) );
  AND4_X1 U7939 ( .A1(n9002), .A2(n9001), .A3(n9000), .A4(n8999), .ZN(n11996)
         );
  NAND2_X1 U7940 ( .A1(n11124), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n6855) );
  AOI22_X1 U7941 ( .A1(n11190), .A2(n11191), .B1(P3_REG1_REG_8__SCAN_IN), .B2(
        n10428), .ZN(n10182) );
  NOR2_X1 U7942 ( .A1(n6638), .A2(n11783), .ZN(n6982) );
  NAND2_X1 U7943 ( .A1(n11849), .A2(n6642), .ZN(n12653) );
  NAND2_X1 U7944 ( .A1(n7444), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7443) );
  OAI211_X1 U7945 ( .C1(n11846), .C2(n6835), .A(P3_REG1_REG_13__SCAN_IN), .B(
        n6832), .ZN(n12649) );
  NAND2_X1 U7946 ( .A1(n6837), .A2(n6635), .ZN(n6835) );
  AND2_X1 U7947 ( .A1(n6834), .A2(n6837), .ZN(n6833) );
  NAND2_X1 U7948 ( .A1(n12689), .A2(n10193), .ZN(n12706) );
  AND2_X1 U7949 ( .A1(n7431), .A2(n7429), .ZN(n12708) );
  AND2_X1 U7950 ( .A1(n12709), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7430) );
  INV_X1 U7951 ( .A(n7363), .ZN(n7360) );
  NAND2_X1 U7952 ( .A1(n7363), .A2(n7364), .ZN(n7362) );
  NOR2_X1 U7953 ( .A1(n12821), .A2(n7413), .ZN(n7412) );
  INV_X1 U7954 ( .A(n9266), .ZN(n7413) );
  NOR2_X1 U7955 ( .A1(n12254), .A2(n7852), .ZN(n7851) );
  INV_X1 U7956 ( .A(n12250), .ZN(n7852) );
  NAND2_X1 U7957 ( .A1(n12852), .A2(n12251), .ZN(n9152) );
  INV_X1 U7958 ( .A(n12860), .ZN(n12889) );
  AND4_X1 U7959 ( .A1(n9047), .A2(n9046), .A3(n9045), .A4(n9044), .ZN(n12943)
         );
  OR2_X1 U7960 ( .A1(n9247), .A2(n9246), .ZN(n9248) );
  INV_X1 U7961 ( .A(n7271), .ZN(n8997) );
  INV_X1 U7962 ( .A(n8973), .ZN(n6703) );
  NOR2_X1 U7963 ( .A1(n12198), .A2(n7877), .ZN(n7876) );
  INV_X1 U7964 ( .A(n12194), .ZN(n7877) );
  AND2_X1 U7965 ( .A1(n12194), .A2(n12195), .ZN(n12326) );
  AOI21_X1 U7966 ( .B1(n8896), .B2(n7847), .A(n6577), .ZN(n7846) );
  INV_X1 U7967 ( .A(n12176), .ZN(n7847) );
  AND4_X1 U7968 ( .A1(n8937), .A2(n8936), .A3(n8935), .A4(n8934), .ZN(n11663)
         );
  NAND2_X1 U7969 ( .A1(n11536), .A2(n7780), .ZN(n11517) );
  NAND2_X1 U7970 ( .A1(n8875), .A2(n12176), .ZN(n11535) );
  AND2_X1 U7971 ( .A1(n12636), .A2(n15656), .ZN(n9279) );
  AND2_X1 U7972 ( .A1(n9144), .A2(n9143), .ZN(n12489) );
  OR2_X1 U7973 ( .A1(n12245), .A2(n12244), .ZN(n12873) );
  OR2_X1 U7974 ( .A1(n12881), .A2(n12887), .ZN(n12883) );
  AND2_X1 U7975 ( .A1(n12359), .A2(n9287), .ZN(n13052) );
  AOI21_X1 U7976 ( .B1(n7859), .B2(n12984), .A(n7857), .ZN(n7856) );
  INV_X1 U7977 ( .A(n12216), .ZN(n7857) );
  INV_X1 U7978 ( .A(n7859), .ZN(n7858) );
  AND2_X1 U7979 ( .A1(n12208), .A2(n12209), .ZN(n12997) );
  AND2_X2 U7980 ( .A1(n11569), .A2(n9231), .ZN(n9233) );
  AOI21_X1 U7981 ( .B1(n7782), .B2(n7403), .A(n6551), .ZN(n7401) );
  AND2_X1 U7982 ( .A1(n12269), .A2(n10843), .ZN(n15656) );
  AND2_X1 U7983 ( .A1(n10829), .A2(n13224), .ZN(n10865) );
  AND2_X1 U7984 ( .A1(n12269), .A2(n10839), .ZN(n15638) );
  NAND2_X1 U7985 ( .A1(n7267), .A2(n7266), .ZN(n8711) );
  INV_X1 U7986 ( .A(n13253), .ZN(n7266) );
  OAI21_X1 U7987 ( .B1(n12279), .B2(n12278), .A(n12277), .ZN(n13229) );
  NOR2_X1 U7988 ( .A1(n8800), .A2(n7689), .ZN(n7688) );
  INV_X1 U7989 ( .A(n8797), .ZN(n7689) );
  OR2_X1 U7990 ( .A1(n9190), .A2(n8796), .ZN(n8798) );
  OR2_X1 U7991 ( .A1(n8725), .A2(P3_IR_REG_24__SCAN_IN), .ZN(n8698) );
  AOI21_X1 U7992 ( .B1(n7666), .B2(n7668), .A(n6671), .ZN(n7665) );
  INV_X1 U7993 ( .A(n9126), .ZN(n7666) );
  INV_X1 U7994 ( .A(n7668), .ZN(n7667) );
  INV_X1 U7995 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8677) );
  INV_X1 U7996 ( .A(n8691), .ZN(n8723) );
  NOR2_X1 U7997 ( .A1(n9083), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n9067) );
  NAND2_X1 U7998 ( .A1(n9115), .A2(n8786), .ZN(n9127) );
  INV_X1 U7999 ( .A(n7680), .ZN(n7679) );
  OAI21_X1 U8000 ( .B1(n9063), .B2(n7681), .A(n9095), .ZN(n7680) );
  INV_X1 U8001 ( .A(n8782), .ZN(n7681) );
  NAND2_X1 U8002 ( .A1(n9064), .A2(n9063), .ZN(n9066) );
  OR2_X1 U8003 ( .A1(n9051), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n9083) );
  AND2_X1 U8004 ( .A1(n8780), .A2(n8779), .ZN(n9079) );
  INV_X1 U8005 ( .A(n6882), .ZN(n6881) );
  OAI21_X1 U8006 ( .B1(n8777), .B2(n6883), .A(n9079), .ZN(n6882) );
  INV_X1 U8007 ( .A(n8778), .ZN(n6883) );
  NAND2_X1 U8008 ( .A1(n6902), .A2(n6900), .ZN(n8775) );
  AND2_X1 U8009 ( .A1(n6901), .A2(n7656), .ZN(n6900) );
  AOI21_X1 U8010 ( .B1(n6583), .B2(n8770), .A(n7658), .ZN(n7657) );
  INV_X1 U8011 ( .A(n8772), .ZN(n7658) );
  AND2_X1 U8012 ( .A1(n10507), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8771) );
  INV_X1 U8013 ( .A(n8770), .ZN(n7659) );
  NAND2_X1 U8014 ( .A1(n8993), .A2(n8765), .ZN(n8767) );
  AND2_X1 U8015 ( .A1(n8761), .A2(n8760), .ZN(n8964) );
  NAND2_X1 U8016 ( .A1(n8965), .A2(n8964), .ZN(n8967) );
  AND2_X1 U8017 ( .A1(n8758), .A2(n8757), .ZN(n8949) );
  OR2_X1 U8018 ( .A1(n8939), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8951) );
  AND2_X1 U8019 ( .A1(n8756), .A2(n8755), .ZN(n8942) );
  OR2_X1 U8020 ( .A1(n8923), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n8939) );
  INV_X1 U8021 ( .A(n8919), .ZN(n8753) );
  NAND2_X1 U8022 ( .A1(n8731), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8836) );
  NAND2_X1 U8023 ( .A1(n7194), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8293) );
  INV_X1 U8024 ( .A(n8275), .ZN(n7194) );
  OAI22_X1 U8025 ( .A1(n13340), .A2(n13308), .B1(n13307), .B2(n13341), .ZN(
        n13309) );
  INV_X1 U8026 ( .A(n14024), .ZN(n13754) );
  NAND2_X1 U8027 ( .A1(n8051), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8421) );
  INV_X1 U8028 ( .A(n8407), .ZN(n8051) );
  NAND2_X1 U8029 ( .A1(n7065), .A2(n7071), .ZN(n13441) );
  NAND2_X1 U8030 ( .A1(n13457), .A2(n7073), .ZN(n7065) );
  NAND2_X1 U8031 ( .A1(n13441), .A2(n13442), .ZN(n13440) );
  INV_X1 U8032 ( .A(n7061), .ZN(n7060) );
  OAI21_X1 U8033 ( .B1(n7063), .B2(n7062), .A(n12135), .ZN(n7061) );
  OR2_X1 U8034 ( .A1(n8126), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8094) );
  OR2_X1 U8035 ( .A1(n8375), .A2(n8374), .ZN(n8388) );
  NAND2_X1 U8036 ( .A1(n13433), .A2(n13432), .ZN(n13467) );
  NAND2_X1 U8037 ( .A1(n8612), .A2(n8561), .ZN(n13786) );
  AOI21_X1 U8038 ( .B1(n7478), .B2(n6488), .A(n7477), .ZN(n7476) );
  INV_X1 U8039 ( .A(n13741), .ZN(n7477) );
  AND2_X1 U8040 ( .A1(n7478), .A2(n13708), .ZN(n7262) );
  NAND2_X1 U8041 ( .A1(n8063), .A2(n14363), .ZN(n10254) );
  NOR2_X1 U8042 ( .A1(n8126), .A2(n11027), .ZN(n8129) );
  OAI21_X1 U8043 ( .B1(n13838), .B2(P2_REG1_REG_1__SCAN_IN), .A(n6701), .ZN(
        n13836) );
  NAND2_X1 U8044 ( .A1(n13838), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6701) );
  AOI21_X1 U8045 ( .B1(n15457), .B2(n13868), .A(n13867), .ZN(n13866) );
  INV_X1 U8046 ( .A(n6963), .ZN(n6962) );
  OAI21_X1 U8047 ( .B1(n10591), .B2(n6964), .A(n15472), .ZN(n6963) );
  AOI21_X1 U8048 ( .B1(n6962), .B2(n6964), .A(n6960), .ZN(n6959) );
  INV_X1 U8049 ( .A(n10614), .ZN(n6960) );
  AOI21_X1 U8050 ( .B1(n13883), .B2(P2_REG1_REG_15__SCAN_IN), .A(n7306), .ZN(
        n13895) );
  AND2_X1 U8051 ( .A1(n7308), .A2(n13884), .ZN(n7306) );
  XNOR2_X1 U8052 ( .A(n13933), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n13934) );
  INV_X1 U8053 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7948) );
  INV_X1 U8054 ( .A(n14314), .ZN(n13946) );
  NAND2_X1 U8055 ( .A1(n8515), .A2(n8514), .ZN(n13955) );
  NOR2_X1 U8056 ( .A1(n8493), .A2(n6763), .ZN(n6762) );
  INV_X1 U8057 ( .A(n8492), .ZN(n6763) );
  AND2_X1 U8058 ( .A1(n13993), .A2(n8606), .ZN(n8493) );
  NAND2_X1 U8059 ( .A1(n8605), .A2(n8600), .ZN(n14000) );
  OR2_X1 U8060 ( .A1(n14008), .A2(n13986), .ZN(n8600) );
  AND2_X1 U8061 ( .A1(n8076), .A2(n8075), .ZN(n14012) );
  NOR2_X1 U8062 ( .A1(n7560), .A2(n6746), .ZN(n6745) );
  AND2_X1 U8063 ( .A1(n13757), .A2(n13755), .ZN(n6746) );
  AOI21_X1 U8064 ( .B1(n7559), .B2(n7561), .A(n6538), .ZN(n7558) );
  NAND2_X1 U8065 ( .A1(n14053), .A2(n14052), .ZN(n14051) );
  NAND2_X1 U8066 ( .A1(n6466), .A2(n14055), .ZN(n14054) );
  AND2_X1 U8067 ( .A1(n7313), .A2(n6591), .ZN(n7506) );
  OR2_X1 U8068 ( .A1(n14081), .A2(n7312), .ZN(n7313) );
  NAND2_X1 U8069 ( .A1(n8595), .A2(n8596), .ZN(n7312) );
  NAND2_X1 U8070 ( .A1(n14080), .A2(n8428), .ZN(n14065) );
  OR2_X1 U8071 ( .A1(n14098), .A2(n8596), .ZN(n7508) );
  NAND2_X1 U8072 ( .A1(n8397), .A2(n6471), .ZN(n7305) );
  NAND2_X1 U8073 ( .A1(n7305), .A2(n7304), .ZN(n14080) );
  AND2_X1 U8074 ( .A1(n14081), .A2(n8414), .ZN(n7304) );
  INV_X1 U8075 ( .A(n13300), .ZN(n14181) );
  NAND2_X1 U8076 ( .A1(n14110), .A2(n14111), .ZN(n8397) );
  AND2_X1 U8077 ( .A1(n7546), .A2(n8330), .ZN(n7545) );
  OR2_X1 U8078 ( .A1(n8356), .A2(n8355), .ZN(n8358) );
  AND2_X1 U8079 ( .A1(n6791), .A2(n7509), .ZN(n6790) );
  NAND2_X1 U8080 ( .A1(n6587), .A2(n8583), .ZN(n7509) );
  NAND2_X1 U8081 ( .A1(n6460), .A2(n8577), .ZN(n6791) );
  INV_X1 U8082 ( .A(n6460), .ZN(n6792) );
  INV_X1 U8083 ( .A(n7552), .ZN(n7550) );
  NAND2_X1 U8084 ( .A1(n7555), .A2(n6533), .ZN(n7554) );
  NAND2_X1 U8085 ( .A1(n6484), .A2(n8282), .ZN(n7555) );
  NAND2_X1 U8086 ( .A1(n8579), .A2(n8578), .ZN(n8581) );
  AOI21_X1 U8087 ( .B1(n7492), .B2(n7490), .A(n6517), .ZN(n7489) );
  NAND2_X1 U8088 ( .A1(n6774), .A2(n6772), .ZN(n6778) );
  INV_X1 U8089 ( .A(n8575), .ZN(n7490) );
  XNOR2_X1 U8090 ( .A(n13585), .B(n13820), .ZN(n13772) );
  NAND2_X1 U8091 ( .A1(n6739), .A2(n8267), .ZN(n11813) );
  OR2_X1 U8092 ( .A1(n11414), .A2(n7299), .ZN(n7298) );
  NAND2_X1 U8093 ( .A1(n6774), .A2(n6775), .ZN(n11865) );
  OAI21_X1 U8094 ( .B1(n11410), .B2(n11414), .A(n6568), .ZN(n11701) );
  NAND2_X1 U8095 ( .A1(n11701), .A2(n13766), .ZN(n11700) );
  AOI22_X1 U8096 ( .A1(n15566), .A2(n13826), .B1(n13827), .B2(n15545), .ZN(
        n7485) );
  OR2_X1 U8097 ( .A1(n15562), .A2(n15826), .ZN(n15563) );
  NAND2_X1 U8098 ( .A1(n6771), .A2(n8178), .ZN(n11352) );
  INV_X1 U8099 ( .A(n8177), .ZN(n8178) );
  NAND2_X1 U8100 ( .A1(n7543), .A2(n7542), .ZN(n6771) );
  NAND2_X1 U8101 ( .A1(n7544), .A2(n8140), .ZN(n11208) );
  NAND2_X1 U8102 ( .A1(n11295), .A2(n8139), .ZN(n8140) );
  INV_X1 U8103 ( .A(n8110), .ZN(n7544) );
  INV_X1 U8104 ( .A(n13827), .ZN(n15544) );
  AND3_X1 U8105 ( .A1(n13512), .A2(n7237), .A3(n15533), .ZN(n11217) );
  AND2_X1 U8106 ( .A1(n13507), .A2(n13503), .ZN(n12371) );
  NOR2_X1 U8107 ( .A1(n13507), .A2(n7237), .ZN(n11297) );
  NAND2_X1 U8108 ( .A1(n14181), .A2(n13936), .ZN(n10742) );
  AND2_X1 U8109 ( .A1(n8653), .A2(n11018), .ZN(n10734) );
  INV_X1 U8110 ( .A(n13952), .ZN(n13789) );
  NOR2_X1 U8111 ( .A1(n14209), .A2(n7326), .ZN(n7325) );
  AND2_X1 U8112 ( .A1(n14210), .A2(n15525), .ZN(n7326) );
  NAND2_X1 U8113 ( .A1(n8291), .A2(n8290), .ZN(n13590) );
  INV_X1 U8114 ( .A(n15826), .ZN(n15566) );
  INV_X1 U8115 ( .A(n8118), .ZN(n8125) );
  AND2_X1 U8116 ( .A1(n11861), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10298) );
  XNOR2_X1 U8117 ( .A(n8060), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8063) );
  NAND2_X1 U8118 ( .A1(n14357), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8060) );
  AND2_X1 U8119 ( .A1(n7912), .A2(n8032), .ZN(n6795) );
  NOR2_X1 U8120 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n7912) );
  AND4_X1 U8121 ( .A1(n6949), .A2(n8539), .A3(n8031), .A4(n8032), .ZN(n6948)
         );
  AND2_X1 U8122 ( .A1(n8285), .A2(n7913), .ZN(n6946) );
  NAND2_X1 U8123 ( .A1(n8401), .A2(n8400), .ZN(n8556) );
  NAND2_X1 U8124 ( .A1(n6949), .A2(n8163), .ZN(n8346) );
  INV_X1 U8125 ( .A(n7893), .ZN(n7892) );
  OAI21_X1 U8126 ( .B1(n9494), .B2(n11437), .A(n9493), .ZN(n7893) );
  OR2_X1 U8127 ( .A1(n9572), .A2(n9573), .ZN(n7248) );
  NAND2_X1 U8128 ( .A1(n6988), .A2(n6989), .ZN(n10300) );
  AND2_X1 U8129 ( .A1(n6990), .A2(n7214), .ZN(n6988) );
  INV_X1 U8130 ( .A(n10904), .ZN(n7214) );
  AND2_X1 U8131 ( .A1(n6996), .A2(n14390), .ZN(n6995) );
  OR2_X1 U8132 ( .A1(n14461), .A2(n6997), .ZN(n6996) );
  NAND2_X1 U8133 ( .A1(n14404), .A2(n9733), .ZN(n14460) );
  NAND2_X1 U8134 ( .A1(n9736), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9756) );
  INV_X1 U8135 ( .A(n9737), .ZN(n9736) );
  NAND2_X1 U8136 ( .A1(n11589), .A2(n7911), .ZN(n7910) );
  AND2_X1 U8137 ( .A1(n9565), .A2(n9531), .ZN(n7911) );
  OR2_X1 U8138 ( .A1(n9649), .A2(n7906), .ZN(n7905) );
  AND2_X1 U8139 ( .A1(n9650), .A2(n7907), .ZN(n7906) );
  NAND2_X1 U8140 ( .A1(n14380), .A2(n9610), .ZN(n7907) );
  INV_X1 U8141 ( .A(n14438), .ZN(n7901) );
  NOR2_X1 U8142 ( .A1(n7947), .A2(n12397), .ZN(n7220) );
  NAND2_X1 U8143 ( .A1(n6722), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9636) );
  INV_X1 U8144 ( .A(n6722), .ZN(n9634) );
  NAND2_X1 U8145 ( .A1(n10121), .A2(n10123), .ZN(n7748) );
  AND4_X1 U8146 ( .A1(n9519), .A2(n9518), .A3(n9517), .A4(n9516), .ZN(n11983)
         );
  NOR2_X1 U8147 ( .A1(n15173), .A2(n15171), .ZN(n9339) );
  OAI21_X1 U8148 ( .B1(n14568), .B2(n10489), .A(n10472), .ZN(n10536) );
  OR2_X1 U8149 ( .A1(n10643), .A2(n6607), .ZN(n7009) );
  AND2_X1 U8150 ( .A1(n10703), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7337) );
  NAND2_X1 U8151 ( .A1(n7009), .A2(n7008), .ZN(n10700) );
  INV_X1 U8152 ( .A(n10646), .ZN(n7008) );
  NAND2_X1 U8153 ( .A1(n14576), .A2(n6697), .ZN(n11326) );
  OR2_X1 U8154 ( .A1(n14585), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6697) );
  NAND2_X1 U8155 ( .A1(n11718), .A2(n7340), .ZN(n14597) );
  OR2_X1 U8156 ( .A1(n11721), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7340) );
  NOR2_X1 U8157 ( .A1(n14612), .A2(n14594), .ZN(n7014) );
  NAND2_X1 U8158 ( .A1(n9867), .A2(n9866), .ZN(n9939) );
  INV_X1 U8159 ( .A(n15009), .ZN(n14656) );
  NAND2_X1 U8160 ( .A1(n14716), .A2(n14749), .ZN(n14753) );
  OAI21_X1 U8161 ( .B1(n14778), .B2(n7711), .A(n7709), .ZN(n14738) );
  NAND2_X1 U8162 ( .A1(n14714), .A2(n14719), .ZN(n14752) );
  NAND2_X1 U8163 ( .A1(n14757), .A2(n14772), .ZN(n14756) );
  NAND2_X1 U8164 ( .A1(n14758), .A2(n14903), .ZN(n14760) );
  NOR2_X1 U8165 ( .A1(n7728), .A2(n14818), .ZN(n7727) );
  INV_X1 U8166 ( .A(n14682), .ZN(n7728) );
  INV_X1 U8167 ( .A(n14680), .ZN(n7722) );
  NOR2_X1 U8168 ( .A1(n14884), .A2(n7730), .ZN(n7729) );
  INV_X1 U8169 ( .A(n14678), .ZN(n7730) );
  NAND2_X1 U8170 ( .A1(n7143), .A2(n7141), .ZN(n14900) );
  NOR2_X1 U8171 ( .A1(n7142), .A2(n14697), .ZN(n7141) );
  INV_X1 U8172 ( .A(n14677), .ZN(n7142) );
  AND2_X1 U8173 ( .A1(n9845), .A2(n15167), .ZN(n14903) );
  NAND2_X1 U8174 ( .A1(n14676), .A2(n14675), .ZN(n14918) );
  AND2_X1 U8175 ( .A1(n9700), .A2(n9699), .ZN(n14922) );
  INV_X1 U8176 ( .A(n14982), .ZN(n14931) );
  AOI21_X1 U8177 ( .B1(n6929), .B2(n6927), .A(n6926), .ZN(n6925) );
  INV_X1 U8178 ( .A(n6933), .ZN(n6932) );
  OAI21_X1 U8179 ( .B1(n7349), .B2(n12063), .A(n12029), .ZN(n6933) );
  INV_X1 U8180 ( .A(n12043), .ZN(n12046) );
  INV_X1 U8181 ( .A(n7118), .ZN(n7122) );
  NAND2_X1 U8182 ( .A1(n11103), .A2(n11102), .ZN(n11107) );
  NAND2_X1 U8183 ( .A1(n7736), .A2(n9465), .ZN(n11310) );
  INV_X1 U8184 ( .A(n9464), .ZN(n7736) );
  INV_X1 U8185 ( .A(n14903), .ZN(n14980) );
  NAND2_X1 U8186 ( .A1(n9693), .A2(n9692), .ZN(n15076) );
  AND2_X1 U8187 ( .A1(n9410), .A2(n9409), .ZN(n15373) );
  AND2_X1 U8188 ( .A1(n9809), .A2(n9808), .ZN(n10391) );
  XNOR2_X1 U8189 ( .A(n9916), .B(n9915), .ZN(n12454) );
  NAND2_X1 U8190 ( .A1(n9912), .A2(n9911), .ZN(n9916) );
  NOR2_X1 U8191 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n7138) );
  XNOR2_X1 U8192 ( .A(n8524), .B(n8523), .ZN(n12457) );
  NAND2_X1 U8193 ( .A1(n9341), .A2(n9326), .ZN(n9824) );
  NAND2_X1 U8194 ( .A1(n8016), .A2(SI_22_), .ZN(n8460) );
  AND2_X1 U8195 ( .A1(n8443), .A2(n8460), .ZN(n9734) );
  OR2_X1 U8196 ( .A1(n8417), .A2(n7311), .ZN(n8430) );
  NAND2_X1 U8197 ( .A1(n9578), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9597) );
  NAND2_X1 U8198 ( .A1(n7251), .A2(n9495), .ZN(n9520) );
  NAND2_X1 U8199 ( .A1(n8136), .A2(n9431), .ZN(n8119) );
  OR2_X1 U8200 ( .A1(n10381), .A2(n13858), .ZN(n7242) );
  NOR2_X1 U8201 ( .A1(n7460), .A2(n10777), .ZN(n7459) );
  INV_X1 U8202 ( .A(n10771), .ZN(n7460) );
  AND2_X1 U8203 ( .A1(n11281), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n6686) );
  INV_X1 U8204 ( .A(n11287), .ZN(n6687) );
  INV_X1 U8205 ( .A(n11286), .ZN(n6688) );
  AOI21_X1 U8206 ( .B1(n7448), .B2(n7454), .A(n6561), .ZN(n7445) );
  AND2_X1 U8207 ( .A1(n11009), .A2(n11008), .ZN(n7241) );
  NAND2_X1 U8208 ( .A1(n9101), .A2(n9100), .ZN(n12910) );
  NAND2_X1 U8209 ( .A1(n11163), .A2(n11162), .ZN(n11167) );
  INV_X1 U8210 ( .A(n12593), .ZN(n12626) );
  NOR2_X1 U8211 ( .A1(n7406), .A2(n6508), .ZN(n6684) );
  NOR2_X1 U8212 ( .A1(n7404), .A2(n10417), .ZN(n7406) );
  INV_X1 U8213 ( .A(n13036), .ZN(n12618) );
  NAND2_X1 U8214 ( .A1(n7833), .A2(n6560), .ZN(n7203) );
  INV_X1 U8215 ( .A(n7842), .ZN(n7832) );
  NAND2_X1 U8216 ( .A1(n12508), .A2(n12469), .ZN(n12624) );
  NAND2_X1 U8217 ( .A1(n10842), .A2(n15588), .ZN(n12631) );
  AOI21_X1 U8218 ( .B1(n6823), .B2(n7623), .A(n6822), .ZN(n6820) );
  AND2_X1 U8219 ( .A1(n7621), .A2(n7622), .ZN(n6823) );
  NAND2_X1 U8220 ( .A1(n6585), .A2(n12363), .ZN(n6822) );
  NOR2_X1 U8221 ( .A1(n7626), .A2(n7625), .ZN(n7622) );
  NAND2_X1 U8222 ( .A1(n12308), .A2(n6824), .ZN(n6819) );
  NOR2_X1 U8223 ( .A1(n12342), .A2(n12357), .ZN(n6824) );
  NAND2_X1 U8224 ( .A1(n9161), .A2(n9160), .ZN(n12637) );
  INV_X1 U8225 ( .A(n13050), .ZN(n12861) );
  INV_X1 U8226 ( .A(n11996), .ZN(n12999) );
  INV_X1 U8227 ( .A(n13119), .ZN(n12642) );
  NOR2_X1 U8228 ( .A1(n10829), .A2(n12154), .ZN(n12647) );
  OAI211_X1 U8229 ( .C1(n7644), .C2(n10139), .A(n10173), .B(n7643), .ZN(n10172) );
  NAND2_X1 U8230 ( .A1(n7645), .A2(n7646), .ZN(n7644) );
  NAND2_X1 U8231 ( .A1(n10139), .A2(n6531), .ZN(n7643) );
  NAND2_X1 U8232 ( .A1(n10935), .A2(n6497), .ZN(n7389) );
  OAI21_X1 U8233 ( .B1(n6498), .B2(n7386), .A(n7385), .ZN(n11123) );
  INV_X1 U8234 ( .A(n7390), .ZN(n7386) );
  XNOR2_X1 U8235 ( .A(n12747), .B(n12748), .ZN(n6875) );
  NAND2_X1 U8236 ( .A1(n7188), .A2(n6874), .ZN(n6873) );
  NOR2_X1 U8237 ( .A1(n6658), .A2(n7189), .ZN(n7188) );
  NAND2_X1 U8238 ( .A1(n12751), .A2(n12752), .ZN(n6874) );
  INV_X1 U8239 ( .A(n12749), .ZN(n7189) );
  OR2_X1 U8240 ( .A1(n12746), .A2(n7649), .ZN(n7393) );
  NAND2_X1 U8241 ( .A1(n12744), .A2(n7650), .ZN(n7649) );
  NAND2_X1 U8242 ( .A1(n6673), .A2(n7651), .ZN(n7650) );
  AOI21_X1 U8243 ( .B1(n12751), .B2(n12343), .A(n7653), .ZN(n7652) );
  NAND2_X1 U8244 ( .A1(n10197), .A2(n12526), .ZN(n7653) );
  XNOR2_X1 U8245 ( .A(n10194), .B(n10200), .ZN(n7654) );
  NOR2_X1 U8246 ( .A1(n15601), .A2(n11514), .ZN(n13010) );
  INV_X1 U8247 ( .A(n9279), .ZN(n7865) );
  NAND2_X1 U8248 ( .A1(n9192), .A2(n9191), .ZN(n13034) );
  NAND2_X1 U8249 ( .A1(n9165), .A2(n9164), .ZN(n13061) );
  NAND2_X1 U8250 ( .A1(n9117), .A2(n9116), .ZN(n13073) );
  NAND2_X1 U8251 ( .A1(n7407), .A2(n12294), .ZN(n9117) );
  INV_X1 U8252 ( .A(n10965), .ZN(n7407) );
  NAND2_X1 U8253 ( .A1(n9088), .A2(n9087), .ZN(n13088) );
  OR2_X1 U8254 ( .A1(n10564), .A2(n7404), .ZN(n9088) );
  NAND2_X1 U8255 ( .A1(n9041), .A2(n9040), .ZN(n13100) );
  NOR2_X1 U8256 ( .A1(n11396), .A2(n11395), .ZN(n12991) );
  OR2_X1 U8257 ( .A1(n8947), .A2(n8946), .ZN(n13127) );
  NOR2_X1 U8258 ( .A1(n10429), .A2(n7404), .ZN(n8946) );
  OR2_X1 U8259 ( .A1(n12300), .A2(n11529), .ZN(n8867) );
  INV_X1 U8260 ( .A(n15601), .ZN(n15599) );
  NAND2_X1 U8261 ( .A1(n13136), .A2(n15676), .ZN(n7421) );
  INV_X1 U8262 ( .A(n13136), .ZN(n6681) );
  XNOR2_X1 U8263 ( .A(n12786), .B(n12785), .ZN(n13140) );
  NAND2_X1 U8264 ( .A1(n12274), .A2(n12273), .ZN(n13139) );
  NAND2_X1 U8265 ( .A1(n9131), .A2(n9130), .ZN(n13168) );
  NAND2_X1 U8266 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n8802), .ZN(n7201) );
  NAND2_X1 U8267 ( .A1(n8803), .A2(P3_IR_REG_28__SCAN_IN), .ZN(n7202) );
  XNOR2_X1 U8268 ( .A(n8861), .B(n8860), .ZN(n10423) );
  NAND2_X1 U8269 ( .A1(n12448), .A2(n10248), .ZN(n8498) );
  INV_X1 U8270 ( .A(n13581), .ZN(n12099) );
  NOR2_X1 U8271 ( .A1(n7519), .A2(n7934), .ZN(n7518) );
  INV_X1 U8272 ( .A(n11773), .ZN(n7519) );
  NAND2_X1 U8273 ( .A1(n8306), .A2(n8305), .ZN(n14296) );
  NAND2_X1 U8274 ( .A1(n8386), .A2(n8385), .ZN(n13648) );
  NAND2_X1 U8275 ( .A1(n10741), .A2(n15503), .ZN(n13479) );
  OR2_X1 U8276 ( .A1(n13475), .A2(n8530), .ZN(n8069) );
  NAND2_X1 U8277 ( .A1(n10585), .A2(n13846), .ZN(n13845) );
  NAND2_X1 U8278 ( .A1(n13848), .A2(n6683), .ZN(n15458) );
  OR2_X1 U8279 ( .A1(n13851), .A2(n10568), .ZN(n6683) );
  OAI21_X1 U8280 ( .B1(n13935), .B2(n15445), .A(n7292), .ZN(n7291) );
  NAND2_X1 U8281 ( .A1(n13934), .A2(n15470), .ZN(n7292) );
  OAI21_X1 U8282 ( .B1(n7948), .B2(n13938), .A(n13937), .ZN(n7287) );
  AND2_X1 U8283 ( .A1(n6952), .A2(n14181), .ZN(n13939) );
  XNOR2_X1 U8284 ( .A(n6953), .B(n13943), .ZN(n6952) );
  NAND2_X1 U8285 ( .A1(n7301), .A2(n8492), .ZN(n13982) );
  NAND2_X1 U8286 ( .A1(n7330), .A2(n7328), .ZN(n14208) );
  AOI21_X1 U8287 ( .B1(n13811), .B2(n14190), .A(n7329), .ZN(n7328) );
  NAND2_X1 U8288 ( .A1(n7331), .A2(n15556), .ZN(n7330) );
  NOR2_X1 U8289 ( .A1(n13986), .A2(n15495), .ZN(n7329) );
  INV_X1 U8290 ( .A(n8088), .ZN(n8091) );
  NAND2_X1 U8291 ( .A1(n14355), .A2(n10248), .ZN(n10252) );
  OAI21_X1 U8292 ( .B1(n10275), .B2(n6738), .A(n6737), .ZN(n6736) );
  NOR2_X1 U8293 ( .A1(n13960), .A2(n7939), .ZN(n8623) );
  AOI21_X1 U8294 ( .B1(n13951), .B2(n13950), .A(n13789), .ZN(n6735) );
  NOR2_X1 U8295 ( .A1(n10277), .A2(n10276), .ZN(n10279) );
  INV_X1 U8296 ( .A(n13974), .ZN(n14318) );
  OR2_X1 U8297 ( .A1(n13981), .A2(n14310), .ZN(n6808) );
  OR2_X1 U8298 ( .A1(n10323), .A2(n8123), .ZN(n7566) );
  INV_X1 U8299 ( .A(n8100), .ZN(n7567) );
  CLKBUF_X1 U8300 ( .A(n13791), .Z(n11137) );
  INV_X1 U8301 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10314) );
  NAND2_X1 U8302 ( .A1(n9498), .A2(n9497), .ZN(n15389) );
  NAND2_X1 U8303 ( .A1(n14451), .A2(n9595), .ZN(n14379) );
  NAND2_X1 U8304 ( .A1(n9753), .A2(n9752), .ZN(n15051) );
  AND4_X1 U8305 ( .A1(n9387), .A2(n9386), .A3(n9385), .A4(n9384), .ZN(n12071)
         );
  AND2_X1 U8306 ( .A1(n14491), .A2(n14982), .ZN(n14478) );
  NAND2_X1 U8307 ( .A1(n9449), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7701) );
  AND2_X1 U8308 ( .A1(n9712), .A2(n9711), .ZN(n14869) );
  NAND2_X1 U8309 ( .A1(n11930), .A2(n6998), .ZN(n14415) );
  NOR2_X1 U8310 ( .A1(n14413), .A2(n6999), .ZN(n6998) );
  INV_X1 U8311 ( .A(n7248), .ZN(n6999) );
  AND2_X1 U8312 ( .A1(n9799), .A2(n9798), .ZN(n14812) );
  OR2_X1 U8313 ( .A1(n14801), .A2(n9876), .ZN(n9799) );
  NAND2_X1 U8314 ( .A1(n9771), .A2(n9770), .ZN(n15046) );
  INV_X1 U8315 ( .A(n14494), .ZN(n14479) );
  OAI211_X1 U8316 ( .C1(n10320), .C2(n9907), .A(n9453), .B(n9452), .ZN(n10657)
         );
  INV_X1 U8317 ( .A(n14741), .ZN(n14783) );
  NAND2_X1 U8318 ( .A1(n7889), .A2(n7222), .ZN(n7221) );
  NAND2_X1 U8319 ( .A1(n14389), .A2(n7887), .ZN(n7222) );
  INV_X1 U8320 ( .A(n7890), .ZN(n7887) );
  OR2_X1 U8321 ( .A1(n15168), .A2(n9907), .ZN(n9909) );
  NAND2_X1 U8322 ( .A1(n9841), .A2(n9840), .ZN(n14800) );
  INV_X1 U8323 ( .A(n14812), .ZN(n14711) );
  NAND2_X1 U8324 ( .A1(n9762), .A2(n9761), .ZN(n14856) );
  OR2_X1 U8325 ( .A1(n14836), .A2(n9876), .ZN(n9762) );
  OR2_X1 U8326 ( .A1(n9353), .A2(n7183), .ZN(n9503) );
  NAND4_X1 U8327 ( .A1(n9417), .A2(n9416), .A3(n9415), .A4(n9414), .ZN(n14508)
         );
  NAND2_X1 U8328 ( .A1(n6918), .A2(n6917), .ZN(n9435) );
  NAND2_X1 U8329 ( .A1(n9443), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6918) );
  AND3_X1 U8330 ( .A1(n9429), .A2(n9427), .A3(n9428), .ZN(n6917) );
  NAND2_X1 U8331 ( .A1(n10448), .A2(n10447), .ZN(n14551) );
  OAI21_X1 U8332 ( .B1(n10546), .B2(n10541), .A(n10452), .ZN(n10544) );
  NOR2_X1 U8333 ( .A1(n10453), .A2(n10454), .ZN(n10527) );
  NOR2_X1 U8334 ( .A1(n14592), .A2(n14591), .ZN(n14596) );
  INV_X1 U8335 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n14648) );
  AOI21_X1 U8336 ( .B1(n6689), .B2(n15270), .A(n9940), .ZN(n7016) );
  INV_X1 U8337 ( .A(n7334), .ZN(n6689) );
  NAND2_X1 U8338 ( .A1(n7333), .A2(n6677), .ZN(n7018) );
  INV_X1 U8339 ( .A(n6678), .ZN(n6677) );
  NAND2_X1 U8340 ( .A1(n7334), .A2(n15270), .ZN(n7333) );
  OAI21_X1 U8341 ( .B1(n14646), .B2(n11724), .A(n7335), .ZN(n6678) );
  NAND2_X1 U8342 ( .A1(n9523), .A2(n9522), .ZN(n15397) );
  AND2_X1 U8343 ( .A1(n9402), .A2(n9401), .ZN(n11250) );
  OAI21_X1 U8344 ( .B1(n7709), .B2(n6728), .A(n6576), .ZN(n6727) );
  OAI21_X1 U8345 ( .B1(n14724), .B2(n15422), .A(n15015), .ZN(n6916) );
  INV_X2 U8346 ( .A(n15424), .ZN(n15425) );
  NAND3_X1 U8347 ( .A1(n9309), .A2(n6453), .A3(n6452), .ZN(n9347) );
  NAND2_X1 U8348 ( .A1(n10390), .A2(n7457), .ZN(n7164) );
  NAND2_X1 U8349 ( .A1(n15234), .A2(n15233), .ZN(n15239) );
  NAND3_X1 U8350 ( .A1(n7162), .A2(n15225), .A3(n7161), .ZN(n15234) );
  INV_X1 U8351 ( .A(n15231), .ZN(n7161) );
  MUX2_X1 U8352 ( .A(n9990), .B(n9989), .S(n10991), .Z(n9991) );
  NAND2_X1 U8353 ( .A1(n10001), .A2(n6521), .ZN(n7741) );
  INV_X1 U8354 ( .A(n10003), .ZN(n7739) );
  NAND2_X1 U8355 ( .A1(n7226), .A2(n13529), .ZN(n13538) );
  INV_X1 U8356 ( .A(n10007), .ZN(n10008) );
  OR2_X1 U8357 ( .A1(n10019), .A2(n7752), .ZN(n7750) );
  INV_X1 U8358 ( .A(n10018), .ZN(n7752) );
  OR2_X1 U8359 ( .A1(n13544), .A2(n13546), .ZN(n7225) );
  NAND2_X1 U8360 ( .A1(n6870), .A2(n12172), .ZN(n6869) );
  NAND2_X1 U8361 ( .A1(n6582), .A2(n12269), .ZN(n7618) );
  OR2_X1 U8362 ( .A1(n12170), .A2(n15590), .ZN(n7620) );
  AND2_X1 U8363 ( .A1(n7618), .A2(n7619), .ZN(n6868) );
  NAND2_X1 U8364 ( .A1(n7617), .A2(n12269), .ZN(n7616) );
  INV_X1 U8365 ( .A(n12174), .ZN(n7617) );
  OAI21_X1 U8366 ( .B1(n7751), .B2(n6574), .A(n7027), .ZN(n7033) );
  OR2_X1 U8367 ( .A1(n13556), .A2(n7480), .ZN(n7479) );
  NAND2_X1 U8368 ( .A1(n6717), .A2(n6716), .ZN(n7169) );
  INV_X1 U8369 ( .A(n13555), .ZN(n7480) );
  AOI211_X1 U8370 ( .C1(n12186), .C2(n12185), .A(n12184), .B(n12183), .ZN(
        n12193) );
  OAI21_X1 U8371 ( .B1(n10072), .B2(n10071), .A(n10070), .ZN(n10081) );
  NAND2_X1 U8372 ( .A1(n15071), .A2(n10082), .ZN(n10084) );
  NAND2_X1 U8373 ( .A1(n6814), .A2(n12214), .ZN(n6813) );
  OAI21_X1 U8374 ( .B1(n12207), .B2(n6816), .A(n6815), .ZN(n6814) );
  INV_X1 U8375 ( .A(n12215), .ZN(n6815) );
  NAND2_X1 U8376 ( .A1(n6712), .A2(n6711), .ZN(n13588) );
  AOI21_X1 U8377 ( .B1(n6463), .B2(n7484), .A(n6578), .ZN(n6711) );
  AND2_X1 U8378 ( .A1(n6506), .A2(n13577), .ZN(n7484) );
  OR2_X1 U8379 ( .A1(n13638), .A2(n13610), .ZN(n13623) );
  AOI21_X1 U8380 ( .B1(n6812), .B2(n6810), .A(n12952), .ZN(n12225) );
  NOR2_X1 U8381 ( .A1(n6811), .A2(n12966), .ZN(n6810) );
  NAND2_X1 U8382 ( .A1(n6813), .A2(n6695), .ZN(n6812) );
  INV_X1 U8383 ( .A(n12218), .ZN(n6811) );
  AOI21_X1 U8384 ( .B1(n7611), .B2(n6514), .A(n12884), .ZN(n6864) );
  NAND2_X1 U8385 ( .A1(n7043), .A2(n7042), .ZN(n10098) );
  AOI21_X1 U8386 ( .B1(n6451), .B2(n7046), .A(n6472), .ZN(n7042) );
  AOI21_X1 U8387 ( .B1(n7469), .B2(n7471), .A(n7468), .ZN(n7467) );
  INV_X1 U8388 ( .A(n13654), .ZN(n7468) );
  NAND2_X1 U8389 ( .A1(n7105), .A2(n7103), .ZN(n7099) );
  INV_X1 U8390 ( .A(n7105), .ZN(n8011) );
  NOR2_X1 U8391 ( .A1(n7583), .A2(n6507), .ZN(n7582) );
  INV_X1 U8392 ( .A(n7588), .ZN(n7583) );
  AOI21_X1 U8393 ( .B1(n6860), .B2(n6862), .A(n6584), .ZN(n6859) );
  NOR2_X1 U8394 ( .A1(n12859), .A2(n7609), .ZN(n7608) );
  INV_X1 U8395 ( .A(n12249), .ZN(n7609) );
  INV_X1 U8396 ( .A(n12252), .ZN(n7606) );
  NAND2_X1 U8397 ( .A1(n7037), .A2(n10987), .ZN(n7036) );
  INV_X1 U8398 ( .A(n9941), .ZN(n7037) );
  NOR2_X1 U8399 ( .A1(n8014), .A2(n10964), .ZN(n7588) );
  INV_X1 U8400 ( .A(n8432), .ZN(n8014) );
  OR2_X1 U8401 ( .A1(n8002), .A2(n7081), .ZN(n7080) );
  NAND4_X1 U8402 ( .A1(n6696), .A2(n6695), .A3(n6694), .A4(n6450), .ZN(n12334)
         );
  INV_X1 U8403 ( .A(n12887), .ZN(n6693) );
  OR2_X1 U8404 ( .A1(n9242), .A2(n12966), .ZN(n9244) );
  INV_X1 U8405 ( .A(n12321), .ZN(n12322) );
  INV_X1 U8406 ( .A(n8761), .ZN(n7675) );
  INV_X1 U8407 ( .A(n7674), .ZN(n7673) );
  OAI21_X1 U8408 ( .B1(n8964), .B2(n7675), .A(n8979), .ZN(n7674) );
  INV_X1 U8409 ( .A(n8756), .ZN(n6898) );
  INV_X1 U8410 ( .A(n13669), .ZN(n7168) );
  NAND2_X1 U8411 ( .A1(n13790), .A2(n7208), .ZN(n7199) );
  INV_X1 U8412 ( .A(n13731), .ZN(n7208) );
  OAI22_X1 U8413 ( .A1(n13729), .A2(n13728), .B1(n13727), .B2(n13726), .ZN(
        n13731) );
  AND2_X1 U8414 ( .A1(n6505), .A2(n8598), .ZN(n6766) );
  AND2_X1 U8415 ( .A1(n15485), .A2(n7488), .ZN(n15487) );
  NAND2_X1 U8416 ( .A1(n7049), .A2(n7048), .ZN(n10115) );
  AOI21_X1 U8417 ( .B1(n6465), .B2(n7052), .A(n6566), .ZN(n7048) );
  CLKBUF_X1 U8418 ( .A(n10085), .Z(n10082) );
  INV_X1 U8419 ( .A(n12014), .ZN(n7706) );
  INV_X1 U8420 ( .A(n8494), .ZN(n7601) );
  NAND2_X1 U8421 ( .A1(n8431), .A2(n6547), .ZN(n7102) );
  NAND2_X1 U8422 ( .A1(n8007), .A2(n8006), .ZN(n7319) );
  INV_X1 U8423 ( .A(n7994), .ZN(n7598) );
  INV_X1 U8424 ( .A(n7987), .ZN(n7094) );
  NAND2_X1 U8425 ( .A1(n7984), .A2(n10416), .ZN(n7987) );
  OAI21_X1 U8426 ( .B1(n6443), .B2(n10326), .A(n7207), .ZN(n7961) );
  NAND2_X1 U8427 ( .A1(n6443), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7207) );
  INV_X1 U8428 ( .A(n12498), .ZN(n7836) );
  OR2_X1 U8429 ( .A1(n12615), .A2(n7842), .ZN(n7841) );
  INV_X1 U8430 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n15804) );
  OAI211_X1 U8431 ( .C1(n12262), .C2(n6846), .A(n6844), .B(n6842), .ZN(n12268)
         );
  NOR2_X1 U8432 ( .A1(n6848), .A2(n6847), .ZN(n6846) );
  NAND2_X1 U8433 ( .A1(n6588), .A2(n6848), .ZN(n6844) );
  NAND2_X1 U8434 ( .A1(n7440), .A2(n10814), .ZN(n10818) );
  NAND2_X1 U8435 ( .A1(n10179), .A2(n10178), .ZN(n10811) );
  NAND2_X1 U8436 ( .A1(n6980), .A2(n11126), .ZN(n6978) );
  INV_X1 U8437 ( .A(n7434), .ZN(n7433) );
  NOR2_X1 U8438 ( .A1(n7435), .A2(n11539), .ZN(n6980) );
  NAND2_X1 U8439 ( .A1(n10221), .A2(n11198), .ZN(n7384) );
  INV_X1 U8440 ( .A(n11610), .ZN(n6985) );
  NAND2_X1 U8441 ( .A1(n6473), .A2(n6668), .ZN(n7376) );
  INV_X1 U8442 ( .A(n11459), .ZN(n7378) );
  NAND2_X1 U8443 ( .A1(n6826), .A2(n6825), .ZN(n10187) );
  INV_X1 U8444 ( .A(n6827), .ZN(n6826) );
  OAI21_X1 U8445 ( .B1(n7255), .B2(n10186), .A(n6647), .ZN(n6827) );
  INV_X1 U8446 ( .A(n6836), .ZN(n6834) );
  NAND2_X1 U8447 ( .A1(n12669), .A2(n10235), .ZN(n10192) );
  NAND2_X1 U8448 ( .A1(n12674), .A2(n10237), .ZN(n10238) );
  INV_X1 U8449 ( .A(n10242), .ZN(n7370) );
  NOR2_X1 U8450 ( .A1(n7369), .A2(n12716), .ZN(n7361) );
  NAND2_X1 U8451 ( .A1(n7639), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n7638) );
  NAND2_X1 U8452 ( .A1(n9206), .A2(n9205), .ZN(n9214) );
  OR2_X1 U8453 ( .A1(n13034), .A2(n13043), .ZN(n12260) );
  NAND2_X1 U8454 ( .A1(n7170), .A2(n9155), .ZN(n9182) );
  NOR2_X1 U8455 ( .A1(n9027), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7272) );
  NAND2_X1 U8456 ( .A1(n9233), .A2(n7401), .ZN(n7397) );
  AND2_X1 U8457 ( .A1(n9230), .A2(n12320), .ZN(n7417) );
  INV_X1 U8458 ( .A(n10849), .ZN(n12163) );
  NAND2_X1 U8459 ( .A1(n12887), .A2(n12241), .ZN(n7883) );
  OR2_X1 U8460 ( .A1(n12910), .A2(n12638), .ZN(n12237) );
  NAND2_X1 U8461 ( .A1(n11920), .A2(n9235), .ZN(n7786) );
  NOR2_X1 U8462 ( .A1(n12205), .A2(n7874), .ZN(n7873) );
  INV_X1 U8463 ( .A(n12200), .ZN(n7874) );
  OR2_X1 U8464 ( .A1(n12316), .A2(n8728), .ZN(n8816) );
  INV_X1 U8465 ( .A(n8799), .ZN(n7686) );
  INV_X1 U8466 ( .A(n7688), .ZN(n7683) );
  AOI21_X1 U8467 ( .B1(n7665), .B2(n7667), .A(n7663), .ZN(n7662) );
  INV_X1 U8468 ( .A(n6904), .ZN(n6903) );
  OAI21_X1 U8469 ( .B1(n7670), .B2(n8992), .A(n7657), .ZN(n6904) );
  NAND2_X1 U8470 ( .A1(n6903), .A2(n8992), .ZN(n6901) );
  INV_X1 U8471 ( .A(n8766), .ZN(n7660) );
  AOI21_X1 U8472 ( .B1(n7673), .B2(n7675), .A(n7671), .ZN(n7670) );
  INV_X1 U8473 ( .A(n8763), .ZN(n7671) );
  NOR2_X1 U8474 ( .A1(n6898), .A2(n6895), .ZN(n6894) );
  INV_X1 U8475 ( .A(n8754), .ZN(n6895) );
  OAI21_X1 U8476 ( .B1(n8942), .B2(n6898), .A(n8949), .ZN(n6897) );
  OAI21_X1 U8477 ( .B1(n8744), .B2(n6892), .A(n8747), .ZN(n6891) );
  INV_X1 U8478 ( .A(n6891), .ZN(n6889) );
  NAND2_X1 U8479 ( .A1(n6976), .A2(n8860), .ZN(n8907) );
  INV_X1 U8480 ( .A(n8859), .ZN(n6976) );
  NAND2_X1 U8481 ( .A1(n10313), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8737) );
  AOI21_X1 U8482 ( .B1(n11683), .B2(n11621), .A(n11617), .ZN(n11619) );
  OR2_X1 U8483 ( .A1(n13725), .A2(n13724), .ZN(n7579) );
  OR2_X1 U8484 ( .A1(n13670), .A2(n13682), .ZN(n6726) );
  INV_X1 U8485 ( .A(n7196), .ZN(n8324) );
  OR2_X1 U8486 ( .A1(n13720), .A2(n13719), .ZN(n8612) );
  NOR2_X1 U8487 ( .A1(n14217), .A2(n14047), .ZN(n6956) );
  INV_X1 U8488 ( .A(n8597), .ZN(n7505) );
  AOI21_X1 U8489 ( .B1(n6790), .B2(n6792), .A(n6553), .ZN(n6789) );
  NAND2_X1 U8490 ( .A1(n7196), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8356) );
  NOR2_X1 U8491 ( .A1(n14166), .A2(n14184), .ZN(n7925) );
  NOR2_X1 U8492 ( .A1(n7491), .A2(n6773), .ZN(n6772) );
  INV_X1 U8493 ( .A(n6775), .ZN(n6773) );
  INV_X1 U8494 ( .A(n7492), .ZN(n7491) );
  AND2_X1 U8495 ( .A1(n7493), .A2(n13772), .ZN(n7492) );
  NAND2_X1 U8496 ( .A1(n8576), .A2(n8575), .ZN(n7493) );
  NAND2_X1 U8497 ( .A1(n6485), .A2(n7299), .ZN(n7295) );
  NAND2_X1 U8498 ( .A1(n11177), .A2(n11178), .ZN(n11176) );
  OR2_X1 U8499 ( .A1(n10250), .A2(n10316), .ZN(n8152) );
  OR2_X1 U8500 ( .A1(n8262), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n8270) );
  OR2_X1 U8501 ( .A1(n8346), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n8213) );
  NAND2_X1 U8502 ( .A1(n7897), .A2(n7896), .ZN(n7895) );
  INV_X1 U8503 ( .A(n11431), .ZN(n7897) );
  INV_X1 U8504 ( .A(n9467), .ZN(n6731) );
  NOR2_X1 U8505 ( .A1(n9538), .A2(n9537), .ZN(n6730) );
  NOR2_X1 U8506 ( .A1(n9602), .A2(n11344), .ZN(n6722) );
  AND3_X1 U8507 ( .A1(n9963), .A2(n14772), .A3(n6509), .ZN(n9936) );
  AOI22_X1 U8508 ( .A1(n12422), .A2(n14994), .B1(n9436), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n9437) );
  NAND2_X1 U8509 ( .A1(n7129), .A2(n14793), .ZN(n7128) );
  AND2_X1 U8510 ( .A1(n6532), .A2(n14700), .ZN(n14701) );
  NAND2_X1 U8511 ( .A1(n7704), .A2(n7134), .ZN(n7133) );
  INV_X1 U8512 ( .A(n7704), .ZN(n7135) );
  NOR2_X1 U8513 ( .A1(n14692), .A2(n15103), .ZN(n7756) );
  INV_X1 U8514 ( .A(n7929), .ZN(n7696) );
  INV_X1 U8515 ( .A(n14663), .ZN(n7707) );
  NAND2_X1 U8516 ( .A1(n14666), .A2(n14665), .ZN(n12031) );
  NOR2_X1 U8517 ( .A1(n7352), .A2(n12063), .ZN(n6935) );
  NAND2_X1 U8518 ( .A1(n6730), .A2(n9349), .ZN(n9382) );
  AND2_X1 U8519 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_REG3_REG_11__SCAN_IN), 
        .ZN(n9349) );
  INV_X1 U8520 ( .A(n11240), .ZN(n7725) );
  NAND2_X1 U8521 ( .A1(n6731), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9413) );
  XNOR2_X1 U8522 ( .A(n7698), .B(n14512), .ZN(n11066) );
  INV_X1 U8523 ( .A(n10973), .ZN(n9943) );
  OR2_X1 U8524 ( .A1(n14885), .A2(n15066), .ZN(n14871) );
  INV_X1 U8525 ( .A(n7760), .ZN(n7759) );
  AND2_X1 U8526 ( .A1(n11050), .A2(n11513), .ZN(n9942) );
  AND2_X1 U8527 ( .A1(n7576), .A2(n7089), .ZN(n7084) );
  INV_X1 U8528 ( .A(n7575), .ZN(n7085) );
  INV_X1 U8529 ( .A(n8070), .ZN(n7089) );
  NOR2_X1 U8530 ( .A1(n8025), .A2(SI_25_), .ZN(n7087) );
  INV_X1 U8531 ( .A(n9824), .ZN(n9360) );
  NOR2_X1 U8532 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n9359) );
  NAND2_X1 U8533 ( .A1(n9369), .A2(n9612), .ZN(n7041) );
  INV_X1 U8534 ( .A(n7983), .ZN(n7569) );
  OAI21_X1 U8535 ( .B1(n6443), .B2(n10317), .A(n7205), .ZN(n8148) );
  NAND2_X1 U8536 ( .A1(n6442), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7205) );
  NAND2_X1 U8537 ( .A1(n11739), .A2(n11740), .ZN(n11973) );
  AOI21_X1 U8538 ( .B1(n7453), .B2(n7451), .A(n7449), .ZN(n7448) );
  INV_X1 U8539 ( .A(n11730), .ZN(n7449) );
  NAND2_X1 U8540 ( .A1(n11973), .A2(n11972), .ZN(n15189) );
  INV_X1 U8541 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n8912) );
  INV_X1 U8542 ( .A(n7170), .ZN(n9168) );
  XNOR2_X1 U8543 ( .A(n12463), .B(n15615), .ZN(n11160) );
  AND4_X1 U8544 ( .A1(n11794), .A2(n11796), .A3(n11638), .A4(n11637), .ZN(
        n11639) );
  NAND2_X1 U8545 ( .A1(n7810), .A2(n11651), .ZN(n11749) );
  INV_X1 U8546 ( .A(n7825), .ZN(n7824) );
  NAND2_X1 U8547 ( .A1(n7823), .A2(n7825), .ZN(n7822) );
  INV_X1 U8548 ( .A(n7827), .ZN(n7823) );
  XNOR2_X1 U8549 ( .A(n10845), .B(n12494), .ZN(n6764) );
  XNOR2_X1 U8550 ( .A(n12463), .B(n15585), .ZN(n11007) );
  NAND2_X1 U8551 ( .A1(n6799), .A2(n12479), .ZN(n12605) );
  INV_X1 U8552 ( .A(n12607), .ZN(n6799) );
  NAND2_X1 U8553 ( .A1(n8877), .A2(n8876), .ZN(n8898) );
  INV_X1 U8554 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8876) );
  INV_X1 U8555 ( .A(n8878), .ZN(n8877) );
  NAND2_X1 U8556 ( .A1(n7270), .A2(n7269), .ZN(n8913) );
  INV_X1 U8557 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n7269) );
  INV_X1 U8558 ( .A(n8898), .ZN(n7270) );
  INV_X1 U8559 ( .A(n10835), .ZN(n12365) );
  AND2_X1 U8560 ( .A1(n12310), .A2(n6601), .ZN(n7661) );
  NAND2_X1 U8561 ( .A1(n12821), .A2(n7259), .ZN(n7258) );
  INV_X1 U8562 ( .A(n12312), .ZN(n7626) );
  NAND2_X1 U8563 ( .A1(n12341), .A2(n12349), .ZN(n7625) );
  OAI21_X1 U8564 ( .B1(n12342), .B2(n12314), .A(n12313), .ZN(n12318) );
  INV_X1 U8565 ( .A(n12311), .ZN(n12314) );
  NAND2_X1 U8566 ( .A1(n12270), .A2(n7235), .ZN(n7621) );
  NOR2_X1 U8567 ( .A1(n12275), .A2(n7236), .ZN(n7235) );
  INV_X1 U8568 ( .A(n12268), .ZN(n12270) );
  NAND2_X1 U8569 ( .A1(n12536), .A2(n12269), .ZN(n7236) );
  AND2_X1 U8570 ( .A1(n12306), .A2(n12305), .ZN(n12352) );
  NAND2_X1 U8571 ( .A1(n7776), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7775) );
  NAND2_X1 U8572 ( .A1(n7438), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10174) );
  INV_X1 U8573 ( .A(n7632), .ZN(n10813) );
  XNOR2_X1 U8574 ( .A(n10146), .B(n6979), .ZN(n11126) );
  NAND2_X1 U8575 ( .A1(n10213), .A2(n10825), .ZN(n7390) );
  NAND2_X1 U8576 ( .A1(n11126), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n11125) );
  XNOR2_X1 U8577 ( .A(n7437), .B(n7436), .ZN(n11035) );
  NAND2_X1 U8578 ( .A1(n6851), .A2(n6850), .ZN(n7641) );
  AOI21_X1 U8579 ( .B1(n7630), .B2(n6852), .A(n6580), .ZN(n6851) );
  NAND2_X1 U8580 ( .A1(n11124), .A2(n6853), .ZN(n6850) );
  OR2_X1 U8581 ( .A1(n7382), .A2(n7381), .ZN(n7380) );
  INV_X1 U8582 ( .A(n7384), .ZN(n7381) );
  AOI21_X1 U8583 ( .B1(n11033), .B2(n6455), .A(n7383), .ZN(n7382) );
  INV_X1 U8584 ( .A(n11192), .ZN(n7383) );
  NOR2_X1 U8585 ( .A1(n7427), .A2(n11466), .ZN(n7426) );
  NAND2_X1 U8586 ( .A1(n10150), .A2(n6985), .ZN(n6983) );
  NAND2_X1 U8587 ( .A1(n7375), .A2(n7373), .ZN(n11601) );
  NOR2_X1 U8588 ( .A1(n7376), .A2(n7374), .ZN(n7373) );
  INV_X1 U8589 ( .A(n11603), .ZN(n7374) );
  AND2_X1 U8590 ( .A1(n7375), .A2(n7372), .ZN(n11602) );
  INV_X1 U8591 ( .A(n7376), .ZN(n7372) );
  XNOR2_X1 U8592 ( .A(n10187), .B(n11783), .ZN(n11789) );
  NAND2_X1 U8593 ( .A1(n6646), .A2(n11840), .ZN(n11842) );
  NAND2_X1 U8594 ( .A1(n12653), .A2(n6641), .ZN(n12673) );
  NAND2_X1 U8595 ( .A1(n12673), .A2(n7371), .ZN(n12674) );
  AND2_X1 U8596 ( .A1(n12676), .A2(n12672), .ZN(n7371) );
  NAND2_X1 U8597 ( .A1(n7441), .A2(n12665), .ZN(n12663) );
  NAND2_X1 U8598 ( .A1(n12649), .A2(n10190), .ZN(n12670) );
  NAND2_X1 U8599 ( .A1(n11845), .A2(n7629), .ZN(n10189) );
  NAND2_X1 U8600 ( .A1(n12670), .A2(n12671), .ZN(n12669) );
  XNOR2_X1 U8601 ( .A(n10192), .B(n10157), .ZN(n12690) );
  INV_X1 U8602 ( .A(n7637), .ZN(n7636) );
  NAND2_X1 U8603 ( .A1(n7655), .A2(n10164), .ZN(n7651) );
  INV_X1 U8604 ( .A(n12791), .ZN(n9269) );
  NAND2_X1 U8605 ( .A1(n7849), .A2(n12259), .ZN(n6885) );
  AND2_X1 U8606 ( .A1(n12260), .A2(n12263), .ZN(n12815) );
  AOI21_X1 U8607 ( .B1(n7412), .B2(n7411), .A(n6563), .ZN(n7410) );
  INV_X1 U8608 ( .A(n7272), .ZN(n9042) );
  INV_X1 U8609 ( .A(n8958), .ZN(n8957) );
  NAND2_X1 U8610 ( .A1(n7268), .A2(n8912), .ZN(n8931) );
  INV_X1 U8611 ( .A(n8913), .ZN(n7268) );
  NAND2_X1 U8612 ( .A1(n6705), .A2(n6704), .ZN(n8958) );
  INV_X1 U8613 ( .A(n8931), .ZN(n6705) );
  INV_X1 U8614 ( .A(n11450), .ZN(n7419) );
  INV_X1 U8615 ( .A(n12327), .ZN(n11526) );
  NAND2_X1 U8616 ( .A1(n12163), .A2(n12368), .ZN(n12267) );
  NAND2_X1 U8617 ( .A1(n9152), .A2(n12250), .ZN(n12829) );
  NAND2_X1 U8618 ( .A1(n12237), .A2(n12238), .ZN(n12900) );
  NAND2_X1 U8619 ( .A1(n9241), .A2(n9240), .ZN(n12962) );
  AOI21_X1 U8620 ( .B1(n7871), .B2(n7873), .A(n7870), .ZN(n7869) );
  INV_X1 U8621 ( .A(n7873), .ZN(n7872) );
  INV_X1 U8622 ( .A(n7876), .ZN(n7871) );
  NAND2_X1 U8623 ( .A1(n7782), .A2(n7400), .ZN(n12118) );
  NAND2_X1 U8624 ( .A1(n11919), .A2(n9236), .ZN(n12119) );
  NAND2_X1 U8625 ( .A1(n9233), .A2(n7402), .ZN(n7400) );
  AND2_X1 U8626 ( .A1(n11956), .A2(n9235), .ZN(n11921) );
  NAND2_X1 U8627 ( .A1(n8874), .A2(n8873), .ZN(n7424) );
  INV_X1 U8628 ( .A(n15651), .ZN(n15637) );
  OR2_X1 U8629 ( .A1(n10966), .A2(n10840), .ZN(n10835) );
  NOR2_X1 U8630 ( .A1(n9285), .A2(n9290), .ZN(n10859) );
  NOR2_X1 U8631 ( .A1(n9291), .A2(n9290), .ZN(n10862) );
  NAND2_X1 U8632 ( .A1(n8708), .A2(n8707), .ZN(n11391) );
  OAI21_X1 U8633 ( .B1(n8798), .B2(n7684), .A(n7682), .ZN(n12279) );
  INV_X1 U8634 ( .A(n7685), .ZN(n7684) );
  AOI21_X1 U8635 ( .B1(n7683), .B2(n7685), .A(n6672), .ZN(n7682) );
  NOR2_X1 U8636 ( .A1(n12271), .A2(n7686), .ZN(n7685) );
  INV_X1 U8637 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7394) );
  INV_X1 U8638 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8694) );
  AND2_X1 U8639 ( .A1(n7817), .A2(n7816), .ZN(n7815) );
  INV_X1 U8640 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7816) );
  NAND2_X1 U8641 ( .A1(n9067), .A2(n7817), .ZN(n8685) );
  NAND2_X1 U8642 ( .A1(n7171), .A2(n12446), .ZN(n6899) );
  NAND2_X1 U8643 ( .A1(n7812), .A2(n7813), .ZN(n8693) );
  NAND2_X1 U8644 ( .A1(n8907), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8889) );
  INV_X1 U8645 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8888) );
  XNOR2_X1 U8646 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .ZN(n6876) );
  NAND2_X1 U8647 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n8838) );
  NAND2_X1 U8648 ( .A1(n7540), .A2(n7538), .ZN(n13329) );
  NOR2_X1 U8649 ( .A1(n13332), .A2(n7539), .ZN(n7538) );
  INV_X1 U8650 ( .A(n13268), .ZN(n7539) );
  NOR2_X1 U8651 ( .A1(n13357), .A2(n7074), .ZN(n7073) );
  INV_X1 U8652 ( .A(n7076), .ZN(n7074) );
  NAND2_X1 U8653 ( .A1(n13288), .A2(n7077), .ZN(n7076) );
  INV_X1 U8654 ( .A(n13289), .ZN(n7077) );
  OR2_X1 U8655 ( .A1(n13457), .A2(n13458), .ZN(n7075) );
  AND2_X1 U8656 ( .A1(n13365), .A2(n7946), .ZN(n13366) );
  NOR2_X1 U8657 ( .A1(n12132), .A2(n7064), .ZN(n7063) );
  INV_X1 U8658 ( .A(n11881), .ZN(n7064) );
  INV_X1 U8659 ( .A(n8293), .ZN(n8048) );
  AND2_X1 U8660 ( .A1(n13489), .A2(n13483), .ZN(n13404) );
  NOR2_X1 U8661 ( .A1(n11473), .A2(n13412), .ZN(n7245) );
  INV_X1 U8662 ( .A(n7930), .ZN(n7054) );
  NOR2_X1 U8663 ( .A1(n11472), .A2(n11471), .ZN(n13412) );
  AOI21_X1 U8664 ( .B1(n7526), .B2(n7528), .A(n6522), .ZN(n7525) );
  NAND2_X1 U8665 ( .A1(n8050), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8407) );
  AND2_X1 U8666 ( .A1(n13280), .A2(n13483), .ZN(n7541) );
  XNOR2_X1 U8667 ( .A(n14210), .B(n13314), .ZN(n13316) );
  NAND2_X1 U8668 ( .A1(n13316), .A2(n13315), .ZN(n13368) );
  OR2_X1 U8669 ( .A1(n13320), .A2(n13396), .ZN(n13468) );
  NOR2_X1 U8670 ( .A1(n7533), .A2(n13301), .ZN(n7529) );
  NAND2_X1 U8671 ( .A1(n8531), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6754) );
  NAND2_X1 U8672 ( .A1(n8208), .A2(n6544), .ZN(n6751) );
  NAND2_X1 U8673 ( .A1(n13836), .A2(n13837), .ZN(n13835) );
  OAI21_X1 U8674 ( .B1(n13866), .B2(n10674), .A(n7303), .ZN(n7302) );
  NOR2_X1 U8675 ( .A1(n10571), .A2(n6513), .ZN(n7303) );
  OAI22_X1 U8676 ( .A1(n10719), .A2(n10718), .B1(n10720), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n10785) );
  OR2_X1 U8677 ( .A1(n8346), .A2(n8347), .ZN(n8288) );
  AND2_X1 U8678 ( .A1(n11380), .A2(n11670), .ZN(n11382) );
  OAI22_X1 U8679 ( .A1(n13895), .A2(n13894), .B1(n13893), .B2(n13892), .ZN(
        n13917) );
  NOR2_X1 U8680 ( .A1(n6968), .A2(n13927), .ZN(n6967) );
  INV_X1 U8681 ( .A(n13909), .ZN(n6968) );
  NOR2_X1 U8682 ( .A1(n6951), .A2(n13946), .ZN(n6950) );
  INV_X1 U8683 ( .A(n7915), .ZN(n6951) );
  INV_X1 U8684 ( .A(n13809), .ZN(n10268) );
  NAND2_X1 U8685 ( .A1(n10285), .A2(n8609), .ZN(n10267) );
  NOR2_X1 U8686 ( .A1(n13786), .A2(n10264), .ZN(n8609) );
  AND2_X1 U8687 ( .A1(n8528), .A2(n8501), .ZN(n13973) );
  OR2_X1 U8688 ( .A1(n10284), .A2(n10283), .ZN(n7935) );
  NAND2_X1 U8689 ( .A1(n13810), .A2(n14190), .ZN(n10287) );
  INV_X1 U8690 ( .A(n7501), .ZN(n13984) );
  AND2_X1 U8691 ( .A1(n7496), .A2(n7502), .ZN(n14001) );
  OR2_X1 U8692 ( .A1(n14019), .A2(n14020), .ZN(n14021) );
  NAND2_X1 U8693 ( .A1(n14058), .A2(n14227), .ZN(n14038) );
  INV_X1 U8694 ( .A(n7919), .ZN(n14085) );
  AND2_X1 U8695 ( .A1(n14193), .A2(n7922), .ZN(n14126) );
  AND2_X1 U8696 ( .A1(n6461), .A2(n7923), .ZN(n7922) );
  NAND2_X1 U8697 ( .A1(n14193), .A2(n6461), .ZN(n14146) );
  NAND2_X1 U8698 ( .A1(n8049), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8375) );
  INV_X1 U8699 ( .A(n8358), .ZN(n8049) );
  NOR2_X1 U8700 ( .A1(n13585), .A2(n13590), .ZN(n6957) );
  INV_X1 U8701 ( .A(n8254), .ZN(n7195) );
  NAND2_X1 U8702 ( .A1(n8047), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8231) );
  INV_X1 U8703 ( .A(n8229), .ZN(n8047) );
  INV_X1 U8704 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8221) );
  AND2_X1 U8705 ( .A1(n11415), .A2(n6516), .ZN(n11873) );
  NAND2_X1 U8706 ( .A1(n11415), .A2(n11588), .ZN(n11695) );
  NAND2_X1 U8707 ( .A1(n11415), .A2(n6467), .ZN(n11763) );
  NAND2_X1 U8708 ( .A1(n11414), .A2(n11413), .ZN(n7297) );
  NAND2_X1 U8709 ( .A1(n6755), .A2(n6753), .ZN(n6752) );
  AOI22_X1 U8710 ( .A1(n8403), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n10576), .B2(
        n10612), .ZN(n6753) );
  OAI211_X1 U8711 ( .C1(n6752), .C2(n13824), .A(n6750), .B(n6748), .ZN(n8571)
         );
  NAND2_X1 U8712 ( .A1(n6752), .A2(n6751), .ZN(n6750) );
  NAND2_X1 U8713 ( .A1(n6752), .A2(n6749), .ZN(n6748) );
  INV_X1 U8714 ( .A(n6754), .ZN(n6749) );
  INV_X1 U8715 ( .A(n8571), .ZN(n11414) );
  NAND2_X1 U8716 ( .A1(n7178), .A2(n15545), .ZN(n15562) );
  INV_X1 U8717 ( .A(n8566), .ZN(n11210) );
  NAND2_X1 U8718 ( .A1(n8138), .A2(n11025), .ZN(n11295) );
  AND2_X1 U8719 ( .A1(n8562), .A2(n14271), .ZN(n6737) );
  NAND2_X1 U8720 ( .A1(n13789), .A2(n13950), .ZN(n6738) );
  NAND2_X1 U8721 ( .A1(n7301), .A2(n6759), .ZN(n6758) );
  INV_X1 U8722 ( .A(n6757), .ZN(n6756) );
  NOR2_X1 U8723 ( .A1(n10283), .A2(n6760), .ZN(n6759) );
  INV_X1 U8724 ( .A(n14105), .ZN(n14256) );
  INV_X1 U8725 ( .A(n15525), .ZN(n15565) );
  AND2_X1 U8726 ( .A1(n11023), .A2(n13743), .ZN(n15525) );
  OR2_X1 U8727 ( .A1(n8658), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n8632) );
  NAND2_X1 U8728 ( .A1(n8332), .A2(n8370), .ZN(n7517) );
  OR2_X1 U8729 ( .A1(n8150), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n8160) );
  INV_X1 U8730 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8731) );
  NAND2_X1 U8731 ( .A1(n14459), .A2(n6690), .ZN(n7886) );
  AND2_X1 U8732 ( .A1(n7889), .A2(n9751), .ZN(n6690) );
  OR2_X1 U8733 ( .A1(n14379), .A2(n14380), .ZN(n14377) );
  NAND2_X1 U8734 ( .A1(n9754), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9773) );
  AND2_X1 U8735 ( .A1(n11589), .A2(n9531), .ZN(n11942) );
  INV_X1 U8736 ( .A(n6986), .ZN(n6990) );
  AND2_X1 U8737 ( .A1(n9510), .A2(n9511), .ZN(n7193) );
  INV_X1 U8738 ( .A(n6720), .ZN(n9792) );
  NAND2_X1 U8739 ( .A1(n6720), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9835) );
  NAND2_X1 U8740 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9467) );
  INV_X1 U8741 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9537) );
  INV_X1 U8742 ( .A(n6730), .ZN(n9553) );
  NAND2_X1 U8743 ( .A1(n6729), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9584) );
  INV_X1 U8744 ( .A(n9382), .ZN(n6729) );
  NAND2_X1 U8745 ( .A1(n9582), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9602) );
  INV_X1 U8746 ( .A(n9584), .ZN(n9582) );
  NAND2_X1 U8747 ( .A1(n6721), .A2(n9672), .ZN(n9694) );
  NAND2_X1 U8748 ( .A1(n12393), .A2(n7891), .ZN(n7890) );
  INV_X1 U8749 ( .A(n7947), .ZN(n7891) );
  NAND2_X1 U8750 ( .A1(n14377), .A2(n9610), .ZN(n14424) );
  OR2_X1 U8751 ( .A1(n9844), .A2(n9823), .ZN(n9829) );
  AND3_X1 U8752 ( .A1(n9620), .A2(n9619), .A3(n9618), .ZN(n14932) );
  AND3_X1 U8753 ( .A1(n9639), .A2(n9638), .A3(n9637), .ZN(n12018) );
  AND4_X1 U8754 ( .A1(n9589), .A2(n9588), .A3(n9587), .A4(n9586), .ZN(n14661)
         );
  AND4_X1 U8755 ( .A1(n9557), .A2(n9556), .A3(n9555), .A4(n9554), .ZN(n11981)
         );
  AND4_X1 U8756 ( .A1(n9543), .A2(n9542), .A3(n9541), .A4(n9540), .ZN(n11832)
         );
  NAND2_X1 U8757 ( .A1(n9444), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7733) );
  INV_X1 U8758 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14513) );
  INV_X1 U8759 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14531) );
  NOR2_X1 U8760 ( .A1(n15271), .A2(n15429), .ZN(n7336) );
  NOR2_X1 U8761 ( .A1(n11316), .A2(n6502), .ZN(n14582) );
  NAND2_X1 U8762 ( .A1(n11325), .A2(n11324), .ZN(n14577) );
  NAND2_X1 U8763 ( .A1(n14577), .A2(n14578), .ZN(n14576) );
  AND2_X1 U8764 ( .A1(n11340), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7341) );
  INV_X1 U8765 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n11344) );
  AOI21_X1 U8766 ( .B1(n14600), .B2(n14599), .A(n6700), .ZN(n14601) );
  AND2_X1 U8767 ( .A1(n14597), .A2(n14598), .ZN(n6700) );
  NAND2_X1 U8768 ( .A1(n14601), .A2(n14602), .ZN(n14610) );
  NAND2_X1 U8769 ( .A1(n11722), .A2(n14598), .ZN(n14590) );
  NAND2_X1 U8770 ( .A1(n7011), .A2(n7263), .ZN(n14639) );
  NAND2_X1 U8771 ( .A1(n7264), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7263) );
  NAND2_X1 U8772 ( .A1(n14622), .A2(n14621), .ZN(n7011) );
  INV_X1 U8773 ( .A(n14625), .ZN(n7264) );
  AND2_X1 U8774 ( .A1(n14644), .A2(n9940), .ZN(n7335) );
  NAND2_X1 U8775 ( .A1(n14637), .A2(n14636), .ZN(n14638) );
  NAND2_X1 U8776 ( .A1(n7110), .A2(n9925), .ZN(n14726) );
  NAND2_X1 U8777 ( .A1(n6719), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n14731) );
  OAI211_X1 U8778 ( .C1(n7110), .C2(n14740), .A(n7107), .B(n7106), .ZN(n14721)
         );
  NAND2_X1 U8779 ( .A1(n7109), .A2(n7108), .ZN(n7106) );
  NAND2_X1 U8780 ( .A1(n7110), .A2(n6468), .ZN(n7107) );
  NOR2_X1 U8781 ( .A1(n14772), .A2(n6943), .ZN(n6942) );
  INV_X1 U8782 ( .A(n14713), .ZN(n6943) );
  OR2_X1 U8783 ( .A1(n6520), .A2(n7938), .ZN(n7697) );
  INV_X1 U8784 ( .A(n15046), .ZN(n14822) );
  NOR2_X2 U8785 ( .A1(n14871), .A2(n14854), .ZN(n14853) );
  INV_X1 U8786 ( .A(n15051), .ZN(n14833) );
  NAND2_X1 U8787 ( .A1(n6733), .A2(n6732), .ZN(n9737) );
  NOR2_X1 U8788 ( .A1(n12384), .A2(n9721), .ZN(n6732) );
  INV_X1 U8789 ( .A(n6733), .ZN(n9722) );
  AND2_X1 U8790 ( .A1(n9744), .A2(n9743), .ZN(n14870) );
  INV_X1 U8791 ( .A(n6920), .ZN(n6919) );
  NAND2_X1 U8792 ( .A1(n14941), .A2(n6923), .ZN(n6922) );
  OAI21_X1 U8793 ( .B1(n6492), .B2(n6921), .A(n14696), .ZN(n6920) );
  AND2_X1 U8794 ( .A1(n9660), .A2(n9659), .ZN(n14921) );
  NAND2_X1 U8795 ( .A1(n12021), .A2(n7756), .ZN(n14946) );
  NOR2_X1 U8796 ( .A1(n14961), .A2(n15103), .ZN(n14960) );
  NAND2_X1 U8797 ( .A1(n14971), .A2(n12030), .ZN(n12033) );
  NAND2_X1 U8798 ( .A1(n12073), .A2(n12014), .ZN(n14979) );
  AND2_X1 U8799 ( .A1(n6504), .A2(n14977), .ZN(n7769) );
  NAND2_X1 U8800 ( .A1(n7712), .A2(n6518), .ZN(n12069) );
  NAND2_X1 U8801 ( .A1(n12010), .A2(n6462), .ZN(n7713) );
  AOI21_X1 U8802 ( .B1(n7351), .B2(n7353), .A(n6554), .ZN(n7349) );
  AND2_X1 U8803 ( .A1(n11824), .A2(n14503), .ZN(n12043) );
  NAND2_X1 U8804 ( .A1(n11825), .A2(n7771), .ZN(n12065) );
  NAND2_X1 U8805 ( .A1(n11825), .A2(n11824), .ZN(n12039) );
  AOI21_X1 U8806 ( .B1(n7346), .B2(n7348), .A(n6557), .ZN(n7344) );
  OR2_X1 U8807 ( .A1(n9500), .A2(n9499), .ZN(n9513) );
  INV_X1 U8808 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9512) );
  OR2_X1 U8809 ( .A1(n9513), .A2(n9512), .ZN(n9538) );
  NAND2_X1 U8810 ( .A1(n7116), .A2(n7114), .ZN(n7726) );
  INV_X1 U8811 ( .A(n7115), .ZN(n7114) );
  OAI21_X1 U8812 ( .B1(n7119), .B2(n6454), .A(n15304), .ZN(n7115) );
  INV_X1 U8813 ( .A(n7119), .ZN(n7113) );
  NAND2_X1 U8814 ( .A1(n11113), .A2(n11250), .ZN(n15314) );
  INV_X1 U8815 ( .A(n11366), .ZN(n11362) );
  AND2_X1 U8816 ( .A1(n7144), .A2(n10993), .ZN(n11363) );
  NAND2_X1 U8817 ( .A1(n11363), .A2(n11362), .ZN(n11361) );
  CLKBUF_X1 U8818 ( .A(n11066), .Z(n7190) );
  NAND2_X1 U8819 ( .A1(n9435), .A2(n14994), .ZN(n11064) );
  NAND2_X1 U8820 ( .A1(n11073), .A2(n14994), .ZN(n10992) );
  INV_X1 U8821 ( .A(n14687), .ZN(n6728) );
  NAND2_X1 U8822 ( .A1(n14844), .A2(n14710), .ZN(n14819) );
  INV_X1 U8823 ( .A(n15406), .ZN(n15418) );
  OAI211_X1 U8824 ( .C1(n9912), .C2(n9865), .A(n9864), .B(n9863), .ZN(n14355)
         );
  XNOR2_X1 U8825 ( .A(n9852), .B(n9851), .ZN(n14361) );
  NAND2_X1 U8826 ( .A1(n8495), .A2(n8494), .ZN(n8508) );
  NAND2_X1 U8827 ( .A1(n7086), .A2(n7083), .ZN(n8028) );
  XNOR2_X1 U8828 ( .A(n9327), .B(P1_IR_REG_24__SCAN_IN), .ZN(n9810) );
  AND2_X1 U8829 ( .A1(n8480), .A2(n8479), .ZN(n12114) );
  NAND2_X1 U8830 ( .A1(n7575), .A2(n7576), .ZN(n7574) );
  XNOR2_X1 U8831 ( .A(n8434), .B(n8433), .ZN(n11707) );
  NAND2_X1 U8832 ( .A1(n7316), .A2(n8006), .ZN(n8399) );
  NAND2_X1 U8833 ( .A1(n7322), .A2(n7321), .ZN(n7316) );
  XNOR2_X1 U8834 ( .A(n8367), .B(n8369), .ZN(n10871) );
  NAND2_X1 U8835 ( .A1(n7082), .A2(n8002), .ZN(n8367) );
  NOR2_X1 U8836 ( .A1(n9368), .A2(n9473), .ZN(n9624) );
  NOR3_X1 U8837 ( .A1(n9368), .A2(n9473), .A3(P1_IR_REG_15__SCAN_IN), .ZN(
        n9627) );
  NAND2_X1 U8838 ( .A1(n7592), .A2(n7994), .ZN(n8345) );
  NAND2_X1 U8839 ( .A1(n7992), .A2(n7599), .ZN(n7592) );
  NAND2_X1 U8840 ( .A1(n7992), .A2(n7991), .ZN(n8316) );
  XNOR2_X1 U8841 ( .A(n9597), .B(P1_IR_REG_13__SCAN_IN), .ZN(n11340) );
  OAI21_X1 U8842 ( .B1(n9376), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9577) );
  NAND2_X1 U8843 ( .A1(n7573), .A2(n7979), .ZN(n8268) );
  NAND2_X1 U8844 ( .A1(n8260), .A2(n7977), .ZN(n7573) );
  INV_X1 U8845 ( .A(n7967), .ZN(n8239) );
  NOR2_X1 U8846 ( .A1(n9406), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n7251) );
  NAND2_X1 U8847 ( .A1(n7024), .A2(n7022), .ZN(n9404) );
  AND2_X1 U8848 ( .A1(n7023), .A2(n9474), .ZN(n7022) );
  INV_X1 U8849 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9474) );
  NAND2_X1 U8850 ( .A1(n9450), .A2(n9303), .ZN(n9319) );
  INV_X1 U8851 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9303) );
  OAI211_X1 U8852 ( .C1(n10371), .C2(n7156), .A(n7153), .B(n7152), .ZN(n10377)
         );
  AND2_X1 U8853 ( .A1(n7154), .A2(n7158), .ZN(n7153) );
  INV_X1 U8854 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14546) );
  NAND2_X1 U8855 ( .A1(n10758), .A2(n10757), .ZN(n10768) );
  XNOR2_X1 U8856 ( .A(n11277), .B(n10776), .ZN(n10777) );
  OAI21_X1 U8857 ( .B1(n11501), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n11500), .ZN(
        n11732) );
  XNOR2_X1 U8858 ( .A(n11636), .B(n12494), .ZN(n11794) );
  OAI21_X1 U8859 ( .B1(n12517), .B2(n7838), .A(n7834), .ZN(n12535) );
  INV_X1 U8860 ( .A(n7802), .ZN(n6800) );
  INV_X1 U8861 ( .A(n12509), .ZN(n7801) );
  NAND2_X1 U8862 ( .A1(n12605), .A2(n12481), .ZN(n12525) );
  OR2_X1 U8863 ( .A1(n7838), .A2(n7831), .ZN(n7828) );
  AND2_X1 U8864 ( .A1(n9151), .A2(n9150), .ZN(n12848) );
  NAND2_X1 U8865 ( .A1(n7096), .A2(n7819), .ZN(n12548) );
  NAND2_X1 U8866 ( .A1(n12605), .A2(n7821), .ZN(n7096) );
  AND4_X1 U8867 ( .A1(n9016), .A2(n9015), .A3(n9014), .A4(n9013), .ZN(n12985)
         );
  NAND2_X1 U8868 ( .A1(n12622), .A2(n12473), .ZN(n12563) );
  NAND2_X1 U8869 ( .A1(n12622), .A2(n7798), .ZN(n12564) );
  NAND2_X1 U8870 ( .A1(n11421), .A2(n11420), .ZN(n11422) );
  NAND2_X1 U8871 ( .A1(n6785), .A2(n6783), .ZN(n12571) );
  AOI21_X1 U8872 ( .B1(n6786), .B2(n6787), .A(n6784), .ZN(n6783) );
  INV_X1 U8873 ( .A(n12572), .ZN(n6784) );
  OAI21_X1 U8874 ( .B1(n12471), .B2(n6787), .A(n6786), .ZN(n12573) );
  NAND2_X1 U8875 ( .A1(n7820), .A2(n7825), .ZN(n12592) );
  NAND2_X1 U8876 ( .A1(n12605), .A2(n7827), .ZN(n7820) );
  OAI21_X1 U8877 ( .B1(n12605), .B2(n7824), .A(n7821), .ZN(n12590) );
  AND4_X1 U8878 ( .A1(n9032), .A2(n9031), .A3(n9030), .A4(n9029), .ZN(n12953)
         );
  NAND2_X1 U8879 ( .A1(n11994), .A2(n11993), .ZN(n7807) );
  INV_X1 U8880 ( .A(n12796), .ZN(n12775) );
  NAND2_X1 U8881 ( .A1(n9199), .A2(n9198), .ZN(n12822) );
  INV_X1 U8882 ( .A(n12848), .ZN(n12875) );
  NAND2_X1 U8883 ( .A1(n9140), .A2(n9139), .ZN(n12860) );
  INV_X1 U8884 ( .A(n13070), .ZN(n12638) );
  INV_X1 U8885 ( .A(n12953), .ZN(n12976) );
  INV_X1 U8886 ( .A(n10174), .ZN(n11142) );
  NAND2_X1 U8887 ( .A1(n7187), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10958) );
  OR2_X1 U8888 ( .A1(n10948), .A2(n13015), .ZN(n10949) );
  NAND2_X1 U8889 ( .A1(n10147), .A2(n11125), .ZN(n11083) );
  INV_X1 U8890 ( .A(n6857), .ZN(n11087) );
  AOI22_X1 U8891 ( .A1(n11081), .A2(n11082), .B1(n10218), .B2(n10217), .ZN(
        n11034) );
  OAI22_X1 U8892 ( .A1(n11032), .A2(n10181), .B1(n7436), .B2(n7640), .ZN(
        n11190) );
  INV_X1 U8893 ( .A(n7641), .ZN(n7640) );
  XNOR2_X1 U8894 ( .A(n10182), .B(n11466), .ZN(n11458) );
  NAND2_X1 U8895 ( .A1(n7377), .A2(n7380), .ZN(n11461) );
  NAND2_X1 U8896 ( .A1(n11034), .A2(n6503), .ZN(n7377) );
  NAND2_X1 U8897 ( .A1(n6984), .A2(n6983), .ZN(n11613) );
  AND2_X1 U8898 ( .A1(n6828), .A2(n7255), .ZN(n11600) );
  NAND2_X1 U8899 ( .A1(n11458), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n6828) );
  NOR2_X1 U8900 ( .A1(n12666), .A2(n7443), .ZN(n12664) );
  NAND2_X1 U8901 ( .A1(n7442), .A2(n7444), .ZN(n12648) );
  OAI211_X1 U8902 ( .C1(n11846), .C2(n6635), .A(n6837), .B(n6831), .ZN(n12650)
         );
  NAND2_X1 U8903 ( .A1(n11846), .A2(n6836), .ZN(n6831) );
  NAND2_X1 U8904 ( .A1(n7432), .A2(n10159), .ZN(n12687) );
  NOR2_X1 U8905 ( .A1(n12687), .A2(n12688), .ZN(n12711) );
  NOR2_X1 U8906 ( .A1(n12695), .A2(n6459), .ZN(n12718) );
  NAND2_X1 U8907 ( .A1(n12708), .A2(n6666), .ZN(n6977) );
  NAND2_X1 U8908 ( .A1(n12695), .A2(n7368), .ZN(n7366) );
  NAND2_X1 U8909 ( .A1(n12299), .A2(n12298), .ZN(n12757) );
  NAND2_X1 U8910 ( .A1(n15601), .A2(n12780), .ZN(n6709) );
  NAND2_X1 U8911 ( .A1(n9266), .A2(n7414), .ZN(n12820) );
  NAND2_X1 U8912 ( .A1(n9265), .A2(n6494), .ZN(n7414) );
  NAND2_X1 U8913 ( .A1(n9175), .A2(n7848), .ZN(n12819) );
  NAND2_X1 U8914 ( .A1(n9152), .A2(n7851), .ZN(n7848) );
  NAND2_X1 U8915 ( .A1(n9265), .A2(n9264), .ZN(n12836) );
  OR2_X1 U8916 ( .A1(n10636), .A2(n7404), .ZN(n9072) );
  AND3_X1 U8917 ( .A1(n9078), .A2(n9077), .A3(n9076), .ZN(n13085) );
  AND3_X1 U8918 ( .A1(n9094), .A2(n9093), .A3(n9092), .ZN(n13091) );
  NAND2_X1 U8919 ( .A1(n9055), .A2(n9054), .ZN(n13094) );
  AND3_X1 U8920 ( .A1(n9061), .A2(n9060), .A3(n9059), .ZN(n13097) );
  AND4_X1 U8921 ( .A1(n8990), .A2(n8989), .A3(n8988), .A4(n8987), .ZN(n13119)
         );
  NAND2_X1 U8922 ( .A1(n7875), .A2(n12200), .ZN(n12117) );
  NAND2_X1 U8923 ( .A1(n8948), .A2(n7876), .ZN(n7875) );
  NAND2_X1 U8924 ( .A1(n8948), .A2(n12194), .ZN(n11918) );
  INV_X1 U8925 ( .A(n9233), .ZN(n11958) );
  INV_X1 U8926 ( .A(n11663), .ZN(n15655) );
  NAND2_X1 U8927 ( .A1(n11517), .A2(n9230), .ZN(n11570) );
  NAND2_X1 U8928 ( .A1(n11535), .A2(n8896), .ZN(n11515) );
  OR2_X1 U8929 ( .A1(n12300), .A2(n11453), .ZN(n8853) );
  NAND2_X1 U8930 ( .A1(n10166), .A2(n7628), .ZN(n8830) );
  AND2_X1 U8931 ( .A1(n10339), .A2(n10419), .ZN(n7628) );
  INV_X1 U8932 ( .A(n7790), .ZN(n7789) );
  INV_X1 U8933 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n15725) );
  NOR2_X1 U8934 ( .A1(n15664), .A2(n15602), .ZN(n7863) );
  NOR2_X1 U8935 ( .A1(n9279), .A2(n6528), .ZN(n7867) );
  INV_X1 U8936 ( .A(n12489), .ZN(n13162) );
  NAND2_X1 U8937 ( .A1(n12241), .A2(n12883), .ZN(n12867) );
  NAND2_X1 U8938 ( .A1(n9026), .A2(n9025), .ZN(n13200) );
  OAI21_X1 U8939 ( .B1(n12982), .B2(n7858), .A(n7856), .ZN(n12961) );
  NAND2_X1 U8940 ( .A1(n9008), .A2(n9007), .ZN(n13206) );
  NAND2_X1 U8941 ( .A1(n7861), .A2(n12213), .ZN(n12975) );
  NAND2_X1 U8942 ( .A1(n12982), .A2(n6694), .ZN(n7861) );
  OR2_X1 U8943 ( .A1(n9233), .A2(n7783), .ZN(n7398) );
  AND2_X1 U8944 ( .A1(n10828), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13224) );
  INV_X1 U8945 ( .A(n13224), .ZN(n12154) );
  INV_X1 U8946 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7884) );
  NAND2_X1 U8947 ( .A1(n7687), .A2(n8799), .ZN(n12272) );
  OAI21_X1 U8948 ( .B1(n9127), .B2(n7667), .A(n7665), .ZN(n9163) );
  NAND2_X1 U8949 ( .A1(n9129), .A2(n8788), .ZN(n9142) );
  NAND2_X1 U8950 ( .A1(n8684), .A2(n8723), .ZN(n11291) );
  OR2_X1 U8951 ( .A1(n9127), .A2(n9126), .ZN(n9128) );
  INV_X1 U8952 ( .A(n9286), .ZN(n12316) );
  OAI21_X1 U8953 ( .B1(n9064), .B2(n7681), .A(n7679), .ZN(n9098) );
  OAI21_X1 U8954 ( .B1(n9050), .B2(n6883), .A(n6881), .ZN(n9082) );
  NAND2_X1 U8955 ( .A1(n6880), .A2(n8778), .ZN(n9080) );
  INV_X1 U8956 ( .A(SI_15_), .ZN(n10503) );
  OAI21_X1 U8957 ( .B1(n8767), .B2(n7659), .A(n7657), .ZN(n9034) );
  INV_X1 U8958 ( .A(SI_12_), .ZN(n10416) );
  INV_X1 U8959 ( .A(SI_11_), .ZN(n10356) );
  NAND2_X1 U8960 ( .A1(n8967), .A2(n8761), .ZN(n8980) );
  INV_X1 U8961 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8969) );
  NOR2_X1 U8962 ( .A1(n7814), .A2(n8859), .ZN(n8968) );
  NAND2_X1 U8963 ( .A1(n8945), .A2(n8756), .ZN(n8950) );
  XNOR2_X1 U8964 ( .A(n8941), .B(n8940), .ZN(n10428) );
  NAND2_X1 U8965 ( .A1(n8751), .A2(n8750), .ZN(n8920) );
  NAND2_X1 U8966 ( .A1(n6890), .A2(n8745), .ZN(n8886) );
  NAND2_X1 U8967 ( .A1(n8872), .A2(n8744), .ZN(n6890) );
  NAND2_X1 U8968 ( .A1(n10139), .A2(n8846), .ZN(n7642) );
  NAND2_X1 U8969 ( .A1(n7540), .A2(n13268), .ZN(n13331) );
  AND2_X1 U8970 ( .A1(n7520), .A2(n7522), .ZN(n11774) );
  AND2_X1 U8971 ( .A1(n11224), .A2(n6519), .ZN(n6458) );
  NAND2_X1 U8972 ( .A1(n7075), .A2(n7076), .ZN(n13358) );
  NAND2_X1 U8973 ( .A1(n13440), .A2(n13296), .ZN(n13389) );
  NAND2_X1 U8974 ( .A1(n7059), .A2(n12131), .ZN(n12134) );
  NAND2_X1 U8975 ( .A1(n11882), .A2(n7063), .ZN(n7059) );
  OAI21_X1 U8976 ( .B1(n11882), .B2(n7062), .A(n7060), .ZN(n12145) );
  AND2_X1 U8977 ( .A1(n7055), .A2(n7053), .ZN(n13414) );
  NOR2_X1 U8978 ( .A1(n11476), .A2(n7054), .ZN(n7053) );
  NAND2_X1 U8979 ( .A1(n6458), .A2(n7245), .ZN(n7055) );
  AOI21_X1 U8980 ( .B1(n11475), .B2(n11474), .A(n13412), .ZN(n11476) );
  OAI211_X2 U8981 ( .C1(n7177), .C2(n10327), .A(n8166), .B(n8165), .ZN(n15826)
         );
  NAND2_X1 U8982 ( .A1(n7537), .A2(n7536), .ZN(n13433) );
  NAND2_X1 U8983 ( .A1(n11626), .A2(n7523), .ZN(n11768) );
  AOI21_X1 U8984 ( .B1(n7060), .B2(n7062), .A(n12144), .ZN(n7057) );
  XNOR2_X1 U8985 ( .A(n13305), .B(n13304), .ZN(n13452) );
  OR2_X1 U8986 ( .A1(n10749), .A2(n13743), .ZN(n13461) );
  NAND2_X1 U8987 ( .A1(n11882), .A2(n11881), .ZN(n12133) );
  OR2_X1 U8988 ( .A1(n8131), .A2(n10569), .ZN(n8093) );
  NAND2_X1 U8989 ( .A1(n10877), .A2(n10876), .ZN(n10878) );
  INV_X1 U8990 ( .A(n13495), .ZN(n13459) );
  NAND2_X1 U8991 ( .A1(n7174), .A2(n13368), .ZN(n13473) );
  NAND2_X1 U8992 ( .A1(n7176), .A2(n7175), .ZN(n7174) );
  INV_X1 U8993 ( .A(n13315), .ZN(n7175) );
  INV_X1 U8994 ( .A(n13316), .ZN(n7176) );
  INV_X1 U8995 ( .A(n13479), .ZN(n13498) );
  INV_X1 U8996 ( .A(n13481), .ZN(n13487) );
  AND2_X1 U8997 ( .A1(n7476), .A2(n8558), .ZN(n7474) );
  NAND2_X1 U8998 ( .A1(n8081), .A2(n8080), .ZN(n14026) );
  NAND2_X1 U8999 ( .A1(n8491), .A2(n8490), .ZN(n14041) );
  OR2_X1 U9000 ( .A1(n14028), .A2(n8530), .ZN(n8491) );
  NAND2_X1 U9001 ( .A1(n8475), .A2(n8474), .ZN(n14024) );
  OAI211_X1 U9002 ( .C1(n13428), .C2(n8530), .A(n8378), .B(n8377), .ZN(n13816)
         );
  OR2_X1 U9003 ( .A1(n8362), .A2(n8361), .ZN(n13818) );
  NAND2_X1 U9004 ( .A1(n6747), .A2(n6754), .ZN(n13824) );
  INV_X1 U9005 ( .A(n6751), .ZN(n6747) );
  NAND4_X1 U9006 ( .A1(n8173), .A2(n8172), .A3(n8171), .A4(n8170), .ZN(n13826)
         );
  OR2_X1 U9007 ( .A1(n7486), .A2(n7056), .ZN(n13827) );
  NOR2_X1 U9008 ( .A1(n8530), .A2(n15502), .ZN(n7056) );
  OR2_X1 U9009 ( .A1(n8126), .A2(n11185), .ZN(n8083) );
  NOR2_X1 U9010 ( .A1(n8129), .A2(n8128), .ZN(n8133) );
  NAND2_X1 U9011 ( .A1(n15455), .A2(n15456), .ZN(n15454) );
  NAND2_X1 U9012 ( .A1(n15458), .A2(n15459), .ZN(n15457) );
  NAND2_X1 U9013 ( .A1(n10592), .A2(n10591), .ZN(n10684) );
  NAND2_X1 U9014 ( .A1(n10684), .A2(n10593), .ZN(n15471) );
  OAI21_X1 U9015 ( .B1(n10592), .B2(n6964), .A(n6962), .ZN(n15469) );
  NAND2_X1 U9016 ( .A1(n6961), .A2(n6959), .ZN(n10595) );
  AOI22_X1 U9017 ( .A1(n10616), .A2(n10617), .B1(P2_REG1_REG_7__SCAN_IN), .B2(
        n10612), .ZN(n10625) );
  NAND2_X1 U9018 ( .A1(n10632), .A2(n6971), .ZN(n10722) );
  NOR2_X1 U9019 ( .A1(n10601), .A2(n6972), .ZN(n6971) );
  INV_X1 U9020 ( .A(n10599), .ZN(n6972) );
  NAND2_X1 U9021 ( .A1(n10722), .A2(n10721), .ZN(n10781) );
  NAND2_X1 U9022 ( .A1(n10722), .A2(n6969), .ZN(n10782) );
  NOR2_X1 U9023 ( .A1(n10780), .A2(n6970), .ZN(n6969) );
  INV_X1 U9024 ( .A(n10721), .ZN(n6970) );
  OR2_X1 U9025 ( .A1(n10726), .A2(n10725), .ZN(n10921) );
  AOI21_X1 U9026 ( .B1(n10723), .B2(P2_REG1_REG_10__SCAN_IN), .A(n10784), .ZN(
        n10913) );
  AND2_X1 U9027 ( .A1(n11267), .A2(n11266), .ZN(n11271) );
  INV_X1 U9028 ( .A(n15444), .ZN(n15470) );
  AND2_X1 U9029 ( .A1(n10605), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15468) );
  OR2_X1 U9030 ( .A1(n13914), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n13932) );
  XNOR2_X1 U9031 ( .A(n13955), .B(n10268), .ZN(n13952) );
  AND2_X1 U9032 ( .A1(n8622), .A2(n13945), .ZN(n13960) );
  XNOR2_X1 U9033 ( .A(n10275), .B(n10274), .ZN(n13969) );
  AOI211_X1 U9034 ( .C1(n13720), .C2(n10273), .A(n15561), .B(n10272), .ZN(
        n13968) );
  AOI21_X1 U9035 ( .B1(n7301), .B2(n6762), .A(n6761), .ZN(n10281) );
  NAND2_X1 U9036 ( .A1(n6740), .A2(n7558), .ZN(n14018) );
  NAND2_X1 U9037 ( .A1(n14054), .A2(n8598), .ZN(n14037) );
  NAND2_X1 U9038 ( .A1(n14051), .A2(n8459), .ZN(n14035) );
  NAND2_X1 U9039 ( .A1(n7503), .A2(n7506), .ZN(n14067) );
  NAND2_X1 U9040 ( .A1(n14098), .A2(n6483), .ZN(n7503) );
  NAND2_X1 U9041 ( .A1(n7508), .A2(n6483), .ZN(n14084) );
  NAND2_X1 U9042 ( .A1(n7508), .A2(n8595), .ZN(n14082) );
  NAND2_X1 U9043 ( .A1(n7310), .A2(n10248), .ZN(n8420) );
  INV_X1 U9044 ( .A(n12447), .ZN(n7310) );
  NAND2_X1 U9045 ( .A1(n7305), .A2(n8414), .ZN(n14078) );
  NAND2_X1 U9046 ( .A1(n8397), .A2(n8396), .ZN(n14096) );
  INV_X1 U9047 ( .A(n13648), .ZN(n14262) );
  INV_X1 U9048 ( .A(n7547), .ZN(n7282) );
  OAI21_X1 U9049 ( .B1(n8579), .B2(n6792), .A(n6790), .ZN(n14159) );
  OAI21_X1 U9050 ( .B1(n11813), .B2(n7550), .A(n7548), .ZN(n14174) );
  NAND2_X1 U9051 ( .A1(n7510), .A2(n7511), .ZN(n14175) );
  NAND2_X1 U9052 ( .A1(n8581), .A2(n6456), .ZN(n7510) );
  NAND2_X1 U9053 ( .A1(n7553), .A2(n7551), .ZN(n14199) );
  INV_X1 U9054 ( .A(n7554), .ZN(n7551) );
  NAND2_X1 U9055 ( .A1(n11813), .A2(n6484), .ZN(n7553) );
  NAND2_X1 U9056 ( .A1(n8581), .A2(n8580), .ZN(n14187) );
  OAI21_X1 U9057 ( .B1(n11813), .B2(n8282), .A(n8281), .ZN(n11894) );
  OAI21_X1 U9058 ( .B1(n11865), .B2(n8576), .A(n8575), .ZN(n11803) );
  OAI21_X1 U9059 ( .B1(n11413), .B2(n7299), .A(n6485), .ZN(n11864) );
  NAND2_X1 U9060 ( .A1(n8265), .A2(n8264), .ZN(n13581) );
  NAND2_X1 U9061 ( .A1(n11700), .A2(n8572), .ZN(n11761) );
  INV_X1 U9062 ( .A(n6752), .ZN(n11588) );
  NAND2_X1 U9063 ( .A1(n6945), .A2(n13515), .ZN(n11183) );
  INV_X1 U9064 ( .A(n13503), .ZN(n7237) );
  NAND2_X1 U9065 ( .A1(n10740), .A2(n15517), .ZN(n15503) );
  AND2_X1 U9066 ( .A1(n15831), .A2(n11137), .ZN(n15484) );
  AND2_X1 U9067 ( .A1(n15831), .A2(n11022), .ZN(n15827) );
  INV_X1 U9068 ( .A(n13535), .ZN(n13531) );
  INV_X1 U9069 ( .A(n14208), .ZN(n7327) );
  INV_X1 U9070 ( .A(n7324), .ZN(n7323) );
  OAI21_X1 U9071 ( .B1(n14211), .B2(n14310), .A(n7325), .ZN(n7324) );
  INV_X1 U9072 ( .A(n14008), .ZN(n14321) );
  NAND2_X1 U9073 ( .A1(n7182), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6803) );
  INV_X1 U9074 ( .A(n14213), .ZN(n6805) );
  INV_X1 U9075 ( .A(n14214), .ZN(n6806) );
  AND2_X1 U9076 ( .A1(n10578), .A2(n10298), .ZN(n15517) );
  NOR2_X1 U9077 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n7483) );
  INV_X1 U9078 ( .A(n6793), .ZN(n8059) );
  XNOR2_X1 U9079 ( .A(n8061), .B(n15801), .ZN(n14363) );
  NAND2_X1 U9080 ( .A1(n6794), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8061) );
  NAND2_X1 U9081 ( .A1(n6793), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6734) );
  XNOR2_X1 U9082 ( .A(n8044), .B(n8043), .ZN(n14366) );
  NAND2_X1 U9083 ( .A1(n8638), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8044) );
  INV_X1 U9084 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11863) );
  AND2_X1 U9085 ( .A1(n8461), .A2(n8447), .ZN(n11907) );
  INV_X1 U9086 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n15733) );
  INV_X1 U9087 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10874) );
  INV_X1 U9088 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10713) );
  INV_X1 U9089 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10558) );
  INV_X1 U9090 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10505) );
  INV_X1 U9091 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10485) );
  INV_X1 U9092 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10412) );
  INV_X1 U9093 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10402) );
  INV_X1 U9094 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10350) );
  INV_X1 U9095 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10334) );
  INV_X1 U9096 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10347) );
  INV_X1 U9097 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10331) );
  INV_X1 U9098 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10327) );
  INV_X1 U9099 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10316) );
  INV_X1 U9100 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10315) );
  INV_X1 U9101 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10313) );
  XNOR2_X1 U9102 ( .A(n8087), .B(n8097), .ZN(n13851) );
  NAND2_X1 U9103 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n7309) );
  NAND2_X1 U9104 ( .A1(n7908), .A2(n9689), .ZN(n14397) );
  NAND2_X1 U9105 ( .A1(n7192), .A2(n9560), .ZN(n7191) );
  NAND2_X1 U9106 ( .A1(n12381), .A2(n9718), .ZN(n14406) );
  NAND2_X1 U9107 ( .A1(n11930), .A2(n7248), .ZN(n14414) );
  NAND2_X1 U9108 ( .A1(n7902), .A2(n7905), .ZN(n14437) );
  AOI21_X1 U9109 ( .B1(n6995), .B2(n6997), .A(n6993), .ZN(n6992) );
  NAND2_X1 U9110 ( .A1(n14460), .A2(n6995), .ZN(n6994) );
  INV_X1 U9111 ( .A(n12396), .ZN(n6993) );
  INV_X1 U9112 ( .A(n14702), .ZN(n15071) );
  AND2_X1 U9113 ( .A1(n9605), .A2(n9604), .ZN(n14981) );
  NAND2_X1 U9114 ( .A1(n9575), .A2(n9574), .ZN(n7213) );
  NAND2_X1 U9115 ( .A1(n7910), .A2(n9570), .ZN(n11932) );
  AOI21_X1 U9116 ( .B1(n10662), .B2(n10663), .A(n9442), .ZN(n10655) );
  AND2_X1 U9117 ( .A1(n7905), .A2(n7901), .ZN(n7900) );
  INV_X1 U9118 ( .A(n14498), .ZN(n14462) );
  OR2_X1 U9119 ( .A1(n10134), .A2(n10133), .ZN(n10136) );
  INV_X1 U9120 ( .A(n14798), .ZN(n14830) );
  INV_X1 U9121 ( .A(n14870), .ZN(n14831) );
  INV_X1 U9122 ( .A(n14921), .ZN(n14500) );
  INV_X1 U9123 ( .A(n14932), .ZN(n14691) );
  INV_X1 U9124 ( .A(n12018), .ZN(n14690) );
  INV_X1 U9125 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10518) );
  NAND2_X1 U9126 ( .A1(n14515), .A2(n14516), .ZN(n14534) );
  NAND2_X1 U9127 ( .A1(n10451), .A2(n10450), .ZN(n15267) );
  NAND2_X1 U9128 ( .A1(n10466), .A2(n10465), .ZN(n15274) );
  OR2_X1 U9129 ( .A1(n10540), .A2(n15435), .ZN(n7338) );
  OAI21_X1 U9130 ( .B1(n10550), .B2(n10478), .A(n10477), .ZN(n10522) );
  INV_X1 U9131 ( .A(n7009), .ZN(n10647) );
  AND2_X1 U9132 ( .A1(n7007), .A2(n7006), .ZN(n11316) );
  INV_X1 U9133 ( .A(n10698), .ZN(n7006) );
  NAND2_X1 U9134 ( .A1(n10700), .A2(n10699), .ZN(n7007) );
  NAND2_X1 U9135 ( .A1(n7021), .A2(n7020), .ZN(n11337) );
  INV_X1 U9136 ( .A(n11320), .ZN(n7020) );
  INV_X1 U9137 ( .A(n11321), .ZN(n7021) );
  AOI21_X1 U9138 ( .B1(n11337), .B2(n11336), .A(n11335), .ZN(n11720) );
  NAND2_X1 U9139 ( .A1(n14596), .A2(n7013), .ZN(n14608) );
  NOR2_X1 U9140 ( .A1(n6657), .A2(n7014), .ZN(n7013) );
  NAND2_X1 U9141 ( .A1(n14608), .A2(n7012), .ZN(n14622) );
  INV_X1 U9142 ( .A(n7014), .ZN(n7012) );
  XNOR2_X1 U9143 ( .A(n14639), .B(n14634), .ZN(n14623) );
  INV_X1 U9144 ( .A(n9939), .ZN(n15004) );
  AND2_X1 U9145 ( .A1(n9918), .A2(n9917), .ZN(n15009) );
  NAND2_X1 U9146 ( .A1(n12457), .A2(n9461), .ZN(n9883) );
  INV_X1 U9147 ( .A(n14753), .ZN(n14751) );
  AOI21_X1 U9148 ( .B1(n14739), .B2(n15359), .A(n7234), .ZN(n7927) );
  INV_X1 U9149 ( .A(n14742), .ZN(n7234) );
  AOI21_X1 U9150 ( .B1(n14762), .B2(n15359), .A(n14761), .ZN(n15029) );
  NAND2_X1 U9151 ( .A1(n14760), .A2(n14759), .ZN(n14761) );
  OAI21_X1 U9152 ( .B1(n14791), .B2(n14793), .A(n7129), .ZN(n14780) );
  NAND2_X1 U9153 ( .A1(n14828), .A2(n14682), .ZN(n14810) );
  NAND2_X1 U9154 ( .A1(n7723), .A2(n7721), .ZN(n14851) );
  NAND2_X1 U9155 ( .A1(n14866), .A2(n14867), .ZN(n7723) );
  NAND2_X1 U9156 ( .A1(n14900), .A2(n14678), .ZN(n14883) );
  OAI21_X1 U9157 ( .B1(n14941), .B2(n6928), .A(n6925), .ZN(n14909) );
  NAND2_X1 U9158 ( .A1(n12033), .A2(n7929), .ZN(n15110) );
  INV_X1 U9159 ( .A(n15116), .ZN(n14977) );
  NAND2_X1 U9160 ( .A1(n7350), .A2(n12028), .ZN(n12038) );
  NAND2_X1 U9161 ( .A1(n12027), .A2(n12026), .ZN(n7350) );
  NAND2_X1 U9162 ( .A1(n11254), .A2(n15303), .ZN(n7345) );
  NAND2_X1 U9163 ( .A1(n7121), .A2(n11108), .ZN(n11238) );
  NAND2_X1 U9164 ( .A1(n11107), .A2(n7122), .ZN(n7121) );
  INV_X1 U9165 ( .A(n14952), .ZN(n15332) );
  OR2_X1 U9166 ( .A1(n14729), .A2(n9940), .ZN(n14952) );
  CLKBUF_X1 U9167 ( .A(n7699), .Z(n15341) );
  NAND2_X1 U9168 ( .A1(n14729), .A2(n14997), .ZN(n14935) );
  INV_X1 U9169 ( .A(n14990), .ZN(n14992) );
  NAND2_X1 U9170 ( .A1(n10392), .A2(n10971), .ZN(n15338) );
  NOR2_X1 U9171 ( .A1(n6939), .A2(n6938), .ZN(n6937) );
  NOR2_X1 U9172 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n6938) );
  NOR2_X1 U9173 ( .A1(n7139), .A2(n7138), .ZN(n7137) );
  NAND2_X1 U9174 ( .A1(n9345), .A2(n9318), .ZN(n7136) );
  OAI21_X1 U9175 ( .B1(n9824), .B2(n9330), .A(n9332), .ZN(n7249) );
  XNOR2_X1 U9176 ( .A(n8465), .B(n8464), .ZN(n11860) );
  INV_X1 U9177 ( .A(n11050), .ZN(n15176) );
  INV_X1 U9178 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11708) );
  INV_X1 U9179 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10715) );
  INV_X1 U9180 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10670) );
  INV_X1 U9181 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10555) );
  XNOR2_X1 U9182 ( .A(n9599), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11721) );
  NAND2_X1 U9183 ( .A1(n9598), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9599) );
  INV_X1 U9184 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10507) );
  XNOR2_X1 U9185 ( .A(n9577), .B(P1_IR_REG_12__SCAN_IN), .ZN(n14585) );
  INV_X1 U9186 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10351) );
  AND2_X1 U9187 ( .A1(n9534), .A2(n9549), .ZN(n10644) );
  INV_X1 U9188 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10335) );
  XNOR2_X1 U9189 ( .A(n7010), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10540) );
  NOR2_X1 U9190 ( .A1(n7251), .A2(n15153), .ZN(n7010) );
  INV_X1 U9191 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10330) );
  INV_X1 U9192 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10322) );
  OAI21_X1 U9193 ( .B1(n8105), .B2(n8104), .A(n8103), .ZN(n8108) );
  OAI21_X1 U9194 ( .B1(n6442), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n8120), .ZN(
        n8121) );
  NAND2_X1 U9195 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n7342) );
  XNOR2_X1 U9196 ( .A(n10770), .B(n10764), .ZN(n15181) );
  XNOR2_X1 U9197 ( .A(n11732), .B(n6685), .ZN(n11730) );
  INV_X1 U9198 ( .A(n11733), .ZN(n6685) );
  NAND2_X1 U9199 ( .A1(n7185), .A2(n11285), .ZN(n11495) );
  NAND2_X1 U9200 ( .A1(n11497), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n11498) );
  AND2_X1 U9201 ( .A1(n15186), .A2(n7462), .ZN(n7463) );
  INV_X1 U9202 ( .A(n15194), .ZN(n7462) );
  NAND2_X1 U9203 ( .A1(n15195), .A2(n15194), .ZN(n7145) );
  INV_X1 U9204 ( .A(n15220), .ZN(n7465) );
  NAND2_X1 U9205 ( .A1(n15221), .A2(n15220), .ZN(n15225) );
  OAI211_X1 U9206 ( .C1(n15239), .C2(n7186), .A(n7149), .B(n7148), .ZN(n15247)
         );
  NAND2_X1 U9207 ( .A1(n7150), .A2(n15246), .ZN(n7149) );
  NOR2_X1 U9208 ( .A1(n15247), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n15249) );
  CLKBUF_X2 U9209 ( .A(n12647), .Z(P3_U3897) );
  NAND2_X1 U9210 ( .A1(n7797), .A2(n11420), .ZN(n11166) );
  XNOR2_X1 U9211 ( .A(n7203), .B(n7839), .ZN(n12621) );
  AOI21_X1 U9212 ( .B1(n6820), .B2(n6819), .A(n6818), .ZN(n6817) );
  INV_X1 U9213 ( .A(n12369), .ZN(n6818) );
  AOI21_X1 U9214 ( .B1(n10935), .B2(n10803), .A(n10802), .ZN(n10805) );
  NAND2_X1 U9215 ( .A1(n7389), .A2(n7388), .ZN(n10809) );
  AOI21_X1 U9216 ( .B1(n6875), .B2(n12692), .A(n6873), .ZN(n12753) );
  NAND2_X1 U9217 ( .A1(n7247), .A2(n7246), .ZN(P3_U3201) );
  AOI21_X1 U9218 ( .B1(n7654), .B2(n12692), .A(n10247), .ZN(n7246) );
  AND3_X1 U9219 ( .A1(n7648), .A2(n7652), .A3(n7393), .ZN(n7247) );
  AOI21_X1 U9220 ( .B1(n6708), .B2(n15599), .A(n6706), .ZN(n12452) );
  OR2_X1 U9221 ( .A1(n12451), .A2(n6707), .ZN(n6706) );
  NAND2_X1 U9222 ( .A1(n7868), .A2(n7865), .ZN(n6708) );
  NAND2_X1 U9223 ( .A1(n7421), .A2(n7420), .ZN(n13029) );
  NAND2_X1 U9224 ( .A1(n15674), .A2(n13027), .ZN(n7420) );
  NAND2_X1 U9225 ( .A1(n12801), .A2(n13115), .ZN(n7232) );
  NAND2_X1 U9226 ( .A1(n6681), .A2(n15666), .ZN(n6680) );
  NAND2_X1 U9227 ( .A1(n12801), .A2(n13217), .ZN(n7231) );
  INV_X1 U9228 ( .A(n7287), .ZN(n7286) );
  NAND2_X1 U9229 ( .A1(n7291), .A2(n11137), .ZN(n7290) );
  NOR2_X1 U9230 ( .A1(n6526), .A2(n7240), .ZN(n7239) );
  NOR2_X1 U9231 ( .A1(n15580), .A2(n10280), .ZN(n7240) );
  AOI21_X1 U9232 ( .B1(n14315), .B2(n15580), .A(n10294), .ZN(n10295) );
  OAI22_X1 U9233 ( .A1(n14318), .A2(n14294), .B1(n15580), .B2(n10293), .ZN(
        n10294) );
  AND2_X1 U9234 ( .A1(n10259), .A2(n7180), .ZN(n7179) );
  NAND2_X1 U9235 ( .A1(n7182), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7180) );
  NAND2_X1 U9236 ( .A1(n8667), .A2(n15571), .ZN(n7494) );
  OAI21_X1 U9237 ( .B1(n10279), .B2(n7182), .A(n7274), .ZN(P2_U3495) );
  NOR2_X1 U9238 ( .A1(n6525), .A2(n7275), .ZN(n7274) );
  NOR2_X1 U9239 ( .A1(n15571), .A2(n10278), .ZN(n7275) );
  OAI21_X1 U9240 ( .B1(n14315), .B2(n7182), .A(n7212), .ZN(n14317) );
  NAND2_X1 U9241 ( .A1(n7182), .A2(n14316), .ZN(n7212) );
  NAND2_X1 U9242 ( .A1(n6804), .A2(n6801), .ZN(P2_U3492) );
  INV_X1 U9243 ( .A(n6802), .ZN(n6801) );
  NAND2_X1 U9244 ( .A1(n14320), .A2(n15571), .ZN(n6804) );
  OAI21_X1 U9245 ( .B1(n14321), .B2(n14350), .A(n6803), .ZN(n6802) );
  XNOR2_X1 U9246 ( .A(n7221), .B(n6500), .ZN(n14485) );
  INV_X1 U9247 ( .A(n6699), .ZN(n6698) );
  OAI21_X1 U9248 ( .B1(n15287), .B2(n14648), .A(n14647), .ZN(n6699) );
  OAI21_X1 U9249 ( .B1(n15025), .B2(n14990), .A(n7355), .ZN(P1_U3266) );
  INV_X1 U9250 ( .A(n7356), .ZN(n7355) );
  OAI21_X1 U9251 ( .B1(n15029), .B2(n15336), .A(n7357), .ZN(n7356) );
  AOI21_X1 U9252 ( .B1(n15026), .B2(n15332), .A(n14773), .ZN(n7357) );
  OR2_X1 U9253 ( .A1(n15017), .A2(n6911), .ZN(n6913) );
  AOI21_X1 U9254 ( .B1(n6446), .B2(n6479), .A(n6649), .ZN(n6910) );
  NAND2_X1 U9255 ( .A1(n15443), .A2(n15359), .ZN(n6911) );
  NAND2_X1 U9256 ( .A1(n6446), .A2(n15402), .ZN(n6912) );
  OR2_X1 U9257 ( .A1(n7163), .A2(n7164), .ZN(n10754) );
  INV_X1 U9258 ( .A(n7458), .ZN(n7163) );
  NAND2_X1 U9259 ( .A1(n7146), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n10779) );
  INV_X1 U9260 ( .A(n7166), .ZN(n7146) );
  AND4_X1 U9261 ( .A1(n12333), .A2(n12997), .A3(n12332), .A4(n12331), .ZN(
        n6450) );
  OAI211_X2 U9262 ( .C1(n10974), .C2(n11710), .A(n7035), .B(n7036), .ZN(n10002) );
  AND2_X1 U9263 ( .A1(n6589), .A2(n7044), .ZN(n6451) );
  NOR2_X1 U9264 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n6452) );
  INV_X2 U9265 ( .A(n6443), .ZN(n10339) );
  NAND2_X1 U9266 ( .A1(n8202), .A2(n10338), .ZN(n8123) );
  INV_X2 U9267 ( .A(n10085), .ZN(n10124) );
  AND2_X1 U9268 ( .A1(n11251), .A2(n15380), .ZN(n6454) );
  INV_X1 U9269 ( .A(n14944), .ZN(n6927) );
  OR2_X1 U9270 ( .A1(n10219), .A2(n10433), .ZN(n6455) );
  OAI211_X1 U9271 ( .C1(n8123), .C2(n10318), .A(n8153), .B(n8152), .ZN(n13762)
         );
  AND2_X1 U9272 ( .A1(n6559), .A2(n8580), .ZN(n6456) );
  INV_X1 U9273 ( .A(n12615), .ZN(n7839) );
  NOR2_X1 U9274 ( .A1(n12323), .A2(n12327), .ZN(n6457) );
  AND2_X1 U9275 ( .A1(n10239), .A2(n10157), .ZN(n6459) );
  AND2_X1 U9276 ( .A1(n8583), .A2(n6456), .ZN(n6460) );
  NAND2_X1 U9277 ( .A1(n8506), .A2(n8505), .ZN(n13811) );
  INV_X1 U9278 ( .A(n8598), .ZN(n6769) );
  INV_X1 U9279 ( .A(n7783), .ZN(n7782) );
  NAND2_X1 U9280 ( .A1(n7784), .A2(n12201), .ZN(n7783) );
  AND2_X1 U9281 ( .A1(n7925), .A2(n7924), .ZN(n6461) );
  AND2_X1 U9282 ( .A1(n15289), .A2(n7714), .ZN(n6462) );
  NOR2_X1 U9283 ( .A1(n6714), .A2(n6713), .ZN(n6463) );
  AND2_X1 U9284 ( .A1(n7928), .A2(n7694), .ZN(n6464) );
  AND2_X1 U9285 ( .A1(n6581), .A2(n7050), .ZN(n6465) );
  NAND2_X1 U9286 ( .A1(n10973), .A2(n10974), .ZN(n9560) );
  NOR2_X1 U9287 ( .A1(n6562), .A2(n7504), .ZN(n6466) );
  NAND2_X1 U9288 ( .A1(n8013), .A2(SI_21_), .ZN(n8431) );
  AND2_X1 U9289 ( .A1(n11588), .A2(n7921), .ZN(n6467) );
  AND2_X1 U9290 ( .A1(n14740), .A2(n9925), .ZN(n6468) );
  AND4_X1 U9291 ( .A1(n6947), .A2(n6946), .A3(n8036), .A4(n8348), .ZN(n6469)
         );
  NAND2_X1 U9292 ( .A1(n8354), .A2(n8353), .ZN(n14166) );
  OR2_X1 U9293 ( .A1(n13623), .A2(n13620), .ZN(n6470) );
  XNOR2_X1 U9294 ( .A(n8008), .B(SI_19_), .ZN(n8398) );
  INV_X1 U9295 ( .A(n7403), .ZN(n7402) );
  NAND2_X1 U9296 ( .A1(n9236), .A2(n9232), .ZN(n7403) );
  INV_X1 U9297 ( .A(n7454), .ZN(n7453) );
  NAND2_X1 U9298 ( .A1(n11498), .A2(n7455), .ZN(n7454) );
  AND2_X1 U9299 ( .A1(n12351), .A2(n12307), .ZN(n12310) );
  INV_X1 U9300 ( .A(n12310), .ZN(n12342) );
  AND2_X1 U9301 ( .A1(n6542), .A2(n8396), .ZN(n6471) );
  INV_X1 U9302 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n14356) );
  INV_X1 U9303 ( .A(n13718), .ZN(n13943) );
  NAND2_X1 U9304 ( .A1(n10252), .A2(n10251), .ZN(n13718) );
  INV_X1 U9305 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7913) );
  INV_X1 U9306 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8058) );
  AND2_X1 U9307 ( .A1(n10094), .A2(n7250), .ZN(n6472) );
  NAND2_X1 U9308 ( .A1(n12394), .A2(n7220), .ZN(n7889) );
  OR2_X1 U9309 ( .A1(n7380), .A2(n7378), .ZN(n6473) );
  AND2_X1 U9310 ( .A1(n13652), .A2(n6594), .ZN(n6474) );
  NAND2_X1 U9311 ( .A1(n9325), .A2(n9324), .ZN(n15121) );
  INV_X1 U9312 ( .A(n15121), .ZN(n7770) );
  AND3_X1 U9313 ( .A1(n6983), .A2(n6638), .A3(n6984), .ZN(n6475) );
  AND2_X1 U9314 ( .A1(n12259), .A2(n12251), .ZN(n6476) );
  AND2_X1 U9315 ( .A1(n7756), .A2(n7755), .ZN(n6477) );
  INV_X1 U9316 ( .A(n8745), .ZN(n6892) );
  NAND2_X1 U9317 ( .A1(n10316), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8745) );
  INV_X1 U9318 ( .A(n8558), .ZN(n13761) );
  AND2_X1 U9319 ( .A1(n11113), .A2(n7759), .ZN(n6478) );
  NOR2_X1 U9320 ( .A1(n15422), .A2(n15440), .ZN(n6479) );
  AOI21_X1 U9321 ( .B1(n8027), .B2(n8494), .A(n6648), .ZN(n7602) );
  INV_X1 U9322 ( .A(n12722), .ZN(n7639) );
  INV_X1 U9323 ( .A(n12716), .ZN(n7368) );
  NAND2_X1 U9324 ( .A1(n7651), .A2(n10199), .ZN(n6480) );
  INV_X1 U9325 ( .A(n10593), .ZN(n6964) );
  AND2_X1 U9326 ( .A1(n7078), .A2(n6941), .ZN(n6481) );
  INV_X1 U9327 ( .A(n12063), .ZN(n7134) );
  NAND2_X1 U9328 ( .A1(n12483), .A2(n13070), .ZN(n6482) );
  NAND2_X1 U9329 ( .A1(n9179), .A2(n9178), .ZN(n13046) );
  INV_X1 U9330 ( .A(n9444), .ZN(n9886) );
  NOR2_X1 U9331 ( .A1(n14081), .A2(n7507), .ZN(n6483) );
  AND2_X1 U9332 ( .A1(n7556), .A2(n8281), .ZN(n6484) );
  INV_X1 U9333 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8149) );
  AND2_X1 U9334 ( .A1(n7298), .A2(n8251), .ZN(n6485) );
  INV_X1 U9335 ( .A(n12030), .ZN(n7695) );
  NAND2_X1 U9336 ( .A1(n6879), .A2(n6877), .ZN(n9064) );
  INV_X1 U9337 ( .A(n13983), .ZN(n7500) );
  OR2_X1 U9338 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10174), .ZN(n6486) );
  AND2_X1 U9339 ( .A1(n7547), .A2(n7545), .ZN(n6487) );
  NAND2_X1 U9340 ( .A1(n13730), .A2(n13723), .ZN(n6488) );
  AND2_X1 U9341 ( .A1(n14687), .A2(n14772), .ZN(n6489) );
  AND2_X1 U9342 ( .A1(n13580), .A2(n13579), .ZN(n6490) );
  AND2_X1 U9343 ( .A1(n7219), .A2(n10270), .ZN(n6491) );
  INV_X1 U9344 ( .A(n11088), .ZN(n6856) );
  AND2_X1 U9345 ( .A1(n15083), .A2(n14902), .ZN(n6492) );
  AND2_X1 U9346 ( .A1(n12294), .A2(n10437), .ZN(n6493) );
  NOR2_X1 U9347 ( .A1(n9267), .A2(n7415), .ZN(n6494) );
  NAND2_X1 U9348 ( .A1(n13508), .A2(n13300), .ZN(n10876) );
  INV_X1 U9349 ( .A(n7352), .ZN(n7351) );
  OAI21_X1 U9350 ( .B1(n12026), .B2(n7353), .A(n12045), .ZN(n7352) );
  AND2_X1 U9351 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_27__SCAN_IN), .ZN(
        n6495) );
  AND2_X1 U9352 ( .A1(n12556), .A2(n7840), .ZN(n6496) );
  AND2_X1 U9353 ( .A1(n10211), .A2(n10803), .ZN(n6497) );
  AND2_X1 U9354 ( .A1(n7388), .A2(n7387), .ZN(n6498) );
  INV_X1 U9355 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n7647) );
  OR3_X1 U9356 ( .A1(n9473), .A2(n9373), .A3(n7041), .ZN(n6499) );
  XOR2_X1 U9357 ( .A(n12404), .B(n12405), .Z(n6500) );
  AND2_X1 U9358 ( .A1(n9317), .A2(n9316), .ZN(n6501) );
  INV_X1 U9359 ( .A(n6721), .ZN(n9675) );
  NOR2_X1 U9360 ( .A1(n9636), .A2(n9616), .ZN(n6721) );
  OAI211_X1 U9361 ( .C1(n9907), .C2(n10343), .A(n7700), .B(n7701), .ZN(n7699)
         );
  NAND2_X1 U9362 ( .A1(n10161), .A2(n10565), .ZN(n7265) );
  INV_X1 U9363 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8678) );
  AND2_X1 U9364 ( .A1(n11317), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6502) );
  AND2_X1 U9365 ( .A1(n6455), .A2(n7384), .ZN(n6503) );
  AND2_X1 U9366 ( .A1(n7771), .A2(n7770), .ZN(n6504) );
  INV_X1 U9367 ( .A(n11494), .ZN(n7451) );
  AND2_X1 U9368 ( .A1(n6483), .A2(n8597), .ZN(n6505) );
  NAND2_X1 U9369 ( .A1(n8248), .A2(n8247), .ZN(n13567) );
  INV_X1 U9370 ( .A(n13567), .ZN(n7921) );
  AND2_X1 U9371 ( .A1(n13576), .A2(n13575), .ZN(n6506) );
  OR2_X1 U9372 ( .A1(n13200), .A2(n12953), .ZN(n12219) );
  INV_X1 U9373 ( .A(n7838), .ZN(n7837) );
  NAND2_X1 U9374 ( .A1(n6496), .A2(n7839), .ZN(n7838) );
  NAND2_X1 U9375 ( .A1(n6931), .A2(n14693), .ZN(n14927) );
  NAND2_X1 U9376 ( .A1(n8220), .A2(n8219), .ZN(n14301) );
  INV_X1 U9377 ( .A(n14301), .ZN(n7920) );
  OR2_X1 U9378 ( .A1(n8019), .A2(n7586), .ZN(n6507) );
  AND2_X1 U9379 ( .A1(n9099), .A2(n10218), .ZN(n6508) );
  INV_X1 U9380 ( .A(n13988), .ZN(n7917) );
  INV_X1 U9381 ( .A(n8605), .ZN(n7499) );
  AND4_X1 U9382 ( .A1(n14752), .A2(n9910), .A3(n14790), .A4(n14779), .ZN(n6509) );
  INV_X1 U9383 ( .A(n14772), .ZN(n7711) );
  AND3_X1 U9384 ( .A1(n14779), .A2(n7128), .A3(n14683), .ZN(n6510) );
  AND4_X1 U9385 ( .A1(n8674), .A2(n8673), .A3(n9022), .A4(n8672), .ZN(n6511)
         );
  OR2_X1 U9386 ( .A1(n14184), .A2(n14191), .ZN(n6512) );
  AND2_X1 U9387 ( .A1(n10680), .A2(n10672), .ZN(n6513) );
  OR2_X1 U9388 ( .A1(n12230), .A2(n12932), .ZN(n6514) );
  NAND2_X1 U9389 ( .A1(n14843), .A2(n14842), .ZN(n14844) );
  AND2_X1 U9390 ( .A1(n13002), .A2(n13119), .ZN(n6515) );
  AND2_X1 U9391 ( .A1(n6467), .A2(n7920), .ZN(n6516) );
  NOR2_X1 U9392 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n8549) );
  INV_X1 U9393 ( .A(n14695), .ZN(n6926) );
  AND2_X1 U9394 ( .A1(n13585), .A2(n11866), .ZN(n6517) );
  AND2_X1 U9395 ( .A1(n12012), .A2(n7713), .ZN(n6518) );
  OR2_X1 U9396 ( .A1(n11226), .A2(n11225), .ZN(n6519) );
  AND2_X1 U9397 ( .A1(n14818), .A2(n14710), .ZN(n6520) );
  AND3_X1 U9398 ( .A1(n10000), .A2(n9998), .A3(n9999), .ZN(n6521) );
  AND2_X1 U9399 ( .A1(n13299), .A2(n13298), .ZN(n6522) );
  AND3_X1 U9400 ( .A1(n9307), .A2(n9308), .A3(n9335), .ZN(n6523) );
  AND2_X1 U9401 ( .A1(n7920), .A2(n13822), .ZN(n6524) );
  INV_X1 U9402 ( .A(n14127), .ZN(n7923) );
  NOR2_X1 U9403 ( .A1(n13966), .A2(n14350), .ZN(n6525) );
  NOR2_X1 U9404 ( .A1(n13966), .A2(n14294), .ZN(n6526) );
  AND2_X1 U9405 ( .A1(n7147), .A2(n15246), .ZN(n6527) );
  INV_X1 U9406 ( .A(n11250), .ZN(n15380) );
  AND2_X1 U9407 ( .A1(n13036), .A2(n15638), .ZN(n6528) );
  INV_X1 U9408 ( .A(n14692), .ZN(n15095) );
  NAND2_X1 U9409 ( .A1(n9615), .A2(n9614), .ZN(n14692) );
  INV_X1 U9410 ( .A(n14184), .ZN(n14351) );
  NAND2_X1 U9411 ( .A1(n8322), .A2(n8321), .ZN(n14184) );
  INV_X1 U9412 ( .A(n14047), .ZN(n14227) );
  NAND2_X1 U9413 ( .A1(n8467), .A2(n8466), .ZN(n14047) );
  NAND2_X2 U9414 ( .A1(n9883), .A2(n9882), .ZN(n14748) );
  AND2_X1 U9415 ( .A1(n7075), .A2(n7073), .ZN(n6529) );
  AND2_X1 U9416 ( .A1(n7414), .A2(n7412), .ZN(n6530) );
  AND2_X1 U9417 ( .A1(n7646), .A2(P3_IR_REG_2__SCAN_IN), .ZN(n6531) );
  INV_X1 U9418 ( .A(n10093), .ZN(n7045) );
  NAND2_X1 U9419 ( .A1(n15058), .A2(n14870), .ZN(n6532) );
  OR2_X1 U9420 ( .A1(n11902), .A2(n12148), .ZN(n6533) );
  INV_X1 U9421 ( .A(n15126), .ZN(n7772) );
  NAND2_X1 U9422 ( .A1(n9379), .A2(n9378), .ZN(n15126) );
  AND2_X1 U9423 ( .A1(n7723), .A2(n14680), .ZN(n6534) );
  AND2_X1 U9424 ( .A1(n7143), .A2(n14677), .ZN(n6535) );
  AND2_X1 U9425 ( .A1(n13789), .A2(n8613), .ZN(n6536) );
  AND2_X1 U9426 ( .A1(n8565), .A2(n8564), .ZN(n6537) );
  NAND2_X1 U9427 ( .A1(n8526), .A2(n8525), .ZN(n13720) );
  INV_X1 U9428 ( .A(n7318), .ZN(n7317) );
  OAI21_X1 U9429 ( .B1(n8398), .B2(n7319), .A(n8010), .ZN(n7318) );
  AND2_X1 U9430 ( .A1(n14047), .A2(n14024), .ZN(n6538) );
  AND2_X1 U9431 ( .A1(n7066), .A2(n7525), .ZN(n6539) );
  OR2_X1 U9432 ( .A1(n12502), .A2(n12822), .ZN(n6540) );
  OR2_X1 U9433 ( .A1(n10131), .A2(n10133), .ZN(n6541) );
  INV_X1 U9434 ( .A(n7560), .ZN(n7559) );
  OAI21_X1 U9435 ( .B1(n14052), .B2(n7561), .A(n8476), .ZN(n7560) );
  OR2_X1 U9436 ( .A1(n14105), .A2(n13814), .ZN(n6542) );
  OR2_X1 U9437 ( .A1(n14321), .A2(n13986), .ZN(n6543) );
  INV_X1 U9438 ( .A(n14073), .ZN(n7918) );
  AND2_X1 U9439 ( .A1(n8207), .A2(n8209), .ZN(n6544) );
  AND2_X1 U9440 ( .A1(n8802), .A2(n7884), .ZN(n6545) );
  AND2_X1 U9441 ( .A1(n7360), .A2(n7366), .ZN(n6546) );
  NAND2_X1 U9442 ( .A1(n8432), .A2(n8416), .ZN(n6547) );
  AND4_X1 U9443 ( .A1(n10060), .A2(n10059), .A3(n10058), .A4(n10057), .ZN(
        n6548) );
  NOR2_X1 U9444 ( .A1(n14296), .A2(n13819), .ZN(n6549) );
  AND2_X1 U9445 ( .A1(n8621), .A2(n8620), .ZN(n6550) );
  INV_X1 U9446 ( .A(n7512), .ZN(n7511) );
  NOR2_X1 U9447 ( .A1(n14197), .A2(n13819), .ZN(n7512) );
  INV_X1 U9448 ( .A(n14740), .ZN(n7109) );
  AND2_X1 U9449 ( .A1(n13122), .A2(n12998), .ZN(n6551) );
  AND2_X1 U9450 ( .A1(n11911), .A2(n12998), .ZN(n6552) );
  NOR2_X1 U9451 ( .A1(n14166), .A2(n8585), .ZN(n6553) );
  NOR2_X1 U9452 ( .A1(n15126), .A2(n14502), .ZN(n6554) );
  NOR2_X1 U9453 ( .A1(n15103), .A2(n14690), .ZN(n6555) );
  NOR2_X1 U9454 ( .A1(n15076), .A2(n14698), .ZN(n6556) );
  NOR2_X1 U9455 ( .A1(n14505), .A2(n15397), .ZN(n6557) );
  NOR2_X1 U9456 ( .A1(n6594), .A2(n13652), .ZN(n6558) );
  OR2_X1 U9457 ( .A1(n14296), .A2(n13775), .ZN(n6559) );
  INV_X1 U9458 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8253) );
  OR2_X1 U9459 ( .A1(n6496), .A2(n7832), .ZN(n6560) );
  AND2_X1 U9460 ( .A1(n7450), .A2(n7452), .ZN(n6561) );
  AND2_X1 U9461 ( .A1(n14098), .A2(n6505), .ZN(n6562) );
  AND2_X1 U9462 ( .A1(n13046), .A2(n13035), .ZN(n6563) );
  INV_X1 U9463 ( .A(n10109), .ZN(n7051) );
  INV_X1 U9464 ( .A(n7557), .ZN(n6761) );
  NAND2_X1 U9465 ( .A1(n14210), .A2(n14004), .ZN(n7557) );
  NAND2_X1 U9466 ( .A1(n7500), .A2(n7501), .ZN(n6564) );
  NAND2_X1 U9467 ( .A1(n7433), .A2(n6978), .ZN(n7437) );
  AND2_X1 U9468 ( .A1(n13548), .A2(n13547), .ZN(n6565) );
  INV_X1 U9469 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8370) );
  NOR2_X1 U9470 ( .A1(n7753), .A2(n10111), .ZN(n6566) );
  AND2_X1 U9471 ( .A1(n12485), .A2(n12908), .ZN(n6567) );
  NAND2_X1 U9472 ( .A1(n11588), .A2(n13824), .ZN(n6568) );
  AND4_X1 U9473 ( .A1(n8036), .A2(n8348), .A3(n8285), .A4(n8058), .ZN(n6569)
         );
  INV_X1 U9474 ( .A(n12010), .ZN(n7716) );
  INV_X1 U9475 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n15801) );
  OR2_X1 U9476 ( .A1(n15373), .A2(n14508), .ZN(n6570) );
  AND2_X1 U9477 ( .A1(n12475), .A2(n12641), .ZN(n6571) );
  OR2_X1 U9478 ( .A1(n10132), .A2(n6541), .ZN(n6572) );
  AND2_X1 U9479 ( .A1(n12815), .A2(n12261), .ZN(n6573) );
  AND2_X1 U9480 ( .A1(n7030), .A2(n7032), .ZN(n6574) );
  AND2_X1 U9481 ( .A1(n15027), .A2(n14783), .ZN(n6575) );
  INV_X1 U9482 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10317) );
  INV_X1 U9483 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10326) );
  INV_X1 U9484 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10346) );
  INV_X1 U9485 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10319) );
  INV_X1 U9486 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10401) );
  INV_X1 U9487 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8043) );
  NAND2_X1 U9488 ( .A1(n14748), .A2(n14686), .ZN(n6576) );
  INV_X1 U9489 ( .A(n8007), .ZN(n7321) );
  NAND2_X1 U9490 ( .A1(n12180), .A2(n12187), .ZN(n6577) );
  INV_X1 U9491 ( .A(n10987), .ZN(n11710) );
  INV_X1 U9492 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10411) );
  INV_X1 U9493 ( .A(n7882), .ZN(n7881) );
  NAND2_X1 U9494 ( .A1(n12248), .A2(n7883), .ZN(n7882) );
  AND2_X1 U9495 ( .A1(n6715), .A2(n6490), .ZN(n6578) );
  NAND2_X1 U9496 ( .A1(n6758), .A2(n6756), .ZN(n10275) );
  NAND2_X1 U9497 ( .A1(n14835), .A2(n14822), .ZN(n14808) );
  INV_X1 U9498 ( .A(n14808), .ZN(n7754) );
  OR2_X1 U9499 ( .A1(n12887), .A2(n6866), .ZN(n6579) );
  NOR2_X1 U9500 ( .A1(n10218), .A2(n15672), .ZN(n6580) );
  OR2_X1 U9501 ( .A1(n10112), .A2(n10110), .ZN(n6581) );
  NAND2_X1 U9502 ( .A1(n12172), .A2(n12161), .ZN(n6582) );
  INV_X1 U9503 ( .A(n8595), .ZN(n7507) );
  INV_X1 U9504 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8846) );
  INV_X1 U9505 ( .A(n6719), .ZN(n9874) );
  NOR2_X1 U9506 ( .A1(n9835), .A2(n9834), .ZN(n6719) );
  OR2_X1 U9507 ( .A1(n8771), .A2(n7660), .ZN(n6583) );
  NAND2_X1 U9508 ( .A1(n14058), .A2(n6956), .ZN(n14007) );
  INV_X1 U9509 ( .A(n10094), .ZN(n7749) );
  NAND2_X1 U9510 ( .A1(n12873), .A2(n12246), .ZN(n6584) );
  NOR2_X1 U9511 ( .A1(n12318), .A2(n12317), .ZN(n6585) );
  OR2_X1 U9512 ( .A1(n7964), .A2(SI_6_), .ZN(n6586) );
  NAND2_X1 U9513 ( .A1(n8091), .A2(n8090), .ZN(n13515) );
  INV_X1 U9514 ( .A(n7104), .ZN(n7103) );
  NAND2_X1 U9515 ( .A1(n8431), .A2(n10964), .ZN(n7104) );
  OR2_X1 U9516 ( .A1(n8582), .A2(n7512), .ZN(n6587) );
  NAND2_X1 U9517 ( .A1(n12395), .A2(n7223), .ZN(n12394) );
  INV_X1 U9518 ( .A(n8398), .ZN(n7320) );
  NAND2_X1 U9519 ( .A1(n12815), .A2(n12259), .ZN(n6588) );
  NAND2_X1 U9520 ( .A1(n7749), .A2(n10095), .ZN(n6589) );
  AND3_X1 U9521 ( .A1(n13061), .A2(n13050), .A3(n12269), .ZN(n6590) );
  NAND2_X1 U9522 ( .A1(n14092), .A2(n13659), .ZN(n6591) );
  OR2_X1 U9523 ( .A1(n13660), .A2(n13661), .ZN(n6592) );
  OR2_X1 U9524 ( .A1(n9456), .A2(n9455), .ZN(n6593) );
  AND2_X1 U9525 ( .A1(n13650), .A2(n13649), .ZN(n6594) );
  NAND2_X1 U9526 ( .A1(n8601), .A2(n13999), .ZN(n14020) );
  INV_X1 U9527 ( .A(n14020), .ZN(n6743) );
  AND2_X1 U9528 ( .A1(n14721), .A2(n14719), .ZN(n6595) );
  AND2_X1 U9529 ( .A1(n6885), .A2(n6884), .ZN(n6596) );
  OR2_X1 U9530 ( .A1(n11744), .A2(n12998), .ZN(n12204) );
  INV_X1 U9531 ( .A(n12204), .ZN(n7870) );
  OR2_X1 U9532 ( .A1(n13557), .A2(n13555), .ZN(n6597) );
  XNOR2_X1 U9533 ( .A(n14092), .B(n13659), .ZN(n14081) );
  OR2_X1 U9534 ( .A1(n6565), .A2(n13550), .ZN(n6598) );
  OR2_X1 U9535 ( .A1(n7993), .A2(SI_14_), .ZN(n6599) );
  AND2_X1 U9536 ( .A1(n7856), .A2(n12219), .ZN(n6600) );
  AND2_X1 U9537 ( .A1(n12341), .A2(n12771), .ZN(n6601) );
  AND3_X1 U9538 ( .A1(n8092), .A2(n8095), .A3(n8094), .ZN(n6602) );
  AND3_X1 U9539 ( .A1(n12171), .A2(n12162), .A3(n10853), .ZN(n6603) );
  AND2_X1 U9540 ( .A1(n7819), .A2(n12486), .ZN(n6604) );
  AND2_X1 U9541 ( .A1(n13034), .A2(n12822), .ZN(n6605) );
  AND2_X1 U9542 ( .A1(n9941), .A2(n11513), .ZN(n6606) );
  AND2_X1 U9543 ( .A1(n10644), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6607) );
  OR2_X1 U9544 ( .A1(n15518), .A2(n13761), .ZN(n13300) );
  AND2_X1 U9545 ( .A1(n12637), .A2(n9154), .ZN(n6608) );
  INV_X1 U9546 ( .A(n9751), .ZN(n6997) );
  AND2_X1 U9547 ( .A1(n8370), .A2(n8550), .ZN(n6609) );
  OR2_X1 U9548 ( .A1(n12618), .A2(n12801), .ZN(n6610) );
  AND2_X1 U9549 ( .A1(n7320), .A2(n8006), .ZN(n6611) );
  INV_X1 U9550 ( .A(n9230), .ZN(n7779) );
  INV_X1 U9551 ( .A(n7571), .ZN(n7570) );
  NOR2_X1 U9552 ( .A1(n8269), .A2(n7572), .ZN(n7571) );
  AND2_X1 U9553 ( .A1(n7523), .A2(n7521), .ZN(n6612) );
  NAND2_X1 U9554 ( .A1(n14217), .A2(n14041), .ZN(n6613) );
  INV_X1 U9555 ( .A(n15628), .ZN(n12645) );
  NAND2_X1 U9556 ( .A1(n14073), .A2(n13501), .ZN(n6614) );
  AND2_X1 U9557 ( .A1(n12591), .A2(n7822), .ZN(n7821) );
  AND2_X1 U9558 ( .A1(n7283), .A2(n13758), .ZN(n6615) );
  OR2_X1 U9559 ( .A1(n14763), .A2(n14748), .ZN(n6616) );
  AND2_X1 U9560 ( .A1(n8753), .A2(n8750), .ZN(n6617) );
  AND2_X1 U9561 ( .A1(n9702), .A2(n9689), .ZN(n6618) );
  OR2_X1 U9562 ( .A1(n10106), .A2(n10104), .ZN(n6619) );
  OR2_X1 U9563 ( .A1(n10123), .A2(n10121), .ZN(n6620) );
  OR2_X1 U9564 ( .A1(n10020), .A2(n10018), .ZN(n6621) );
  NAND2_X1 U9565 ( .A1(n12324), .A2(n12182), .ZN(n6622) );
  AND2_X1 U9566 ( .A1(n7841), .A2(n6540), .ZN(n6623) );
  AND2_X1 U9567 ( .A1(n7465), .A2(n15211), .ZN(n6624) );
  INV_X1 U9568 ( .A(n7130), .ZN(n7129) );
  NOR2_X1 U9569 ( .A1(n15040), .A2(n14711), .ZN(n7130) );
  OR2_X1 U9570 ( .A1(n13683), .A2(n7227), .ZN(n6625) );
  AND2_X1 U9571 ( .A1(n6497), .A2(n7390), .ZN(n6626) );
  AND2_X1 U9572 ( .A1(n13684), .A2(n6726), .ZN(n6627) );
  OAI21_X1 U9573 ( .B1(n6769), .B2(n14055), .A(n8599), .ZN(n6768) );
  AND2_X1 U9574 ( .A1(n7080), .A2(n8005), .ZN(n6628) );
  NAND2_X1 U9575 ( .A1(n12533), .A2(n12618), .ZN(n6629) );
  NAND2_X1 U9576 ( .A1(n13535), .A2(n15496), .ZN(n8141) );
  NOR2_X1 U9577 ( .A1(n7938), .A2(n14829), .ZN(n6630) );
  NOR2_X1 U9578 ( .A1(n10136), .A2(n10135), .ZN(n6631) );
  NAND2_X1 U9579 ( .A1(n14212), .A2(n14271), .ZN(n6632) );
  INV_X1 U9580 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8802) );
  AND2_X1 U9581 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_5__SCAN_IN), 
        .ZN(n6633) );
  INV_X1 U9582 ( .A(n8004), .ZN(n7081) );
  NAND2_X1 U9583 ( .A1(n10327), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8748) );
  INV_X1 U9584 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n10360) );
  INV_X1 U9585 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9310) );
  XNOR2_X1 U9586 ( .A(n15250), .B(n15245), .ZN(n15246) );
  INV_X1 U9587 ( .A(n15246), .ZN(n7186) );
  OR2_X1 U9588 ( .A1(n12337), .A2(n6691), .ZN(n6634) );
  INV_X1 U9589 ( .A(n15329), .ZN(n11113) );
  INV_X1 U9590 ( .A(n12884), .ZN(n6867) );
  INV_X1 U9591 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6966) );
  NAND2_X1 U9592 ( .A1(n11208), .A2(n8141), .ZN(n15480) );
  NAND2_X1 U9593 ( .A1(n7629), .A2(n6841), .ZN(n6635) );
  NAND2_X1 U9594 ( .A1(n12069), .A2(n12063), .ZN(n12073) );
  NAND2_X1 U9595 ( .A1(n14193), .A2(n7925), .ZN(n14145) );
  OAI21_X1 U9596 ( .B1(n12073), .B2(n7707), .A(n7704), .ZN(n14942) );
  NAND2_X1 U9597 ( .A1(n11415), .A2(n6958), .ZN(n6636) );
  NAND2_X1 U9598 ( .A1(n14193), .A2(n14351), .ZN(n6637) );
  NAND2_X1 U9599 ( .A1(n7297), .A2(n8210), .ZN(n11693) );
  NAND2_X1 U9600 ( .A1(n8042), .A2(n8626), .ZN(n8630) );
  NAND2_X1 U9601 ( .A1(n6905), .A2(n9154), .ZN(n13056) );
  NAND2_X1 U9602 ( .A1(n6770), .A2(n8195), .ZN(n11413) );
  NAND2_X1 U9603 ( .A1(n7345), .A2(n11255), .ZN(n11821) );
  NAND2_X1 U9604 ( .A1(n7401), .A2(n7398), .ZN(n12996) );
  NAND2_X1 U9605 ( .A1(n11607), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6638) );
  NAND2_X1 U9606 ( .A1(n8570), .A2(n8569), .ZN(n11410) );
  NAND2_X1 U9607 ( .A1(n6778), .A2(n7489), .ZN(n11895) );
  NAND2_X1 U9608 ( .A1(n11107), .A2(n11106), .ZN(n15319) );
  NAND2_X1 U9609 ( .A1(n7726), .A2(n11240), .ZN(n11828) );
  NAND2_X1 U9610 ( .A1(n7807), .A2(n11999), .ZN(n12466) );
  AND2_X1 U9611 ( .A1(n6985), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n6639) );
  INV_X1 U9612 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8687) );
  INV_X1 U9613 ( .A(n10233), .ZN(n6841) );
  AND2_X1 U9614 ( .A1(n11749), .A2(n11746), .ZN(n6640) );
  AND2_X1 U9615 ( .A1(n8539), .A2(n8031), .ZN(n8625) );
  AND2_X1 U9616 ( .A1(n12651), .A2(n12652), .ZN(n6641) );
  AND2_X1 U9617 ( .A1(n11850), .A2(n11848), .ZN(n6642) );
  OR3_X1 U9618 ( .A1(n9368), .A2(n9473), .A3(n7041), .ZN(n6643) );
  INV_X1 U9619 ( .A(n9925), .ZN(n7108) );
  INV_X1 U9620 ( .A(n7758), .ZN(n15313) );
  NAND2_X1 U9621 ( .A1(n11113), .A2(n7761), .ZN(n7758) );
  INV_X1 U9622 ( .A(n7768), .ZN(n14972) );
  NAND2_X1 U9623 ( .A1(n11825), .A2(n6504), .ZN(n7768) );
  NOR2_X1 U9624 ( .A1(n15290), .A2(n15289), .ZN(n15288) );
  NAND2_X1 U9625 ( .A1(n10151), .A2(n11840), .ZN(n6644) );
  NAND2_X1 U9626 ( .A1(n9204), .A2(n9203), .ZN(n12801) );
  AND2_X1 U9627 ( .A1(n8509), .A2(SI_27_), .ZN(n6645) );
  INV_X1 U9628 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9369) );
  AND2_X1 U9629 ( .A1(n10151), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n6646) );
  OR2_X1 U9630 ( .A1(n10185), .A2(n10184), .ZN(n6647) );
  AND2_X1 U9631 ( .A1(n8507), .A2(n13249), .ZN(n6648) );
  AND2_X1 U9632 ( .A1(n15440), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6649) );
  NOR2_X1 U9633 ( .A1(P3_REG0_REG_28__SCAN_IN), .A2(n15666), .ZN(n6650) );
  AND2_X1 U9634 ( .A1(n14126), .A2(n14262), .ZN(n14099) );
  INV_X1 U9635 ( .A(n7442), .ZN(n12666) );
  OR2_X1 U9636 ( .A1(n10154), .A2(n10233), .ZN(n7442) );
  INV_X1 U9637 ( .A(n8416), .ZN(n7311) );
  INV_X2 U9638 ( .A(n15664), .ZN(n15666) );
  OR2_X1 U9639 ( .A1(n15666), .A2(n13137), .ZN(n6651) );
  NOR2_X1 U9640 ( .A1(n15288), .A2(n7945), .ZN(n6652) );
  AND2_X1 U9641 ( .A1(n11536), .A2(n9229), .ZN(n6653) );
  NOR2_X1 U9642 ( .A1(n11841), .A2(n13001), .ZN(n6654) );
  AND2_X1 U9643 ( .A1(n6639), .A2(n10354), .ZN(n6655) );
  OR2_X1 U9644 ( .A1(n11672), .A2(n14292), .ZN(n6656) );
  INV_X1 U9645 ( .A(n15571), .ZN(n7182) );
  INV_X1 U9646 ( .A(n11432), .ZN(n7896) );
  INV_X1 U9647 ( .A(n15676), .ZN(n15674) );
  AND3_X2 U9648 ( .A1(n8730), .A2(n11390), .A3(n8729), .ZN(n15676) );
  OR2_X1 U9649 ( .A1(n10575), .A2(n10603), .ZN(n15493) );
  INV_X1 U9650 ( .A(n15493), .ZN(n14190) );
  AND2_X1 U9651 ( .A1(n14612), .A2(n14594), .ZN(n6657) );
  AND2_X2 U9652 ( .A1(n11396), .A2(n15588), .ZN(n15601) );
  AND2_X1 U9653 ( .A1(n15581), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n6658) );
  INV_X1 U9654 ( .A(n11137), .ZN(n13936) );
  AND2_X2 U9655 ( .A1(n10734), .A2(n8661), .ZN(n15580) );
  AND2_X1 U9656 ( .A1(n10581), .A2(n14366), .ZN(n15475) );
  NAND2_X1 U9657 ( .A1(n8336), .A2(n8335), .ZN(n14341) );
  INV_X1 U9658 ( .A(n14341), .ZN(n7924) );
  INV_X1 U9659 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6907) );
  AND2_X1 U9660 ( .A1(n12744), .A2(n6480), .ZN(n6659) );
  NAND2_X1 U9661 ( .A1(n9655), .A2(n9654), .ZN(n15088) );
  INV_X1 U9662 ( .A(n15088), .ZN(n7755) );
  INV_X1 U9663 ( .A(n12131), .ZN(n7062) );
  INV_X1 U9664 ( .A(n15389), .ZN(n7762) );
  INV_X1 U9665 ( .A(n15481), .ZN(n7178) );
  AND2_X1 U9666 ( .A1(n10241), .A2(n12722), .ZN(n6660) );
  NAND2_X1 U9667 ( .A1(n10855), .A2(n10857), .ZN(n10892) );
  AND2_X1 U9668 ( .A1(n13512), .A2(n7237), .ZN(n6661) );
  AND2_X1 U9669 ( .A1(n10632), .A2(n10599), .ZN(n6662) );
  AND2_X1 U9670 ( .A1(n12705), .A2(n10565), .ZN(n6663) );
  NAND2_X1 U9671 ( .A1(n11083), .A2(n11084), .ZN(n6664) );
  AND2_X1 U9672 ( .A1(n6857), .A2(n6856), .ZN(n6665) );
  AND2_X1 U9673 ( .A1(n12736), .A2(n10160), .ZN(n6666) );
  NOR2_X1 U9674 ( .A1(n7370), .A2(n12736), .ZN(n7369) );
  AND2_X1 U9675 ( .A1(n10974), .A2(n9941), .ZN(n6667) );
  NAND2_X1 U9676 ( .A1(n10224), .A2(n11466), .ZN(n6668) );
  NOR2_X1 U9677 ( .A1(n7177), .A2(n12455), .ZN(n6669) );
  AND2_X1 U9678 ( .A1(n6498), .A2(n7389), .ZN(n6670) );
  AND2_X1 U9679 ( .A1(n11909), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6671) );
  AND2_X1 U9680 ( .A1(n12458), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6672) );
  OR2_X1 U9681 ( .A1(n7655), .A2(n10164), .ZN(n6673) );
  INV_X1 U9682 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7455) );
  NOR2_X1 U9683 ( .A1(n7638), .A2(n12736), .ZN(n6674) );
  INV_X1 U9684 ( .A(n7934), .ZN(n7522) );
  INV_X1 U9685 ( .A(SI_22_), .ZN(n7586) );
  INV_X1 U9686 ( .A(n13884), .ZN(n7307) );
  INV_X1 U9687 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7003) );
  XNOR2_X1 U9688 ( .A(n8688), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12343) );
  INV_X1 U9689 ( .A(n12343), .ZN(n12357) );
  INV_X1 U9690 ( .A(n14598), .ZN(n7339) );
  AND2_X1 U9691 ( .A1(n7458), .A2(n10390), .ZN(n6675) );
  INV_X1 U9692 ( .A(n9940), .ZN(n14817) );
  AND2_X1 U9693 ( .A1(n10144), .A2(n10815), .ZN(n6676) );
  INV_X1 U9694 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7457) );
  INV_X1 U9695 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n6704) );
  INV_X1 U9696 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n6702) );
  INV_X1 U9697 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7005) );
  INV_X1 U9698 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7183) );
  XNOR2_X1 U9699 ( .A(n7641), .B(n10433), .ZN(n11032) );
  INV_X1 U9700 ( .A(n10433), .ZN(n7436) );
  NAND2_X1 U9701 ( .A1(n7630), .A2(n11130), .ZN(n6854) );
  INV_X1 U9702 ( .A(n11130), .ZN(n6979) );
  INV_X1 U9703 ( .A(n7369), .ZN(n7364) );
  OR2_X1 U9704 ( .A1(n15017), .A2(n15400), .ZN(n6914) );
  NAND2_X1 U9705 ( .A1(n14900), .A2(n7729), .ZN(n14881) );
  NAND2_X1 U9706 ( .A1(n14828), .A2(n7727), .ZN(n14815) );
  NAND2_X1 U9707 ( .A1(n7769), .A2(n11825), .ZN(n14973) );
  INV_X1 U9708 ( .A(n9435), .ZN(n11073) );
  INV_X2 U9710 ( .A(n9319), .ZN(n7024) );
  NOR2_X1 U9711 ( .A1(n10497), .A2(n10496), .ZN(n10546) );
  NAND2_X1 U9712 ( .A1(n14565), .A2(n14566), .ZN(n14564) );
  NAND2_X1 U9713 ( .A1(n10705), .A2(n10704), .ZN(n11325) );
  NAND2_X1 U9714 ( .A1(n11341), .A2(n11342), .ZN(n11718) );
  OAI21_X1 U9715 ( .B1(n14626), .B2(n14625), .A(n14624), .ZN(n14635) );
  NAND2_X1 U9716 ( .A1(n6679), .A2(n6698), .ZN(P1_U3262) );
  NAND2_X1 U9717 ( .A1(n7018), .A2(n7015), .ZN(n6679) );
  NOR2_X1 U9718 ( .A1(n15264), .A2(n7336), .ZN(n14565) );
  NOR2_X1 U9719 ( .A1(n11339), .A2(n7341), .ZN(n11341) );
  NOR2_X1 U9720 ( .A1(n10702), .A2(n7337), .ZN(n10705) );
  OAI21_X1 U9721 ( .B1(n12853), .B2(n9259), .A(n9262), .ZN(n7773) );
  NOR2_X1 U9722 ( .A1(n12768), .A2(n12770), .ZN(n7423) );
  NAND3_X1 U9723 ( .A1(n6680), .A2(n13141), .A3(n6651), .ZN(P3_U3456) );
  NAND2_X1 U9724 ( .A1(n7409), .A2(n7410), .ZN(n12814) );
  NAND3_X1 U9725 ( .A1(n6682), .A2(n7290), .A3(n7286), .ZN(P2_U3233) );
  NAND2_X1 U9726 ( .A1(n7288), .A2(n13936), .ZN(n6682) );
  NOR3_X1 U9727 ( .A1(n11260), .A2(n11259), .A3(n11262), .ZN(n11373) );
  NAND2_X1 U9728 ( .A1(n7864), .A2(n7862), .ZN(n9294) );
  NAND4_X2 U9729 ( .A1(n7184), .A2(n7813), .A3(n7812), .A4(n6511), .ZN(n8701)
         );
  NAND2_X1 U9730 ( .A1(n7228), .A2(n7412), .ZN(n7409) );
  NAND2_X1 U9731 ( .A1(n7155), .A2(n7157), .ZN(n7154) );
  NAND2_X1 U9732 ( .A1(n7162), .A2(n15225), .ZN(n15232) );
  NAND3_X1 U9733 ( .A1(n15239), .A2(n7186), .A3(n15238), .ZN(n7148) );
  AOI21_X2 U9734 ( .B1(n6688), .B2(n6687), .A(n6686), .ZN(n11499) );
  OAI21_X1 U9735 ( .B1(n10527), .B2(n10525), .A(n10526), .ZN(n10639) );
  NAND2_X1 U9736 ( .A1(n10544), .A2(n7338), .ZN(n10453) );
  NAND2_X1 U9737 ( .A1(n14453), .A2(n14452), .ZN(n14451) );
  NAND2_X1 U9738 ( .A1(n9666), .A2(n9665), .ZN(n14469) );
  NOR2_X1 U9739 ( .A1(n9487), .A2(n10301), .ZN(n9490) );
  INV_X4 U9740 ( .A(n9801), .ZN(n12422) );
  INV_X1 U9741 ( .A(n9312), .ZN(n7139) );
  NOR3_X1 U9742 ( .A1(n12809), .A2(n12339), .A3(n7258), .ZN(n12340) );
  NOR2_X4 U9743 ( .A1(n14796), .A2(n15033), .ZN(n14781) );
  INV_X1 U9744 ( .A(n12984), .ZN(n6694) );
  INV_X1 U9745 ( .A(n12974), .ZN(n6695) );
  INV_X1 U9746 ( .A(n12952), .ZN(n6696) );
  NAND2_X1 U9747 ( .A1(n13329), .A2(n13272), .ZN(n13484) );
  NAND2_X1 U9748 ( .A1(n7058), .A2(n7057), .ZN(n13261) );
  INV_X1 U9749 ( .A(n7524), .ZN(n7523) );
  NAND2_X2 U9750 ( .A1(n8202), .A2(n10339), .ZN(n10250) );
  NAND2_X1 U9751 ( .A1(n7562), .A2(n15774), .ZN(n7603) );
  INV_X1 U9752 ( .A(n14867), .ZN(n7719) );
  OAI21_X1 U9753 ( .B1(n14866), .B2(n7720), .A(n7717), .ZN(n14827) );
  INV_X4 U9754 ( .A(n10339), .ZN(n10338) );
  OAI211_X1 U9755 ( .C1(n15444), .C2(n13934), .A(n7289), .B(n15465), .ZN(n7288) );
  XNOR2_X1 U9756 ( .A(n7308), .B(n7307), .ZN(n13883) );
  AOI22_X1 U9757 ( .A1(n13928), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n13926), 
        .B2(n13927), .ZN(n13930) );
  XNOR2_X1 U9758 ( .A(n13925), .B(n13927), .ZN(n13928) );
  INV_X1 U9759 ( .A(n7302), .ZN(n10676) );
  OAI21_X1 U9760 ( .B1(n11674), .B2(n11673), .A(n6656), .ZN(n7308) );
  NAND2_X1 U9761 ( .A1(n13935), .A2(n15475), .ZN(n7289) );
  NAND2_X1 U9762 ( .A1(n9010), .A2(n9009), .ZN(n9027) );
  NOR2_X2 U9763 ( .A1(n8985), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7271) );
  INV_X1 U9764 ( .A(n9134), .ZN(n9133) );
  NAND2_X1 U9765 ( .A1(n9120), .A2(n9134), .ZN(n12891) );
  NAND2_X1 U9766 ( .A1(n9118), .A2(n15793), .ZN(n9134) );
  NOR2_X2 U9767 ( .A1(n9056), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9074) );
  NAND2_X1 U9768 ( .A1(n6603), .A2(n12161), .ZN(n8850) );
  NAND2_X1 U9769 ( .A1(n7866), .A2(n7789), .ZN(n7788) );
  NAND2_X1 U9770 ( .A1(n7788), .A2(n7787), .ZN(n9282) );
  NAND2_X2 U9771 ( .A1(n9112), .A2(n12237), .ZN(n12881) );
  NAND2_X1 U9772 ( .A1(n7855), .A2(n7853), .ZN(n12950) );
  NAND2_X1 U9773 ( .A1(n12793), .A2(n9269), .ZN(n7233) );
  OAI21_X2 U9774 ( .B1(n12881), .B2(n7882), .A(n7878), .ZN(n12852) );
  NAND2_X1 U9775 ( .A1(n12161), .A2(n12171), .ZN(n15590) );
  AOI21_X1 U9776 ( .B1(n12929), .B2(n9257), .A(n7931), .ZN(n12853) );
  NAND2_X1 U9777 ( .A1(n6710), .A2(n6709), .ZN(n12789) );
  NAND2_X1 U9778 ( .A1(n13136), .A2(n15599), .ZN(n6710) );
  NAND2_X1 U9779 ( .A1(n13578), .A2(n6463), .ZN(n6712) );
  AOI21_X1 U9780 ( .B1(n13588), .B2(n13587), .A(n13586), .ZN(n13594) );
  NAND3_X1 U9781 ( .A1(n7224), .A2(n7466), .A3(n6598), .ZN(n6717) );
  NAND2_X1 U9782 ( .A1(n14731), .A2(n9875), .ZN(n14766) );
  NAND3_X1 U9783 ( .A1(n7932), .A2(n13658), .A3(n6592), .ZN(n6723) );
  NAND2_X1 U9784 ( .A1(n6725), .A2(n6627), .ZN(n13709) );
  NAND3_X1 U9785 ( .A1(n7167), .A2(n6625), .A3(n7482), .ZN(n6725) );
  NAND2_X1 U9786 ( .A1(n6731), .A2(n6633), .ZN(n9500) );
  NAND2_X2 U9787 ( .A1(n14366), .A2(n8615), .ZN(n8202) );
  NAND3_X1 U9788 ( .A1(n7295), .A2(n7296), .A3(n8266), .ZN(n6739) );
  NAND2_X1 U9789 ( .A1(n6744), .A2(n6745), .ZN(n6740) );
  NAND3_X1 U9790 ( .A1(n6745), .A2(n6744), .A3(n14020), .ZN(n6741) );
  NAND2_X1 U9791 ( .A1(n10345), .A2(n10248), .ZN(n6755) );
  NAND2_X1 U9792 ( .A1(n6764), .A2(n15592), .ZN(n10891) );
  AOI21_X1 U9793 ( .B1(n6766), .B2(n14098), .A(n6768), .ZN(n6765) );
  NAND4_X1 U9794 ( .A1(n11163), .A2(n6782), .A3(n7797), .A4(n11423), .ZN(n6781) );
  NAND3_X1 U9795 ( .A1(n11163), .A2(n6782), .A3(n7797), .ZN(n11421) );
  NAND2_X1 U9796 ( .A1(n11010), .A2(n7241), .ZN(n11163) );
  NAND2_X1 U9797 ( .A1(n12471), .A2(n6786), .ZN(n6785) );
  NAND2_X1 U9798 ( .A1(n8579), .A2(n6790), .ZN(n6788) );
  NAND2_X1 U9799 ( .A1(n6788), .A2(n6789), .ZN(n14123) );
  NAND4_X1 U9800 ( .A1(n6795), .A2(n8040), .A3(n8625), .A4(n8041), .ZN(n6793)
         );
  NAND4_X1 U9801 ( .A1(n6569), .A2(n8040), .A3(n8625), .A4(n6795), .ZN(n6794)
         );
  NOR2_X2 U9802 ( .A1(n8162), .A2(n8284), .ZN(n8040) );
  NAND2_X1 U9803 ( .A1(n12607), .A2(n7821), .ZN(n6796) );
  NAND3_X1 U9804 ( .A1(n6806), .A2(n6632), .A3(n6805), .ZN(n14320) );
  OAI21_X1 U9805 ( .B1(n7285), .B2(n7547), .A(n6615), .ZN(n7280) );
  NAND3_X1 U9806 ( .A1(n6808), .A2(n13972), .A3(n13977), .ZN(n14315) );
  NAND2_X1 U9807 ( .A1(n12364), .A2(n12363), .ZN(n6821) );
  NAND2_X1 U9808 ( .A1(n6821), .A2(n6817), .ZN(P3_U3296) );
  NAND2_X1 U9809 ( .A1(n11458), .A2(n6829), .ZN(n6825) );
  NAND2_X1 U9810 ( .A1(n11846), .A2(n6833), .ZN(n6832) );
  NAND2_X1 U9811 ( .A1(n11846), .A2(n11847), .ZN(n11845) );
  NAND2_X1 U9812 ( .A1(n6855), .A2(n6854), .ZN(n6857) );
  NAND2_X1 U9813 ( .A1(n7612), .A2(n6860), .ZN(n6858) );
  NAND2_X1 U9814 ( .A1(n6858), .A2(n6859), .ZN(n7610) );
  INV_X4 U9815 ( .A(n8938), .ZN(n9099) );
  NAND2_X2 U9816 ( .A1(n8938), .A2(n10338), .ZN(n9038) );
  NAND2_X1 U9817 ( .A1(n12169), .A2(n7619), .ZN(n6870) );
  NAND2_X1 U9818 ( .A1(n7620), .A2(n6868), .ZN(n6872) );
  NAND2_X1 U9819 ( .A1(n6869), .A2(n7618), .ZN(n6871) );
  NAND3_X1 U9820 ( .A1(n6872), .A2(n7615), .A3(n6871), .ZN(n12186) );
  NAND2_X1 U9821 ( .A1(n8732), .A2(n6876), .ZN(n8734) );
  XNOR2_X1 U9822 ( .A(n6876), .B(n8836), .ZN(n10441) );
  NAND2_X1 U9823 ( .A1(n9050), .A2(n6881), .ZN(n6879) );
  NAND3_X1 U9824 ( .A1(n9175), .A2(n6476), .A3(n12852), .ZN(n6884) );
  NAND3_X1 U9825 ( .A1(n6885), .A2(n12260), .A3(n6884), .ZN(n9200) );
  OAI21_X1 U9826 ( .B1(n6891), .B2(n8745), .A(n8748), .ZN(n6887) );
  NAND2_X1 U9827 ( .A1(n8872), .A2(n6889), .ZN(n6888) );
  NAND2_X1 U9828 ( .A1(n6893), .A2(n6896), .ZN(n8759) );
  NAND2_X1 U9829 ( .A1(n8922), .A2(n6894), .ZN(n6893) );
  NAND2_X1 U9830 ( .A1(n8785), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8786) );
  NAND2_X1 U9831 ( .A1(n6899), .A2(n8786), .ZN(n9113) );
  NAND2_X1 U9832 ( .A1(n7672), .A2(n6903), .ZN(n6902) );
  NAND2_X1 U9833 ( .A1(n7672), .A2(n7670), .ZN(n8993) );
  NAND2_X1 U9834 ( .A1(n6905), .A2(n6608), .ZN(n12253) );
  NAND2_X1 U9835 ( .A1(n11817), .A2(n12294), .ZN(n6905) );
  NAND2_X1 U9836 ( .A1(n6906), .A2(n11366), .ZN(n10978) );
  XNOR2_X1 U9837 ( .A(n6906), .B(n11366), .ZN(n15353) );
  NAND2_X1 U9838 ( .A1(n10976), .A2(n10975), .ZN(n6906) );
  OAI211_X1 U9839 ( .C1(n6915), .C2(n15440), .A(n6913), .B(n6910), .ZN(
        P1_U3557) );
  NAND2_X1 U9840 ( .A1(n6481), .A2(n14724), .ZN(n15016) );
  NAND3_X1 U9841 ( .A1(n6915), .A2(n6914), .A3(n6912), .ZN(n15133) );
  NAND2_X1 U9842 ( .A1(n14941), .A2(n14944), .ZN(n6931) );
  INV_X1 U9843 ( .A(n6929), .ZN(n6928) );
  NAND2_X1 U9844 ( .A1(n12027), .A2(n6935), .ZN(n6934) );
  NAND2_X1 U9845 ( .A1(n6934), .A2(n6932), .ZN(n14971) );
  NAND2_X1 U9846 ( .A1(n6936), .A2(n7349), .ZN(n12064) );
  NAND2_X1 U9847 ( .A1(n12027), .A2(n7351), .ZN(n6936) );
  NAND3_X1 U9848 ( .A1(n9312), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_IR_REG_29__SCAN_IN), .ZN(n6940) );
  NAND3_X1 U9849 ( .A1(n9309), .A2(n6453), .A3(n9310), .ZN(n9312) );
  NAND3_X1 U9850 ( .A1(n14777), .A2(n6942), .A3(n6595), .ZN(n6941) );
  NAND2_X1 U9851 ( .A1(n14777), .A2(n14713), .ZN(n14771) );
  NAND2_X1 U9852 ( .A1(n6944), .A2(n15289), .ZN(n11823) );
  XNOR2_X1 U9853 ( .A(n6944), .B(n15289), .ZN(n15411) );
  NAND2_X1 U9854 ( .A1(n7343), .A2(n7344), .ZN(n6944) );
  INV_X1 U9855 ( .A(n6661), .ZN(n6945) );
  NAND2_X1 U9856 ( .A1(n6948), .A2(n6469), .ZN(n8638) );
  INV_X1 U9857 ( .A(n8284), .ZN(n6947) );
  INV_X1 U9858 ( .A(n8162), .ZN(n6949) );
  AND2_X2 U9859 ( .A1(n8041), .A2(n8040), .ZN(n8332) );
  AND2_X1 U9860 ( .A1(n8625), .A2(n8032), .ZN(n8042) );
  NAND2_X1 U9861 ( .A1(n7917), .A2(n7915), .ZN(n13945) );
  NAND2_X1 U9862 ( .A1(n7917), .A2(n6950), .ZN(n6953) );
  INV_X1 U9863 ( .A(n6953), .ZN(n13944) );
  NAND3_X1 U9864 ( .A1(n11415), .A2(n6958), .A3(n11809), .ZN(n11807) );
  NAND3_X1 U9865 ( .A1(n11415), .A2(n6958), .A3(n6957), .ZN(n14194) );
  NAND2_X1 U9866 ( .A1(n10592), .A2(n6962), .ZN(n6961) );
  NOR2_X1 U9867 ( .A1(n14356), .A2(n8548), .ZN(n8553) );
  NAND2_X1 U9868 ( .A1(n8096), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8087) );
  NAND2_X1 U9869 ( .A1(n8150), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8099) );
  NAND2_X1 U9870 ( .A1(n7515), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8544) );
  OAI21_X1 U9871 ( .B1(n8160), .B2(P2_IR_REG_4__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8161) );
  NAND2_X1 U9872 ( .A1(n8658), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8660) );
  NAND2_X1 U9873 ( .A1(n8545), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8542) );
  NAND2_X1 U9874 ( .A1(n8245), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8246) );
  NAND2_X1 U9875 ( .A1(n8632), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8633) );
  NAND2_X1 U9876 ( .A1(n8634), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8629) );
  OAI21_X1 U9877 ( .B1(n8270), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8271) );
  NAND2_X1 U9878 ( .A1(n13912), .A2(n13931), .ZN(n13914) );
  NAND2_X1 U9879 ( .A1(n13910), .A2(n6967), .ZN(n13931) );
  NAND2_X1 U9880 ( .A1(n13910), .A2(n13909), .ZN(n13911) );
  NAND2_X1 U9881 ( .A1(n11377), .A2(n11376), .ZN(n11379) );
  NAND2_X1 U9882 ( .A1(n11377), .A2(n6973), .ZN(n11670) );
  AND2_X4 U9883 ( .A1(n7438), .A2(n7439), .ZN(n10139) );
  NAND2_X1 U9884 ( .A1(n12708), .A2(n10160), .ZN(n10161) );
  NAND2_X1 U9885 ( .A1(n10146), .A2(n11130), .ZN(n10147) );
  NAND2_X1 U9886 ( .A1(n11462), .A2(n6639), .ZN(n6984) );
  OAI21_X1 U9887 ( .B1(n6983), .B2(n11783), .A(n6981), .ZN(n10152) );
  AOI21_X1 U9888 ( .B1(n11462), .B2(n6655), .A(n6982), .ZN(n6981) );
  NAND2_X1 U9889 ( .A1(n11462), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n11611) );
  INV_X1 U9890 ( .A(n10654), .ZN(n6991) );
  OAI21_X1 U9891 ( .B1(n10654), .B2(n6987), .A(n6593), .ZN(n6986) );
  INV_X1 U9892 ( .A(n9442), .ZN(n6987) );
  NAND2_X1 U9893 ( .A1(n6989), .A2(n6990), .ZN(n10903) );
  NAND3_X1 U9894 ( .A1(n6991), .A2(n10663), .A3(n10662), .ZN(n6989) );
  NAND2_X1 U9895 ( .A1(n14460), .A2(n14461), .ZN(n14459) );
  NAND2_X1 U9896 ( .A1(n15158), .A2(n7004), .ZN(n7000) );
  OAI21_X1 U9897 ( .B1(n7001), .B2(n15158), .A(n7000), .ZN(n9424) );
  INV_X1 U9898 ( .A(n15162), .ZN(n9351) );
  AND2_X1 U9899 ( .A1(n9352), .A2(n15162), .ZN(n9444) );
  OAI21_X1 U9900 ( .B1(n15162), .B2(n7003), .A(n7002), .ZN(n7001) );
  NAND2_X1 U9901 ( .A1(n15162), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7002) );
  NAND2_X1 U9902 ( .A1(n15162), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n7004) );
  NAND2_X1 U9903 ( .A1(n9309), .A2(n6453), .ZN(n9317) );
  NAND2_X1 U9904 ( .A1(n7017), .A2(n7016), .ZN(n7015) );
  NAND2_X1 U9905 ( .A1(n14646), .A2(n15277), .ZN(n7017) );
  INV_X1 U9906 ( .A(n9404), .ZN(n9321) );
  INV_X1 U9907 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7023) );
  OAI21_X1 U9908 ( .B1(n7750), .B2(n7032), .A(n7034), .ZN(n7031) );
  INV_X1 U9909 ( .A(n10022), .ZN(n7032) );
  NAND2_X1 U9910 ( .A1(n7033), .A2(n10061), .ZN(n7218) );
  INV_X1 U9911 ( .A(n10021), .ZN(n7034) );
  NAND2_X1 U9912 ( .A1(n6606), .A2(n10974), .ZN(n7035) );
  NAND4_X1 U9913 ( .A1(n7040), .A2(n7039), .A3(n7038), .A4(n10137), .ZN(
        P1_U3242) );
  NAND3_X1 U9914 ( .A1(n7732), .A2(n7731), .A3(n6631), .ZN(n7038) );
  OR2_X1 U9915 ( .A1(n7732), .A2(n6572), .ZN(n7040) );
  NAND2_X1 U9916 ( .A1(n10092), .A2(n6451), .ZN(n7043) );
  NAND2_X1 U9917 ( .A1(n10108), .A2(n6465), .ZN(n7049) );
  NOR2_X2 U9918 ( .A1(n13414), .A2(n11480), .ZN(n11620) );
  NAND2_X1 U9919 ( .A1(n8113), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8095) );
  NAND2_X1 U9920 ( .A1(n11882), .A2(n7060), .ZN(n7058) );
  OR3_X2 U9921 ( .A1(n13457), .A2(n7527), .A3(n7070), .ZN(n7069) );
  OR2_X1 U9922 ( .A1(n14723), .A2(n14722), .ZN(n7078) );
  NAND3_X1 U9923 ( .A1(n7591), .A2(n8004), .A3(n7589), .ZN(n7079) );
  NAND2_X1 U9924 ( .A1(n7591), .A2(n7589), .ZN(n7082) );
  NAND2_X1 U9925 ( .A1(n7079), .A2(n6628), .ZN(n8380) );
  NAND3_X1 U9926 ( .A1(n7575), .A2(n7576), .A3(n8477), .ZN(n8480) );
  NAND3_X1 U9927 ( .A1(n7086), .A2(n7083), .A3(n7602), .ZN(n7090) );
  AOI21_X1 U9928 ( .B1(n7576), .B2(n7088), .A(n7087), .ZN(n7086) );
  NOR2_X1 U9929 ( .A1(n8070), .A2(n8477), .ZN(n7088) );
  NAND2_X1 U9930 ( .A1(n8480), .A2(n7576), .ZN(n8071) );
  NAND3_X1 U9931 ( .A1(n7092), .A2(n7976), .A3(n7571), .ZN(n7091) );
  NAND2_X1 U9932 ( .A1(n7315), .A2(n7098), .ZN(n7097) );
  NAND2_X1 U9933 ( .A1(n7105), .A2(n10964), .ZN(n8415) );
  AND4_X2 U9934 ( .A1(n9306), .A2(n7024), .A3(n9304), .A4(n9305), .ZN(n9309)
         );
  INV_X1 U9935 ( .A(n9309), .ZN(n9343) );
  OAI21_X1 U9936 ( .B1(n11107), .B2(n7113), .A(n7112), .ZN(n15302) );
  AOI21_X1 U9937 ( .B1(n7118), .B2(n7119), .A(n6454), .ZN(n7112) );
  NAND2_X1 U9938 ( .A1(n7117), .A2(n11107), .ZN(n7116) );
  NAND3_X1 U9939 ( .A1(n14779), .A2(n7128), .A3(n7130), .ZN(n7124) );
  NAND2_X1 U9940 ( .A1(n6510), .A2(n14815), .ZN(n7125) );
  NAND2_X1 U9941 ( .A1(n14791), .A2(n7129), .ZN(n7126) );
  NAND2_X2 U9942 ( .A1(n7126), .A2(n7127), .ZN(n14778) );
  NAND3_X1 U9943 ( .A1(n7132), .A2(n14673), .A3(n7131), .ZN(n14926) );
  NAND3_X1 U9944 ( .A1(n7702), .A2(n7133), .A3(n7135), .ZN(n7131) );
  NAND3_X1 U9945 ( .A1(n12069), .A2(n7133), .A3(n7702), .ZN(n7132) );
  NAND2_X2 U9946 ( .A1(n10407), .A2(n10338), .ZN(n9425) );
  NAND2_X2 U9947 ( .A1(n15167), .A2(n14651), .ZN(n10407) );
  INV_X1 U9948 ( .A(n14512), .ZN(n10991) );
  OAI21_X1 U9949 ( .B1(n6441), .B2(n14512), .A(n10992), .ZN(n7144) );
  NAND2_X1 U9950 ( .A1(n7145), .A2(n15198), .ZN(n15196) );
  NAND2_X1 U9951 ( .A1(n15239), .A2(n15238), .ZN(n7147) );
  INV_X1 U9952 ( .A(n15238), .ZN(n7150) );
  NAND2_X1 U9953 ( .A1(n10371), .A2(n7151), .ZN(n7152) );
  NAND2_X1 U9954 ( .A1(n10371), .A2(n10370), .ZN(n7160) );
  INV_X1 U9955 ( .A(n10370), .ZN(n7155) );
  INV_X1 U9956 ( .A(n7157), .ZN(n7156) );
  NAND2_X1 U9957 ( .A1(n7160), .A2(n10359), .ZN(n10361) );
  NAND2_X1 U9958 ( .A1(n7159), .A2(n10360), .ZN(n7158) );
  INV_X1 U9959 ( .A(n10359), .ZN(n7159) );
  NAND2_X1 U9960 ( .A1(n10778), .A2(n10777), .ZN(n7165) );
  OR2_X1 U9961 ( .A1(n13564), .A2(n13563), .ZN(n13570) );
  NAND2_X1 U9962 ( .A1(n7169), .A2(n7479), .ZN(n13562) );
  OAI22_X1 U9963 ( .A1(n13594), .A2(n13593), .B1(n13615), .B2(n13614), .ZN(
        n13647) );
  AOI21_X1 U9964 ( .B1(n13664), .B2(n13663), .A(n13662), .ZN(n7481) );
  OAI21_X1 U9965 ( .B1(n13668), .B2(n13667), .A(n7168), .ZN(n7167) );
  NAND2_X1 U9966 ( .A1(n8957), .A2(n8956), .ZN(n8973) );
  NAND2_X1 U9967 ( .A1(n9074), .A2(n9073), .ZN(n9091) );
  NAND2_X1 U9968 ( .A1(n9133), .A2(n9132), .ZN(n9145) );
  INV_X2 U9969 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n15680) );
  NAND2_X1 U9970 ( .A1(n7271), .A2(n15765), .ZN(n9011) );
  INV_X1 U9971 ( .A(n9011), .ZN(n9010) );
  NAND2_X1 U9972 ( .A1(n7272), .A2(n15703), .ZN(n9056) );
  NAND2_X1 U9973 ( .A1(n9200), .A2(n12263), .ZN(n12790) );
  INV_X1 U9974 ( .A(n9175), .ZN(n7850) );
  AOI21_X1 U9975 ( .B1(n12792), .B2(n12782), .A(n12346), .ZN(n12356) );
  NAND2_X1 U9976 ( .A1(n12871), .A2(n12870), .ZN(n9261) );
  NAND2_X1 U9977 ( .A1(n9260), .A2(n12887), .ZN(n12871) );
  NAND2_X1 U9978 ( .A1(n9066), .A2(n8782), .ZN(n9096) );
  INV_X1 U9979 ( .A(n8785), .ZN(n7171) );
  NAND2_X1 U9980 ( .A1(n7229), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7691) );
  NAND2_X1 U9981 ( .A1(n8734), .A2(n8733), .ZN(n8845) );
  NAND2_X1 U9982 ( .A1(n8742), .A2(n8741), .ZN(n8872) );
  NAND2_X1 U9983 ( .A1(n8751), .A2(n6617), .ZN(n8922) );
  XNOR2_X1 U9984 ( .A(n9153), .B(n12115), .ZN(n11817) );
  NAND2_X1 U9985 ( .A1(n12795), .A2(n9269), .ZN(n12794) );
  INV_X1 U9986 ( .A(n12380), .ZN(n7408) );
  NAND2_X1 U9987 ( .A1(n7494), .A2(n8668), .ZN(P2_U3496) );
  NOR2_X1 U9988 ( .A1(n7423), .A2(n12778), .ZN(n7422) );
  OAI21_X1 U9989 ( .B1(n8260), .B2(n7570), .A(n7568), .ZN(n8283) );
  NAND2_X1 U9990 ( .A1(n15183), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7185) );
  NAND2_X1 U9991 ( .A1(n7463), .A2(n7464), .ZN(n15198) );
  NAND2_X1 U9992 ( .A1(n7894), .A2(n7892), .ZN(n11504) );
  NAND2_X1 U9993 ( .A1(n10128), .A2(n10127), .ZN(n7731) );
  NAND2_X1 U9994 ( .A1(n10129), .A2(n10130), .ZN(n7732) );
  NAND2_X1 U9995 ( .A1(n13264), .A2(n13263), .ZN(n7540) );
  OAI211_X1 U9997 ( .C1(SI_2_), .C2(n8089), .A(n7954), .B(n8102), .ZN(n8147)
         );
  NAND2_X1 U9998 ( .A1(n7953), .A2(n7952), .ZN(n8102) );
  NAND2_X1 U9999 ( .A1(n8023), .A2(n11820), .ZN(n7575) );
  NAND2_X1 U10000 ( .A1(n8380), .A2(n6611), .ZN(n7315) );
  NAND2_X1 U10001 ( .A1(n7534), .A2(n13321), .ZN(n7533) );
  INV_X1 U10002 ( .A(n7533), .ZN(n7531) );
  NAND2_X1 U10003 ( .A1(n13322), .A2(n7535), .ZN(n7534) );
  NAND2_X1 U10004 ( .A1(n7181), .A2(n7179), .ZN(P2_U3498) );
  OR2_X1 U10005 ( .A1(n10260), .A2(n7182), .ZN(n7181) );
  XNOR2_X1 U10006 ( .A(n13742), .B(n8614), .ZN(n8557) );
  NAND2_X1 U10007 ( .A1(n11650), .A2(n11649), .ZN(n11653) );
  NAND2_X1 U10008 ( .A1(n7693), .A2(n7692), .ZN(n14941) );
  NAND2_X1 U10009 ( .A1(n15198), .A2(n15197), .ZN(n15199) );
  NAND2_X1 U10010 ( .A1(n10958), .A2(n6486), .ZN(n10930) );
  INV_X1 U10011 ( .A(n10956), .ZN(n7187) );
  NAND2_X1 U10012 ( .A1(n7257), .A2(n10565), .ZN(n7256) );
  NAND2_X1 U10013 ( .A1(n11626), .A2(n6612), .ZN(n7520) );
  NAND2_X1 U10014 ( .A1(n7197), .A2(n7530), .ZN(n13470) );
  NAND2_X1 U10015 ( .A1(n11620), .A2(n7244), .ZN(n11626) );
  NAND2_X1 U10016 ( .A1(n7520), .A2(n7518), .ZN(n11882) );
  OAI21_X1 U10017 ( .B1(n13309), .B2(n7532), .A(n7531), .ZN(n7530) );
  NAND3_X1 U10018 ( .A1(n8147), .A2(n8146), .A3(n7958), .ZN(n7198) );
  NAND2_X1 U10019 ( .A1(n7929), .A2(n7695), .ZN(n7694) );
  NAND2_X1 U10020 ( .A1(n14794), .A2(n14793), .ZN(n14792) );
  NAND2_X1 U10021 ( .A1(n14775), .A2(n14774), .ZN(n14777) );
  NAND2_X1 U10022 ( .A1(n7354), .A2(n7697), .ZN(n14794) );
  NAND2_X1 U10023 ( .A1(n13489), .A2(n7541), .ZN(n13287) );
  NAND2_X1 U10024 ( .A1(n11253), .A2(n11252), .ZN(n15303) );
  NAND2_X1 U10025 ( .A1(n10978), .A2(n10977), .ZN(n11306) );
  NAND2_X1 U10026 ( .A1(n10690), .A2(n7191), .ZN(n10663) );
  INV_X1 U10027 ( .A(n10687), .ZN(n7192) );
  NAND2_X1 U10028 ( .A1(n9439), .A2(n10687), .ZN(n10690) );
  AND2_X1 U10029 ( .A1(n9313), .A2(n15706), .ZN(n9341) );
  AOI21_X1 U10030 ( .B1(n11504), .B2(n11503), .A(n7193), .ZN(n11591) );
  OR2_X1 U10031 ( .A1(n13641), .A2(n13606), .ZN(n13638) );
  NOR2_X1 U10032 ( .A1(n13646), .A2(n6474), .ZN(n7473) );
  NAND2_X1 U10033 ( .A1(n7529), .A2(n13303), .ZN(n7197) );
  NAND3_X1 U10034 ( .A1(n7578), .A2(n13790), .A3(n7577), .ZN(n13730) );
  NAND2_X1 U10035 ( .A1(n7198), .A2(n7960), .ZN(n8238) );
  NAND2_X1 U10036 ( .A1(n7199), .A2(n13730), .ZN(n13735) );
  INV_X1 U10037 ( .A(n7829), .ZN(n12538) );
  INV_X4 U10038 ( .A(n7404), .ZN(n12294) );
  NAND2_X1 U10039 ( .A1(n14371), .A2(n10248), .ZN(n8073) );
  NAND2_X1 U10040 ( .A1(n8022), .A2(n8021), .ZN(n8024) );
  NAND2_X1 U10041 ( .A1(n7972), .A2(n7971), .ZN(n8211) );
  NAND2_X1 U10042 ( .A1(n7211), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7210) );
  NAND2_X2 U10043 ( .A1(n7204), .A2(n8045), .ZN(n14210) );
  NAND2_X1 U10044 ( .A1(n7276), .A2(n10248), .ZN(n7204) );
  NAND2_X1 U10045 ( .A1(n7446), .A2(n7445), .ZN(n11969) );
  INV_X1 U10046 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7206) );
  NAND2_X1 U10047 ( .A1(n7243), .A2(n7242), .ZN(n10389) );
  XNOR2_X2 U10048 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n10370) );
  NAND2_X1 U10049 ( .A1(n7209), .A2(n8119), .ZN(n7953) );
  NAND2_X1 U10050 ( .A1(n7951), .A2(n7210), .ZN(n7209) );
  INV_X1 U10051 ( .A(n6442), .ZN(n7211) );
  OAI21_X1 U10052 ( .B1(n13983), .B2(n7502), .A(n7498), .ZN(n7497) );
  NAND2_X1 U10053 ( .A1(n14415), .A2(n7213), .ZN(n14453) );
  NAND2_X1 U10055 ( .A1(n10089), .A2(n10090), .ZN(n10092) );
  NAND2_X1 U10056 ( .A1(n7218), .A2(n6548), .ZN(n7217) );
  NAND3_X1 U10057 ( .A1(n10267), .A2(n10266), .A3(n15556), .ZN(n7219) );
  INV_X1 U10058 ( .A(n10265), .ZN(n10285) );
  NAND2_X1 U10059 ( .A1(n8604), .A2(n13998), .ZN(n7254) );
  NAND2_X1 U10060 ( .A1(n7579), .A2(n13733), .ZN(n7577) );
  AOI21_X1 U10061 ( .B1(n13665), .B2(n13666), .A(n7481), .ZN(n13668) );
  NAND3_X1 U10062 ( .A1(n7225), .A2(n13542), .A3(n13543), .ZN(n7224) );
  NAND3_X1 U10063 ( .A1(n13524), .A2(n13523), .A3(n13522), .ZN(n7226) );
  INV_X4 U10064 ( .A(n12494), .ZN(n12463) );
  AND2_X4 U10065 ( .A1(n7794), .A2(n10851), .ZN(n12494) );
  NAND2_X1 U10066 ( .A1(n8705), .A2(n13258), .ZN(n7267) );
  AOI21_X1 U10067 ( .B1(n12743), .B2(n7265), .A(n12742), .ZN(n12746) );
  NOR2_X1 U10068 ( .A1(n10150), .A2(n7426), .ZN(n11462) );
  NAND2_X1 U10069 ( .A1(n11789), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n11788) );
  AOI21_X1 U10070 ( .B1(n7657), .B2(n7659), .A(n9033), .ZN(n7656) );
  INV_X1 U10071 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n8086) );
  INV_X1 U10072 ( .A(n13670), .ZN(n7227) );
  OAI211_X1 U10073 ( .C1(n12706), .C2(n7636), .A(n7634), .B(n7633), .ZN(n12728) );
  NAND2_X2 U10074 ( .A1(n15608), .A2(n15585), .ZN(n12171) );
  AOI21_X1 U10075 ( .B1(n13570), .B2(n13569), .A(n13568), .ZN(n13572) );
  NAND2_X1 U10076 ( .A1(n13709), .A2(n7262), .ZN(n7475) );
  INV_X1 U10077 ( .A(n8791), .ZN(n7229) );
  NAND2_X1 U10078 ( .A1(n12268), .A2(n6610), .ZN(n12264) );
  INV_X1 U10079 ( .A(n9265), .ZN(n7228) );
  NAND2_X1 U10080 ( .A1(n7610), .A2(n7608), .ZN(n7607) );
  NAND2_X1 U10081 ( .A1(n15840), .A2(n15839), .ZN(n7243) );
  OAI21_X2 U10082 ( .B1(n12800), .B2(n15644), .A(n12799), .ZN(n13030) );
  OAI21_X1 U10083 ( .B1(n7851), .B2(n7850), .A(n12821), .ZN(n7849) );
  INV_X1 U10084 ( .A(n7347), .ZN(n7346) );
  NAND2_X1 U10085 ( .A1(n14843), .A2(n6630), .ZN(n7354) );
  INV_X1 U10086 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7230) );
  NAND2_X1 U10087 ( .A1(n13144), .A2(n7231), .ZN(P3_U3454) );
  NAND2_X1 U10088 ( .A1(n13033), .A2(n7232), .ZN(P3_U3486) );
  AOI21_X2 U10089 ( .B1(n10300), .B2(n9490), .A(n7933), .ZN(n11433) );
  NAND2_X1 U10090 ( .A1(n7908), .A2(n6618), .ZN(n14398) );
  NAND2_X1 U10091 ( .A1(n9996), .A2(n10994), .ZN(n11366) );
  NOR2_X2 U10092 ( .A1(n13742), .A2(n13791), .ZN(n13499) );
  NAND2_X1 U10093 ( .A1(n13008), .A2(n12165), .ZN(n12162) );
  AOI21_X1 U10094 ( .B1(n7607), .B2(n7605), .A(n6590), .ZN(n12258) );
  NAND2_X1 U10095 ( .A1(n7278), .A2(n7586), .ZN(n8443) );
  NAND2_X1 U10096 ( .A1(n14398), .A2(n9705), .ZN(n12383) );
  NAND2_X1 U10097 ( .A1(n7919), .A2(n7918), .ZN(n14068) );
  INV_X1 U10098 ( .A(n8016), .ZN(n7278) );
  INV_X1 U10099 ( .A(n15168), .ZN(n7276) );
  NAND2_X1 U10100 ( .A1(n8443), .A2(n7277), .ZN(n8022) );
  NAND2_X1 U10101 ( .A1(n6491), .A2(n7273), .ZN(n10277) );
  OAI21_X1 U10102 ( .B1(n10279), .B2(n15578), .A(n7239), .ZN(P2_U3527) );
  NAND2_X1 U10103 ( .A1(n10893), .A2(n10894), .ZN(n11010) );
  NAND2_X1 U10104 ( .A1(n7808), .A2(n7809), .ZN(n11991) );
  NAND2_X2 U10105 ( .A1(n8938), .A2(n10339), .ZN(n7404) );
  INV_X1 U10106 ( .A(n9366), .ZN(n9305) );
  NAND2_X1 U10107 ( .A1(n14709), .A2(n14708), .ZN(n14843) );
  NAND2_X1 U10108 ( .A1(n10156), .A2(n10501), .ZN(n10159) );
  NAND2_X1 U10109 ( .A1(n13470), .A2(n13366), .ZN(n13377) );
  NAND2_X1 U10110 ( .A1(n12710), .A2(n12709), .ZN(n7431) );
  NOR2_X1 U10111 ( .A1(n11195), .A2(n11196), .ZN(n11194) );
  NOR2_X2 U10112 ( .A1(n7497), .A2(n7253), .ZN(n10282) );
  NAND2_X1 U10113 ( .A1(n10183), .A2(n11466), .ZN(n7255) );
  NAND2_X1 U10114 ( .A1(n7902), .A2(n7900), .ZN(n9666) );
  NAND2_X1 U10115 ( .A1(n8767), .A2(n8766), .ZN(n9003) );
  NAND2_X1 U10116 ( .A1(n9435), .A2(n9434), .ZN(n9438) );
  XNOR2_X2 U10117 ( .A(n9451), .B(P1_IR_REG_2__SCAN_IN), .ZN(n14537) );
  NAND2_X1 U10118 ( .A1(n7664), .A2(n7662), .ZN(n8790) );
  AND2_X2 U10119 ( .A1(n8703), .A2(n7792), .ZN(n8806) );
  NAND4_X1 U10120 ( .A1(n12326), .A2(n15583), .A3(n12327), .A4(n12328), .ZN(
        n12329) );
  NAND2_X1 U10121 ( .A1(n7926), .A2(n7661), .ZN(n12344) );
  INV_X1 U10122 ( .A(n7979), .ZN(n7572) );
  INV_X1 U10123 ( .A(n13968), .ZN(n7273) );
  OAI21_X1 U10124 ( .B1(n7284), .B2(n7280), .A(n13759), .ZN(n14110) );
  OAI22_X1 U10125 ( .A1(n7282), .A2(n7281), .B1(n8366), .B2(n8365), .ZN(n14133) );
  NAND2_X1 U10126 ( .A1(n7545), .A2(n7283), .ZN(n7281) );
  INV_X1 U10127 ( .A(n8365), .ZN(n7283) );
  NAND2_X1 U10128 ( .A1(n7293), .A2(n11295), .ZN(n7294) );
  NAND2_X1 U10129 ( .A1(n6485), .A2(n11413), .ZN(n7296) );
  XNOR2_X1 U10130 ( .A(n8086), .B(n7309), .ZN(n13838) );
  OAI21_X1 U10131 ( .B1(n7506), .B2(n7505), .A(n6614), .ZN(n7504) );
  NAND2_X1 U10132 ( .A1(n7327), .A2(n7323), .ZN(n14319) );
  NAND2_X1 U10133 ( .A1(n6564), .A2(n7332), .ZN(n7331) );
  NAND2_X1 U10134 ( .A1(n13984), .A2(n13983), .ZN(n7332) );
  AOI21_X1 U10135 ( .B1(n15267), .B2(n15266), .A(n15265), .ZN(n15264) );
  MUX2_X1 U10136 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10446), .S(n14517), .Z(
        n14515) );
  XNOR2_X2 U10137 ( .A(n7342), .B(P1_IR_REG_1__SCAN_IN), .ZN(n14517) );
  NAND2_X1 U10138 ( .A1(n15303), .A2(n7346), .ZN(n7343) );
  NOR2_X2 U10139 ( .A1(n14770), .A2(n7358), .ZN(n15025) );
  NAND2_X1 U10140 ( .A1(n7362), .A2(n7359), .ZN(n10243) );
  NAND2_X1 U10141 ( .A1(n12695), .A2(n7361), .ZN(n7359) );
  NAND2_X1 U10142 ( .A1(n7366), .A2(n7367), .ZN(n12732) );
  INV_X1 U10143 ( .A(n12733), .ZN(n7365) );
  NAND2_X1 U10144 ( .A1(n11034), .A2(n7379), .ZN(n7375) );
  OAI21_X1 U10145 ( .B1(n11034), .B2(n11033), .A(n6455), .ZN(n11193) );
  NAND2_X1 U10146 ( .A1(n10935), .A2(n6626), .ZN(n7385) );
  MUX2_X1 U10147 ( .A(n13015), .B(n10955), .S(n13246), .Z(n10201) );
  NAND2_X4 U10148 ( .A1(n8807), .A2(n7391), .ZN(n13246) );
  NOR2_X1 U10149 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_27__SCAN_IN), 
        .ZN(n7392) );
  INV_X2 U10150 ( .A(n8701), .ZN(n8703) );
  NAND3_X1 U10151 ( .A1(n6511), .A2(n8683), .A3(n8682), .ZN(n8695) );
  NAND2_X1 U10152 ( .A1(n7397), .A2(n7399), .ZN(n9239) );
  NAND2_X1 U10153 ( .A1(n7408), .A2(n12294), .ZN(n9131) );
  NAND2_X1 U10154 ( .A1(n7777), .A2(n7416), .ZN(n11569) );
  NAND3_X1 U10155 ( .A1(n7418), .A2(n7417), .A3(n9228), .ZN(n7416) );
  NAND3_X1 U10156 ( .A1(n7418), .A2(n9228), .A3(n12320), .ZN(n11536) );
  AND2_X1 U10157 ( .A1(n9228), .A2(n7418), .ZN(n11537) );
  NAND2_X1 U10158 ( .A1(n10151), .A2(n6654), .ZN(n7425) );
  NAND3_X1 U10159 ( .A1(n7432), .A2(n10159), .A3(n7430), .ZN(n7429) );
  NAND2_X1 U10160 ( .A1(n10158), .A2(n10157), .ZN(n7432) );
  AND2_X2 U10161 ( .A1(n10139), .A2(n7811), .ZN(n7812) );
  NAND3_X1 U10162 ( .A1(n10144), .A2(n10815), .A3(P3_REG2_REG_3__SCAN_IN), 
        .ZN(n10795) );
  NAND2_X1 U10163 ( .A1(n10795), .A2(n10815), .ZN(n7440) );
  NAND2_X1 U10164 ( .A1(n7442), .A2(n7443), .ZN(n7441) );
  NAND2_X1 U10165 ( .A1(n10154), .A2(n10233), .ZN(n7444) );
  NAND2_X1 U10166 ( .A1(n11495), .A2(n7447), .ZN(n7446) );
  NAND2_X1 U10167 ( .A1(n11495), .A2(n11494), .ZN(n7456) );
  INV_X1 U10168 ( .A(n11498), .ZN(n7452) );
  NAND2_X1 U10169 ( .A1(n7456), .A2(n11498), .ZN(n11731) );
  XNOR2_X2 U10170 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n10366) );
  NAND2_X1 U10171 ( .A1(n15181), .A2(n15182), .ZN(n7461) );
  NAND2_X1 U10172 ( .A1(n7461), .A2(n10771), .ZN(n10778) );
  NAND2_X1 U10173 ( .A1(n7464), .A2(n15186), .ZN(n15195) );
  NAND2_X1 U10174 ( .A1(n15212), .A2(n6624), .ZN(n15224) );
  NAND2_X1 U10175 ( .A1(n15212), .A2(n15211), .ZN(n15221) );
  OAI21_X1 U10176 ( .B1(n13647), .B2(n7472), .A(n7471), .ZN(n13657) );
  NAND2_X1 U10177 ( .A1(n7470), .A2(n7467), .ZN(n13658) );
  NAND3_X1 U10178 ( .A1(n13647), .A2(n7471), .A3(n13656), .ZN(n7470) );
  NAND2_X1 U10179 ( .A1(n7475), .A2(n7476), .ZN(n13753) );
  NAND2_X1 U10180 ( .A1(n7475), .A2(n7474), .ZN(n13803) );
  NOR2_X1 U10181 ( .A1(n13562), .A2(n13561), .ZN(n13563) );
  NAND2_X1 U10182 ( .A1(n13668), .A2(n13667), .ZN(n7482) );
  NAND2_X1 U10183 ( .A1(n8059), .A2(n7483), .ZN(n14357) );
  NAND2_X1 U10184 ( .A1(n7487), .A2(n7485), .ZN(n8568) );
  NAND3_X1 U10185 ( .A1(n8142), .A2(n8143), .A3(n8144), .ZN(n7486) );
  NAND3_X1 U10186 ( .A1(n15488), .A2(n15487), .A3(n15551), .ZN(n7487) );
  NAND2_X1 U10187 ( .A1(n8566), .A2(n8565), .ZN(n7488) );
  NAND2_X1 U10188 ( .A1(n11176), .A2(n6537), .ZN(n15488) );
  INV_X1 U10189 ( .A(n11895), .ZN(n8579) );
  NAND2_X1 U10190 ( .A1(n13998), .A2(n8604), .ZN(n7496) );
  INV_X1 U10191 ( .A(n8603), .ZN(n7502) );
  NAND2_X1 U10192 ( .A1(n8332), .A2(n7514), .ZN(n7515) );
  NAND2_X1 U10193 ( .A1(n7517), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8371) );
  AOI21_X1 U10194 ( .B1(n7517), .B2(n8553), .A(n7516), .ZN(n8554) );
  AND2_X1 U10195 ( .A1(n8551), .A2(n8552), .ZN(n7516) );
  OAI21_X1 U10196 ( .B1(n11628), .B2(n11627), .A(n11625), .ZN(n7524) );
  NAND2_X1 U10197 ( .A1(n13303), .A2(n13302), .ZN(n7537) );
  INV_X1 U10198 ( .A(n13309), .ZN(n7536) );
  NAND2_X1 U10199 ( .A1(n8110), .A2(n8141), .ZN(n7542) );
  NAND3_X1 U10200 ( .A1(n7548), .A2(n7550), .A3(n6512), .ZN(n7546) );
  NAND3_X1 U10201 ( .A1(n7563), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n7562) );
  NAND3_X1 U10202 ( .A1(n7581), .A2(n7579), .A3(n7580), .ZN(n7578) );
  OAI21_X1 U10203 ( .B1(n7587), .B2(n6507), .A(n7584), .ZN(n8020) );
  OAI21_X1 U10204 ( .B1(n7992), .B2(n7596), .A(n7593), .ZN(n8331) );
  NAND2_X1 U10205 ( .A1(n7992), .A2(n7593), .ZN(n7591) );
  NAND3_X1 U10206 ( .A1(n7604), .A2(n7603), .A3(n7949), .ZN(n9431) );
  AOI21_X1 U10207 ( .B1(n13803), .B2(n7944), .A(n13802), .ZN(n13804) );
  XNOR2_X1 U10208 ( .A(n8108), .B(n8107), .ZN(n10323) );
  AOI21_X1 U10209 ( .B1(n10289), .B2(n15556), .A(n10288), .ZN(n13972) );
  NAND2_X1 U10210 ( .A1(n7623), .A2(n7621), .ZN(n12308) );
  NAND2_X1 U10211 ( .A1(n12265), .A2(n7624), .ZN(n7623) );
  OAI21_X1 U10212 ( .B1(n12266), .B2(n12267), .A(n12783), .ZN(n7627) );
  NAND2_X1 U10213 ( .A1(n12706), .A2(n12705), .ZN(n12704) );
  NAND2_X1 U10214 ( .A1(n12706), .A2(n6663), .ZN(n7633) );
  AOI21_X1 U10215 ( .B1(n7637), .B2(n7635), .A(n6674), .ZN(n7634) );
  AND2_X1 U10216 ( .A1(n7638), .A2(n12736), .ZN(n7637) );
  NAND2_X1 U10217 ( .A1(n12746), .A2(n6659), .ZN(n7648) );
  INV_X1 U10218 ( .A(n10199), .ZN(n7655) );
  NAND2_X1 U10219 ( .A1(n9127), .A2(n7665), .ZN(n7664) );
  NAND2_X1 U10220 ( .A1(n8965), .A2(n7673), .ZN(n7672) );
  NAND2_X1 U10221 ( .A1(n9064), .A2(n7679), .ZN(n7678) );
  NAND2_X1 U10222 ( .A1(n8798), .A2(n7688), .ZN(n7687) );
  NAND2_X1 U10223 ( .A1(n8798), .A2(n8797), .ZN(n9202) );
  NAND2_X1 U10224 ( .A1(n7691), .A2(n8792), .ZN(n9153) );
  NAND2_X1 U10225 ( .A1(n7691), .A2(n7690), .ZN(n9177) );
  NAND2_X1 U10226 ( .A1(n8792), .A2(n12115), .ZN(n7690) );
  NAND2_X1 U10227 ( .A1(n9177), .A2(n8793), .ZN(n8795) );
  NAND2_X1 U10228 ( .A1(n14971), .A2(n6464), .ZN(n7693) );
  NAND2_X1 U10229 ( .A1(n9669), .A2(n14517), .ZN(n7700) );
  NAND2_X2 U10230 ( .A1(n10407), .A2(n10339), .ZN(n9907) );
  INV_X1 U10231 ( .A(n14778), .ZN(n7708) );
  NAND2_X1 U10232 ( .A1(n15290), .A2(n7715), .ZN(n7712) );
  NAND2_X1 U10233 ( .A1(n7726), .A2(n7724), .ZN(n11831) );
  NAND2_X1 U10234 ( .A1(n11310), .A2(n10980), .ZN(n10996) );
  AND2_X1 U10235 ( .A1(n9459), .A2(n7735), .ZN(n7734) );
  NAND2_X1 U10236 ( .A1(n10006), .A2(n10007), .ZN(n10005) );
  NAND3_X1 U10237 ( .A1(n7742), .A2(n7740), .A3(n7741), .ZN(n7738) );
  NAND2_X1 U10238 ( .A1(n10003), .A2(n7744), .ZN(n7740) );
  OAI21_X1 U10239 ( .B1(n9995), .B2(n9994), .A(n9993), .ZN(n7742) );
  NAND3_X1 U10240 ( .A1(n10103), .A2(n10102), .A3(n6619), .ZN(n7745) );
  NAND2_X1 U10241 ( .A1(n7745), .A2(n7746), .ZN(n10108) );
  NAND3_X1 U10242 ( .A1(n10120), .A2(n10119), .A3(n6620), .ZN(n7747) );
  NAND2_X1 U10243 ( .A1(n7747), .A2(n7748), .ZN(n10125) );
  NAND2_X1 U10244 ( .A1(n10098), .A2(n10099), .ZN(n10097) );
  NAND3_X1 U10245 ( .A1(n10016), .A2(n10017), .A3(n6621), .ZN(n7751) );
  NAND2_X1 U10246 ( .A1(n12021), .A2(n6477), .ZN(n14929) );
  NAND2_X1 U10247 ( .A1(n7757), .A2(n11113), .ZN(n15298) );
  NAND2_X1 U10248 ( .A1(n7764), .A2(n14781), .ZN(n7766) );
  NAND2_X2 U10249 ( .A1(n13238), .A2(n8821), .ZN(n12300) );
  NAND2_X1 U10250 ( .A1(n15674), .A2(n9218), .ZN(n7787) );
  NAND2_X1 U10251 ( .A1(n8703), .A2(n7791), .ZN(n8818) );
  NAND2_X1 U10252 ( .A1(n8703), .A2(n8702), .ZN(n8805) );
  OAI21_X1 U10253 ( .B1(n11994), .B2(n7804), .A(n7802), .ZN(n12510) );
  AOI21_X1 U10254 ( .B1(n7802), .B2(n7804), .A(n7801), .ZN(n7800) );
  INV_X1 U10255 ( .A(n11653), .ZN(n7810) );
  NAND2_X1 U10256 ( .A1(n11653), .A2(n11746), .ZN(n7808) );
  NAND3_X1 U10257 ( .A1(n7813), .A2(n7812), .A3(n6511), .ZN(n9051) );
  NAND4_X1 U10258 ( .A1(n8670), .A2(n8671), .A3(n8669), .A4(n8891), .ZN(n7814)
         );
  NAND2_X1 U10259 ( .A1(n9067), .A2(n7815), .ZN(n7818) );
  NAND2_X1 U10260 ( .A1(n9067), .A2(n8678), .ZN(n9070) );
  OAI211_X1 U10261 ( .C1(n12517), .C2(n7828), .A(n7830), .B(n6629), .ZN(n7829)
         );
  OAI21_X1 U10262 ( .B1(n12517), .B2(n12499), .A(n12498), .ZN(n12555) );
  NAND3_X1 U10263 ( .A1(n12517), .A2(n7842), .A3(n12498), .ZN(n7833) );
  NAND2_X1 U10264 ( .A1(n12500), .A2(n13051), .ZN(n7842) );
  OAI21_X1 U10265 ( .B1(n8875), .B2(n7845), .A(n7846), .ZN(n11567) );
  NAND2_X1 U10266 ( .A1(n7844), .A2(n7843), .ZN(n8930) );
  NAND2_X1 U10267 ( .A1(n8875), .A2(n7846), .ZN(n7843) );
  AOI21_X1 U10268 ( .B1(n7846), .B2(n7845), .A(n6622), .ZN(n7844) );
  INV_X1 U10269 ( .A(n8896), .ZN(n7845) );
  NAND2_X1 U10270 ( .A1(n13012), .A2(n10896), .ZN(n12161) );
  NAND2_X1 U10271 ( .A1(n12162), .A2(n10853), .ZN(n15584) );
  NAND2_X1 U10272 ( .A1(n12982), .A2(n6600), .ZN(n7855) );
  NAND3_X1 U10273 ( .A1(n7856), .A2(n7858), .A3(n12219), .ZN(n7854) );
  NAND3_X1 U10274 ( .A1(n12453), .A2(n7866), .A3(n15666), .ZN(n7864) );
  NAND2_X2 U10275 ( .A1(n8806), .A2(n6545), .ZN(n13232) );
  XNOR2_X2 U10276 ( .A(n7885), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8821) );
  NAND2_X2 U10277 ( .A1(n13232), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7885) );
  NAND2_X1 U10278 ( .A1(n7886), .A2(n7888), .ZN(n12408) );
  NAND3_X1 U10279 ( .A1(n11433), .A2(n9491), .A3(n7895), .ZN(n7894) );
  NAND2_X1 U10280 ( .A1(n14379), .A2(n7903), .ZN(n7902) );
  NOR2_X1 U10281 ( .A1(n13955), .A2(n13974), .ZN(n7914) );
  NOR2_X1 U10282 ( .A1(n13988), .A2(n13974), .ZN(n10292) );
  NOR2_X2 U10283 ( .A1(n14068), .A2(n14059), .ZN(n14058) );
  INV_X1 U10284 ( .A(n13518), .ZN(n13521) );
  XNOR2_X1 U10285 ( .A(n12344), .B(n12357), .ZN(n12362) );
  OAI21_X1 U10286 ( .B1(n13753), .B2(n13752), .A(n13751), .ZN(n13806) );
  NAND2_X1 U10287 ( .A1(n13753), .A2(n13750), .ZN(n13751) );
  INV_X1 U10288 ( .A(n9919), .ZN(n9930) );
  NAND2_X1 U10289 ( .A1(n8667), .A2(n15580), .ZN(n8663) );
  NAND2_X1 U10290 ( .A1(n10285), .A2(n7935), .ZN(n10289) );
  NAND2_X1 U10291 ( .A1(n8111), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8117) );
  NAND2_X1 U10292 ( .A1(n8111), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8084) );
  INV_X1 U10293 ( .A(n8563), .ZN(n8138) );
  INV_X1 U10294 ( .A(n11367), .ZN(n10983) );
  NAND2_X1 U10295 ( .A1(n10983), .A2(n15356), .ZN(n10984) );
  INV_X1 U10296 ( .A(n15344), .ZN(n15328) );
  OR2_X1 U10297 ( .A1(n15344), .A2(n14817), .ZN(n11044) );
  XNOR2_X1 U10298 ( .A(n14688), .B(n14717), .ZN(n15017) );
  INV_X1 U10299 ( .A(n13954), .ZN(n8624) );
  INV_X1 U10300 ( .A(n8063), .ZN(n12456) );
  INV_X1 U10301 ( .A(n8806), .ZN(n8807) );
  AOI21_X1 U10302 ( .B1(n9271), .B2(n12536), .A(n13052), .ZN(n9281) );
  INV_X1 U10303 ( .A(n10300), .ZN(n10902) );
  INV_X1 U10304 ( .A(n8821), .ZN(n12461) );
  NAND2_X1 U10305 ( .A1(n10849), .A2(n11291), .ZN(n15651) );
  AOI211_X1 U10306 ( .C1(n13946), .C2(n13945), .A(n15561), .B(n13944), .ZN(
        n14205) );
  OAI22_X1 U10307 ( .A1(n10250), .A2(n10313), .B1(n8202), .B2(n13851), .ZN(
        n8088) );
  OAI22_X1 U10308 ( .A1(n10250), .A2(n10315), .B1(n8202), .B2(n15452), .ZN(
        n8100) );
  AND3_X1 U10309 ( .A1(n13989), .A2(n14181), .A3(n13988), .ZN(n14209) );
  NAND2_X1 U10310 ( .A1(n14011), .A2(n13993), .ZN(n13988) );
  CLKBUF_X3 U10311 ( .A(n13530), .Z(n13738) );
  AND4_X1 U10312 ( .A1(n12348), .A2(n12536), .A3(n12340), .A4(n12791), .ZN(
        n7926) );
  AND2_X1 U10313 ( .A1(n14959), .A2(n14957), .ZN(n7928) );
  AND2_X1 U10314 ( .A1(n12031), .A2(n12032), .ZN(n7929) );
  XNOR2_X1 U10315 ( .A(n11478), .B(n11477), .ZN(n7930) );
  NAND2_X1 U10316 ( .A1(n9256), .A2(n9255), .ZN(n7931) );
  NAND2_X1 U10317 ( .A1(n13657), .A2(n13655), .ZN(n7932) );
  NAND2_X2 U10318 ( .A1(n11020), .A2(n15503), .ZN(n15831) );
  OR2_X1 U10319 ( .A1(n15006), .A2(n15005), .ZN(n15440) );
  AND2_X1 U10320 ( .A1(n9489), .A2(n9488), .ZN(n7933) );
  AND2_X1 U10321 ( .A1(n11772), .A2(n11771), .ZN(n7934) );
  OR2_X1 U10322 ( .A1(n15025), .A2(n15422), .ZN(n7936) );
  AND2_X1 U10323 ( .A1(n7991), .A2(n7990), .ZN(n7937) );
  AND2_X1 U10324 ( .A1(n14822), .A2(n14798), .ZN(n7938) );
  INV_X1 U10325 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10173) );
  INV_X1 U10326 ( .A(n9313), .ZN(n9345) );
  AND2_X1 U10327 ( .A1(n13955), .A2(n15525), .ZN(n7939) );
  NAND2_X1 U10328 ( .A1(n13952), .A2(n15556), .ZN(n7940) );
  AND2_X1 U10329 ( .A1(n7987), .A2(n7986), .ZN(n7941) );
  AND2_X1 U10330 ( .A1(n8002), .A2(n8001), .ZN(n7942) );
  NAND2_X1 U10331 ( .A1(n15496), .A2(n13531), .ZN(n15485) );
  AND2_X1 U10332 ( .A1(n13811), .A2(n14188), .ZN(n7943) );
  AND3_X1 U10333 ( .A1(n13801), .A2(n13936), .A3(n13792), .ZN(n7944) );
  AND2_X1 U10334 ( .A1(n11987), .A2(n11832), .ZN(n7945) );
  AND2_X1 U10335 ( .A1(n13368), .A2(n13371), .ZN(n7946) );
  NOR2_X1 U10336 ( .A1(n15664), .A2(n15651), .ZN(n13217) );
  AND2_X1 U10337 ( .A1(n15676), .A2(n15637), .ZN(n13115) );
  NOR2_X1 U10338 ( .A1(n12400), .A2(n12399), .ZN(n7947) );
  NAND2_X1 U10339 ( .A1(n13530), .A2(n13515), .ZN(n13516) );
  INV_X1 U10340 ( .A(n13519), .ZN(n13520) );
  NAND2_X1 U10341 ( .A1(n10011), .A2(n10010), .ZN(n10015) );
  NAND2_X1 U10342 ( .A1(n14869), .A2(n10124), .ZN(n10083) );
  NAND2_X1 U10343 ( .A1(n10084), .A2(n10083), .ZN(n10087) );
  INV_X1 U10344 ( .A(n12854), .ZN(n9258) );
  NAND2_X1 U10345 ( .A1(n12855), .A2(n9258), .ZN(n9259) );
  INV_X1 U10346 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9307) );
  INV_X1 U10347 ( .A(n11654), .ZN(n11651) );
  NAND2_X1 U10348 ( .A1(n7639), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n10160) );
  INV_X1 U10349 ( .A(n12326), .ZN(n9232) );
  AND2_X1 U10350 ( .A1(n8612), .A2(n15556), .ZN(n8613) );
  NAND2_X1 U10351 ( .A1(n8586), .A2(n14122), .ZN(n8587) );
  AND2_X1 U10352 ( .A1(n14699), .A2(n14884), .ZN(n14700) );
  NAND2_X1 U10353 ( .A1(n10949), .A2(n10141), .ZN(n10937) );
  NAND2_X1 U10354 ( .A1(n6475), .A2(n11783), .ZN(n10151) );
  INV_X1 U10355 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8307) );
  NOR2_X1 U10356 ( .A1(n8588), .A2(n8587), .ZN(n8589) );
  INV_X1 U10357 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n15765) );
  OAI22_X1 U10358 ( .A1(n10250), .A2(n10314), .B1(n8202), .B2(n13838), .ZN(
        n8118) );
  INV_X1 U10359 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8037) );
  AND2_X1 U10360 ( .A1(n10303), .A2(n10302), .ZN(n9487) );
  INV_X1 U10361 ( .A(n11943), .ZN(n9563) );
  XNOR2_X1 U10362 ( .A(n9945), .B(n9948), .ZN(n9946) );
  INV_X1 U10363 ( .A(n9756), .ZN(n9754) );
  INV_X1 U10364 ( .A(n15417), .ZN(n11824) );
  NAND2_X1 U10365 ( .A1(n7999), .A2(n10553), .ZN(n8002) );
  INV_X1 U10366 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8956) );
  INV_X1 U10367 ( .A(n12625), .ZN(n12470) );
  INV_X1 U10368 ( .A(n10501), .ZN(n10157) );
  INV_X1 U10369 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8672) );
  INV_X1 U10370 ( .A(n13301), .ZN(n13302) );
  NAND2_X1 U10371 ( .A1(n13732), .A2(n13733), .ZN(n13734) );
  NOR2_X1 U10372 ( .A1(n10254), .A2(n8127), .ZN(n8128) );
  INV_X1 U10373 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n15703) );
  INV_X1 U10374 ( .A(n10742), .ZN(n10740) );
  INV_X1 U10375 ( .A(n9593), .ZN(n9594) );
  INV_X1 U10376 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9499) );
  NAND2_X1 U10377 ( .A1(n9608), .A2(n9609), .ZN(n9610) );
  NAND2_X1 U10378 ( .A1(n14880), .A2(n14701), .ZN(n14709) );
  NAND2_X1 U10379 ( .A1(n9315), .A2(n9314), .ZN(n9316) );
  NAND2_X1 U10380 ( .A1(n7980), .A2(n10356), .ZN(n7983) );
  INV_X1 U10381 ( .A(n10865), .ZN(n10840) );
  INV_X1 U10382 ( .A(n12908), .ZN(n12528) );
  INV_X1 U10383 ( .A(n12822), .ZN(n13043) );
  OAI21_X1 U10384 ( .B1(n10947), .B2(n10173), .A(n10172), .ZN(n10931) );
  INV_X1 U10385 ( .A(n12637), .ZN(n13058) );
  INV_X1 U10386 ( .A(n15638), .ZN(n15652) );
  OR2_X1 U10387 ( .A1(n15601), .A2(n15652), .ZN(n12989) );
  AND2_X1 U10388 ( .A1(n8817), .A2(n8816), .ZN(n15644) );
  INV_X1 U10389 ( .A(n15656), .ZN(n15642) );
  INV_X1 U10390 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8702) );
  NAND2_X1 U10391 ( .A1(n8691), .A2(n8694), .ZN(n8725) );
  NAND2_X1 U10392 ( .A1(n10335), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8756) );
  INV_X1 U10393 ( .A(n14041), .ZN(n13400) );
  OR2_X1 U10394 ( .A1(n10605), .A2(P2_U3088), .ZN(n10604) );
  INV_X1 U10395 ( .A(n14210), .ZN(n13993) );
  OR2_X1 U10396 ( .A1(n14138), .A2(n14152), .ZN(n14140) );
  INV_X1 U10397 ( .A(n14191), .ZN(n14160) );
  INV_X1 U10398 ( .A(n15484), .ZN(n15829) );
  OR2_X1 U10399 ( .A1(n14370), .A2(n8636), .ZN(n8640) );
  INV_X1 U10400 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n14417) );
  NAND2_X1 U10401 ( .A1(n14800), .A2(n14982), .ZN(n14759) );
  NAND2_X1 U10402 ( .A1(n11823), .A2(n11822), .ZN(n12027) );
  INV_X2 U10403 ( .A(n12411), .ZN(n12425) );
  NAND2_X1 U10404 ( .A1(n10972), .A2(n10971), .ZN(n14997) );
  NAND2_X1 U10405 ( .A1(n8429), .A2(n8415), .ZN(n8417) );
  INV_X1 U10406 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9320) );
  INV_X1 U10407 ( .A(n12634), .ZN(n12589) );
  OR2_X1 U10408 ( .A1(n12300), .A2(n8822), .ZN(n8825) );
  INV_X1 U10409 ( .A(n12755), .ZN(n12675) );
  INV_X1 U10410 ( .A(n12750), .ZN(n12692) );
  INV_X1 U10411 ( .A(n12815), .ZN(n12809) );
  NAND2_X1 U10412 ( .A1(n10841), .A2(n11394), .ZN(n15588) );
  INV_X1 U10413 ( .A(n12804), .ZN(n13004) );
  AND2_X1 U10414 ( .A1(n15602), .A2(n15676), .ZN(n13049) );
  AND3_X1 U10415 ( .A1(n9285), .A2(n9291), .A3(n8727), .ZN(n11390) );
  AND2_X1 U10416 ( .A1(n15644), .A2(n15659), .ZN(n13138) );
  INV_X1 U10417 ( .A(n13052), .ZN(n15611) );
  AND2_X1 U10418 ( .A1(n8763), .A2(n8762), .ZN(n8979) );
  INV_X1 U10419 ( .A(n13491), .ZN(n13474) );
  AND2_X1 U10420 ( .A1(n11232), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13495) );
  OR2_X1 U10421 ( .A1(n8131), .A2(n8179), .ZN(n8187) );
  NOR2_X1 U10422 ( .A1(n10914), .A2(n10915), .ZN(n11260) );
  INV_X1 U10423 ( .A(n11268), .ZN(n11375) );
  NOR2_X1 U10424 ( .A1(n10604), .A2(n10603), .ZN(n15447) );
  INV_X1 U10425 ( .A(n15495), .ZN(n14188) );
  XNOR2_X1 U10426 ( .A(n13825), .B(n14307), .ZN(n13765) );
  INV_X1 U10427 ( .A(n14350), .ZN(n10258) );
  NAND2_X2 U10428 ( .A1(n13748), .A2(n8611), .ZN(n15556) );
  INV_X1 U10429 ( .A(n14271), .ZN(n14310) );
  AND2_X1 U10430 ( .A1(n8640), .A2(n8654), .ZN(n15509) );
  AND2_X1 U10431 ( .A1(n9833), .A2(n9830), .ZN(n14496) );
  INV_X1 U10432 ( .A(n14645), .ZN(n15270) );
  AND2_X1 U10433 ( .A1(n10515), .A2(n10479), .ZN(n15277) );
  OR2_X1 U10434 ( .A1(n10971), .A2(n11837), .ZN(n10457) );
  AND2_X1 U10435 ( .A1(n9845), .A2(n10511), .ZN(n14982) );
  NAND2_X1 U10436 ( .A1(n10989), .A2(n10988), .ZN(n15359) );
  INV_X1 U10437 ( .A(n15311), .ZN(n14995) );
  NAND2_X1 U10438 ( .A1(n9811), .A2(n10393), .ZN(n15005) );
  INV_X1 U10439 ( .A(n15359), .ZN(n15400) );
  INV_X1 U10440 ( .A(n15402), .ZN(n15422) );
  NAND2_X1 U10441 ( .A1(n15305), .A2(n15393), .ZN(n15402) );
  AND2_X1 U10442 ( .A1(n10296), .A2(n10397), .ZN(n10971) );
  NAND2_X1 U10443 ( .A1(n9321), .A2(n9320), .ZN(n9406) );
  AND2_X1 U10444 ( .A1(n10196), .A2(n10195), .ZN(n15581) );
  INV_X1 U10445 ( .A(n12631), .ZN(n12610) );
  NAND2_X1 U10446 ( .A1(n10866), .A2(n10865), .ZN(n12634) );
  INV_X1 U10447 ( .A(n12352), .ZN(n12760) );
  INV_X1 U10448 ( .A(n13051), .ZN(n13035) );
  INV_X1 U10449 ( .A(n13091), .ZN(n12640) );
  INV_X1 U10450 ( .A(n13010), .ZN(n13007) );
  INV_X1 U10451 ( .A(n13049), .ZN(n13118) );
  INV_X1 U10452 ( .A(n13151), .ZN(n13220) );
  AND2_X1 U10453 ( .A1(n9293), .A2(n9292), .ZN(n15664) );
  OR2_X1 U10454 ( .A1(n12155), .A2(n12154), .ZN(n12156) );
  INV_X1 U10455 ( .A(SI_16_), .ZN(n10553) );
  INV_X1 U10456 ( .A(SI_13_), .ZN(n10510) );
  OR2_X1 U10457 ( .A1(n13461), .A2(n15493), .ZN(n13491) );
  OR3_X1 U10458 ( .A1(n10749), .A2(n10736), .A3(n15525), .ZN(n13481) );
  INV_X1 U10459 ( .A(n15475), .ZN(n15445) );
  INV_X1 U10460 ( .A(n15447), .ZN(n15465) );
  INV_X1 U10461 ( .A(n15827), .ZN(n15504) );
  AND2_X1 U10462 ( .A1(n14080), .A2(n14079), .ZN(n14251) );
  NAND2_X1 U10463 ( .A1(n15831), .A2(n11351), .ZN(n14200) );
  NAND2_X1 U10464 ( .A1(n13718), .A2(n14280), .ZN(n10262) );
  INV_X1 U10465 ( .A(n14092), .ZN(n14335) );
  INV_X1 U10466 ( .A(n14166), .ZN(n14346) );
  INV_X1 U10467 ( .A(n15571), .ZN(n15569) );
  AND2_X2 U10468 ( .A1(n8666), .A2(n8665), .ZN(n15571) );
  INV_X1 U10469 ( .A(n15510), .ZN(n15511) );
  INV_X1 U10470 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10669) );
  INV_X1 U10471 ( .A(n15076), .ZN(n14899) );
  XNOR2_X1 U10472 ( .A(n9806), .B(n9805), .ZN(n9850) );
  NAND2_X1 U10473 ( .A1(n10658), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14494) );
  NAND2_X1 U10474 ( .A1(n9828), .A2(n9827), .ZN(n14498) );
  NAND2_X1 U10475 ( .A1(n9934), .A2(n9933), .ZN(n14740) );
  INV_X1 U10476 ( .A(n14869), .ZN(n14904) );
  INV_X1 U10477 ( .A(n11981), .ZN(n14503) );
  OR2_X1 U10478 ( .A1(n15336), .A2(n15400), .ZN(n14970) );
  OR2_X1 U10479 ( .A1(n15336), .A2(n14910), .ZN(n14990) );
  NOR2_X1 U10480 ( .A1(n15006), .A2(n11048), .ZN(n15149) );
  INV_X1 U10481 ( .A(n15149), .ZN(n15424) );
  AND2_X1 U10482 ( .A1(n10404), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10397) );
  INV_X1 U10483 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10872) );
  INV_X1 U10484 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10487) );
  INV_X1 U10485 ( .A(n10295), .ZN(P2_U3526) );
  INV_X1 U10486 ( .A(n14525), .ZN(P1_U4016) );
  OAI21_X1 U10487 ( .B1(n9850), .B2(n14498), .A(n9849), .ZN(P1_U3225) );
  MUX2_X1 U10488 ( .A(n10322), .B(n10315), .S(n6442), .Z(n7955) );
  INV_X1 U10489 ( .A(SI_3_), .ZN(n10422) );
  NAND2_X1 U10490 ( .A1(n7955), .A2(n10422), .ZN(n7954) );
  AND2_X1 U10491 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n7949) );
  AND2_X1 U10492 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7950) );
  NAND2_X1 U10493 ( .A1(n6442), .A2(n7950), .ZN(n8136) );
  INV_X1 U10494 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10342) );
  AOI21_X1 U10495 ( .B1(n6443), .B2(P1_DATAO_REG_1__SCAN_IN), .A(SI_1_), .ZN(
        n7951) );
  NAND2_X1 U10496 ( .A1(n6443), .A2(n10314), .ZN(n8120) );
  OAI211_X1 U10497 ( .C1(P2_DATAO_REG_1__SCAN_IN), .C2(n6442), .A(n8120), .B(
        SI_1_), .ZN(n7952) );
  NAND2_X1 U10498 ( .A1(n8089), .A2(SI_2_), .ZN(n8103) );
  NAND2_X1 U10499 ( .A1(n8103), .A2(n10422), .ZN(n7956) );
  INV_X1 U10500 ( .A(n7955), .ZN(n8106) );
  NAND2_X1 U10501 ( .A1(n7956), .A2(n8106), .ZN(n8146) );
  AND2_X1 U10502 ( .A1(SI_2_), .A2(SI_3_), .ZN(n7957) );
  NAND2_X1 U10503 ( .A1(n8089), .A2(n7957), .ZN(n8145) );
  NAND2_X1 U10504 ( .A1(n8148), .A2(SI_4_), .ZN(n8156) );
  AND2_X1 U10505 ( .A1(n8145), .A2(n8156), .ZN(n7958) );
  NOR2_X1 U10506 ( .A1(n8148), .A2(SI_4_), .ZN(n7959) );
  NOR2_X1 U10507 ( .A1(n8158), .A2(n7959), .ZN(n7960) );
  NAND2_X1 U10508 ( .A1(n7965), .A2(SI_7_), .ZN(n8241) );
  INV_X1 U10509 ( .A(n8241), .ZN(n7962) );
  MUX2_X1 U10510 ( .A(n10330), .B(n10331), .S(n6442), .Z(n8189) );
  INV_X1 U10511 ( .A(n8189), .ZN(n7964) );
  NAND2_X1 U10512 ( .A1(n7964), .A2(SI_6_), .ZN(n8198) );
  NAND2_X1 U10513 ( .A1(n7961), .A2(SI_5_), .ZN(n8188) );
  NAND2_X1 U10514 ( .A1(n8198), .A2(n8188), .ZN(n8236) );
  NOR2_X1 U10515 ( .A1(n7962), .A2(n8236), .ZN(n7963) );
  NAND2_X1 U10516 ( .A1(n8238), .A2(n7963), .ZN(n7969) );
  MUX2_X1 U10517 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n6443), .Z(n7970) );
  XNOR2_X1 U10518 ( .A(n7970), .B(SI_8_), .ZN(n8243) );
  AOI21_X1 U10519 ( .B1(n7967), .B2(n8241), .A(n8243), .ZN(n7968) );
  NAND2_X1 U10520 ( .A1(n7969), .A2(n7968), .ZN(n7972) );
  NAND2_X1 U10521 ( .A1(n7970), .A2(SI_8_), .ZN(n7971) );
  MUX2_X1 U10522 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n6443), .Z(n7974) );
  XNOR2_X1 U10523 ( .A(n7974), .B(SI_9_), .ZN(n8212) );
  INV_X1 U10524 ( .A(n8212), .ZN(n7973) );
  NAND2_X1 U10525 ( .A1(n8211), .A2(n7973), .ZN(n7976) );
  NAND2_X1 U10526 ( .A1(n7974), .A2(SI_9_), .ZN(n7975) );
  XNOR2_X1 U10527 ( .A(n7978), .B(SI_10_), .ZN(n8261) );
  INV_X1 U10528 ( .A(n8261), .ZN(n7977) );
  NAND2_X1 U10529 ( .A1(n7978), .A2(SI_10_), .ZN(n7979) );
  INV_X1 U10530 ( .A(n7980), .ZN(n7981) );
  NAND2_X1 U10531 ( .A1(n7981), .A2(SI_11_), .ZN(n7982) );
  NAND2_X1 U10532 ( .A1(n7983), .A2(n7982), .ZN(n8269) );
  MUX2_X1 U10533 ( .A(n10487), .B(n10485), .S(n6442), .Z(n7984) );
  INV_X1 U10534 ( .A(n7984), .ZN(n7985) );
  NAND2_X1 U10535 ( .A1(n7985), .A2(SI_12_), .ZN(n7986) );
  MUX2_X1 U10536 ( .A(n10507), .B(n10505), .S(n10338), .Z(n7988) );
  INV_X1 U10537 ( .A(n7988), .ZN(n7989) );
  NAND2_X1 U10538 ( .A1(n7989), .A2(SI_13_), .ZN(n7990) );
  MUX2_X1 U10539 ( .A(n10555), .B(n10558), .S(n10338), .Z(n8317) );
  NAND2_X1 U10540 ( .A1(n7993), .A2(SI_14_), .ZN(n7994) );
  MUX2_X1 U10541 ( .A(n10670), .B(n10669), .S(n10338), .Z(n7995) );
  INV_X1 U10542 ( .A(n7995), .ZN(n7996) );
  NAND2_X1 U10543 ( .A1(n7996), .A2(SI_15_), .ZN(n7997) );
  MUX2_X1 U10544 ( .A(n10715), .B(n10713), .S(n10338), .Z(n7999) );
  INV_X1 U10545 ( .A(n7999), .ZN(n8000) );
  NAND2_X1 U10546 ( .A1(n8000), .A2(SI_16_), .ZN(n8001) );
  MUX2_X1 U10547 ( .A(n10872), .B(n10874), .S(n6443), .Z(n8368) );
  INV_X1 U10548 ( .A(n8368), .ZN(n8003) );
  NAND2_X1 U10549 ( .A1(n8003), .A2(SI_17_), .ZN(n8004) );
  INV_X1 U10550 ( .A(SI_17_), .ZN(n10566) );
  NAND2_X1 U10551 ( .A1(n8368), .A2(n10566), .ZN(n8005) );
  MUX2_X1 U10552 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n10338), .Z(n8381) );
  NOR2_X1 U10553 ( .A1(n8381), .A2(SI_18_), .ZN(n8007) );
  NAND2_X1 U10554 ( .A1(n8381), .A2(SI_18_), .ZN(n8006) );
  MUX2_X1 U10555 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n10338), .Z(n8008) );
  INV_X1 U10556 ( .A(n8008), .ZN(n8009) );
  INV_X1 U10557 ( .A(SI_19_), .ZN(n10716) );
  NAND2_X1 U10558 ( .A1(n8009), .A2(n10716), .ZN(n8010) );
  MUX2_X1 U10559 ( .A(n11708), .B(n15733), .S(n10338), .Z(n8012) );
  INV_X1 U10560 ( .A(SI_21_), .ZN(n12379) );
  INV_X1 U10561 ( .A(SI_20_), .ZN(n10964) );
  MUX2_X1 U10562 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n10338), .Z(n8416) );
  INV_X1 U10563 ( .A(n8012), .ZN(n8013) );
  MUX2_X1 U10564 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n10338), .Z(n8444) );
  INV_X1 U10565 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8015) );
  MUX2_X1 U10566 ( .A(n8015), .B(n11863), .S(n10338), .Z(n8017) );
  INV_X1 U10567 ( .A(SI_23_), .ZN(n11559) );
  NAND2_X1 U10568 ( .A1(n8017), .A2(n11559), .ZN(n8463) );
  INV_X1 U10569 ( .A(n8463), .ZN(n8019) );
  INV_X1 U10570 ( .A(n8017), .ZN(n8018) );
  NAND2_X1 U10571 ( .A1(n8018), .A2(SI_23_), .ZN(n8462) );
  INV_X1 U10572 ( .A(n8020), .ZN(n8021) );
  INV_X1 U10573 ( .A(n8024), .ZN(n8023) );
  INV_X1 U10574 ( .A(SI_24_), .ZN(n11820) );
  MUX2_X1 U10575 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n10338), .Z(n8477) );
  MUX2_X1 U10576 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n10338), .Z(n8025) );
  XNOR2_X1 U10577 ( .A(n8025), .B(SI_25_), .ZN(n8070) );
  MUX2_X1 U10578 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n10338), .Z(n8026) );
  OAI21_X1 U10579 ( .B1(SI_26_), .B2(n8026), .A(n8494), .ZN(n8027) );
  NAND2_X1 U10580 ( .A1(n8028), .A2(n8027), .ZN(n8029) );
  INV_X1 U10581 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8034) );
  NAND4_X1 U10582 ( .A1(n8097), .A2(n8098), .A3(n8149), .A4(n8037), .ZN(n8162)
         );
  NAND4_X1 U10583 ( .A1(n8216), .A2(n8214), .A3(n8039), .A4(n8038), .ZN(n8284)
         );
  INV_X1 U10584 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14368) );
  OR2_X1 U10585 ( .A1(n7177), .A2(n14368), .ZN(n8045) );
  INV_X1 U10586 ( .A(n8182), .ZN(n8046) );
  OR2_X2 U10587 ( .A1(n8231), .A2(n8221), .ZN(n8254) );
  INV_X1 U10588 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8355) );
  INV_X1 U10589 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8374) );
  INV_X1 U10590 ( .A(n8388), .ZN(n8050) );
  INV_X1 U10591 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13446) );
  OR2_X2 U10592 ( .A1(n8421), .A2(n13446), .ZN(n8452) );
  NAND2_X1 U10593 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .ZN(n8052) );
  OR2_X2 U10594 ( .A1(n8452), .A2(n8052), .ZN(n8468) );
  INV_X1 U10595 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8074) );
  INV_X1 U10596 ( .A(n8076), .ZN(n8055) );
  INV_X1 U10597 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8056) );
  NAND2_X1 U10598 ( .A1(n8076), .A2(n8056), .ZN(n8057) );
  NAND2_X1 U10599 ( .A1(n8500), .A2(n8057), .ZN(n13475) );
  INV_X1 U10600 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8066) );
  OR2_X2 U10601 ( .A1(n8063), .A2(n14363), .ZN(n8131) );
  NAND2_X1 U10602 ( .A1(n8531), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8065) );
  NAND2_X1 U10603 ( .A1(n8532), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8064) );
  OAI211_X1 U10604 ( .C1(n8066), .C2(n8535), .A(n8065), .B(n8064), .ZN(n8067)
         );
  INV_X1 U10605 ( .A(n8067), .ZN(n8068) );
  NAND2_X2 U10606 ( .A1(n8069), .A2(n8068), .ZN(n14004) );
  XNOR2_X1 U10607 ( .A(n8071), .B(n8070), .ZN(n14371) );
  INV_X1 U10608 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n14373) );
  OR2_X1 U10609 ( .A1(n7177), .A2(n14373), .ZN(n8072) );
  NAND2_X1 U10610 ( .A1(n8485), .A2(n8074), .ZN(n8075) );
  NAND2_X1 U10611 ( .A1(n14012), .A2(n8112), .ZN(n8081) );
  INV_X1 U10612 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n15747) );
  NAND2_X1 U10613 ( .A1(n8531), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8078) );
  NAND2_X1 U10614 ( .A1(n8532), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8077) );
  OAI211_X1 U10615 ( .C1(n15747), .C2(n8535), .A(n8078), .B(n8077), .ZN(n8079)
         );
  INV_X1 U10616 ( .A(n8079), .ZN(n8080) );
  NAND2_X1 U10617 ( .A1(n8113), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8085) );
  INV_X1 U10618 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11185) );
  INV_X1 U10619 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10568) );
  OR2_X1 U10620 ( .A1(n8131), .A2(n10568), .ZN(n8082) );
  NAND2_X1 U10621 ( .A1(n13832), .A2(n8086), .ZN(n8096) );
  INV_X1 U10622 ( .A(SI_2_), .ZN(n10430) );
  XNOR2_X1 U10623 ( .A(n8089), .B(n10430), .ZN(n8101) );
  XNOR2_X1 U10624 ( .A(n8102), .B(n8101), .ZN(n10320) );
  OR2_X1 U10625 ( .A1(n8123), .A2(n10320), .ZN(n8090) );
  NAND2_X1 U10626 ( .A1(n13829), .A2(n15533), .ZN(n8564) );
  NAND2_X1 U10627 ( .A1(n11210), .A2(n8564), .ZN(n11179) );
  NAND2_X1 U10628 ( .A1(n11298), .A2(n15533), .ZN(n11205) );
  INV_X1 U10629 ( .A(n11205), .ZN(n8109) );
  INV_X1 U10630 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11216) );
  NAND2_X1 U10631 ( .A1(n8111), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8092) );
  INV_X1 U10632 ( .A(n8096), .ZN(n8163) );
  NAND2_X1 U10633 ( .A1(n8163), .A2(n8097), .ZN(n8150) );
  XNOR2_X1 U10634 ( .A(n8099), .B(n8098), .ZN(n15452) );
  INV_X1 U10635 ( .A(n8101), .ZN(n8105) );
  INV_X1 U10636 ( .A(n8102), .ZN(n8104) );
  XNOR2_X1 U10637 ( .A(n8106), .B(n10422), .ZN(n8107) );
  OAI21_X1 U10638 ( .B1(n11179), .B2(n8109), .A(n13763), .ZN(n8110) );
  INV_X1 U10639 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10567) );
  OR2_X1 U10640 ( .A1(n8131), .A2(n10567), .ZN(n8116) );
  INV_X1 U10641 ( .A(n8126), .ZN(n8112) );
  NAND2_X1 U10642 ( .A1(n8112), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8115) );
  NAND2_X1 U10643 ( .A1(n8113), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8114) );
  XNOR2_X1 U10644 ( .A(n8119), .B(SI_1_), .ZN(n8122) );
  XNOR2_X1 U10645 ( .A(n8122), .B(n8121), .ZN(n10343) );
  OR2_X1 U10646 ( .A1(n8123), .A2(n10343), .ZN(n8124) );
  NAND2_X2 U10647 ( .A1(n8125), .A2(n8124), .ZN(n15524) );
  XNOR2_X1 U10648 ( .A(n13508), .B(n15524), .ZN(n8563) );
  NAND2_X1 U10649 ( .A1(n8111), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8134) );
  INV_X1 U10650 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11027) );
  INV_X1 U10651 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n8127) );
  INV_X1 U10652 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n8130) );
  OR2_X1 U10653 ( .A1(n8131), .A2(n8130), .ZN(n8132) );
  NAND3_X2 U10654 ( .A1(n8134), .A2(n8133), .A3(n8132), .ZN(n13507) );
  NAND2_X1 U10655 ( .A1(n6443), .A2(SI_0_), .ZN(n8135) );
  NAND2_X1 U10656 ( .A1(n8135), .A2(n8731), .ZN(n8137) );
  AND2_X1 U10657 ( .A1(n8136), .A2(n8137), .ZN(n14376) );
  MUX2_X1 U10658 ( .A(P2_IR_REG_0__SCAN_IN), .B(n14376), .S(n8202), .Z(n13503)
         );
  INV_X1 U10659 ( .A(n12371), .ZN(n11025) );
  INV_X1 U10660 ( .A(n13508), .ZN(n10882) );
  INV_X1 U10661 ( .A(n15524), .ZN(n13512) );
  NAND2_X1 U10662 ( .A1(n10882), .A2(n13512), .ZN(n11174) );
  AND2_X1 U10663 ( .A1(n11205), .A2(n11174), .ZN(n8139) );
  NAND2_X1 U10664 ( .A1(n8111), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8144) );
  INV_X1 U10665 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10589) );
  OR2_X1 U10666 ( .A1(n10254), .A2(n10589), .ZN(n8143) );
  OR2_X1 U10667 ( .A1(n8131), .A2(n15576), .ZN(n8142) );
  XNOR2_X1 U10668 ( .A(P2_REG3_REG_3__SCAN_IN), .B(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n15502) );
  NAND3_X1 U10669 ( .A1(n8147), .A2(n8146), .A3(n8145), .ZN(n8155) );
  INV_X1 U10670 ( .A(SI_4_), .ZN(n10435) );
  XNOR2_X1 U10671 ( .A(n8148), .B(n10435), .ZN(n8154) );
  XNOR2_X1 U10672 ( .A(n8155), .B(n8154), .ZN(n10318) );
  NAND2_X1 U10673 ( .A1(n8160), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8151) );
  OR2_X1 U10674 ( .A1(n8202), .A2(n13861), .ZN(n8153) );
  NAND2_X1 U10675 ( .A1(n8155), .A2(n8154), .ZN(n8157) );
  NAND2_X1 U10676 ( .A1(n8157), .A2(n8156), .ZN(n8159) );
  XNOR2_X1 U10677 ( .A(n8158), .B(n8159), .ZN(n10325) );
  NAND2_X1 U10678 ( .A1(n10248), .A2(n10325), .ZN(n8166) );
  MUX2_X1 U10679 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8161), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n8164) );
  NAND2_X1 U10680 ( .A1(n8164), .A2(n8346), .ZN(n10680) );
  OR2_X1 U10681 ( .A1(n8202), .A2(n10680), .ZN(n8165) );
  NAND2_X1 U10682 ( .A1(n8113), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8173) );
  INV_X1 U10683 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10672) );
  OR2_X1 U10684 ( .A1(n8131), .A2(n10672), .ZN(n8172) );
  INV_X1 U10685 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8168) );
  NAND2_X1 U10686 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n8167) );
  NAND2_X1 U10687 ( .A1(n8168), .A2(n8167), .ZN(n8169) );
  NAND2_X1 U10688 ( .A1(n8182), .A2(n8169), .ZN(n13416) );
  OR2_X1 U10689 ( .A1(n8530), .A2(n13416), .ZN(n8171) );
  NAND2_X1 U10690 ( .A1(n8111), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8170) );
  AOI22_X1 U10691 ( .A1(n13827), .A2(n13762), .B1(n15826), .B2(n13826), .ZN(
        n8174) );
  AOI21_X1 U10692 ( .B1(n15545), .B2(n15544), .A(n15494), .ZN(n8176) );
  NAND3_X1 U10693 ( .A1(n15494), .A2(n15544), .A3(n15545), .ZN(n8175) );
  OAI21_X1 U10694 ( .B1(n8176), .B2(n15826), .A(n8175), .ZN(n8177) );
  INV_X1 U10695 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n8179) );
  NAND2_X1 U10696 ( .A1(n8111), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8186) );
  INV_X1 U10697 ( .A(n8180), .ZN(n8205) );
  INV_X1 U10698 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8181) );
  NAND2_X1 U10699 ( .A1(n8182), .A2(n8181), .ZN(n8183) );
  NAND2_X1 U10700 ( .A1(n8205), .A2(n8183), .ZN(n11486) );
  OR2_X1 U10701 ( .A1(n8530), .A2(n11486), .ZN(n8185) );
  INV_X1 U10702 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11357) );
  OR2_X1 U10703 ( .A1(n10254), .A2(n11357), .ZN(n8184) );
  NAND4_X1 U10704 ( .A1(n8187), .A2(n8186), .A3(n8185), .A4(n8184), .ZN(n13825) );
  NAND2_X1 U10705 ( .A1(n8238), .A2(n8188), .ZN(n8197) );
  XNOR2_X1 U10706 ( .A(n8189), .B(SI_6_), .ZN(n8196) );
  INV_X1 U10707 ( .A(n8196), .ZN(n8190) );
  XNOR2_X1 U10708 ( .A(n8197), .B(n8190), .ZN(n10329) );
  NAND2_X1 U10709 ( .A1(n10329), .A2(n10248), .ZN(n8194) );
  NAND2_X1 U10710 ( .A1(n8346), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8192) );
  INV_X1 U10711 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8191) );
  XNOR2_X1 U10712 ( .A(n8192), .B(n8191), .ZN(n15464) );
  OR2_X1 U10713 ( .A1(n8202), .A2(n15464), .ZN(n8193) );
  INV_X1 U10714 ( .A(n13765), .ZN(n11354) );
  INV_X1 U10715 ( .A(n13825), .ZN(n11582) );
  INV_X1 U10716 ( .A(n14307), .ZN(n13554) );
  NAND2_X1 U10717 ( .A1(n11582), .A2(n13554), .ZN(n8195) );
  NAND2_X1 U10718 ( .A1(n8197), .A2(n8196), .ZN(n8199) );
  NAND2_X1 U10719 ( .A1(n8199), .A2(n8198), .ZN(n8201) );
  XNOR2_X1 U10720 ( .A(n8201), .B(n8200), .ZN(n10345) );
  NAND2_X1 U10721 ( .A1(n8213), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8203) );
  XNOR2_X1 U10722 ( .A(n8203), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10612) );
  NAND2_X1 U10723 ( .A1(n8111), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8209) );
  INV_X1 U10724 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8204) );
  NAND2_X1 U10725 ( .A1(n8205), .A2(n8204), .ZN(n8206) );
  NAND2_X1 U10726 ( .A1(n8229), .A2(n8206), .ZN(n11583) );
  OR2_X1 U10727 ( .A1(n8530), .A2(n11583), .ZN(n8208) );
  INV_X1 U10728 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11412) );
  OR2_X1 U10729 ( .A1(n10254), .A2(n11412), .ZN(n8207) );
  INV_X1 U10730 ( .A(n13824), .ZN(n11487) );
  NAND2_X1 U10731 ( .A1(n11487), .A2(n11588), .ZN(n8210) );
  XNOR2_X1 U10732 ( .A(n8211), .B(n8212), .ZN(n10349) );
  NAND2_X1 U10733 ( .A1(n10349), .A2(n10248), .ZN(n8220) );
  INV_X1 U10734 ( .A(n8213), .ZN(n8215) );
  INV_X1 U10735 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n8214) );
  NAND2_X1 U10736 ( .A1(n8215), .A2(n8214), .ZN(n8245) );
  INV_X1 U10737 ( .A(n8245), .ZN(n8217) );
  NAND2_X1 U10738 ( .A1(n8217), .A2(n8216), .ZN(n8262) );
  NAND2_X1 U10739 ( .A1(n8262), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8218) );
  XNOR2_X1 U10740 ( .A(n8218), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10720) );
  AOI22_X1 U10741 ( .A1(n8403), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n10576), 
        .B2(n10720), .ZN(n8219) );
  NAND2_X1 U10742 ( .A1(n8532), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8227) );
  NAND2_X1 U10743 ( .A1(n8111), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8226) );
  NAND2_X1 U10744 ( .A1(n8231), .A2(n8221), .ZN(n8222) );
  NAND2_X1 U10745 ( .A1(n8254), .A2(n8222), .ZN(n11764) );
  OR2_X1 U10746 ( .A1(n8530), .A2(n11764), .ZN(n8225) );
  INV_X1 U10747 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n8223) );
  OR2_X1 U10748 ( .A1(n8131), .A2(n8223), .ZN(n8224) );
  NAND4_X1 U10749 ( .A1(n8227), .A2(n8226), .A3(n8225), .A4(n8224), .ZN(n13822) );
  NAND2_X1 U10750 ( .A1(n8531), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8235) );
  NAND2_X1 U10751 ( .A1(n8532), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8234) );
  INV_X1 U10752 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8228) );
  NAND2_X1 U10753 ( .A1(n8229), .A2(n8228), .ZN(n8230) );
  NAND2_X1 U10754 ( .A1(n8231), .A2(n8230), .ZN(n11697) );
  OR2_X1 U10755 ( .A1(n8530), .A2(n11697), .ZN(n8233) );
  INV_X1 U10756 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15719) );
  OR2_X1 U10757 ( .A1(n8535), .A2(n15719), .ZN(n8232) );
  INV_X1 U10758 ( .A(n8236), .ZN(n8237) );
  NAND2_X1 U10759 ( .A1(n8238), .A2(n8237), .ZN(n8240) );
  NAND2_X1 U10760 ( .A1(n8240), .A2(n8239), .ZN(n8242) );
  NAND2_X1 U10761 ( .A1(n8242), .A2(n8241), .ZN(n8244) );
  XNOR2_X1 U10762 ( .A(n8244), .B(n8243), .ZN(n10333) );
  NAND2_X1 U10763 ( .A1(n10333), .A2(n10248), .ZN(n8248) );
  XNOR2_X1 U10764 ( .A(n8246), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10627) );
  AOI22_X1 U10765 ( .A1(n8403), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n10576), 
        .B2(n10627), .ZN(n8247) );
  OAI22_X1 U10766 ( .A1(n14301), .A2(n13822), .B1(n13823), .B2(n13567), .ZN(
        n8252) );
  NAND2_X1 U10767 ( .A1(n13823), .A2(n13567), .ZN(n11758) );
  INV_X1 U10768 ( .A(n13822), .ZN(n11867) );
  NAND2_X1 U10769 ( .A1(n11758), .A2(n11867), .ZN(n8250) );
  AND2_X1 U10770 ( .A1(n13822), .A2(n13823), .ZN(n8249) );
  AOI22_X1 U10771 ( .A1(n8250), .A2(n14301), .B1(n8249), .B2(n13567), .ZN(
        n8251) );
  NAND2_X1 U10772 ( .A1(n8111), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8259) );
  NAND2_X1 U10773 ( .A1(n8531), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8258) );
  NAND2_X1 U10774 ( .A1(n8254), .A2(n8253), .ZN(n8255) );
  NAND2_X1 U10775 ( .A1(n8275), .A2(n8255), .ZN(n11871) );
  OR2_X1 U10776 ( .A1(n8530), .A2(n11871), .ZN(n8257) );
  INV_X1 U10777 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11872) );
  OR2_X1 U10778 ( .A1(n10254), .A2(n11872), .ZN(n8256) );
  NAND4_X1 U10779 ( .A1(n8259), .A2(n8258), .A3(n8257), .A4(n8256), .ZN(n13821) );
  XNOR2_X1 U10780 ( .A(n8260), .B(n8261), .ZN(n10400) );
  NAND2_X1 U10781 ( .A1(n10400), .A2(n10248), .ZN(n8265) );
  NAND2_X1 U10782 ( .A1(n8270), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8263) );
  XNOR2_X1 U10783 ( .A(n8263), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10723) );
  AOI22_X1 U10784 ( .A1(n8403), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n10576), 
        .B2(n10723), .ZN(n8264) );
  OR2_X1 U10785 ( .A1(n13821), .A2(n13581), .ZN(n8266) );
  NAND2_X1 U10786 ( .A1(n13581), .A2(n13821), .ZN(n8267) );
  XNOR2_X1 U10787 ( .A(n8268), .B(n8269), .ZN(n10409) );
  NAND2_X1 U10788 ( .A1(n10409), .A2(n10248), .ZN(n8273) );
  XNOR2_X1 U10789 ( .A(n8271), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10917) );
  AOI22_X1 U10790 ( .A1(n8403), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n10576), 
        .B2(n10917), .ZN(n8272) );
  NAND2_X1 U10791 ( .A1(n8532), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8280) );
  NAND2_X1 U10792 ( .A1(n8111), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8279) );
  INV_X1 U10793 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8274) );
  NAND2_X1 U10794 ( .A1(n8275), .A2(n8274), .ZN(n8276) );
  NAND2_X1 U10795 ( .A1(n8293), .A2(n8276), .ZN(n11886) );
  OR2_X1 U10796 ( .A1(n8530), .A2(n11886), .ZN(n8278) );
  INV_X1 U10797 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10910) );
  OR2_X1 U10798 ( .A1(n8131), .A2(n10910), .ZN(n8277) );
  NAND4_X1 U10799 ( .A1(n8280), .A2(n8279), .A3(n8278), .A4(n8277), .ZN(n13820) );
  AND2_X1 U10800 ( .A1(n13585), .A2(n13820), .ZN(n8282) );
  OR2_X1 U10801 ( .A1(n13585), .A2(n13820), .ZN(n8281) );
  XNOR2_X1 U10802 ( .A(n8283), .B(n7941), .ZN(n10484) );
  NAND2_X1 U10803 ( .A1(n10484), .A2(n10248), .ZN(n8291) );
  NAND2_X1 U10804 ( .A1(n6947), .A2(n8285), .ZN(n8347) );
  NAND2_X1 U10805 ( .A1(n8288), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8286) );
  MUX2_X1 U10806 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8286), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n8287) );
  INV_X1 U10807 ( .A(n8287), .ZN(n8289) );
  NOR2_X1 U10808 ( .A1(n8288), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n8303) );
  NOR2_X1 U10809 ( .A1(n8289), .A2(n8303), .ZN(n11258) );
  AOI22_X1 U10810 ( .A1(n8403), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n10576), 
        .B2(n11258), .ZN(n8290) );
  NAND2_X1 U10811 ( .A1(n8531), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8298) );
  NAND2_X1 U10812 ( .A1(n8111), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8297) );
  INV_X1 U10813 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8292) );
  NAND2_X1 U10814 ( .A1(n8293), .A2(n8292), .ZN(n8294) );
  NAND2_X1 U10815 ( .A1(n8308), .A2(n8294), .ZN(n12140) );
  OR2_X1 U10816 ( .A1(n8530), .A2(n12140), .ZN(n8296) );
  INV_X1 U10817 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11899) );
  OR2_X1 U10818 ( .A1(n10254), .A2(n11899), .ZN(n8295) );
  NAND4_X1 U10819 ( .A1(n8298), .A2(n8297), .A3(n8296), .A4(n8295), .ZN(n14189) );
  INV_X1 U10820 ( .A(n13590), .ZN(n11902) );
  INV_X1 U10821 ( .A(n14189), .ZN(n12148) );
  XNOR2_X1 U10822 ( .A(n8299), .B(n7937), .ZN(n10504) );
  NAND2_X1 U10823 ( .A1(n10504), .A2(n10248), .ZN(n8306) );
  INV_X1 U10824 ( .A(n8303), .ZN(n8300) );
  NAND2_X1 U10825 ( .A1(n8300), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8301) );
  MUX2_X1 U10826 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8301), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n8304) );
  NAND2_X1 U10827 ( .A1(n8303), .A2(n8302), .ZN(n8319) );
  NAND2_X1 U10828 ( .A1(n8304), .A2(n8319), .ZN(n11268) );
  AOI22_X1 U10829 ( .A1(n8403), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n10576), 
        .B2(n11375), .ZN(n8305) );
  NAND2_X1 U10830 ( .A1(n8531), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8314) );
  NAND2_X1 U10831 ( .A1(n8532), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8313) );
  NAND2_X1 U10832 ( .A1(n8308), .A2(n8307), .ZN(n8309) );
  NAND2_X1 U10833 ( .A1(n8324), .A2(n8309), .ZN(n12146) );
  OR2_X1 U10834 ( .A1(n8530), .A2(n12146), .ZN(n8312) );
  INV_X1 U10835 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8310) );
  OR2_X1 U10836 ( .A1(n8535), .A2(n8310), .ZN(n8311) );
  NAND4_X1 U10837 ( .A1(n8314), .A2(n8313), .A3(n8312), .A4(n8311), .ZN(n13819) );
  AND2_X1 U10838 ( .A1(n14296), .A2(n13819), .ZN(n8315) );
  XNOR2_X1 U10839 ( .A(n8317), .B(SI_14_), .ZN(n8318) );
  NAND2_X1 U10840 ( .A1(n10554), .A2(n10248), .ZN(n8322) );
  NAND2_X1 U10841 ( .A1(n8319), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8320) );
  XNOR2_X1 U10842 ( .A(n8320), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11378) );
  AOI22_X1 U10843 ( .A1(n8403), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n10576), 
        .B2(n11378), .ZN(n8321) );
  NAND2_X1 U10844 ( .A1(n8531), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8329) );
  NAND2_X1 U10845 ( .A1(n8532), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8328) );
  INV_X1 U10846 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8323) );
  NAND2_X1 U10847 ( .A1(n8324), .A2(n8323), .ZN(n8325) );
  NAND2_X1 U10848 ( .A1(n8356), .A2(n8325), .ZN(n13333) );
  OR2_X1 U10849 ( .A1(n8530), .A2(n13333), .ZN(n8327) );
  INV_X1 U10850 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14348) );
  OR2_X1 U10851 ( .A1(n8535), .A2(n14348), .ZN(n8326) );
  NAND4_X1 U10852 ( .A1(n8329), .A2(n8328), .A3(n8327), .A4(n8326), .ZN(n14191) );
  NAND2_X1 U10853 ( .A1(n14184), .A2(n14191), .ZN(n8330) );
  XNOR2_X1 U10854 ( .A(n8331), .B(n7942), .ZN(n10712) );
  NAND2_X1 U10855 ( .A1(n10712), .A2(n10248), .ZN(n8336) );
  INV_X1 U10856 ( .A(n8626), .ZN(n8333) );
  NAND2_X1 U10857 ( .A1(n8333), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8334) );
  XNOR2_X1 U10858 ( .A(n8334), .B(P2_IR_REG_16__SCAN_IN), .ZN(n13885) );
  AOI22_X1 U10859 ( .A1(n8403), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n10576), 
        .B2(n13885), .ZN(n8335) );
  INV_X1 U10860 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8343) );
  INV_X1 U10861 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8337) );
  NAND2_X1 U10862 ( .A1(n8358), .A2(n8337), .ZN(n8338) );
  NAND2_X1 U10863 ( .A1(n8375), .A2(n8338), .ZN(n14143) );
  OR2_X1 U10864 ( .A1(n14143), .A2(n8530), .ZN(n8342) );
  NAND2_X1 U10865 ( .A1(n8531), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8340) );
  NAND2_X1 U10866 ( .A1(n8532), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8339) );
  AND2_X1 U10867 ( .A1(n8340), .A2(n8339), .ZN(n8341) );
  OAI211_X1 U10868 ( .C1(n8535), .C2(n8343), .A(n8342), .B(n8341), .ZN(n13817)
         );
  INV_X1 U10869 ( .A(n13817), .ZN(n14161) );
  NOR2_X1 U10870 ( .A1(n14341), .A2(n14161), .ZN(n8591) );
  INV_X1 U10871 ( .A(n8591), .ZN(n14124) );
  NAND2_X1 U10872 ( .A1(n14341), .A2(n14161), .ZN(n8586) );
  NAND2_X1 U10873 ( .A1(n14124), .A2(n8586), .ZN(n14152) );
  XNOR2_X1 U10874 ( .A(n8345), .B(n8344), .ZN(n10668) );
  NAND2_X1 U10875 ( .A1(n10668), .A2(n10248), .ZN(n8354) );
  INV_X1 U10876 ( .A(n8346), .ZN(n8350) );
  INV_X1 U10877 ( .A(n8347), .ZN(n8349) );
  NAND3_X1 U10878 ( .A1(n8350), .A2(n8349), .A3(n8348), .ZN(n8351) );
  NAND2_X1 U10879 ( .A1(n8351), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8352) );
  XNOR2_X1 U10880 ( .A(n8352), .B(P2_IR_REG_15__SCAN_IN), .ZN(n13884) );
  AOI22_X1 U10881 ( .A1(n8403), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n10576), 
        .B2(n13884), .ZN(n8353) );
  NAND2_X1 U10882 ( .A1(n8356), .A2(n8355), .ZN(n8357) );
  NAND2_X1 U10883 ( .A1(n8358), .A2(n8357), .ZN(n13490) );
  NAND2_X1 U10884 ( .A1(n8531), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8359) );
  OAI21_X1 U10885 ( .B1(n13490), .B2(n8530), .A(n8359), .ZN(n8362) );
  INV_X1 U10886 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n14344) );
  NAND2_X1 U10887 ( .A1(n8532), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8360) );
  OAI21_X1 U10888 ( .B1(n8535), .B2(n14344), .A(n8360), .ZN(n8361) );
  OR2_X1 U10889 ( .A1(n14166), .A2(n13818), .ZN(n14151) );
  AND2_X1 U10890 ( .A1(n14152), .A2(n14151), .ZN(n8366) );
  NAND3_X1 U10891 ( .A1(n14152), .A2(n14166), .A3(n13818), .ZN(n8364) );
  NAND2_X1 U10892 ( .A1(n14341), .A2(n13817), .ZN(n8363) );
  NAND2_X1 U10893 ( .A1(n8364), .A2(n8363), .ZN(n8365) );
  XNOR2_X1 U10894 ( .A(n8368), .B(SI_17_), .ZN(n8369) );
  NAND2_X1 U10895 ( .A1(n10871), .A2(n10248), .ZN(n8373) );
  XNOR2_X1 U10896 ( .A(n8371), .B(P2_IR_REG_17__SCAN_IN), .ZN(n13915) );
  AOI22_X1 U10897 ( .A1(n8403), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n10576), 
        .B2(n13915), .ZN(n8372) );
  NAND2_X1 U10898 ( .A1(n8375), .A2(n8374), .ZN(n8376) );
  NAND2_X1 U10899 ( .A1(n8388), .A2(n8376), .ZN(n13428) );
  AOI22_X1 U10900 ( .A1(n8111), .A2(P2_REG0_REG_17__SCAN_IN), .B1(n8532), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n8378) );
  NAND2_X1 U10901 ( .A1(n8531), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8377) );
  NAND2_X1 U10902 ( .A1(n14127), .A2(n13816), .ZN(n13758) );
  OR2_X1 U10903 ( .A1(n14127), .A2(n13816), .ZN(n13759) );
  INV_X1 U10904 ( .A(SI_18_), .ZN(n10638) );
  NAND2_X1 U10905 ( .A1(n8380), .A2(n10638), .ZN(n8379) );
  OAI21_X1 U10906 ( .B1(n8380), .B2(n10638), .A(n8379), .ZN(n8382) );
  XNOR2_X1 U10907 ( .A(n8382), .B(n8381), .ZN(n11060) );
  NAND2_X1 U10908 ( .A1(n11060), .A2(n10248), .ZN(n8386) );
  INV_X1 U10909 ( .A(n8401), .ZN(n8383) );
  NAND2_X1 U10910 ( .A1(n8383), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8384) );
  XNOR2_X1 U10911 ( .A(n8384), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13927) );
  AOI22_X1 U10912 ( .A1(n8403), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n10576), 
        .B2(n13927), .ZN(n8385) );
  INV_X1 U10913 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8387) );
  NAND2_X1 U10914 ( .A1(n8388), .A2(n8387), .ZN(n8389) );
  NAND2_X1 U10915 ( .A1(n8407), .A2(n8389), .ZN(n14115) );
  OR2_X1 U10916 ( .A1(n14115), .A2(n8530), .ZN(n8395) );
  INV_X1 U10917 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8392) );
  NAND2_X1 U10918 ( .A1(n8532), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8391) );
  NAND2_X1 U10919 ( .A1(n8531), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8390) );
  OAI211_X1 U10920 ( .C1(n8392), .C2(n8535), .A(n8391), .B(n8390), .ZN(n8393)
         );
  INV_X1 U10921 ( .A(n8393), .ZN(n8394) );
  NAND2_X1 U10922 ( .A1(n8395), .A2(n8394), .ZN(n13815) );
  INV_X1 U10923 ( .A(n13815), .ZN(n13651) );
  XNOR2_X1 U10924 ( .A(n13648), .B(n13651), .ZN(n14111) );
  OR2_X1 U10925 ( .A1(n13648), .A2(n13815), .ZN(n8396) );
  XNOR2_X1 U10926 ( .A(n8399), .B(n8398), .ZN(n11135) );
  NAND2_X1 U10927 ( .A1(n11135), .A2(n10248), .ZN(n8405) );
  INV_X1 U10928 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8400) );
  NAND2_X1 U10929 ( .A1(n8556), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8402) );
  INV_X1 U10930 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8547) );
  XNOR2_X1 U10931 ( .A(n8402), .B(n8547), .ZN(n13791) );
  AOI22_X1 U10932 ( .A1(n8403), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n10576), 
        .B2(n13936), .ZN(n8404) );
  INV_X1 U10933 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8406) );
  NAND2_X1 U10934 ( .A1(n8407), .A2(n8406), .ZN(n8408) );
  NAND2_X1 U10935 ( .A1(n8421), .A2(n8408), .ZN(n14102) );
  OR2_X1 U10936 ( .A1(n14102), .A2(n8530), .ZN(n8413) );
  INV_X1 U10937 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13929) );
  NAND2_X1 U10938 ( .A1(n8111), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8410) );
  NAND2_X1 U10939 ( .A1(n8532), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8409) );
  OAI211_X1 U10940 ( .C1(n8131), .C2(n13929), .A(n8410), .B(n8409), .ZN(n8411)
         );
  INV_X1 U10941 ( .A(n8411), .ZN(n8412) );
  NAND2_X1 U10942 ( .A1(n8413), .A2(n8412), .ZN(n13814) );
  NAND2_X1 U10943 ( .A1(n14105), .A2(n13814), .ZN(n8414) );
  NAND2_X1 U10944 ( .A1(n8417), .A2(n7311), .ZN(n8418) );
  INV_X1 U10945 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n12446) );
  OR2_X1 U10946 ( .A1(n7177), .A2(n12446), .ZN(n8419) );
  NAND2_X1 U10947 ( .A1(n8421), .A2(n13446), .ZN(n8422) );
  NAND2_X1 U10948 ( .A1(n8452), .A2(n8422), .ZN(n14088) );
  OR2_X1 U10949 ( .A1(n14088), .A2(n8530), .ZN(n8427) );
  INV_X1 U10950 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n14332) );
  NAND2_X1 U10951 ( .A1(n8531), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8424) );
  NAND2_X1 U10952 ( .A1(n8532), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8423) );
  OAI211_X1 U10953 ( .C1(n14332), .C2(n8535), .A(n8424), .B(n8423), .ZN(n8425)
         );
  INV_X1 U10954 ( .A(n8425), .ZN(n8426) );
  NAND2_X1 U10955 ( .A1(n8427), .A2(n8426), .ZN(n13813) );
  INV_X1 U10956 ( .A(n13813), .ZN(n13659) );
  INV_X1 U10957 ( .A(n14081), .ZN(n14077) );
  NAND2_X1 U10958 ( .A1(n14335), .A2(n13659), .ZN(n8428) );
  NAND2_X1 U10959 ( .A1(n8430), .A2(n8429), .ZN(n8434) );
  NAND2_X1 U10960 ( .A1(n8432), .A2(n8431), .ZN(n8433) );
  NAND2_X1 U10961 ( .A1(n11707), .A2(n10248), .ZN(n8436) );
  OR2_X1 U10962 ( .A1(n7177), .A2(n15733), .ZN(n8435) );
  NAND2_X2 U10963 ( .A1(n8436), .A2(n8435), .ZN(n14073) );
  XNOR2_X1 U10964 ( .A(n8452), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n14070) );
  NAND2_X1 U10965 ( .A1(n14070), .A2(n8112), .ZN(n8442) );
  INV_X1 U10966 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8439) );
  NAND2_X1 U10967 ( .A1(n8532), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8438) );
  NAND2_X1 U10968 ( .A1(n8531), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8437) );
  OAI211_X1 U10969 ( .C1(n8439), .C2(n8535), .A(n8438), .B(n8437), .ZN(n8440)
         );
  INV_X1 U10970 ( .A(n8440), .ZN(n8441) );
  NAND2_X1 U10971 ( .A1(n8442), .A2(n8441), .ZN(n13812) );
  NOR2_X1 U10972 ( .A1(n14073), .A2(n13812), .ZN(n13757) );
  NAND2_X1 U10973 ( .A1(n14073), .A2(n13812), .ZN(n13755) );
  NAND2_X1 U10974 ( .A1(n9734), .A2(n8444), .ZN(n8461) );
  INV_X1 U10975 ( .A(n9734), .ZN(n8446) );
  INV_X1 U10976 ( .A(n8444), .ZN(n8445) );
  NAND2_X1 U10977 ( .A1(n8446), .A2(n8445), .ZN(n8447) );
  NAND2_X1 U10978 ( .A1(n11907), .A2(n10248), .ZN(n8449) );
  INV_X1 U10979 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11909) );
  OR2_X1 U10980 ( .A1(n7177), .A2(n11909), .ZN(n8448) );
  INV_X1 U10981 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8451) );
  INV_X1 U10982 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8450) );
  OAI21_X1 U10983 ( .B1(n8452), .B2(n8451), .A(n8450), .ZN(n8453) );
  AND2_X1 U10984 ( .A1(n8468), .A2(n8453), .ZN(n14060) );
  NAND2_X1 U10985 ( .A1(n14060), .A2(n8112), .ZN(n8458) );
  INV_X1 U10986 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n14325) );
  NAND2_X1 U10987 ( .A1(n8531), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8455) );
  NAND2_X1 U10988 ( .A1(n8532), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8454) );
  OAI211_X1 U10989 ( .C1(n14325), .C2(n8535), .A(n8455), .B(n8454), .ZN(n8456)
         );
  INV_X1 U10990 ( .A(n8456), .ZN(n8457) );
  NAND2_X1 U10991 ( .A1(n8458), .A2(n8457), .ZN(n14039) );
  XNOR2_X1 U10992 ( .A(n14059), .B(n14039), .ZN(n14055) );
  INV_X1 U10993 ( .A(n14055), .ZN(n14052) );
  NAND2_X1 U10994 ( .A1(n14059), .A2(n14039), .ZN(n8459) );
  NAND2_X1 U10995 ( .A1(n8461), .A2(n8460), .ZN(n8465) );
  NAND2_X1 U10996 ( .A1(n8463), .A2(n8462), .ZN(n8464) );
  NAND2_X1 U10997 ( .A1(n11860), .A2(n10248), .ZN(n8467) );
  OR2_X1 U10998 ( .A1(n7177), .A2(n11863), .ZN(n8466) );
  INV_X1 U10999 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n15749) );
  NAND2_X1 U11000 ( .A1(n8468), .A2(n15749), .ZN(n8469) );
  NAND2_X1 U11001 ( .A1(n8483), .A2(n8469), .ZN(n14043) );
  OR2_X1 U11002 ( .A1(n14043), .A2(n8530), .ZN(n8475) );
  INV_X1 U11003 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8472) );
  NAND2_X1 U11004 ( .A1(n8531), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8471) );
  NAND2_X1 U11005 ( .A1(n8532), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8470) );
  OAI211_X1 U11006 ( .C1(n8472), .C2(n8535), .A(n8471), .B(n8470), .ZN(n8473)
         );
  INV_X1 U11007 ( .A(n8473), .ZN(n8474) );
  OR2_X1 U11008 ( .A1(n14047), .A2(n14024), .ZN(n8476) );
  INV_X1 U11009 ( .A(n8477), .ZN(n8478) );
  NAND2_X1 U11010 ( .A1(n7574), .A2(n8478), .ZN(n8479) );
  NAND2_X1 U11011 ( .A1(n12114), .A2(n10248), .ZN(n8482) );
  INV_X1 U11012 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12127) );
  OR2_X1 U11013 ( .A1(n7177), .A2(n12127), .ZN(n8481) );
  INV_X1 U11014 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13434) );
  NAND2_X1 U11015 ( .A1(n8483), .A2(n13434), .ZN(n8484) );
  NAND2_X1 U11016 ( .A1(n8485), .A2(n8484), .ZN(n14028) );
  INV_X1 U11017 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8488) );
  NAND2_X1 U11018 ( .A1(n8531), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8487) );
  NAND2_X1 U11019 ( .A1(n8532), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8486) );
  OAI211_X1 U11020 ( .C1(n8488), .C2(n8535), .A(n8487), .B(n8486), .ZN(n8489)
         );
  INV_X1 U11021 ( .A(n8489), .ZN(n8490) );
  OR2_X1 U11022 ( .A1(n14217), .A2(n13400), .ZN(n8601) );
  NAND2_X1 U11023 ( .A1(n14217), .A2(n13400), .ZN(n13999) );
  MUX2_X1 U11024 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n10338), .Z(n8509) );
  XNOR2_X1 U11025 ( .A(n8509), .B(SI_27_), .ZN(n8496) );
  INV_X1 U11026 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14364) );
  OR2_X1 U11027 ( .A1(n7177), .A2(n14364), .ZN(n8497) );
  INV_X1 U11028 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8499) );
  NAND2_X1 U11029 ( .A1(n8500), .A2(n8499), .ZN(n8501) );
  NAND2_X1 U11030 ( .A1(n13973), .A2(n8112), .ZN(n8506) );
  INV_X1 U11031 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n14316) );
  NAND2_X1 U11032 ( .A1(n8531), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8503) );
  NAND2_X1 U11033 ( .A1(n8532), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8502) );
  OAI211_X1 U11034 ( .C1(n14316), .C2(n8535), .A(n8503), .B(n8502), .ZN(n8504)
         );
  INV_X1 U11035 ( .A(n8504), .ZN(n8505) );
  INV_X1 U11036 ( .A(n8509), .ZN(n8507) );
  INV_X1 U11037 ( .A(SI_27_), .ZN(n13249) );
  INV_X1 U11038 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n15165) );
  INV_X1 U11039 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n12458) );
  MUX2_X1 U11040 ( .A(n15165), .B(n12458), .S(n10338), .Z(n8510) );
  INV_X1 U11041 ( .A(SI_28_), .ZN(n13242) );
  NAND2_X1 U11042 ( .A1(n8510), .A2(n13242), .ZN(n8513) );
  INV_X1 U11043 ( .A(n8510), .ZN(n8511) );
  NAND2_X1 U11044 ( .A1(n8511), .A2(SI_28_), .ZN(n8512) );
  NAND2_X1 U11045 ( .A1(n8513), .A2(n8512), .ZN(n8523) );
  INV_X1 U11046 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15163) );
  INV_X1 U11047 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14362) );
  MUX2_X1 U11048 ( .A(n15163), .B(n14362), .S(n6442), .Z(n9857) );
  XNOR2_X1 U11049 ( .A(n9857), .B(SI_29_), .ZN(n9851) );
  NAND2_X1 U11050 ( .A1(n14361), .A2(n10248), .ZN(n8515) );
  OR2_X1 U11051 ( .A1(n7177), .A2(n14362), .ZN(n8514) );
  INV_X1 U11052 ( .A(n8528), .ZN(n8516) );
  NAND2_X1 U11053 ( .A1(n8516), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n13958) );
  OR2_X1 U11054 ( .A1(n13958), .A2(n8530), .ZN(n8522) );
  INV_X1 U11055 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8519) );
  NAND2_X1 U11056 ( .A1(n8531), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8518) );
  NAND2_X1 U11057 ( .A1(n8532), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8517) );
  OAI211_X1 U11058 ( .C1(n8519), .C2(n8535), .A(n8518), .B(n8517), .ZN(n8520)
         );
  INV_X1 U11059 ( .A(n8520), .ZN(n8521) );
  NAND2_X1 U11060 ( .A1(n12457), .A2(n10248), .ZN(n8526) );
  OR2_X1 U11061 ( .A1(n7177), .A2(n12458), .ZN(n8525) );
  INV_X1 U11062 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8527) );
  NAND2_X1 U11063 ( .A1(n8528), .A2(n8527), .ZN(n8529) );
  NAND2_X1 U11064 ( .A1(n13958), .A2(n8529), .ZN(n13382) );
  INV_X1 U11065 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n10278) );
  NAND2_X1 U11066 ( .A1(n8531), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8534) );
  NAND2_X1 U11067 ( .A1(n8532), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8533) );
  OAI211_X1 U11068 ( .C1(n10278), .C2(n8535), .A(n8534), .B(n8533), .ZN(n8536)
         );
  INV_X1 U11069 ( .A(n8536), .ZN(n8537) );
  NAND2_X2 U11070 ( .A1(n8538), .A2(n8537), .ZN(n13810) );
  NAND2_X1 U11071 ( .A1(n13720), .A2(n13810), .ZN(n13950) );
  INV_X1 U11072 ( .A(n8539), .ZN(n8540) );
  INV_X1 U11073 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8543) );
  NAND2_X1 U11074 ( .A1(n8544), .A2(n8543), .ZN(n8545) );
  INV_X1 U11075 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8541) );
  XNOR2_X2 U11076 ( .A(n8542), .B(n8541), .ZN(n8559) );
  INV_X1 U11077 ( .A(n8559), .ZN(n8614) );
  OR2_X1 U11078 ( .A1(n8544), .A2(n8543), .ZN(n8546) );
  INV_X1 U11079 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8548) );
  NAND2_X1 U11080 ( .A1(n8548), .A2(n8547), .ZN(n8555) );
  INV_X1 U11081 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8550) );
  NAND3_X1 U11082 ( .A1(n8549), .A2(P2_IR_REG_20__SCAN_IN), .A3(n8550), .ZN(
        n8552) );
  XNOR2_X1 U11083 ( .A(P2_IR_REG_31__SCAN_IN), .B(P2_IR_REG_20__SCAN_IN), .ZN(
        n8551) );
  OAI21_X2 U11084 ( .B1(n8556), .B2(n8555), .A(n8554), .ZN(n8558) );
  NAND2_X1 U11085 ( .A1(n8557), .A2(n11137), .ZN(n10737) );
  NOR2_X1 U11086 ( .A1(n11137), .A2(n13761), .ZN(n8560) );
  NAND2_X1 U11087 ( .A1(n8560), .A2(n8559), .ZN(n15528) );
  NAND2_X1 U11088 ( .A1(n15501), .A2(n15528), .ZN(n14271) );
  NAND2_X1 U11089 ( .A1(n13720), .A2(n13719), .ZN(n8561) );
  NAND3_X1 U11090 ( .A1(n13789), .A2(n10274), .A3(n13950), .ZN(n8562) );
  NAND2_X1 U11091 ( .A1(n10275), .A2(n13786), .ZN(n13951) );
  NAND2_X1 U11092 ( .A1(n8563), .A2(n11297), .ZN(n11177) );
  NAND2_X1 U11093 ( .A1(n10882), .A2(n15524), .ZN(n11178) );
  NAND2_X1 U11094 ( .A1(n13828), .A2(n13535), .ZN(n8565) );
  NAND2_X1 U11095 ( .A1(n15544), .A2(n13762), .ZN(n15551) );
  NAND2_X1 U11096 ( .A1(n15494), .A2(n15826), .ZN(n8567) );
  NAND2_X1 U11097 ( .A1(n8568), .A2(n8567), .ZN(n11353) );
  NAND2_X1 U11098 ( .A1(n11353), .A2(n13765), .ZN(n8570) );
  NAND2_X1 U11099 ( .A1(n11582), .A2(n14307), .ZN(n8569) );
  XNOR2_X1 U11100 ( .A(n13823), .B(n13567), .ZN(n13766) );
  NAND2_X1 U11101 ( .A1(n7921), .A2(n13823), .ZN(n8572) );
  NAND2_X1 U11102 ( .A1(n11867), .A2(n14301), .ZN(n8573) );
  INV_X1 U11103 ( .A(n13821), .ZN(n8574) );
  NOR2_X1 U11104 ( .A1(n13581), .A2(n8574), .ZN(n8576) );
  NAND2_X1 U11105 ( .A1(n13581), .A2(n8574), .ZN(n8575) );
  INV_X1 U11106 ( .A(n13820), .ZN(n11866) );
  AND2_X1 U11107 ( .A1(n13590), .A2(n12148), .ZN(n8577) );
  INV_X1 U11108 ( .A(n8577), .ZN(n8578) );
  OR2_X1 U11109 ( .A1(n13590), .A2(n12148), .ZN(n8580) );
  INV_X1 U11110 ( .A(n13819), .ZN(n13775) );
  INV_X1 U11111 ( .A(n14296), .ZN(n14197) );
  AND2_X1 U11112 ( .A1(n14184), .A2(n14160), .ZN(n8582) );
  OR2_X1 U11113 ( .A1(n14184), .A2(n14160), .ZN(n8583) );
  INV_X1 U11114 ( .A(n13818), .ZN(n8585) );
  INV_X1 U11115 ( .A(n13816), .ZN(n8584) );
  NAND2_X1 U11116 ( .A1(n14127), .A2(n8584), .ZN(n8590) );
  INV_X1 U11117 ( .A(n8590), .ZN(n8588) );
  NAND2_X1 U11118 ( .A1(n14166), .A2(n8585), .ZN(n14122) );
  NAND2_X1 U11119 ( .A1(n14123), .A2(n8589), .ZN(n8593) );
  AOI22_X1 U11120 ( .A1(n8591), .A2(n8590), .B1(n7923), .B2(n13816), .ZN(n8592) );
  NAND2_X1 U11121 ( .A1(n8593), .A2(n8592), .ZN(n14112) );
  NOR2_X1 U11122 ( .A1(n13648), .A2(n13651), .ZN(n8594) );
  INV_X1 U11123 ( .A(n13814), .ZN(n13653) );
  AND2_X1 U11124 ( .A1(n14105), .A2(n13653), .ZN(n8596) );
  OR2_X1 U11125 ( .A1(n14105), .A2(n13653), .ZN(n8595) );
  INV_X1 U11126 ( .A(n13812), .ZN(n13501) );
  OR2_X1 U11127 ( .A1(n14073), .A2(n13501), .ZN(n8597) );
  INV_X1 U11128 ( .A(n14059), .ZN(n14327) );
  NAND2_X1 U11129 ( .A1(n14327), .A2(n14039), .ZN(n8598) );
  NAND2_X1 U11130 ( .A1(n14047), .A2(n13754), .ZN(n8599) );
  NAND2_X1 U11131 ( .A1(n14008), .A2(n13986), .ZN(n8605) );
  OR2_X1 U11132 ( .A1(n14047), .A2(n13754), .ZN(n13997) );
  NAND2_X1 U11133 ( .A1(n8601), .A2(n13997), .ZN(n8602) );
  NOR2_X1 U11134 ( .A1(n14000), .A2(n8602), .ZN(n8604) );
  NOR2_X1 U11135 ( .A1(n14000), .A2(n13999), .ZN(n8603) );
  OAI21_X2 U11136 ( .B1(n14210), .B2(n8606), .A(n8607), .ZN(n13983) );
  INV_X1 U11137 ( .A(n8607), .ZN(n8608) );
  NOR2_X2 U11138 ( .A1(n10282), .A2(n13785), .ZN(n10265) );
  AND2_X1 U11139 ( .A1(n13974), .A2(n13985), .ZN(n10264) );
  OR2_X1 U11140 ( .A1(n8559), .A2(n13791), .ZN(n13748) );
  NAND2_X1 U11141 ( .A1(n13761), .A2(n8610), .ZN(n8611) );
  NAND4_X1 U11142 ( .A1(n13952), .A2(n13966), .A3(n13810), .A4(n15556), .ZN(
        n8621) );
  NAND2_X1 U11143 ( .A1(n8614), .A2(n8610), .ZN(n10575) );
  OR2_X1 U11144 ( .A1(n10575), .A2(n8615), .ZN(n15495) );
  INV_X1 U11145 ( .A(n8615), .ZN(n10603) );
  INV_X1 U11146 ( .A(P2_B_REG_SCAN_IN), .ZN(n13794) );
  NOR2_X1 U11147 ( .A1(n14366), .A2(n13794), .ZN(n8616) );
  NOR2_X1 U11148 ( .A1(n15493), .A2(n8616), .ZN(n10257) );
  INV_X1 U11149 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n14206) );
  NAND2_X1 U11150 ( .A1(n8111), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8619) );
  INV_X1 U11151 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8617) );
  OR2_X1 U11152 ( .A1(n10254), .A2(n8617), .ZN(n8618) );
  OAI211_X1 U11153 ( .C1(n8131), .C2(n14206), .A(n8619), .B(n8618), .ZN(n13808) );
  AOI22_X1 U11154 ( .A1(n13810), .A2(n14188), .B1(n10257), .B2(n13808), .ZN(
        n8620) );
  NAND2_X1 U11155 ( .A1(n11217), .A2(n13535), .ZN(n15481) );
  NOR2_X4 U11156 ( .A1(n15563), .A2(n14307), .ZN(n11415) );
  INV_X1 U11157 ( .A(n13585), .ZN(n11809) );
  NAND2_X1 U11158 ( .A1(n14099), .A2(n14256), .ZN(n14100) );
  AOI21_X1 U11159 ( .B1(n10271), .B2(n13955), .A(n15561), .ZN(n8622) );
  INV_X1 U11160 ( .A(n15518), .ZN(n11023) );
  NAND2_X1 U11161 ( .A1(n11137), .A2(n8558), .ZN(n13743) );
  NAND2_X1 U11162 ( .A1(n8626), .A2(n8625), .ZN(n8658) );
  INV_X1 U11163 ( .A(n8632), .ZN(n8628) );
  INV_X1 U11164 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8627) );
  NAND2_X1 U11165 ( .A1(n8628), .A2(n8627), .ZN(n8634) );
  MUX2_X1 U11166 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8629), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8631) );
  AND2_X1 U11167 ( .A1(n8631), .A2(n8630), .ZN(n14370) );
  MUX2_X1 U11168 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8633), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8635) );
  NAND2_X1 U11169 ( .A1(n8635), .A2(n8634), .ZN(n12128) );
  XOR2_X1 U11170 ( .A(P2_B_REG_SCAN_IN), .B(n12128), .Z(n8636) );
  NAND2_X1 U11171 ( .A1(n8630), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8637) );
  MUX2_X1 U11172 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8637), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8639) );
  NAND2_X1 U11173 ( .A1(n8639), .A2(n8638), .ZN(n14369) );
  INV_X1 U11174 ( .A(n14369), .ZN(n8654) );
  INV_X1 U11175 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15512) );
  NAND2_X1 U11176 ( .A1(n15509), .A2(n15512), .ZN(n8642) );
  NAND2_X1 U11177 ( .A1(n12128), .A2(n14369), .ZN(n8641) );
  NAND2_X1 U11178 ( .A1(n8642), .A2(n8641), .ZN(n15513) );
  INV_X1 U11179 ( .A(n15513), .ZN(n8653) );
  NOR4_X1 U11180 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n8646) );
  NOR4_X1 U11181 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n8645) );
  NOR4_X1 U11182 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8644) );
  NOR4_X1 U11183 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n8643) );
  NAND4_X1 U11184 ( .A1(n8646), .A2(n8645), .A3(n8644), .A4(n8643), .ZN(n8652)
         );
  NOR2_X1 U11185 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .ZN(
        n8650) );
  NOR4_X1 U11186 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n8649) );
  NOR4_X1 U11187 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n8648) );
  NOR4_X1 U11188 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n8647) );
  NAND4_X1 U11189 ( .A1(n8650), .A2(n8649), .A3(n8648), .A4(n8647), .ZN(n8651)
         );
  OAI21_X1 U11190 ( .B1(n8652), .B2(n8651), .A(n15509), .ZN(n11018) );
  INV_X1 U11191 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15515) );
  NAND2_X1 U11192 ( .A1(n15509), .A2(n15515), .ZN(n8656) );
  OR2_X1 U11193 ( .A1(n14370), .A2(n8654), .ZN(n8655) );
  NAND2_X1 U11194 ( .A1(n8656), .A2(n8655), .ZN(n15516) );
  NAND2_X1 U11195 ( .A1(n15516), .A2(n10742), .ZN(n8664) );
  NOR2_X1 U11196 ( .A1(n12128), .A2(n14369), .ZN(n8657) );
  NAND2_X1 U11197 ( .A1(n14370), .A2(n8657), .ZN(n10578) );
  INV_X1 U11198 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8659) );
  XNOR2_X1 U11199 ( .A(n8660), .B(n8659), .ZN(n11861) );
  NAND2_X1 U11200 ( .A1(n13743), .A2(n8610), .ZN(n13711) );
  OR2_X1 U11201 ( .A1(n13711), .A2(n8559), .ZN(n10747) );
  NAND2_X1 U11202 ( .A1(n15517), .A2(n10747), .ZN(n13798) );
  NOR2_X1 U11203 ( .A1(n8664), .A2(n13798), .ZN(n8661) );
  NAND2_X1 U11204 ( .A1(n15578), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8662) );
  NAND2_X1 U11205 ( .A1(n8663), .A2(n8662), .ZN(P2_U3528) );
  INV_X1 U11206 ( .A(n13798), .ZN(n11017) );
  AND3_X1 U11207 ( .A1(n11018), .A2(n11017), .A3(n15513), .ZN(n8666) );
  INV_X1 U11208 ( .A(n8664), .ZN(n8665) );
  NAND2_X1 U11209 ( .A1(n15569), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8668) );
  INV_X1 U11210 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8675) );
  XNOR2_X2 U11211 ( .A(n8676), .B(n8675), .ZN(n10849) );
  NAND4_X1 U11212 ( .A1(n8679), .A2(n8687), .A3(n8678), .A4(n8677), .ZN(n8681)
         );
  OAI21_X1 U11213 ( .B1(n9083), .B2(n8681), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n8680) );
  MUX2_X1 U11214 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8680), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n8684) );
  INV_X1 U11215 ( .A(n8681), .ZN(n8683) );
  NAND2_X1 U11216 ( .A1(n8685), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8686) );
  NAND2_X1 U11217 ( .A1(n9070), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8688) );
  NAND2_X1 U11218 ( .A1(n12357), .A2(n12368), .ZN(n8728) );
  OAI21_X1 U11219 ( .B1(n15651), .B2(n9286), .A(n8728), .ZN(n8689) );
  NAND2_X1 U11220 ( .A1(n12316), .A2(n12357), .ZN(n9288) );
  NAND2_X1 U11221 ( .A1(n8689), .A2(n9288), .ZN(n8690) );
  NAND2_X1 U11222 ( .A1(n8690), .A2(n12267), .ZN(n8709) );
  NAND2_X1 U11223 ( .A1(n8698), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8692) );
  MUX2_X1 U11224 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8692), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8696) );
  NAND2_X1 U11225 ( .A1(n8696), .A2(n8701), .ZN(n13258) );
  NAND2_X1 U11226 ( .A1(n8725), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8697) );
  MUX2_X1 U11227 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8697), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8699) );
  XNOR2_X1 U11228 ( .A(n11818), .B(P3_B_REG_SCAN_IN), .ZN(n8705) );
  NAND2_X1 U11229 ( .A1(n8701), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8700) );
  MUX2_X1 U11230 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8700), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n8704) );
  NAND2_X1 U11231 ( .A1(n8704), .A2(n8805), .ZN(n13253) );
  INV_X1 U11232 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8706) );
  NAND2_X1 U11233 ( .A1(n12155), .A2(n8706), .ZN(n8708) );
  NAND2_X1 U11234 ( .A1(n13258), .A2(n13253), .ZN(n8707) );
  NAND2_X1 U11235 ( .A1(n8709), .A2(n11391), .ZN(n8730) );
  NAND2_X1 U11236 ( .A1(n11818), .A2(n13253), .ZN(n8710) );
  OR2_X1 U11237 ( .A1(n11391), .A2(n10848), .ZN(n9285) );
  NAND2_X1 U11238 ( .A1(n10848), .A2(n11391), .ZN(n9291) );
  NOR4_X1 U11239 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_27__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_13__SCAN_IN), .ZN(n15686) );
  NOR2_X1 U11240 ( .A1(P3_D_REG_8__SCAN_IN), .A2(P3_D_REG_7__SCAN_IN), .ZN(
        n8714) );
  NOR4_X1 U11241 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_19__SCAN_IN), .ZN(n8713) );
  NOR4_X1 U11242 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_17__SCAN_IN), .ZN(n8712) );
  NAND4_X1 U11243 ( .A1(n15686), .A2(n8714), .A3(n8713), .A4(n8712), .ZN(n8720) );
  NOR4_X1 U11244 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n8718) );
  NOR4_X1 U11245 ( .A1(P3_D_REG_18__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_21__SCAN_IN), .ZN(n8717) );
  NOR4_X1 U11246 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_2__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_4__SCAN_IN), .ZN(n8716) );
  NOR4_X1 U11247 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_3__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n8715) );
  NAND4_X1 U11248 ( .A1(n8718), .A2(n8717), .A3(n8716), .A4(n8715), .ZN(n8719)
         );
  OAI21_X1 U11249 ( .B1(n8720), .B2(n8719), .A(n12155), .ZN(n9284) );
  INV_X1 U11250 ( .A(n13258), .ZN(n8722) );
  NOR2_X1 U11251 ( .A1(n11818), .A2(n13253), .ZN(n8721) );
  NAND2_X1 U11252 ( .A1(n8722), .A2(n8721), .ZN(n10829) );
  NAND2_X1 U11253 ( .A1(n8723), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8724) );
  MUX2_X1 U11254 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8724), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n8726) );
  NAND2_X1 U11255 ( .A1(n8726), .A2(n8725), .ZN(n10828) );
  AND2_X1 U11256 ( .A1(n9284), .A2(n10865), .ZN(n8727) );
  INV_X1 U11257 ( .A(n9288), .ZN(n8814) );
  OR2_X1 U11258 ( .A1(n12267), .A2(n8814), .ZN(n10830) );
  NAND2_X1 U11259 ( .A1(n12267), .A2(n8816), .ZN(n11387) );
  NAND2_X1 U11260 ( .A1(n10830), .A2(n11387), .ZN(n11388) );
  INV_X1 U11261 ( .A(n11391), .ZN(n13225) );
  NAND2_X1 U11262 ( .A1(n11388), .A2(n13225), .ZN(n8729) );
  INV_X1 U11263 ( .A(n13115), .ZN(n9283) );
  INV_X1 U11264 ( .A(n8836), .ZN(n8732) );
  NAND2_X1 U11265 ( .A1(n10314), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8733) );
  NAND2_X1 U11266 ( .A1(n10319), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8735) );
  NAND2_X1 U11267 ( .A1(n8737), .A2(n8735), .ZN(n8844) );
  INV_X1 U11268 ( .A(n8844), .ZN(n8736) );
  NAND2_X1 U11269 ( .A1(n8845), .A2(n8736), .ZN(n8738) );
  NAND2_X1 U11270 ( .A1(n8738), .A2(n8737), .ZN(n8857) );
  NAND2_X1 U11271 ( .A1(n10322), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8739) );
  NAND2_X1 U11272 ( .A1(n8741), .A2(n8739), .ZN(n8858) );
  INV_X1 U11273 ( .A(n8858), .ZN(n8740) );
  NAND2_X1 U11274 ( .A1(n8857), .A2(n8740), .ZN(n8742) );
  NAND2_X1 U11275 ( .A1(n10317), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8743) );
  NAND2_X1 U11276 ( .A1(n8745), .A2(n8743), .ZN(n8871) );
  INV_X1 U11277 ( .A(n8871), .ZN(n8744) );
  NAND2_X1 U11278 ( .A1(n10326), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8746) );
  NAND2_X1 U11279 ( .A1(n8748), .A2(n8746), .ZN(n8887) );
  INV_X1 U11280 ( .A(n8887), .ZN(n8747) );
  NAND2_X1 U11281 ( .A1(n10330), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8749) );
  NAND2_X1 U11282 ( .A1(n8906), .A2(n8749), .ZN(n8751) );
  NAND2_X1 U11283 ( .A1(n10331), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8750) );
  NAND2_X1 U11284 ( .A1(n10347), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8752) );
  NAND2_X1 U11285 ( .A1(n8754), .A2(n8752), .ZN(n8919) );
  NAND2_X1 U11286 ( .A1(n10334), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U11287 ( .A1(n10351), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8758) );
  NAND2_X1 U11288 ( .A1(n10350), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8757) );
  NAND2_X1 U11289 ( .A1(n8759), .A2(n8758), .ZN(n8965) );
  NAND2_X1 U11290 ( .A1(n10401), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8761) );
  NAND2_X1 U11291 ( .A1(n10402), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8760) );
  NAND2_X1 U11292 ( .A1(n10411), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8763) );
  NAND2_X1 U11293 ( .A1(n10412), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8762) );
  NAND2_X1 U11294 ( .A1(n10487), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8766) );
  NAND2_X1 U11295 ( .A1(n10485), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8764) );
  NAND2_X1 U11296 ( .A1(n8766), .A2(n8764), .ZN(n8992) );
  INV_X1 U11297 ( .A(n8992), .ZN(n8765) );
  NAND2_X1 U11298 ( .A1(n10555), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8772) );
  NAND2_X1 U11299 ( .A1(n10558), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8768) );
  NAND2_X1 U11300 ( .A1(n8772), .A2(n8768), .ZN(n9020) );
  AND2_X1 U11301 ( .A1(n10505), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n8769) );
  NOR2_X1 U11302 ( .A1(n9020), .A2(n8769), .ZN(n8770) );
  NAND2_X1 U11303 ( .A1(n10670), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8774) );
  NAND2_X1 U11304 ( .A1(n10669), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8773) );
  NAND2_X1 U11305 ( .A1(n8774), .A2(n8773), .ZN(n9033) );
  NAND2_X1 U11306 ( .A1(n8775), .A2(n8774), .ZN(n9050) );
  NAND2_X1 U11307 ( .A1(n10715), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8778) );
  NAND2_X1 U11308 ( .A1(n10713), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8776) );
  NAND2_X1 U11309 ( .A1(n8778), .A2(n8776), .ZN(n9049) );
  INV_X1 U11310 ( .A(n9049), .ZN(n8777) );
  NAND2_X1 U11311 ( .A1(n10872), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8780) );
  NAND2_X1 U11312 ( .A1(n10874), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8779) );
  INV_X1 U11313 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11061) );
  NAND2_X1 U11314 ( .A1(n11061), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8782) );
  INV_X1 U11315 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11063) );
  NAND2_X1 U11316 ( .A1(n11063), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8781) );
  AND2_X1 U11317 ( .A1(n8782), .A2(n8781), .ZN(n9063) );
  INV_X1 U11318 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11138) );
  NAND2_X1 U11319 ( .A1(n11138), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8784) );
  INV_X1 U11320 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11136) );
  NAND2_X1 U11321 ( .A1(n11136), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8783) );
  AND2_X1 U11322 ( .A1(n8784), .A2(n8783), .ZN(n9095) );
  NAND2_X1 U11323 ( .A1(n11708), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8788) );
  NAND2_X1 U11324 ( .A1(n15733), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8787) );
  AND2_X1 U11325 ( .A1(n8788), .A2(n8787), .ZN(n9126) );
  XNOR2_X1 U11326 ( .A(n11909), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n9141) );
  XNOR2_X1 U11327 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n9162) );
  NAND2_X1 U11328 ( .A1(n11863), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8789) );
  NAND2_X1 U11329 ( .A1(n8790), .A2(n8789), .ZN(n8791) );
  NAND2_X1 U11330 ( .A1(n8791), .A2(n12127), .ZN(n8792) );
  NAND2_X1 U11331 ( .A1(n14373), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8793) );
  INV_X1 U11332 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n15175) );
  NAND2_X1 U11333 ( .A1(n15175), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8794) );
  NAND2_X1 U11334 ( .A1(n8795), .A2(n8794), .ZN(n9190) );
  INV_X1 U11335 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15170) );
  AND2_X1 U11336 ( .A1(n15170), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8796) );
  NAND2_X1 U11337 ( .A1(n14368), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8797) );
  AND2_X1 U11338 ( .A1(n14364), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8800) );
  INV_X1 U11339 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n12449) );
  NAND2_X1 U11340 ( .A1(n12449), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8799) );
  XNOR2_X1 U11341 ( .A(n15165), .B(P1_DATAO_REG_28__SCAN_IN), .ZN(n8801) );
  XNOR2_X1 U11342 ( .A(n12272), .B(n8801), .ZN(n13241) );
  OR2_X1 U11343 ( .A1(n8806), .A2(n7647), .ZN(n8803) );
  NAND2_X1 U11344 ( .A1(n13241), .A2(n12294), .ZN(n8809) );
  INV_X4 U11345 ( .A(n9038), .ZN(n12297) );
  NAND2_X1 U11346 ( .A1(n12297), .A2(SI_28_), .ZN(n8808) );
  NAND2_X1 U11347 ( .A1(n10849), .A2(n12316), .ZN(n8810) );
  NAND2_X1 U11348 ( .A1(n8810), .A2(n11291), .ZN(n8813) );
  OAI21_X1 U11349 ( .B1(n9286), .B2(n11291), .A(n12343), .ZN(n8811) );
  NAND2_X1 U11350 ( .A1(n8811), .A2(n10849), .ZN(n8812) );
  NAND2_X1 U11351 ( .A1(n8813), .A2(n8812), .ZN(n10858) );
  AND2_X1 U11352 ( .A1(n15651), .A2(n8814), .ZN(n8815) );
  NAND2_X1 U11353 ( .A1(n10858), .A2(n8815), .ZN(n8817) );
  NAND2_X1 U11354 ( .A1(n12316), .A2(n12343), .ZN(n15586) );
  OR2_X1 U11355 ( .A1(n15586), .A2(n12368), .ZN(n15659) );
  NAND2_X1 U11356 ( .A1(n8818), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8819) );
  MUX2_X1 U11357 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8819), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n8820) );
  NAND2_X1 U11358 ( .A1(n6447), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8827) );
  AND2_X2 U11359 ( .A1(n12461), .A2(n8823), .ZN(n8851) );
  NAND2_X1 U11360 ( .A1(n8851), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8826) );
  INV_X1 U11361 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n8822) );
  NAND2_X1 U11362 ( .A1(n6448), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8824) );
  NAND4_X2 U11363 ( .A1(n8827), .A2(n8826), .A3(n8825), .A4(n8824), .ZN(n15605) );
  INV_X1 U11364 ( .A(n15605), .ZN(n8831) );
  INV_X1 U11365 ( .A(SI_0_), .ZN(n10421) );
  NAND2_X1 U11366 ( .A1(n10443), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8828) );
  NAND2_X1 U11367 ( .A1(n8836), .A2(n8828), .ZN(n10419) );
  NAND2_X1 U11368 ( .A1(n9099), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n8829) );
  NAND2_X1 U11369 ( .A1(n8831), .A2(n11397), .ZN(n13008) );
  NAND2_X1 U11370 ( .A1(n8897), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8835) );
  NAND2_X1 U11371 ( .A1(n8851), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8834) );
  INV_X1 U11372 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n8832) );
  OR2_X1 U11373 ( .A1(n8880), .A2(n8832), .ZN(n8833) );
  INV_X1 U11374 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n13015) );
  INV_X1 U11375 ( .A(SI_1_), .ZN(n8837) );
  NAND2_X1 U11376 ( .A1(n15592), .A2(n13014), .ZN(n12165) );
  NAND2_X1 U11378 ( .A1(n9058), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8843) );
  NAND2_X1 U11379 ( .A1(n6448), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8842) );
  INV_X1 U11380 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n8839) );
  OR2_X1 U11381 ( .A1(n8880), .A2(n8839), .ZN(n8841) );
  INV_X1 U11382 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10203) );
  OR2_X1 U11383 ( .A1(n12300), .A2(n10203), .ZN(n8840) );
  NAND2_X1 U11384 ( .A1(n12297), .A2(n10430), .ZN(n8849) );
  XNOR2_X1 U11385 ( .A(n8845), .B(n8844), .ZN(n10431) );
  NAND2_X1 U11386 ( .A1(n12294), .A2(n10431), .ZN(n8848) );
  NAND2_X1 U11387 ( .A1(n9099), .A2(n10947), .ZN(n8847) );
  INV_X1 U11388 ( .A(n15585), .ZN(n10896) );
  NAND2_X1 U11389 ( .A1(n8850), .A2(n12171), .ZN(n11449) );
  NAND2_X1 U11390 ( .A1(n9058), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8856) );
  NAND2_X1 U11391 ( .A1(n6449), .A2(n15680), .ZN(n8855) );
  INV_X1 U11392 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n8852) );
  OR2_X1 U11393 ( .A1(n8880), .A2(n8852), .ZN(n8854) );
  INV_X1 U11394 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11453) );
  NAND2_X1 U11395 ( .A1(n12297), .A2(n10422), .ZN(n8864) );
  XNOR2_X1 U11396 ( .A(n8857), .B(n8858), .ZN(n10424) );
  NAND2_X1 U11397 ( .A1(n12294), .A2(n10424), .ZN(n8863) );
  NAND2_X1 U11398 ( .A1(n8859), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8861) );
  INV_X1 U11399 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8860) );
  NAND2_X1 U11400 ( .A1(n9099), .A2(n10423), .ZN(n8862) );
  NAND2_X1 U11401 ( .A1(n15591), .A2(n15615), .ZN(n12174) );
  INV_X1 U11402 ( .A(n15615), .ZN(n11011) );
  NAND2_X1 U11403 ( .A1(n15620), .A2(n11011), .ZN(n12172) );
  AND2_X2 U11404 ( .A1(n12174), .A2(n12172), .ZN(n12323) );
  NAND2_X1 U11405 ( .A1(n11449), .A2(n12323), .ZN(n11448) );
  NAND2_X1 U11406 ( .A1(n11448), .A2(n12174), .ZN(n11523) );
  NAND2_X1 U11407 ( .A1(n9058), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8870) );
  NAND2_X1 U11408 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8865) );
  NAND2_X1 U11409 ( .A1(n8878), .A2(n8865), .ZN(n11530) );
  NAND2_X1 U11410 ( .A1(n6449), .A2(n11530), .ZN(n8869) );
  INV_X1 U11411 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n8866) );
  OR2_X1 U11412 ( .A1(n8880), .A2(n8866), .ZN(n8868) );
  INV_X1 U11413 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11529) );
  XNOR2_X1 U11414 ( .A(n8872), .B(n8871), .ZN(n10437) );
  NAND2_X1 U11415 ( .A1(n9099), .A2(n10436), .ZN(n8873) );
  INV_X1 U11416 ( .A(n15619), .ZN(n11170) );
  NAND2_X1 U11417 ( .A1(n11170), .A2(n12645), .ZN(n12175) );
  NAND2_X1 U11418 ( .A1(n9058), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8885) );
  NAND2_X1 U11419 ( .A1(n8878), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8879) );
  NAND2_X1 U11420 ( .A1(n8898), .A2(n8879), .ZN(n11540) );
  NAND2_X1 U11421 ( .A1(n6449), .A2(n11540), .ZN(n8884) );
  INV_X1 U11422 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n8881) );
  OR2_X1 U11423 ( .A1(n8880), .A2(n8881), .ZN(n8883) );
  INV_X1 U11424 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11539) );
  OR2_X1 U11425 ( .A1(n12300), .A2(n11539), .ZN(n8882) );
  INV_X1 U11426 ( .A(SI_5_), .ZN(n10425) );
  NAND2_X1 U11427 ( .A1(n12297), .A2(n10425), .ZN(n8895) );
  XNOR2_X1 U11428 ( .A(n8886), .B(n8887), .ZN(n10426) );
  NAND2_X1 U11429 ( .A1(n12294), .A2(n10426), .ZN(n8894) );
  NAND2_X1 U11430 ( .A1(n8889), .A2(n8888), .ZN(n8890) );
  NAND2_X1 U11431 ( .A1(n8890), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8892) );
  XNOR2_X1 U11432 ( .A(n8892), .B(n8891), .ZN(n11130) );
  NAND2_X1 U11433 ( .A1(n9099), .A2(n11130), .ZN(n8893) );
  NAND2_X1 U11434 ( .A1(n15623), .A2(n11541), .ZN(n12180) );
  INV_X1 U11435 ( .A(n11541), .ZN(n15627) );
  NAND2_X1 U11436 ( .A1(n15639), .A2(n15627), .ZN(n12181) );
  INV_X1 U11437 ( .A(n12320), .ZN(n8896) );
  NAND2_X1 U11438 ( .A1(n9058), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8904) );
  NAND2_X1 U11439 ( .A1(n8898), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8899) );
  NAND2_X1 U11440 ( .A1(n8913), .A2(n8899), .ZN(n11546) );
  NAND2_X1 U11441 ( .A1(n6448), .A2(n11546), .ZN(n8903) );
  INV_X1 U11442 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n8900) );
  OR2_X1 U11443 ( .A1(n8880), .A2(n8900), .ZN(n8902) );
  INV_X1 U11444 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11518) );
  OR2_X1 U11445 ( .A1(n12300), .A2(n11518), .ZN(n8901) );
  AND4_X2 U11446 ( .A1(n8904), .A2(n8903), .A3(n8902), .A4(n8901), .ZN(n15653)
         );
  XNOR2_X1 U11447 ( .A(n10330), .B(P1_DATAO_REG_6__SCAN_IN), .ZN(n8905) );
  XNOR2_X1 U11448 ( .A(n8906), .B(n8905), .ZN(n10417) );
  NAND2_X1 U11449 ( .A1(n12297), .A2(SI_6_), .ZN(n8911) );
  INV_X1 U11450 ( .A(n8907), .ZN(n8909) );
  NOR2_X1 U11451 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n8908) );
  NAND2_X1 U11452 ( .A1(n8909), .A2(n8908), .ZN(n8923) );
  NAND2_X1 U11453 ( .A1(n8923), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8910) );
  XNOR2_X1 U11454 ( .A(n8910), .B(P3_IR_REG_6__SCAN_IN), .ZN(n10218) );
  NAND2_X1 U11455 ( .A1(n15653), .A2(n15636), .ZN(n12187) );
  NAND2_X1 U11456 ( .A1(n8851), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8918) );
  NAND2_X1 U11457 ( .A1(n9273), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8917) );
  NAND2_X1 U11458 ( .A1(n8913), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8914) );
  NAND2_X1 U11459 ( .A1(n8931), .A2(n8914), .ZN(n11666) );
  NAND2_X1 U11460 ( .A1(n6449), .A2(n11666), .ZN(n8916) );
  NAND2_X1 U11461 ( .A1(n7776), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8915) );
  NAND4_X1 U11462 ( .A1(n8918), .A2(n8917), .A3(n8916), .A4(n8915), .ZN(n12644) );
  NAND2_X1 U11463 ( .A1(n8920), .A2(n8919), .ZN(n8921) );
  NAND2_X1 U11464 ( .A1(n8922), .A2(n8921), .ZN(n10434) );
  NAND2_X1 U11465 ( .A1(n12294), .A2(n10434), .ZN(n8927) );
  NAND2_X1 U11466 ( .A1(n8939), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8925) );
  INV_X1 U11467 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8924) );
  XNOR2_X1 U11468 ( .A(n8925), .B(n8924), .ZN(n10433) );
  NAND2_X1 U11469 ( .A1(n9099), .A2(n10433), .ZN(n8926) );
  OAI211_X1 U11470 ( .C1(n9038), .C2(SI_7_), .A(n8927), .B(n8926), .ZN(n15650)
         );
  XNOR2_X1 U11471 ( .A(n12644), .B(n15650), .ZN(n11636) );
  INV_X1 U11472 ( .A(n11636), .ZN(n12324) );
  INV_X2 U11473 ( .A(n15653), .ZN(n15630) );
  INV_X1 U11474 ( .A(n15636), .ZN(n8928) );
  INV_X1 U11475 ( .A(n12644), .ZN(n15643) );
  INV_X1 U11476 ( .A(n15650), .ZN(n12188) );
  NAND2_X1 U11477 ( .A1(n15643), .A2(n12188), .ZN(n8929) );
  NAND2_X1 U11478 ( .A1(n8930), .A2(n8929), .ZN(n11955) );
  NAND2_X1 U11479 ( .A1(n9058), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8937) );
  NAND2_X1 U11480 ( .A1(n8931), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8932) );
  NAND2_X1 U11481 ( .A1(n8958), .A2(n8932), .ZN(n11962) );
  NAND2_X1 U11482 ( .A1(n6449), .A2(n11962), .ZN(n8936) );
  INV_X1 U11483 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n8933) );
  OR2_X1 U11484 ( .A1(n8880), .A2(n8933), .ZN(n8935) );
  INV_X1 U11485 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11961) );
  OR2_X1 U11486 ( .A1(n12300), .A2(n11961), .ZN(n8934) );
  INV_X1 U11487 ( .A(SI_8_), .ZN(n10427) );
  NAND2_X1 U11488 ( .A1(n8951), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8941) );
  INV_X1 U11489 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8940) );
  OAI22_X1 U11490 ( .A1(n9038), .A2(n10427), .B1(n10166), .B2(n10428), .ZN(
        n8947) );
  OR2_X1 U11491 ( .A1(n8943), .A2(n8942), .ZN(n8944) );
  NAND2_X1 U11492 ( .A1(n8945), .A2(n8944), .ZN(n10429) );
  NAND2_X1 U11493 ( .A1(n11663), .A2(n13127), .ZN(n12194) );
  INV_X1 U11494 ( .A(n13127), .ZN(n9234) );
  NAND2_X1 U11495 ( .A1(n15655), .A2(n9234), .ZN(n12195) );
  XNOR2_X1 U11496 ( .A(n8950), .B(n8949), .ZN(n10340) );
  NAND2_X1 U11497 ( .A1(n10340), .A2(n12294), .ZN(n8955) );
  INV_X1 U11498 ( .A(SI_9_), .ZN(n10341) );
  OAI21_X1 U11499 ( .B1(n8951), .B2(P3_IR_REG_8__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8953) );
  INV_X1 U11500 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8952) );
  XNOR2_X1 U11501 ( .A(n8953), .B(n8952), .ZN(n11466) );
  AOI22_X1 U11502 ( .A1(n12297), .A2(n10341), .B1(n9099), .B2(n11466), .ZN(
        n8954) );
  NAND2_X1 U11503 ( .A1(n9273), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8963) );
  NAND2_X1 U11504 ( .A1(n7776), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8962) );
  NAND2_X1 U11505 ( .A1(n8958), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n8959) );
  NAND2_X1 U11506 ( .A1(n8973), .A2(n8959), .ZN(n11922) );
  NAND2_X1 U11507 ( .A1(n6449), .A2(n11922), .ZN(n8961) );
  NAND2_X1 U11508 ( .A1(n9058), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8960) );
  NOR2_X1 U11509 ( .A1(n12057), .A2(n12643), .ZN(n12198) );
  NAND2_X1 U11510 ( .A1(n12057), .A2(n12643), .ZN(n12200) );
  OR2_X1 U11511 ( .A1(n8965), .A2(n8964), .ZN(n8966) );
  NAND2_X1 U11512 ( .A1(n8967), .A2(n8966), .ZN(n10439) );
  NAND2_X1 U11513 ( .A1(n10439), .A2(n12294), .ZN(n8972) );
  INV_X1 U11514 ( .A(SI_10_), .ZN(n10438) );
  OR2_X1 U11515 ( .A1(n8968), .A2(n7647), .ZN(n8970) );
  XNOR2_X1 U11516 ( .A(n8970), .B(n8969), .ZN(n11607) );
  AOI22_X1 U11517 ( .A1(n12297), .A2(n10438), .B1(n9099), .B2(n11607), .ZN(
        n8971) );
  NAND2_X1 U11518 ( .A1(n8972), .A2(n8971), .ZN(n11744) );
  NAND2_X1 U11519 ( .A1(n9058), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8978) );
  NAND2_X1 U11520 ( .A1(n9273), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8977) );
  NAND2_X1 U11521 ( .A1(n8973), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8974) );
  NAND2_X1 U11522 ( .A1(n8985), .A2(n8974), .ZN(n12120) );
  NAND2_X1 U11523 ( .A1(n6448), .A2(n12120), .ZN(n8976) );
  NAND2_X1 U11524 ( .A1(n7776), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8975) );
  NAND2_X1 U11525 ( .A1(n11744), .A2(n12998), .ZN(n9237) );
  INV_X1 U11526 ( .A(n9237), .ZN(n12205) );
  XNOR2_X1 U11527 ( .A(n8980), .B(n8979), .ZN(n10355) );
  NAND2_X1 U11528 ( .A1(n10355), .A2(n12294), .ZN(n8984) );
  NAND2_X1 U11529 ( .A1(n8693), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8981) );
  MUX2_X1 U11530 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8981), .S(
        P3_IR_REG_11__SCAN_IN), .Z(n8982) );
  OR2_X1 U11531 ( .A1(n8693), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n9005) );
  NAND2_X1 U11532 ( .A1(n8982), .A2(n9005), .ZN(n10354) );
  AOI22_X1 U11533 ( .A1(n12297), .A2(n10356), .B1(n9099), .B2(n10354), .ZN(
        n8983) );
  NAND2_X1 U11534 ( .A1(n8984), .A2(n8983), .ZN(n13002) );
  NAND2_X1 U11535 ( .A1(n9058), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8990) );
  NAND2_X1 U11536 ( .A1(n8985), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8986) );
  NAND2_X1 U11537 ( .A1(n8997), .A2(n8986), .ZN(n13003) );
  NAND2_X1 U11538 ( .A1(n6449), .A2(n13003), .ZN(n8989) );
  INV_X1 U11539 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n13215) );
  OR2_X1 U11540 ( .A1(n8880), .A2(n13215), .ZN(n8988) );
  INV_X1 U11541 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n13001) );
  OR2_X1 U11542 ( .A1(n12300), .A2(n13001), .ZN(n8987) );
  NAND2_X1 U11543 ( .A1(n13002), .A2(n12642), .ZN(n12209) );
  XNOR2_X1 U11544 ( .A(n8993), .B(n8992), .ZN(n10414) );
  NAND2_X1 U11545 ( .A1(n10414), .A2(n12294), .ZN(n8996) );
  NAND2_X1 U11546 ( .A1(n9005), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8994) );
  XNOR2_X1 U11547 ( .A(n8994), .B(P3_IR_REG_12__SCAN_IN), .ZN(n10230) );
  AOI22_X1 U11548 ( .A1(n12297), .A2(SI_12_), .B1(n9099), .B2(n10230), .ZN(
        n8995) );
  NAND2_X1 U11549 ( .A1(n8996), .A2(n8995), .ZN(n13111) );
  NAND2_X1 U11550 ( .A1(n8997), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8998) );
  NAND2_X1 U11551 ( .A1(n9011), .A2(n8998), .ZN(n12987) );
  NAND2_X1 U11552 ( .A1(n6449), .A2(n12987), .ZN(n9002) );
  NAND2_X1 U11553 ( .A1(n9058), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n9001) );
  INV_X1 U11554 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n13211) );
  OR2_X1 U11555 ( .A1(n8880), .A2(n13211), .ZN(n9000) );
  INV_X1 U11556 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n10153) );
  OR2_X1 U11557 ( .A1(n12300), .A2(n10153), .ZN(n8999) );
  OR2_X1 U11558 ( .A1(n13111), .A2(n11996), .ZN(n12212) );
  NAND2_X1 U11559 ( .A1(n13111), .A2(n11996), .ZN(n12213) );
  NAND2_X1 U11560 ( .A1(n12212), .A2(n12213), .ZN(n12984) );
  NAND2_X1 U11561 ( .A1(n9003), .A2(n10507), .ZN(n9018) );
  OR2_X1 U11562 ( .A1(n9003), .A2(n10507), .ZN(n9004) );
  NAND2_X1 U11563 ( .A1(n9018), .A2(n9004), .ZN(n9019) );
  XNOR2_X1 U11564 ( .A(n9019), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n10508) );
  NAND2_X1 U11565 ( .A1(n10508), .A2(n12294), .ZN(n9008) );
  NOR2_X1 U11566 ( .A1(n9005), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n9023) );
  OR2_X1 U11567 ( .A1(n9023), .A2(n7647), .ZN(n9006) );
  XNOR2_X1 U11568 ( .A(n9006), .B(P3_IR_REG_13__SCAN_IN), .ZN(n10233) );
  AOI22_X1 U11569 ( .A1(n12297), .A2(SI_13_), .B1(n9099), .B2(n10233), .ZN(
        n9007) );
  INV_X1 U11570 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n9009) );
  NAND2_X1 U11571 ( .A1(n9011), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9012) );
  NAND2_X1 U11572 ( .A1(n9027), .A2(n9012), .ZN(n12979) );
  NAND2_X1 U11573 ( .A1(n6449), .A2(n12979), .ZN(n9016) );
  NAND2_X1 U11574 ( .A1(n9058), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n9015) );
  INV_X1 U11575 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n13205) );
  OR2_X1 U11576 ( .A1(n8880), .A2(n13205), .ZN(n9014) );
  INV_X1 U11577 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12978) );
  OR2_X1 U11578 ( .A1(n12300), .A2(n12978), .ZN(n9013) );
  NAND2_X1 U11579 ( .A1(n13206), .A2(n12985), .ZN(n12217) );
  INV_X1 U11580 ( .A(n12217), .ZN(n9017) );
  OAI21_X1 U11581 ( .B1(n9019), .B2(n10505), .A(n9018), .ZN(n9021) );
  XNOR2_X1 U11582 ( .A(n9021), .B(n9020), .ZN(n10559) );
  NAND2_X1 U11583 ( .A1(n10559), .A2(n12294), .ZN(n9026) );
  NAND2_X1 U11584 ( .A1(n9023), .A2(n9022), .ZN(n9035) );
  NAND2_X1 U11585 ( .A1(n9035), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9024) );
  XNOR2_X1 U11586 ( .A(n9024), .B(P3_IR_REG_14__SCAN_IN), .ZN(n10560) );
  AOI22_X1 U11587 ( .A1(n12297), .A2(SI_14_), .B1(n9099), .B2(n10560), .ZN(
        n9025) );
  NAND2_X1 U11588 ( .A1(n9058), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9032) );
  NAND2_X1 U11589 ( .A1(n9027), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9028) );
  NAND2_X1 U11590 ( .A1(n9042), .A2(n9028), .ZN(n12971) );
  NAND2_X1 U11591 ( .A1(n6448), .A2(n12971), .ZN(n9031) );
  INV_X1 U11592 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13199) );
  OR2_X1 U11593 ( .A1(n8880), .A2(n13199), .ZN(n9030) );
  INV_X1 U11594 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12970) );
  OR2_X1 U11595 ( .A1(n12300), .A2(n12970), .ZN(n9029) );
  NAND2_X1 U11596 ( .A1(n13200), .A2(n12953), .ZN(n12220) );
  XNOR2_X1 U11597 ( .A(n9034), .B(n9033), .ZN(n10500) );
  NAND2_X1 U11598 ( .A1(n10500), .A2(n12294), .ZN(n9041) );
  OAI21_X1 U11599 ( .B1(n9035), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9036) );
  MUX2_X1 U11600 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9036), .S(
        P3_IR_REG_15__SCAN_IN), .Z(n9037) );
  NAND2_X1 U11601 ( .A1(n9037), .A2(n9051), .ZN(n10501) );
  OAI22_X1 U11602 ( .A1(n9038), .A2(n10503), .B1(n10166), .B2(n10501), .ZN(
        n9039) );
  INV_X1 U11603 ( .A(n9039), .ZN(n9040) );
  NAND2_X1 U11604 ( .A1(n9042), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9043) );
  NAND2_X1 U11605 ( .A1(n9056), .A2(n9043), .ZN(n12955) );
  NAND2_X1 U11606 ( .A1(n12955), .A2(n6449), .ZN(n9047) );
  NAND2_X1 U11607 ( .A1(n9273), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9046) );
  NAND2_X1 U11608 ( .A1(n7776), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n9045) );
  NAND2_X1 U11609 ( .A1(n9058), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n9044) );
  OR2_X1 U11610 ( .A1(n13100), .A2(n12943), .ZN(n12221) );
  NAND2_X1 U11611 ( .A1(n13100), .A2(n12943), .ZN(n12229) );
  NAND2_X1 U11612 ( .A1(n12221), .A2(n12229), .ZN(n12952) );
  NAND2_X1 U11613 ( .A1(n12950), .A2(n6696), .ZN(n9048) );
  NAND2_X1 U11614 ( .A1(n9048), .A2(n12229), .ZN(n12940) );
  XNOR2_X1 U11615 ( .A(n9050), .B(n9049), .ZN(n10551) );
  NAND2_X1 U11616 ( .A1(n10551), .A2(n12294), .ZN(n9055) );
  NAND2_X1 U11617 ( .A1(n9051), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9052) );
  MUX2_X1 U11618 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9052), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n9053) );
  AND2_X1 U11619 ( .A1(n9053), .A2(n9083), .ZN(n12722) );
  AOI22_X1 U11620 ( .A1(n12297), .A2(SI_16_), .B1(n9099), .B2(n12722), .ZN(
        n9054) );
  NAND2_X1 U11621 ( .A1(n9056), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9057) );
  NAND2_X1 U11622 ( .A1(n9089), .A2(n9057), .ZN(n12945) );
  NAND2_X1 U11623 ( .A1(n12945), .A2(n6448), .ZN(n9061) );
  AOI22_X1 U11624 ( .A1(n9058), .A2(P3_REG1_REG_16__SCAN_IN), .B1(n9273), .B2(
        P3_REG0_REG_16__SCAN_IN), .ZN(n9060) );
  NAND2_X1 U11625 ( .A1(n7776), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n9059) );
  NAND2_X1 U11626 ( .A1(n13094), .A2(n13097), .ZN(n12228) );
  NAND2_X1 U11627 ( .A1(n12222), .A2(n12228), .ZN(n12941) );
  INV_X1 U11628 ( .A(n12941), .ZN(n12336) );
  NAND2_X1 U11629 ( .A1(n12940), .A2(n12336), .ZN(n9062) );
  OR2_X1 U11630 ( .A1(n9064), .A2(n9063), .ZN(n9065) );
  NAND2_X1 U11631 ( .A1(n9066), .A2(n9065), .ZN(n10636) );
  INV_X1 U11632 ( .A(n9067), .ZN(n9085) );
  NAND2_X1 U11633 ( .A1(n9085), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9068) );
  MUX2_X1 U11634 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9068), .S(
        P3_IR_REG_18__SCAN_IN), .Z(n9069) );
  AND2_X1 U11635 ( .A1(n9070), .A2(n9069), .ZN(n12752) );
  AOI22_X1 U11636 ( .A1(n12297), .A2(SI_18_), .B1(n9099), .B2(n12752), .ZN(
        n9071) );
  NAND2_X1 U11637 ( .A1(n9072), .A2(n9071), .ZN(n12924) );
  INV_X1 U11638 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n9073) );
  NAND2_X1 U11639 ( .A1(n9091), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9075) );
  NAND2_X1 U11640 ( .A1(n9102), .A2(n9075), .ZN(n12917) );
  NAND2_X1 U11641 ( .A1(n12917), .A2(n6448), .ZN(n9078) );
  AOI22_X1 U11642 ( .A1(n8851), .A2(P3_REG1_REG_18__SCAN_IN), .B1(n9273), .B2(
        P3_REG0_REG_18__SCAN_IN), .ZN(n9077) );
  NAND2_X1 U11643 ( .A1(n7776), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9076) );
  NAND2_X1 U11644 ( .A1(n12924), .A2(n13085), .ZN(n12232) );
  OR2_X1 U11645 ( .A1(n9080), .A2(n9079), .ZN(n9081) );
  NAND2_X1 U11646 ( .A1(n9082), .A2(n9081), .ZN(n10564) );
  NAND2_X1 U11647 ( .A1(n9083), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9084) );
  MUX2_X1 U11648 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9084), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n9086) );
  NAND2_X1 U11649 ( .A1(n9086), .A2(n9085), .ZN(n10565) );
  INV_X1 U11650 ( .A(n10565), .ZN(n12736) );
  AOI22_X1 U11651 ( .A1(n12297), .A2(SI_17_), .B1(n9099), .B2(n12736), .ZN(
        n9087) );
  NAND2_X1 U11652 ( .A1(n9089), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9090) );
  NAND2_X1 U11653 ( .A1(n9091), .A2(n9090), .ZN(n12935) );
  NAND2_X1 U11654 ( .A1(n12935), .A2(n6449), .ZN(n9094) );
  AOI22_X1 U11655 ( .A1(n9273), .A2(P3_REG0_REG_17__SCAN_IN), .B1(n7776), .B2(
        P3_REG2_REG_17__SCAN_IN), .ZN(n9093) );
  NAND2_X1 U11656 ( .A1(n8851), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n9092) );
  NAND2_X1 U11657 ( .A1(n13088), .A2(n13091), .ZN(n12159) );
  NAND2_X1 U11658 ( .A1(n12232), .A2(n12159), .ZN(n9111) );
  OR2_X1 U11659 ( .A1(n9096), .A2(n9095), .ZN(n9097) );
  NAND2_X1 U11660 ( .A1(n9098), .A2(n9097), .ZN(n10717) );
  NAND2_X1 U11661 ( .A1(n10717), .A2(n12294), .ZN(n9101) );
  AOI22_X1 U11662 ( .A1(n12297), .A2(n10716), .B1(n9099), .B2(n12357), .ZN(
        n9100) );
  NOR2_X2 U11663 ( .A1(n9102), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9118) );
  INV_X1 U11664 ( .A(n9118), .ZN(n9119) );
  NAND2_X1 U11665 ( .A1(n9102), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9103) );
  NAND2_X1 U11666 ( .A1(n9119), .A2(n9103), .ZN(n12911) );
  NAND2_X1 U11667 ( .A1(n12911), .A2(n6449), .ZN(n9108) );
  INV_X1 U11668 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13076) );
  NAND2_X1 U11669 ( .A1(n9273), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9105) );
  NAND2_X1 U11670 ( .A1(n7776), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n9104) );
  OAI211_X1 U11671 ( .C1(n13076), .C2(n9276), .A(n9105), .B(n9104), .ZN(n9106)
         );
  INV_X1 U11672 ( .A(n9106), .ZN(n9107) );
  NAND2_X1 U11673 ( .A1(n12910), .A2(n12638), .ZN(n12238) );
  OR2_X1 U11674 ( .A1(n13088), .A2(n13091), .ZN(n9251) );
  INV_X1 U11675 ( .A(n9251), .ZN(n9109) );
  NAND2_X1 U11676 ( .A1(n12232), .A2(n9109), .ZN(n12235) );
  OR2_X1 U11677 ( .A1(n12924), .A2(n13085), .ZN(n12898) );
  AND3_X1 U11678 ( .A1(n12238), .A2(n12235), .A3(n12898), .ZN(n9110) );
  NAND2_X1 U11679 ( .A1(n9113), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9114) );
  NAND2_X1 U11680 ( .A1(n9115), .A2(n9114), .ZN(n10965) );
  NAND2_X1 U11681 ( .A1(n12297), .A2(SI_20_), .ZN(n9116) );
  INV_X1 U11682 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n15793) );
  NAND2_X1 U11683 ( .A1(n9119), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9120) );
  NAND2_X1 U11684 ( .A1(n12891), .A2(n6449), .ZN(n9125) );
  INV_X1 U11685 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13074) );
  NAND2_X1 U11686 ( .A1(n7776), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n9122) );
  NAND2_X1 U11687 ( .A1(n9273), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n9121) );
  OAI211_X1 U11688 ( .C1(n9276), .C2(n13074), .A(n9122), .B(n9121), .ZN(n9123)
         );
  INV_X1 U11689 ( .A(n9123), .ZN(n9124) );
  NAND2_X1 U11690 ( .A1(n13073), .A2(n12528), .ZN(n12242) );
  NAND2_X1 U11691 ( .A1(n9129), .A2(n9128), .ZN(n12380) );
  NAND2_X1 U11692 ( .A1(n12297), .A2(SI_21_), .ZN(n9130) );
  INV_X1 U11693 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n9132) );
  NAND2_X1 U11694 ( .A1(n9134), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9135) );
  NAND2_X1 U11695 ( .A1(n9145), .A2(n9135), .ZN(n12878) );
  NAND2_X1 U11696 ( .A1(n12878), .A2(n6449), .ZN(n9140) );
  INV_X1 U11697 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13067) );
  NAND2_X1 U11698 ( .A1(n7776), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n9137) );
  NAND2_X1 U11699 ( .A1(n9273), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n9136) );
  OAI211_X1 U11700 ( .C1(n9276), .C2(n13067), .A(n9137), .B(n9136), .ZN(n9138)
         );
  INV_X1 U11701 ( .A(n9138), .ZN(n9139) );
  NAND2_X1 U11702 ( .A1(n13168), .A2(n12889), .ZN(n12248) );
  OR2_X1 U11703 ( .A1(n13168), .A2(n12889), .ZN(n12247) );
  XNOR2_X1 U11704 ( .A(n9142), .B(n9141), .ZN(n11293) );
  NAND2_X1 U11705 ( .A1(n11293), .A2(n12294), .ZN(n9144) );
  NAND2_X1 U11706 ( .A1(n12297), .A2(SI_22_), .ZN(n9143) );
  NAND2_X1 U11707 ( .A1(n9145), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9146) );
  NAND2_X1 U11708 ( .A1(n9166), .A2(n9146), .ZN(n12864) );
  NAND2_X1 U11709 ( .A1(n12864), .A2(n6448), .ZN(n9151) );
  INV_X1 U11710 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13064) );
  NAND2_X1 U11711 ( .A1(n9273), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n9148) );
  NAND2_X1 U11712 ( .A1(n7776), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n9147) );
  OAI211_X1 U11713 ( .C1(n9276), .C2(n13064), .A(n9148), .B(n9147), .ZN(n9149)
         );
  INV_X1 U11714 ( .A(n9149), .ZN(n9150) );
  NAND2_X1 U11715 ( .A1(n13162), .A2(n12848), .ZN(n12251) );
  INV_X1 U11716 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12115) );
  NAND2_X1 U11717 ( .A1(n12297), .A2(SI_24_), .ZN(n9154) );
  INV_X1 U11718 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n9155) );
  NAND2_X1 U11719 ( .A1(n9168), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9156) );
  NAND2_X1 U11720 ( .A1(n9182), .A2(n9156), .ZN(n12832) );
  NAND2_X1 U11721 ( .A1(n12832), .A2(n6448), .ZN(n9161) );
  INV_X1 U11722 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n15677) );
  NAND2_X1 U11723 ( .A1(n7776), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n9158) );
  NAND2_X1 U11724 ( .A1(n9273), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n9157) );
  OAI211_X1 U11725 ( .C1(n9276), .C2(n15677), .A(n9158), .B(n9157), .ZN(n9159)
         );
  INV_X1 U11726 ( .A(n9159), .ZN(n9160) );
  XNOR2_X1 U11727 ( .A(n9163), .B(n9162), .ZN(n11557) );
  NAND2_X1 U11728 ( .A1(n11557), .A2(n12294), .ZN(n9165) );
  NAND2_X1 U11729 ( .A1(n12297), .A2(SI_23_), .ZN(n9164) );
  NAND2_X1 U11730 ( .A1(n9166), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9167) );
  NAND2_X1 U11731 ( .A1(n9168), .A2(n9167), .ZN(n12843) );
  NAND2_X1 U11732 ( .A1(n12843), .A2(n6449), .ZN(n9173) );
  INV_X1 U11733 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13062) );
  NAND2_X1 U11734 ( .A1(n7776), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n9170) );
  NAND2_X1 U11735 ( .A1(n9273), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n9169) );
  OAI211_X1 U11736 ( .C1(n9276), .C2(n13062), .A(n9170), .B(n9169), .ZN(n9171)
         );
  INV_X1 U11737 ( .A(n9171), .ZN(n9172) );
  OR2_X1 U11738 ( .A1(n13061), .A2(n13050), .ZN(n12830) );
  NAND2_X1 U11739 ( .A1(n12253), .A2(n12830), .ZN(n12254) );
  NAND3_X1 U11740 ( .A1(n12253), .A2(n13050), .A3(n13061), .ZN(n9174) );
  NAND2_X1 U11741 ( .A1(n13056), .A2(n13058), .ZN(n12255) );
  AND2_X1 U11742 ( .A1(n9174), .A2(n12255), .ZN(n9175) );
  XNOR2_X1 U11743 ( .A(n14373), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n9176) );
  XNOR2_X1 U11744 ( .A(n9177), .B(n9176), .ZN(n13255) );
  NAND2_X1 U11745 ( .A1(n13255), .A2(n12294), .ZN(n9179) );
  NAND2_X1 U11746 ( .A1(n12297), .A2(SI_25_), .ZN(n9178) );
  INV_X1 U11747 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n9180) );
  NAND2_X1 U11748 ( .A1(n9182), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9183) );
  NAND2_X1 U11749 ( .A1(n9193), .A2(n9183), .ZN(n12823) );
  NAND2_X1 U11750 ( .A1(n12823), .A2(n6449), .ZN(n9188) );
  INV_X1 U11751 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n15679) );
  NAND2_X1 U11752 ( .A1(n9058), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9185) );
  NAND2_X1 U11753 ( .A1(n7776), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9184) );
  OAI211_X1 U11754 ( .C1(n8880), .C2(n15679), .A(n9185), .B(n9184), .ZN(n9186)
         );
  INV_X1 U11755 ( .A(n9186), .ZN(n9187) );
  NAND2_X1 U11756 ( .A1(n13046), .A2(n13051), .ZN(n12259) );
  XNOR2_X1 U11758 ( .A(n15170), .B(P1_DATAO_REG_26__SCAN_IN), .ZN(n9189) );
  XNOR2_X1 U11759 ( .A(n9190), .B(n9189), .ZN(n13251) );
  NAND2_X1 U11760 ( .A1(n13251), .A2(n12294), .ZN(n9192) );
  NAND2_X1 U11761 ( .A1(n12297), .A2(SI_26_), .ZN(n9191) );
  NAND2_X1 U11762 ( .A1(n9193), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9194) );
  NAND2_X1 U11763 ( .A1(n9207), .A2(n9194), .ZN(n12810) );
  NAND2_X1 U11764 ( .A1(n12810), .A2(n6449), .ZN(n9199) );
  INV_X1 U11765 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13041) );
  NAND2_X1 U11766 ( .A1(n7776), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n9196) );
  NAND2_X1 U11767 ( .A1(n9273), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n9195) );
  OAI211_X1 U11768 ( .C1(n9276), .C2(n13041), .A(n9196), .B(n9195), .ZN(n9197)
         );
  INV_X1 U11769 ( .A(n9197), .ZN(n9198) );
  NAND2_X1 U11770 ( .A1(n13034), .A2(n13043), .ZN(n12263) );
  XNOR2_X1 U11771 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n9201) );
  XNOR2_X1 U11772 ( .A(n9202), .B(n9201), .ZN(n13245) );
  NAND2_X1 U11773 ( .A1(n13245), .A2(n12294), .ZN(n9204) );
  NAND2_X1 U11774 ( .A1(n12297), .A2(SI_27_), .ZN(n9203) );
  INV_X1 U11775 ( .A(n9207), .ZN(n9206) );
  INV_X1 U11776 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n9205) );
  NAND2_X1 U11777 ( .A1(n9207), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9208) );
  NAND2_X1 U11778 ( .A1(n9214), .A2(n9208), .ZN(n12802) );
  NAND2_X1 U11779 ( .A1(n12802), .A2(n6449), .ZN(n9213) );
  INV_X1 U11780 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n13032) );
  NAND2_X1 U11781 ( .A1(n9273), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n9210) );
  NAND2_X1 U11782 ( .A1(n7776), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n9209) );
  OAI211_X1 U11783 ( .C1(n13032), .C2(n9276), .A(n9210), .B(n9209), .ZN(n9211)
         );
  INV_X1 U11784 ( .A(n9211), .ZN(n9212) );
  NAND2_X1 U11785 ( .A1(n12801), .A2(n12618), .ZN(n12157) );
  NAND2_X1 U11786 ( .A1(n12792), .A2(n12157), .ZN(n9223) );
  NAND2_X1 U11787 ( .A1(n9214), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9215) );
  NAND2_X1 U11788 ( .A1(n12761), .A2(n9215), .ZN(n12540) );
  NAND2_X1 U11789 ( .A1(n12540), .A2(n6448), .ZN(n9221) );
  INV_X1 U11790 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n9218) );
  NAND2_X1 U11791 ( .A1(n9273), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n9217) );
  NAND2_X1 U11792 ( .A1(n7776), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n9216) );
  OAI211_X1 U11793 ( .C1(n9276), .C2(n9218), .A(n9217), .B(n9216), .ZN(n9219)
         );
  INV_X1 U11794 ( .A(n9219), .ZN(n9220) );
  NAND2_X1 U11795 ( .A1(n12772), .A2(n12796), .ZN(n12158) );
  INV_X1 U11796 ( .A(n12536), .ZN(n9222) );
  NAND2_X1 U11797 ( .A1(n15605), .A2(n11397), .ZN(n13017) );
  NAND2_X1 U11798 ( .A1(n13018), .A2(n13017), .ZN(n9225) );
  NAND2_X1 U11799 ( .A1(n15592), .A2(n10845), .ZN(n9224) );
  NAND2_X1 U11800 ( .A1(n9225), .A2(n9224), .ZN(n15589) );
  NAND2_X1 U11801 ( .A1(n15589), .A2(n15590), .ZN(n9227) );
  NAND2_X1 U11802 ( .A1(n15608), .A2(n10896), .ZN(n9226) );
  NAND2_X1 U11803 ( .A1(n9227), .A2(n9226), .ZN(n11450) );
  AND2_X1 U11804 ( .A1(n15620), .A2(n15615), .ZN(n11524) );
  AOI22_X1 U11805 ( .A1(n11526), .A2(n11524), .B1(n15619), .B2(n12645), .ZN(
        n9228) );
  NAND2_X1 U11806 ( .A1(n15623), .A2(n15627), .ZN(n9229) );
  NAND2_X1 U11807 ( .A1(n12187), .A2(n12182), .ZN(n12321) );
  NAND2_X1 U11808 ( .A1(n15630), .A2(n15636), .ZN(n9230) );
  NAND2_X1 U11809 ( .A1(n12644), .A2(n12188), .ZN(n9231) );
  NAND2_X1 U11810 ( .A1(n11663), .A2(n9234), .ZN(n9235) );
  INV_X1 U11811 ( .A(n12057), .ZN(n11923) );
  NAND2_X1 U11812 ( .A1(n11923), .A2(n12643), .ZN(n9236) );
  NAND2_X1 U11813 ( .A1(n12204), .A2(n9237), .ZN(n12201) );
  INV_X1 U11814 ( .A(n11744), .ZN(n13122) );
  OR2_X1 U11815 ( .A1(n13002), .A2(n13119), .ZN(n9238) );
  NAND2_X1 U11816 ( .A1(n9239), .A2(n9238), .ZN(n12983) );
  NAND2_X1 U11817 ( .A1(n12983), .A2(n12984), .ZN(n9241) );
  NAND2_X1 U11818 ( .A1(n13111), .A2(n12999), .ZN(n9240) );
  NAND2_X1 U11819 ( .A1(n12216), .A2(n12217), .ZN(n12974) );
  NAND2_X1 U11820 ( .A1(n13200), .A2(n12976), .ZN(n9245) );
  INV_X1 U11821 ( .A(n9245), .ZN(n9242) );
  NAND2_X1 U11822 ( .A1(n12219), .A2(n12220), .ZN(n12966) );
  AND2_X1 U11823 ( .A1(n12974), .A2(n9244), .ZN(n9243) );
  NAND2_X1 U11824 ( .A1(n12962), .A2(n9243), .ZN(n9249) );
  INV_X1 U11825 ( .A(n9244), .ZN(n9247) );
  INV_X1 U11826 ( .A(n12985), .ZN(n12967) );
  NAND2_X1 U11827 ( .A1(n13206), .A2(n12967), .ZN(n12963) );
  AND2_X1 U11828 ( .A1(n12963), .A2(n9245), .ZN(n9246) );
  NAND2_X1 U11829 ( .A1(n9249), .A2(n9248), .ZN(n12951) );
  NAND2_X1 U11830 ( .A1(n12951), .A2(n12952), .ZN(n12929) );
  INV_X1 U11831 ( .A(n12943), .ZN(n12968) );
  NAND2_X1 U11832 ( .A1(n13100), .A2(n12968), .ZN(n12928) );
  INV_X1 U11833 ( .A(n13097), .ZN(n12641) );
  NAND2_X1 U11834 ( .A1(n13094), .A2(n12641), .ZN(n12930) );
  NAND2_X1 U11835 ( .A1(n13088), .A2(n12640), .ZN(n9250) );
  AND2_X1 U11836 ( .A1(n12930), .A2(n9250), .ZN(n9253) );
  AND2_X1 U11837 ( .A1(n12928), .A2(n9253), .ZN(n9257) );
  INV_X1 U11838 ( .A(n9250), .ZN(n9252) );
  NAND2_X1 U11839 ( .A1(n9251), .A2(n12159), .ZN(n12932) );
  OR2_X1 U11840 ( .A1(n9252), .A2(n12932), .ZN(n9256) );
  INV_X1 U11841 ( .A(n9253), .ZN(n9254) );
  OR2_X1 U11842 ( .A1(n9254), .A2(n12941), .ZN(n9255) );
  AND2_X1 U11843 ( .A1(n13168), .A2(n12860), .ZN(n12244) );
  NAND2_X1 U11844 ( .A1(n13073), .A2(n12908), .ZN(n12870) );
  OR2_X1 U11845 ( .A1(n12910), .A2(n13070), .ZN(n12886) );
  NAND2_X1 U11846 ( .A1(n12898), .A2(n12232), .ZN(n12884) );
  AND2_X1 U11847 ( .A1(n12886), .A2(n12884), .ZN(n12868) );
  NAND2_X1 U11848 ( .A1(n12870), .A2(n12868), .ZN(n12854) );
  INV_X1 U11849 ( .A(n12244), .ZN(n12855) );
  INV_X1 U11850 ( .A(n13085), .ZN(n12639) );
  OR2_X1 U11851 ( .A1(n12924), .A2(n12639), .ZN(n12901) );
  NAND2_X1 U11852 ( .A1(n12900), .A2(n12901), .ZN(n12885) );
  NAND2_X1 U11853 ( .A1(n12885), .A2(n12886), .ZN(n9260) );
  NAND2_X1 U11854 ( .A1(n9261), .A2(n12243), .ZN(n12856) );
  AOI22_X1 U11855 ( .A1(n12855), .A2(n12856), .B1(n12489), .B2(n12848), .ZN(
        n9262) );
  NAND2_X1 U11856 ( .A1(n13162), .A2(n12875), .ZN(n9263) );
  XNOR2_X1 U11857 ( .A(n13061), .B(n13050), .ZN(n12847) );
  NAND2_X1 U11858 ( .A1(n13061), .A2(n12861), .ZN(n9264) );
  AND2_X1 U11859 ( .A1(n13056), .A2(n12637), .ZN(n9267) );
  OR2_X1 U11860 ( .A1(n13056), .A2(n12637), .ZN(n9266) );
  OR2_X1 U11861 ( .A1(n13034), .A2(n12822), .ZN(n9268) );
  OR2_X1 U11862 ( .A1(n12801), .A2(n13036), .ZN(n9270) );
  NAND2_X1 U11863 ( .A1(n12163), .A2(n9286), .ZN(n12359) );
  NAND2_X1 U11864 ( .A1(n12343), .A2(n12368), .ZN(n9287) );
  INV_X1 U11865 ( .A(n12768), .ZN(n9280) );
  INV_X1 U11866 ( .A(n12761), .ZN(n9272) );
  NAND2_X1 U11867 ( .A1(n9272), .A2(n6449), .ZN(n12306) );
  INV_X1 U11868 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n13027) );
  NAND2_X1 U11869 ( .A1(n9273), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9275) );
  NAND2_X1 U11870 ( .A1(n7776), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9274) );
  OAI211_X1 U11871 ( .C1(n13027), .C2(n9276), .A(n9275), .B(n9274), .ZN(n9277)
         );
  INV_X1 U11872 ( .A(n9277), .ZN(n9278) );
  NAND2_X1 U11873 ( .A1(n12306), .A2(n9278), .ZN(n12636) );
  INV_X1 U11874 ( .A(n13243), .ZN(n12758) );
  INV_X1 U11875 ( .A(n13246), .ZN(n10198) );
  NAND2_X1 U11876 ( .A1(n12758), .A2(n10198), .ZN(n10169) );
  NAND2_X1 U11877 ( .A1(n10169), .A2(n10166), .ZN(n10843) );
  INV_X1 U11878 ( .A(n10843), .ZN(n10839) );
  OAI21_X1 U11879 ( .B1(n9283), .B2(n9295), .A(n9282), .ZN(P3_U3487) );
  INV_X1 U11880 ( .A(n9284), .ZN(n9290) );
  NAND2_X1 U11881 ( .A1(n10849), .A2(n9286), .ZN(n12361) );
  OR2_X1 U11882 ( .A1(n12361), .A2(n9287), .ZN(n10860) );
  OR2_X1 U11883 ( .A1(n12267), .A2(n9288), .ZN(n10966) );
  OAI21_X1 U11884 ( .B1(n10840), .B2(n10860), .A(n10835), .ZN(n9289) );
  NAND2_X1 U11885 ( .A1(n10859), .A2(n9289), .ZN(n9293) );
  NAND3_X1 U11886 ( .A1(n10862), .A2(n10865), .A3(n10858), .ZN(n9292) );
  INV_X1 U11887 ( .A(n13217), .ZN(n9296) );
  INV_X1 U11888 ( .A(n12772), .ZN(n9295) );
  OAI21_X1 U11889 ( .B1(n9296), .B2(n9295), .A(n9294), .ZN(P3_U3455) );
  NOR2_X1 U11890 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n9300) );
  NAND4_X1 U11891 ( .A1(n9300), .A2(n9299), .A3(n9298), .A4(n9297), .ZN(n9367)
         );
  INV_X1 U11892 ( .A(n9367), .ZN(n9306) );
  NAND2_X1 U11893 ( .A1(n9322), .A2(n9377), .ZN(n9366) );
  NOR2_X2 U11894 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9450) );
  NAND2_X1 U11895 ( .A1(n9317), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9311) );
  AND2_X1 U11896 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n9318) );
  NAND3_X1 U11897 ( .A1(n9328), .A2(P1_IR_REG_27__SCAN_IN), .A3(n9335), .ZN(
        n9315) );
  XNOR2_X1 U11898 ( .A(P1_IR_REG_27__SCAN_IN), .B(P1_IR_REG_31__SCAN_IN), .ZN(
        n9314) );
  NAND2_X1 U11899 ( .A1(n10484), .A2(n9461), .ZN(n9325) );
  OR2_X1 U11900 ( .A1(n9322), .A2(n15153), .ZN(n9323) );
  NAND2_X1 U11901 ( .A1(n9533), .A2(n9323), .ZN(n9376) );
  INV_X2 U11902 ( .A(n10407), .ZN(n9669) );
  AOI22_X1 U11903 ( .A1(n14585), .A2(n9669), .B1(P2_DATAO_REG_12__SCAN_IN), 
        .B2(n9924), .ZN(n9324) );
  NAND2_X1 U11904 ( .A1(n9313), .A2(n9328), .ZN(n9334) );
  NOR2_X1 U11905 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n9329) );
  NAND2_X1 U11906 ( .A1(n9334), .A2(n9329), .ZN(n9330) );
  XNOR2_X1 U11907 ( .A(n15153), .B(P1_IR_REG_25__SCAN_IN), .ZN(n9331) );
  NAND2_X1 U11908 ( .A1(n9334), .A2(n9331), .ZN(n9332) );
  NAND2_X1 U11909 ( .A1(n9334), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9333) );
  MUX2_X1 U11910 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9333), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n9338) );
  INV_X1 U11911 ( .A(n9334), .ZN(n9336) );
  NAND2_X1 U11912 ( .A1(n9336), .A2(n9335), .ZN(n9337) );
  NAND2_X1 U11913 ( .A1(n9345), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9340) );
  INV_X1 U11914 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n15706) );
  MUX2_X1 U11915 ( .A(n9340), .B(P1_IR_REG_31__SCAN_IN), .S(n15706), .Z(n9342)
         );
  INV_X1 U11916 ( .A(n9341), .ZN(n9358) );
  NAND2_X1 U11917 ( .A1(n9343), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9344) );
  MUX2_X1 U11918 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9344), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n9346) );
  NAND2_X1 U11919 ( .A1(n9346), .A2(n9345), .ZN(n11513) );
  NAND2_X4 U11920 ( .A1(n10296), .A2(n9943), .ZN(n9801) );
  NAND2_X1 U11921 ( .A1(n9382), .A2(n14417), .ZN(n9350) );
  AND2_X1 U11922 ( .A1(n9584), .A2(n9350), .ZN(n14418) );
  NAND2_X1 U11923 ( .A1(n6445), .A2(n14418), .ZN(n9357) );
  AND2_X4 U11924 ( .A1(n15158), .A2(n9351), .ZN(n9919) );
  NAND2_X1 U11925 ( .A1(n9919), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9356) );
  INV_X2 U11926 ( .A(n9886), .ZN(n9920) );
  NAND2_X1 U11927 ( .A1(n9920), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9355) );
  INV_X4 U11928 ( .A(n9353), .ZN(n9927) );
  NAND2_X1 U11929 ( .A1(n9927), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9354) );
  NAND4_X1 U11930 ( .A1(n9357), .A2(n9356), .A3(n9355), .A4(n9354), .ZN(n14983) );
  INV_X1 U11931 ( .A(n14983), .ZN(n12013) );
  INV_X1 U11932 ( .A(n15344), .ZN(n9363) );
  OAI22_X1 U11933 ( .A1(n7770), .A2(n9801), .B1(n12013), .B2(n9800), .ZN(n9574) );
  NAND2_X1 U11934 ( .A1(n15121), .A2(n12427), .ZN(n9365) );
  NAND2_X1 U11935 ( .A1(n14983), .A2(n12422), .ZN(n9364) );
  NAND2_X1 U11936 ( .A1(n9365), .A2(n9364), .ZN(n9375) );
  OR2_X1 U11937 ( .A1(n9367), .A2(n9366), .ZN(n9368) );
  INV_X1 U11938 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9370) );
  NAND2_X1 U11939 ( .A1(n9371), .A2(n9370), .ZN(n9373) );
  XNOR2_X1 U11940 ( .A(P1_IR_REG_19__SCAN_IN), .B(P1_IR_REG_31__SCAN_IN), .ZN(
        n9372) );
  XNOR2_X1 U11941 ( .A(n9375), .B(n12425), .ZN(n9575) );
  NAND2_X1 U11942 ( .A1(n10409), .A2(n9461), .ZN(n9379) );
  XNOR2_X1 U11943 ( .A(n9377), .B(n9376), .ZN(n11317) );
  AOI22_X1 U11944 ( .A1(n11317), .A2(n9669), .B1(P2_DATAO_REG_11__SCAN_IN), 
        .B2(n9924), .ZN(n9378) );
  INV_X1 U11945 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9381) );
  INV_X1 U11946 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9380) );
  OAI21_X1 U11947 ( .B1(n9553), .B2(n9381), .A(n9380), .ZN(n9383) );
  AND2_X1 U11948 ( .A1(n9383), .A2(n9382), .ZN(n12041) );
  NAND2_X1 U11949 ( .A1(n6445), .A2(n12041), .ZN(n9387) );
  NAND2_X1 U11950 ( .A1(n9919), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n9386) );
  NAND2_X1 U11951 ( .A1(n9927), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n9385) );
  NAND2_X1 U11952 ( .A1(n9920), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9384) );
  NOR2_X1 U11953 ( .A1(n12071), .A2(n9800), .ZN(n9388) );
  AOI21_X1 U11954 ( .B1(n15126), .B2(n12422), .A(n9388), .ZN(n9571) );
  INV_X1 U11955 ( .A(n9571), .ZN(n9573) );
  NAND2_X1 U11956 ( .A1(n15126), .A2(n12427), .ZN(n9390) );
  INV_X1 U11957 ( .A(n12071), .ZN(n14502) );
  NAND2_X1 U11958 ( .A1(n14502), .A2(n12422), .ZN(n9389) );
  NAND2_X1 U11959 ( .A1(n9390), .A2(n9389), .ZN(n9391) );
  XNOR2_X1 U11960 ( .A(n9391), .B(n12425), .ZN(n9572) );
  INV_X1 U11961 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9392) );
  NAND2_X1 U11962 ( .A1(n9413), .A2(n9392), .ZN(n9393) );
  AND2_X1 U11963 ( .A1(n9500), .A2(n9393), .ZN(n11115) );
  NAND2_X1 U11964 ( .A1(n6445), .A2(n11115), .ZN(n9397) );
  NAND2_X1 U11965 ( .A1(n9919), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9396) );
  NAND2_X1 U11966 ( .A1(n9920), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9395) );
  NAND2_X1 U11967 ( .A1(n9927), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9394) );
  NAND4_X1 U11968 ( .A1(n9397), .A2(n9396), .A3(n9395), .A4(n9394), .ZN(n14507) );
  INV_X1 U11969 ( .A(n14507), .ZN(n11251) );
  NAND2_X1 U11970 ( .A1(n10329), .A2(n9461), .ZN(n9402) );
  NAND2_X1 U11971 ( .A1(n9406), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9399) );
  INV_X1 U11972 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9398) );
  XNOR2_X1 U11973 ( .A(n9399), .B(n9398), .ZN(n10495) );
  OAI22_X1 U11974 ( .A1(n9690), .A2(n10330), .B1(n7215), .B2(n10495), .ZN(
        n9400) );
  INV_X1 U11975 ( .A(n9400), .ZN(n9401) );
  OAI22_X1 U11976 ( .A1(n11251), .A2(n9801), .B1(n11250), .B2(n9745), .ZN(
        n9403) );
  XOR2_X1 U11977 ( .A(n12425), .B(n9403), .Z(n11437) );
  NAND2_X1 U11978 ( .A1(n10325), .A2(n9461), .ZN(n9410) );
  NAND2_X1 U11979 ( .A1(n9404), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9405) );
  MUX2_X1 U11980 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9405), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n9407) );
  NAND2_X1 U11981 ( .A1(n9407), .A2(n9406), .ZN(n10471) );
  OAI22_X1 U11982 ( .A1(n9690), .A2(n10326), .B1(n7215), .B2(n10471), .ZN(
        n9408) );
  INV_X1 U11983 ( .A(n9408), .ZN(n9409) );
  INV_X1 U11984 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9411) );
  NAND2_X1 U11985 ( .A1(n9467), .A2(n9411), .ZN(n9412) );
  AND2_X1 U11986 ( .A1(n9413), .A2(n9412), .ZN(n15325) );
  NAND2_X1 U11987 ( .A1(n6445), .A2(n15325), .ZN(n9417) );
  NAND2_X1 U11988 ( .A1(n9919), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9416) );
  NAND2_X1 U11989 ( .A1(n9927), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9415) );
  NAND2_X1 U11990 ( .A1(n9920), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9414) );
  NAND2_X1 U11991 ( .A1(n14508), .A2(n12422), .ZN(n9418) );
  OAI21_X1 U11992 ( .B1(n15373), .B2(n9745), .A(n9418), .ZN(n9419) );
  XNOR2_X1 U11993 ( .A(n9419), .B(n12425), .ZN(n11431) );
  NAND2_X1 U11994 ( .A1(n9434), .A2(n14508), .ZN(n9420) );
  OAI21_X1 U11995 ( .B1(n15373), .B2(n9801), .A(n9420), .ZN(n11432) );
  OR2_X1 U11996 ( .A1(n11250), .A2(n9801), .ZN(n9422) );
  NAND2_X1 U11997 ( .A1(n9434), .A2(n14507), .ZN(n9421) );
  AND2_X1 U11998 ( .A1(n9422), .A2(n9421), .ZN(n11436) );
  INV_X1 U11999 ( .A(n11436), .ZN(n9492) );
  AOI21_X1 U12000 ( .B1(n11431), .B2(n11432), .A(n9492), .ZN(n9494) );
  NAND2_X1 U12001 ( .A1(n9919), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9423) );
  INV_X1 U12002 ( .A(n9425), .ZN(n9449) );
  OAI22_X1 U12003 ( .A1(n10991), .A2(n9800), .B1(n6441), .B2(n9801), .ZN(n9440) );
  OAI22_X1 U12004 ( .A1(n10991), .A2(n9801), .B1(n6441), .B2(n9745), .ZN(n9426) );
  XNOR2_X1 U12005 ( .A(n9426), .B(n9560), .ZN(n9441) );
  XOR2_X1 U12006 ( .A(n9440), .B(n9441), .Z(n10662) );
  NAND2_X1 U12007 ( .A1(n9919), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9429) );
  NAND2_X1 U12008 ( .A1(n9458), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9428) );
  NAND2_X1 U12009 ( .A1(n9444), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9427) );
  OR2_X1 U12010 ( .A1(n11073), .A2(n9801), .ZN(n9433) );
  OAI21_X1 U12011 ( .B1(n6442), .B2(n10421), .A(n10443), .ZN(n9430) );
  AND2_X1 U12012 ( .A1(n9431), .A2(n9430), .ZN(n15178) );
  MUX2_X1 U12013 ( .A(P1_IR_REG_0__SCAN_IN), .B(n15178), .S(n10407), .Z(n14994) );
  INV_X1 U12014 ( .A(n10296), .ZN(n9436) );
  AOI22_X1 U12015 ( .A1(n12427), .A2(n14994), .B1(n9436), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n9432) );
  NAND2_X1 U12016 ( .A1(n9433), .A2(n9432), .ZN(n10687) );
  NAND2_X1 U12017 ( .A1(n9438), .A2(n9437), .ZN(n10688) );
  INV_X1 U12018 ( .A(n10688), .ZN(n9439) );
  NOR2_X1 U12019 ( .A1(n9441), .A2(n9440), .ZN(n9442) );
  NAND2_X1 U12020 ( .A1(n9443), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9448) );
  NAND2_X1 U12021 ( .A1(n9919), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9447) );
  NAND2_X1 U12022 ( .A1(n9458), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9446) );
  NAND2_X1 U12023 ( .A1(n9444), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9445) );
  NAND2_X1 U12024 ( .A1(n9449), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9453) );
  NAND2_X1 U12025 ( .A1(n9669), .A2(n14537), .ZN(n9452) );
  OAI22_X1 U12026 ( .A1(n9892), .A2(n9801), .B1(n9891), .B2(n9745), .ZN(n9454)
         );
  XNOR2_X1 U12027 ( .A(n9454), .B(n9560), .ZN(n9456) );
  OAI22_X1 U12028 ( .A1(n9892), .A2(n9800), .B1(n9891), .B2(n9801), .ZN(n9455)
         );
  XNOR2_X1 U12029 ( .A(n9456), .B(n9455), .ZN(n10654) );
  INV_X1 U12030 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9457) );
  NAND2_X1 U12031 ( .A1(n9443), .A2(n9457), .ZN(n9460) );
  NAND2_X1 U12032 ( .A1(n9458), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9459) );
  INV_X1 U12033 ( .A(n10323), .ZN(n9462) );
  NAND2_X1 U12034 ( .A1(n9462), .A2(n9461), .ZN(n9465) );
  NAND2_X1 U12035 ( .A1(n9319), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9463) );
  XNOR2_X1 U12036 ( .A(n9463), .B(n7023), .ZN(n14553) );
  OAI22_X1 U12037 ( .A1(n9425), .A2(n10322), .B1(n7215), .B2(n14553), .ZN(
        n9464) );
  OAI22_X1 U12038 ( .A1(n10980), .A2(n9801), .B1(n15356), .B2(n9745), .ZN(
        n9466) );
  XNOR2_X1 U12039 ( .A(n9466), .B(n9560), .ZN(n9483) );
  OAI22_X1 U12040 ( .A1(n10980), .A2(n9800), .B1(n15356), .B2(n9801), .ZN(
        n9484) );
  XNOR2_X1 U12041 ( .A(n9483), .B(n9484), .ZN(n10904) );
  OAI21_X1 U12042 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n9467), .ZN(n11002) );
  INV_X1 U12043 ( .A(n11002), .ZN(n9468) );
  NAND2_X1 U12044 ( .A1(n9443), .A2(n9468), .ZN(n9472) );
  NAND2_X1 U12045 ( .A1(n9919), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9471) );
  NAND2_X1 U12046 ( .A1(n9920), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9470) );
  NAND2_X1 U12047 ( .A1(n9927), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9469) );
  NAND2_X1 U12048 ( .A1(n14509), .A2(n12422), .ZN(n9479) );
  NAND2_X1 U12049 ( .A1(n9473), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9475) );
  XNOR2_X1 U12050 ( .A(n9475), .B(n9474), .ZN(n15271) );
  OAI22_X1 U12051 ( .A1(n9690), .A2(n10317), .B1(n7215), .B2(n15271), .ZN(
        n9476) );
  INV_X1 U12052 ( .A(n9476), .ZN(n9477) );
  NAND2_X1 U12053 ( .A1(n12427), .A2(n11104), .ZN(n9478) );
  NAND2_X1 U12054 ( .A1(n9479), .A2(n9478), .ZN(n9480) );
  XNOR2_X1 U12055 ( .A(n9480), .B(n12425), .ZN(n10303) );
  NAND2_X1 U12056 ( .A1(n9434), .A2(n14509), .ZN(n9482) );
  NAND2_X1 U12057 ( .A1(n12422), .A2(n11104), .ZN(n9481) );
  NAND2_X1 U12058 ( .A1(n9482), .A2(n9481), .ZN(n10302) );
  INV_X1 U12059 ( .A(n9483), .ZN(n9486) );
  INV_X1 U12060 ( .A(n9484), .ZN(n9485) );
  NOR2_X1 U12061 ( .A1(n9486), .A2(n9485), .ZN(n10301) );
  INV_X1 U12062 ( .A(n10303), .ZN(n9489) );
  INV_X1 U12063 ( .A(n10302), .ZN(n9488) );
  NAND2_X1 U12064 ( .A1(n11437), .A2(n11436), .ZN(n9491) );
  NAND3_X1 U12065 ( .A1(n11431), .A2(n11432), .A3(n9492), .ZN(n9493) );
  NAND2_X1 U12066 ( .A1(n10345), .A2(n9461), .ZN(n9498) );
  INV_X1 U12067 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9495) );
  OAI22_X1 U12068 ( .A1(n9690), .A2(n10346), .B1(n7215), .B2(n10540), .ZN(
        n9496) );
  INV_X1 U12069 ( .A(n9496), .ZN(n9497) );
  NAND2_X1 U12070 ( .A1(n15389), .A2(n12427), .ZN(n9507) );
  NAND2_X1 U12071 ( .A1(n9919), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9505) );
  NAND2_X1 U12072 ( .A1(n9500), .A2(n9499), .ZN(n9501) );
  AND2_X1 U12073 ( .A1(n9513), .A2(n9501), .ZN(n15309) );
  NAND2_X1 U12074 ( .A1(n9443), .A2(n15309), .ZN(n9504) );
  NAND2_X1 U12075 ( .A1(n9920), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9502) );
  NAND4_X1 U12076 ( .A1(n9505), .A2(n9504), .A3(n9503), .A4(n9502), .ZN(n14506) );
  NAND2_X1 U12077 ( .A1(n14506), .A2(n12422), .ZN(n9506) );
  NAND2_X1 U12078 ( .A1(n9507), .A2(n9506), .ZN(n9508) );
  XNOR2_X1 U12079 ( .A(n9508), .B(n12425), .ZN(n9510) );
  AOI22_X1 U12080 ( .A1(n15389), .A2(n12422), .B1(n9434), .B2(n14506), .ZN(
        n9509) );
  XNOR2_X1 U12081 ( .A(n9510), .B(n9509), .ZN(n11503) );
  INV_X1 U12082 ( .A(n9509), .ZN(n9511) );
  NAND2_X1 U12083 ( .A1(n9513), .A2(n9512), .ZN(n9514) );
  NAND2_X1 U12084 ( .A1(n9538), .A2(n9514), .ZN(n11598) );
  INV_X1 U12085 ( .A(n11598), .ZN(n9515) );
  NAND2_X1 U12086 ( .A1(n6445), .A2(n9515), .ZN(n9519) );
  NAND2_X1 U12087 ( .A1(n9919), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9518) );
  NAND2_X1 U12088 ( .A1(n9927), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n9517) );
  NAND2_X1 U12089 ( .A1(n9920), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9516) );
  NAND2_X1 U12090 ( .A1(n10333), .A2(n9461), .ZN(n9523) );
  NAND2_X1 U12091 ( .A1(n9520), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9521) );
  XNOR2_X1 U12092 ( .A(n9521), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10524) );
  AOI22_X1 U12093 ( .A1(n9924), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9669), .B2(
        n10524), .ZN(n9522) );
  NAND2_X1 U12094 ( .A1(n15397), .A2(n12427), .ZN(n9524) );
  OAI21_X1 U12095 ( .B1(n11983), .B2(n9801), .A(n9524), .ZN(n9525) );
  XNOR2_X1 U12096 ( .A(n9525), .B(n12425), .ZN(n9529) );
  NAND2_X1 U12097 ( .A1(n15397), .A2(n12422), .ZN(n9527) );
  OR2_X1 U12098 ( .A1(n11983), .A2(n9800), .ZN(n9526) );
  NAND2_X1 U12099 ( .A1(n9527), .A2(n9526), .ZN(n9528) );
  NOR2_X1 U12100 ( .A1(n9529), .A2(n9528), .ZN(n9530) );
  AOI21_X1 U12101 ( .B1(n9529), .B2(n9528), .A(n9530), .ZN(n11590) );
  INV_X1 U12102 ( .A(n9530), .ZN(n9531) );
  NAND2_X1 U12103 ( .A1(n10349), .A2(n9461), .ZN(n9536) );
  INV_X1 U12104 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9532) );
  OR2_X1 U12105 ( .A1(n9533), .A2(n9532), .ZN(n9534) );
  NAND2_X1 U12106 ( .A1(n9533), .A2(n9532), .ZN(n9549) );
  AOI22_X1 U12107 ( .A1(n10644), .A2(n9669), .B1(n9924), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n9535) );
  NAND2_X1 U12108 ( .A1(n9536), .A2(n9535), .ZN(n11987) );
  NAND2_X1 U12109 ( .A1(n11987), .A2(n12427), .ZN(n9545) );
  NAND2_X1 U12110 ( .A1(n9919), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n9543) );
  NAND2_X1 U12111 ( .A1(n9538), .A2(n9537), .ZN(n9539) );
  AND2_X1 U12112 ( .A1(n9553), .A2(n9539), .ZN(n15295) );
  NAND2_X1 U12113 ( .A1(n6445), .A2(n15295), .ZN(n9542) );
  NAND2_X1 U12114 ( .A1(n9927), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9541) );
  NAND2_X1 U12115 ( .A1(n9920), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9540) );
  OR2_X1 U12116 ( .A1(n11832), .A2(n9801), .ZN(n9544) );
  NAND2_X1 U12117 ( .A1(n9545), .A2(n9544), .ZN(n9546) );
  XNOR2_X1 U12118 ( .A(n9546), .B(n12425), .ZN(n11979) );
  NAND2_X1 U12119 ( .A1(n11987), .A2(n12422), .ZN(n9548) );
  OR2_X1 U12120 ( .A1(n11832), .A2(n9800), .ZN(n9547) );
  NAND2_X1 U12121 ( .A1(n9548), .A2(n9547), .ZN(n11941) );
  NOR2_X1 U12122 ( .A1(n11979), .A2(n11941), .ZN(n9564) );
  NAND2_X1 U12123 ( .A1(n10400), .A2(n9461), .ZN(n9552) );
  NAND2_X1 U12124 ( .A1(n9549), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9550) );
  XNOR2_X1 U12125 ( .A(n9550), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10703) );
  AOI22_X1 U12126 ( .A1(n10703), .A2(n9669), .B1(P2_DATAO_REG_10__SCAN_IN), 
        .B2(n9924), .ZN(n9551) );
  NAND2_X1 U12127 ( .A1(n9552), .A2(n9551), .ZN(n15417) );
  NAND2_X1 U12128 ( .A1(n15417), .A2(n12427), .ZN(n9559) );
  XNOR2_X1 U12129 ( .A(n9553), .B(P1_REG3_REG_10__SCAN_IN), .ZN(n11952) );
  NAND2_X1 U12130 ( .A1(n6445), .A2(n11952), .ZN(n9557) );
  NAND2_X1 U12131 ( .A1(n9919), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9556) );
  NAND2_X1 U12132 ( .A1(n9920), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9555) );
  NAND2_X1 U12133 ( .A1(n9927), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n9554) );
  NAND2_X1 U12134 ( .A1(n14503), .A2(n12422), .ZN(n9558) );
  NAND2_X1 U12135 ( .A1(n9559), .A2(n9558), .ZN(n9561) );
  INV_X1 U12136 ( .A(n9560), .ZN(n12411) );
  XNOR2_X1 U12137 ( .A(n9561), .B(n12411), .ZN(n11945) );
  NOR2_X1 U12138 ( .A1(n11981), .A2(n9800), .ZN(n9562) );
  AOI21_X1 U12139 ( .B1(n15417), .B2(n12422), .A(n9562), .ZN(n11944) );
  NAND2_X1 U12140 ( .A1(n11945), .A2(n11944), .ZN(n11943) );
  NOR2_X1 U12141 ( .A1(n9564), .A2(n9563), .ZN(n9565) );
  INV_X1 U12142 ( .A(n11944), .ZN(n9566) );
  AOI21_X1 U12143 ( .B1(n11979), .B2(n11941), .A(n9566), .ZN(n9568) );
  NAND3_X1 U12144 ( .A1(n11979), .A2(n11941), .A3(n9566), .ZN(n9567) );
  OAI21_X1 U12145 ( .B1(n9568), .B2(n11945), .A(n9567), .ZN(n9569) );
  INV_X1 U12146 ( .A(n9569), .ZN(n9570) );
  XOR2_X1 U12147 ( .A(n9571), .B(n9572), .Z(n11933) );
  XNOR2_X1 U12148 ( .A(n9575), .B(n9574), .ZN(n14413) );
  NAND2_X1 U12149 ( .A1(n10504), .A2(n9461), .ZN(n9581) );
  INV_X1 U12150 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9576) );
  NAND2_X1 U12151 ( .A1(n9577), .A2(n9576), .ZN(n9578) );
  NOR2_X1 U12152 ( .A1(n9690), .A2(n10507), .ZN(n9579) );
  AOI21_X1 U12153 ( .B1(n11340), .B2(n9669), .A(n9579), .ZN(n9580) );
  INV_X1 U12154 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9583) );
  NAND2_X1 U12155 ( .A1(n9584), .A2(n9583), .ZN(n9585) );
  AND2_X1 U12156 ( .A1(n9602), .A2(n9585), .ZN(n14975) );
  NAND2_X1 U12157 ( .A1(n6445), .A2(n14975), .ZN(n9589) );
  NAND2_X1 U12158 ( .A1(n9919), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9588) );
  NAND2_X1 U12159 ( .A1(n9920), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9587) );
  NAND2_X1 U12160 ( .A1(n9927), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n9586) );
  OAI22_X1 U12161 ( .A1(n14977), .A2(n9745), .B1(n14661), .B2(n9801), .ZN(
        n9590) );
  XNOR2_X1 U12162 ( .A(n9590), .B(n12425), .ZN(n9592) );
  NOR2_X1 U12163 ( .A1(n14661), .A2(n9800), .ZN(n9591) );
  AOI21_X1 U12164 ( .B1(n15116), .B2(n12422), .A(n9591), .ZN(n9593) );
  XNOR2_X1 U12165 ( .A(n9592), .B(n9593), .ZN(n14452) );
  NAND2_X1 U12166 ( .A1(n9592), .A2(n9594), .ZN(n9595) );
  NAND2_X1 U12167 ( .A1(n10554), .A2(n9461), .ZN(n9601) );
  INV_X1 U12168 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9596) );
  NAND2_X1 U12169 ( .A1(n9597), .A2(n9596), .ZN(n9598) );
  AOI22_X1 U12170 ( .A1(n11721), .A2(n9669), .B1(P2_DATAO_REG_14__SCAN_IN), 
        .B2(n9924), .ZN(n9600) );
  NAND2_X2 U12171 ( .A1(n9601), .A2(n9600), .ZN(n15107) );
  NAND2_X1 U12172 ( .A1(n9602), .A2(n11344), .ZN(n9603) );
  AND2_X1 U12173 ( .A1(n9634), .A2(n9603), .ZN(n14381) );
  AOI22_X1 U12174 ( .A1(n14381), .A2(n9443), .B1(n9919), .B2(
        P1_REG1_REG_14__SCAN_IN), .ZN(n9605) );
  AOI22_X1 U12175 ( .A1(n9927), .A2(P1_REG0_REG_14__SCAN_IN), .B1(n9920), .B2(
        P1_REG2_REG_14__SCAN_IN), .ZN(n9604) );
  NOR2_X1 U12176 ( .A1(n14981), .A2(n9801), .ZN(n9606) );
  AOI21_X1 U12177 ( .B1(n15107), .B2(n12427), .A(n9606), .ZN(n9607) );
  XNOR2_X1 U12178 ( .A(n9607), .B(n12425), .ZN(n9608) );
  INV_X1 U12179 ( .A(n14981), .ZN(n14689) );
  AOI22_X1 U12180 ( .A1(n15107), .A2(n12422), .B1(n9434), .B2(n14689), .ZN(
        n9609) );
  XNOR2_X1 U12181 ( .A(n9608), .B(n9609), .ZN(n14380) );
  NAND2_X1 U12182 ( .A1(n10712), .A2(n9461), .ZN(n9615) );
  OR2_X1 U12183 ( .A1(n9627), .A2(n15153), .ZN(n9611) );
  XNOR2_X1 U12184 ( .A(n9612), .B(n9611), .ZN(n14612) );
  OAI22_X1 U12185 ( .A1(n9690), .A2(n10715), .B1(n7215), .B2(n14612), .ZN(
        n9613) );
  INV_X1 U12186 ( .A(n9613), .ZN(n9614) );
  NAND2_X1 U12187 ( .A1(n14692), .A2(n12427), .ZN(n9622) );
  INV_X1 U12188 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9616) );
  NAND2_X1 U12189 ( .A1(n9636), .A2(n9616), .ZN(n9617) );
  AND2_X1 U12190 ( .A1(n9675), .A2(n9617), .ZN(n14947) );
  NAND2_X1 U12191 ( .A1(n14947), .A2(n6445), .ZN(n9620) );
  AOI22_X1 U12192 ( .A1(n9927), .A2(P1_REG0_REG_16__SCAN_IN), .B1(n9920), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n9619) );
  NAND2_X1 U12193 ( .A1(n9919), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9618) );
  OR2_X1 U12194 ( .A1(n14932), .A2(n9801), .ZN(n9621) );
  NAND2_X1 U12195 ( .A1(n9622), .A2(n9621), .ZN(n9623) );
  XNOR2_X1 U12196 ( .A(n9623), .B(n12425), .ZN(n14427) );
  AOI22_X1 U12197 ( .A1(n14692), .A2(n12422), .B1(n9434), .B2(n14691), .ZN(
        n14426) );
  INV_X1 U12198 ( .A(n14426), .ZN(n9644) );
  NAND2_X1 U12199 ( .A1(n10668), .A2(n9461), .ZN(n9632) );
  NOR2_X1 U12200 ( .A1(n9624), .A2(n15153), .ZN(n9625) );
  MUX2_X1 U12201 ( .A(n15153), .B(n9625), .S(P1_IR_REG_15__SCAN_IN), .Z(n9626)
         );
  INV_X1 U12202 ( .A(n9626), .ZN(n9629) );
  INV_X1 U12203 ( .A(n9627), .ZN(n9628) );
  NAND2_X1 U12204 ( .A1(n9629), .A2(n9628), .ZN(n14598) );
  OAI22_X1 U12205 ( .A1(n9690), .A2(n10670), .B1(n7215), .B2(n14598), .ZN(
        n9630) );
  INV_X1 U12206 ( .A(n9630), .ZN(n9631) );
  INV_X1 U12207 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9633) );
  NAND2_X1 U12208 ( .A1(n9634), .A2(n9633), .ZN(n9635) );
  NAND2_X1 U12209 ( .A1(n9636), .A2(n9635), .ZN(n14962) );
  INV_X1 U12210 ( .A(n6445), .ZN(n9876) );
  OR2_X1 U12211 ( .A1(n14962), .A2(n9876), .ZN(n9639) );
  AOI22_X1 U12212 ( .A1(n9927), .A2(P1_REG0_REG_15__SCAN_IN), .B1(n9920), .B2(
        P1_REG2_REG_15__SCAN_IN), .ZN(n9638) );
  NAND2_X1 U12213 ( .A1(n9919), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n9637) );
  NOR2_X1 U12214 ( .A1(n12018), .A2(n9800), .ZN(n9640) );
  AOI21_X1 U12215 ( .B1(n15103), .B2(n12422), .A(n9640), .ZN(n9645) );
  INV_X1 U12216 ( .A(n9645), .ZN(n14487) );
  NAND2_X1 U12217 ( .A1(n15103), .A2(n12427), .ZN(n9642) );
  NAND2_X1 U12218 ( .A1(n14690), .A2(n12422), .ZN(n9641) );
  NAND2_X1 U12219 ( .A1(n9642), .A2(n9641), .ZN(n9643) );
  XNOR2_X1 U12220 ( .A(n9643), .B(n12411), .ZN(n14425) );
  INV_X1 U12221 ( .A(n14425), .ZN(n9647) );
  AOI22_X1 U12222 ( .A1(n14427), .A2(n9644), .B1(n14487), .B2(n9647), .ZN(
        n9650) );
  AOI21_X1 U12223 ( .B1(n14425), .B2(n9645), .A(n14426), .ZN(n9648) );
  NAND2_X1 U12224 ( .A1(n14426), .A2(n9645), .ZN(n9646) );
  OAI22_X1 U12225 ( .A1(n9648), .A2(n14427), .B1(n9647), .B2(n9646), .ZN(n9649) );
  NAND2_X1 U12226 ( .A1(n10871), .A2(n9461), .ZN(n9655) );
  NAND2_X1 U12227 ( .A1(n6643), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9651) );
  MUX2_X1 U12228 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9651), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n9652) );
  OR2_X1 U12229 ( .A1(n6643), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n9667) );
  NAND2_X1 U12230 ( .A1(n9652), .A2(n9667), .ZN(n14625) );
  OAI22_X1 U12231 ( .A1(n9690), .A2(n10872), .B1(n14625), .B2(n7215), .ZN(
        n9653) );
  INV_X1 U12232 ( .A(n9653), .ZN(n9654) );
  XNOR2_X1 U12233 ( .A(n9675), .B(P1_REG3_REG_17__SCAN_IN), .ZN(n14934) );
  NAND2_X1 U12234 ( .A1(n14934), .A2(n6445), .ZN(n9660) );
  INV_X1 U12235 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14626) );
  NAND2_X1 U12236 ( .A1(n9920), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9657) );
  NAND2_X1 U12237 ( .A1(n9927), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n9656) );
  OAI211_X1 U12238 ( .C1(n14626), .C2(n9930), .A(n9657), .B(n9656), .ZN(n9658)
         );
  INV_X1 U12239 ( .A(n9658), .ZN(n9659) );
  NOR2_X1 U12240 ( .A1(n14921), .A2(n9801), .ZN(n9661) );
  AOI21_X1 U12241 ( .B1(n15088), .B2(n12427), .A(n9661), .ZN(n9662) );
  XNOR2_X1 U12242 ( .A(n9662), .B(n12425), .ZN(n9664) );
  AOI22_X1 U12243 ( .A1(n15088), .A2(n12422), .B1(n9434), .B2(n14500), .ZN(
        n9663) );
  XNOR2_X1 U12244 ( .A(n9664), .B(n9663), .ZN(n14438) );
  NAND2_X1 U12245 ( .A1(n9664), .A2(n9663), .ZN(n9665) );
  NAND2_X1 U12246 ( .A1(n11060), .A2(n9461), .ZN(n9671) );
  NAND2_X1 U12247 ( .A1(n9667), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9668) );
  XNOR2_X1 U12248 ( .A(n9668), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14640) );
  AOI22_X1 U12249 ( .A1(n9924), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n14640), 
        .B2(n9669), .ZN(n9670) );
  NAND2_X1 U12250 ( .A1(n15083), .A2(n12427), .ZN(n9684) );
  AND2_X1 U12251 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_REG3_REG_18__SCAN_IN), 
        .ZN(n9672) );
  INV_X1 U12252 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9674) );
  INV_X1 U12253 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9673) );
  OAI21_X1 U12254 ( .B1(n9675), .B2(n9674), .A(n9673), .ZN(n9676) );
  NAND2_X1 U12255 ( .A1(n9694), .A2(n9676), .ZN(n14914) );
  OR2_X1 U12256 ( .A1(n14914), .A2(n9876), .ZN(n9682) );
  INV_X1 U12257 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9679) );
  NAND2_X1 U12258 ( .A1(n9920), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9678) );
  NAND2_X1 U12259 ( .A1(n9927), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n9677) );
  OAI211_X1 U12260 ( .C1(n9679), .C2(n9930), .A(n9678), .B(n9677), .ZN(n9680)
         );
  INV_X1 U12261 ( .A(n9680), .ZN(n9681) );
  NAND2_X1 U12262 ( .A1(n9682), .A2(n9681), .ZN(n14902) );
  NAND2_X1 U12263 ( .A1(n14902), .A2(n12422), .ZN(n9683) );
  NAND2_X1 U12264 ( .A1(n9684), .A2(n9683), .ZN(n9685) );
  XNOR2_X1 U12265 ( .A(n9685), .B(n12425), .ZN(n9686) );
  AOI22_X1 U12266 ( .A1(n15083), .A2(n12422), .B1(n9434), .B2(n14902), .ZN(
        n9687) );
  XNOR2_X1 U12267 ( .A(n9686), .B(n9687), .ZN(n14470) );
  INV_X1 U12268 ( .A(n9686), .ZN(n9688) );
  NAND2_X1 U12269 ( .A1(n9688), .A2(n9687), .ZN(n9689) );
  NAND2_X1 U12270 ( .A1(n11135), .A2(n9461), .ZN(n9693) );
  OAI22_X1 U12271 ( .A1(n9690), .A2(n11138), .B1(n7215), .B2(n14817), .ZN(
        n9691) );
  INV_X1 U12272 ( .A(n9691), .ZN(n9692) );
  INV_X1 U12273 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n15744) );
  NAND2_X1 U12274 ( .A1(n9694), .A2(n15744), .ZN(n9695) );
  NAND2_X1 U12275 ( .A1(n9722), .A2(n9695), .ZN(n14896) );
  OR2_X1 U12276 ( .A1(n14896), .A2(n9876), .ZN(n9700) );
  INV_X1 U12277 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n15776) );
  NAND2_X1 U12278 ( .A1(n9919), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n9697) );
  NAND2_X1 U12279 ( .A1(n9920), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n9696) );
  OAI211_X1 U12280 ( .C1(n9353), .C2(n15776), .A(n9697), .B(n9696), .ZN(n9698)
         );
  INV_X1 U12281 ( .A(n9698), .ZN(n9699) );
  OAI22_X1 U12282 ( .A1(n14899), .A2(n9745), .B1(n14922), .B2(n9801), .ZN(
        n9701) );
  XNOR2_X1 U12283 ( .A(n9701), .B(n12425), .ZN(n9704) );
  OAI22_X1 U12284 ( .A1(n14899), .A2(n9801), .B1(n14922), .B2(n9800), .ZN(
        n9703) );
  XNOR2_X1 U12285 ( .A(n9704), .B(n9703), .ZN(n14396) );
  INV_X1 U12286 ( .A(n14396), .ZN(n9702) );
  NAND2_X1 U12287 ( .A1(n9704), .A2(n9703), .ZN(n9705) );
  NAND2_X1 U12288 ( .A1(n9924), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9706) );
  XNOR2_X1 U12289 ( .A(n9722), .B(P1_REG3_REG_20__SCAN_IN), .ZN(n14886) );
  NAND2_X1 U12290 ( .A1(n14886), .A2(n6445), .ZN(n9712) );
  INV_X1 U12291 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9709) );
  NAND2_X1 U12292 ( .A1(n9920), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9708) );
  NAND2_X1 U12293 ( .A1(n9927), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9707) );
  OAI211_X1 U12294 ( .C1(n9709), .C2(n9930), .A(n9708), .B(n9707), .ZN(n9710)
         );
  INV_X1 U12295 ( .A(n9710), .ZN(n9711) );
  OAI22_X1 U12296 ( .A1(n15071), .A2(n9745), .B1(n14869), .B2(n9801), .ZN(
        n9713) );
  XNOR2_X1 U12297 ( .A(n9713), .B(n12425), .ZN(n9715) );
  NOR2_X1 U12298 ( .A1(n14869), .A2(n9800), .ZN(n9714) );
  AOI21_X1 U12299 ( .B1(n14702), .B2(n12422), .A(n9714), .ZN(n9716) );
  XNOR2_X1 U12300 ( .A(n9715), .B(n9716), .ZN(n12382) );
  INV_X1 U12301 ( .A(n9715), .ZN(n9717) );
  OR2_X1 U12302 ( .A1(n9717), .A2(n9716), .ZN(n9718) );
  NAND2_X1 U12303 ( .A1(n11707), .A2(n9461), .ZN(n9720) );
  NAND2_X1 U12304 ( .A1(n9924), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9719) );
  NAND2_X2 U12305 ( .A1(n9720), .A2(n9719), .ZN(n15066) );
  INV_X1 U12306 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n12384) );
  INV_X1 U12307 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9721) );
  OAI21_X1 U12308 ( .B1(n9722), .B2(n12384), .A(n9721), .ZN(n9723) );
  AND2_X1 U12309 ( .A1(n9723), .A2(n9737), .ZN(n14873) );
  NAND2_X1 U12310 ( .A1(n14873), .A2(n6445), .ZN(n9729) );
  INV_X1 U12311 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9726) );
  NAND2_X1 U12312 ( .A1(n9927), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9725) );
  NAND2_X1 U12313 ( .A1(n9920), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9724) );
  OAI211_X1 U12314 ( .C1(n9930), .C2(n9726), .A(n9725), .B(n9724), .ZN(n9727)
         );
  INV_X1 U12315 ( .A(n9727), .ZN(n9728) );
  NAND2_X1 U12316 ( .A1(n9729), .A2(n9728), .ZN(n14855) );
  AOI22_X1 U12317 ( .A1(n15066), .A2(n12427), .B1(n12422), .B2(n14855), .ZN(
        n9730) );
  XNOR2_X1 U12318 ( .A(n9730), .B(n12425), .ZN(n9732) );
  AOI22_X1 U12319 ( .A1(n15066), .A2(n12422), .B1(n9434), .B2(n14855), .ZN(
        n9731) );
  XNOR2_X1 U12320 ( .A(n9732), .B(n9731), .ZN(n14407) );
  NAND2_X1 U12321 ( .A1(n9732), .A2(n9731), .ZN(n9733) );
  NAND2_X1 U12322 ( .A1(n9734), .A2(n10339), .ZN(n9735) );
  XNOR2_X1 U12323 ( .A(n9735), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15177) );
  INV_X1 U12324 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n15766) );
  NAND2_X1 U12325 ( .A1(n9737), .A2(n15766), .ZN(n9738) );
  AND2_X1 U12326 ( .A1(n9756), .A2(n9738), .ZN(n14857) );
  NAND2_X1 U12327 ( .A1(n14857), .A2(n6445), .ZN(n9744) );
  INV_X1 U12328 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9741) );
  NAND2_X1 U12329 ( .A1(n9927), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9740) );
  NAND2_X1 U12330 ( .A1(n9920), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9739) );
  OAI211_X1 U12331 ( .C1(n9741), .C2(n9930), .A(n9740), .B(n9739), .ZN(n9742)
         );
  INV_X1 U12332 ( .A(n9742), .ZN(n9743) );
  OAI22_X1 U12333 ( .A1(n15058), .A2(n9745), .B1(n14870), .B2(n9801), .ZN(
        n9746) );
  XNOR2_X1 U12334 ( .A(n9746), .B(n12425), .ZN(n9748) );
  NOR2_X1 U12335 ( .A1(n14870), .A2(n9800), .ZN(n9747) );
  AOI21_X1 U12336 ( .B1(n14854), .B2(n12422), .A(n9747), .ZN(n9749) );
  XNOR2_X1 U12337 ( .A(n9748), .B(n9749), .ZN(n14461) );
  INV_X1 U12338 ( .A(n9748), .ZN(n9750) );
  NAND2_X1 U12339 ( .A1(n9750), .A2(n9749), .ZN(n9751) );
  NAND2_X1 U12340 ( .A1(n11860), .A2(n9461), .ZN(n9753) );
  NAND2_X1 U12341 ( .A1(n9924), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9752) );
  INV_X1 U12342 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9755) );
  NAND2_X1 U12343 ( .A1(n9756), .A2(n9755), .ZN(n9757) );
  NAND2_X1 U12344 ( .A1(n9773), .A2(n9757), .ZN(n14836) );
  INV_X1 U12345 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n15763) );
  NAND2_X1 U12346 ( .A1(n9919), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n9759) );
  NAND2_X1 U12347 ( .A1(n9920), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9758) );
  OAI211_X1 U12348 ( .C1(n9353), .C2(n15763), .A(n9759), .B(n9758), .ZN(n9760)
         );
  INV_X1 U12349 ( .A(n9760), .ZN(n9761) );
  INV_X1 U12350 ( .A(n14856), .ZN(n14811) );
  OAI22_X1 U12351 ( .A1(n14833), .A2(n9801), .B1(n14811), .B2(n9800), .ZN(
        n9767) );
  NAND2_X1 U12352 ( .A1(n15051), .A2(n12427), .ZN(n9764) );
  NAND2_X1 U12353 ( .A1(n14856), .A2(n12422), .ZN(n9763) );
  NAND2_X1 U12354 ( .A1(n9764), .A2(n9763), .ZN(n9765) );
  XNOR2_X1 U12355 ( .A(n9765), .B(n12425), .ZN(n9766) );
  XOR2_X1 U12356 ( .A(n9767), .B(n9766), .Z(n14390) );
  INV_X1 U12357 ( .A(n9766), .ZN(n9769) );
  INV_X1 U12358 ( .A(n9767), .ZN(n9768) );
  NAND2_X1 U12359 ( .A1(n9769), .A2(n9768), .ZN(n12396) );
  NAND2_X1 U12360 ( .A1(n12114), .A2(n9461), .ZN(n9771) );
  NAND2_X1 U12361 ( .A1(n9924), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9770) );
  INV_X1 U12362 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9772) );
  NAND2_X1 U12363 ( .A1(n9773), .A2(n9772), .ZN(n9774) );
  AND2_X1 U12364 ( .A1(n9792), .A2(n9774), .ZN(n14820) );
  NAND2_X1 U12365 ( .A1(n14820), .A2(n6445), .ZN(n9780) );
  INV_X1 U12366 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9777) );
  NAND2_X1 U12367 ( .A1(n9920), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9776) );
  NAND2_X1 U12368 ( .A1(n9927), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9775) );
  OAI211_X1 U12369 ( .C1(n9777), .C2(n9930), .A(n9776), .B(n9775), .ZN(n9778)
         );
  INV_X1 U12370 ( .A(n9778), .ZN(n9779) );
  OAI22_X1 U12371 ( .A1(n14822), .A2(n9801), .B1(n14798), .B2(n9800), .ZN(
        n9785) );
  NAND2_X1 U12372 ( .A1(n15046), .A2(n12427), .ZN(n9782) );
  NAND2_X1 U12373 ( .A1(n14830), .A2(n12422), .ZN(n9781) );
  NAND2_X1 U12374 ( .A1(n9782), .A2(n9781), .ZN(n9783) );
  XNOR2_X1 U12375 ( .A(n9783), .B(n12425), .ZN(n9784) );
  XOR2_X1 U12376 ( .A(n9785), .B(n9784), .Z(n14445) );
  NAND2_X1 U12377 ( .A1(n14444), .A2(n14445), .ZN(n9788) );
  INV_X1 U12378 ( .A(n9784), .ZN(n9787) );
  INV_X1 U12379 ( .A(n9785), .ZN(n9786) );
  NAND2_X1 U12380 ( .A1(n9787), .A2(n9786), .ZN(n12392) );
  NAND2_X1 U12381 ( .A1(n9788), .A2(n12392), .ZN(n9806) );
  NAND2_X1 U12382 ( .A1(n14371), .A2(n9461), .ZN(n9790) );
  NAND2_X1 U12383 ( .A1(n9924), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9789) );
  INV_X1 U12384 ( .A(n14795), .ZN(n15040) );
  INV_X1 U12385 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9791) );
  NAND2_X1 U12386 ( .A1(n9792), .A2(n9791), .ZN(n9793) );
  NAND2_X1 U12387 ( .A1(n9835), .A2(n9793), .ZN(n14801) );
  INV_X1 U12388 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9796) );
  NAND2_X1 U12389 ( .A1(n9920), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9795) );
  NAND2_X1 U12390 ( .A1(n9927), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9794) );
  OAI211_X1 U12391 ( .C1(n9796), .C2(n9930), .A(n9795), .B(n9794), .ZN(n9797)
         );
  INV_X1 U12392 ( .A(n9797), .ZN(n9798) );
  OAI22_X1 U12393 ( .A1(n15040), .A2(n9801), .B1(n14812), .B2(n9800), .ZN(
        n12389) );
  NAND2_X1 U12394 ( .A1(n14795), .A2(n12427), .ZN(n9803) );
  NAND2_X1 U12395 ( .A1(n14711), .A2(n12422), .ZN(n9802) );
  NAND2_X1 U12396 ( .A1(n9803), .A2(n9802), .ZN(n9804) );
  XNOR2_X1 U12397 ( .A(n9804), .B(n12425), .ZN(n12388) );
  XOR2_X1 U12398 ( .A(n12388), .B(n12389), .Z(n12399) );
  INV_X1 U12399 ( .A(n12399), .ZN(n9805) );
  NAND2_X1 U12400 ( .A1(n15173), .A2(P1_B_REG_SCAN_IN), .ZN(n9807) );
  MUX2_X1 U12401 ( .A(n9807), .B(P1_B_REG_SCAN_IN), .S(n9810), .Z(n9809) );
  INV_X1 U12402 ( .A(n15171), .ZN(n9808) );
  INV_X1 U12403 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10395) );
  NAND2_X1 U12404 ( .A1(n10391), .A2(n10395), .ZN(n9811) );
  INV_X1 U12405 ( .A(n9810), .ZN(n12116) );
  NAND2_X1 U12406 ( .A1(n12116), .A2(n15171), .ZN(n10393) );
  INV_X1 U12407 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10399) );
  NAND2_X1 U12408 ( .A1(n10391), .A2(n10399), .ZN(n9812) );
  NAND2_X1 U12409 ( .A1(n15173), .A2(n15171), .ZN(n10396) );
  NAND2_X1 U12410 ( .A1(n9812), .A2(n10396), .ZN(n11045) );
  OR2_X1 U12411 ( .A1(n15005), .A2(n11045), .ZN(n9844) );
  NOR4_X1 U12412 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n9816) );
  NOR4_X1 U12413 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n9815) );
  NOR4_X1 U12414 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n9814) );
  NOR4_X1 U12415 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n9813) );
  AND4_X1 U12416 ( .A1(n9816), .A2(n9815), .A3(n9814), .A4(n9813), .ZN(n9821)
         );
  NOR2_X1 U12417 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .ZN(
        n15687) );
  NOR4_X1 U12418 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n9819) );
  NOR4_X1 U12419 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n9818) );
  NOR4_X1 U12420 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n9817) );
  AND4_X1 U12421 ( .A1(n15687), .A2(n9819), .A3(n9818), .A4(n9817), .ZN(n9820)
         );
  NAND2_X1 U12422 ( .A1(n9821), .A2(n9820), .ZN(n9822) );
  NAND2_X1 U12423 ( .A1(n10391), .A2(n9822), .ZN(n9843) );
  INV_X1 U12424 ( .A(n9843), .ZN(n9823) );
  INV_X1 U12425 ( .A(n9829), .ZN(n9828) );
  NAND2_X1 U12426 ( .A1(n9824), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9825) );
  XNOR2_X1 U12427 ( .A(n9825), .B(n6907), .ZN(n10404) );
  NAND2_X1 U12428 ( .A1(n15176), .A2(n10987), .ZN(n10406) );
  AND2_X1 U12429 ( .A1(n14817), .A2(n11513), .ZN(n9831) );
  INV_X1 U12430 ( .A(n9831), .ZN(n9826) );
  NAND3_X1 U12431 ( .A1(n9826), .A2(n11050), .A3(n11710), .ZN(n15406) );
  AND3_X1 U12432 ( .A1(n10971), .A2(n10406), .A3(n15406), .ZN(n9827) );
  NAND2_X1 U12433 ( .A1(n9829), .A2(n11044), .ZN(n9833) );
  AND2_X1 U12434 ( .A1(n10971), .A2(n15418), .ZN(n9830) );
  OAI211_X1 U12435 ( .C1(n9831), .C2(n10406), .A(n10296), .B(n10404), .ZN(
        n9842) );
  INV_X1 U12436 ( .A(n9842), .ZN(n9832) );
  NAND2_X1 U12437 ( .A1(n9833), .A2(n9832), .ZN(n10658) );
  INV_X1 U12438 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9834) );
  NAND2_X1 U12439 ( .A1(n9835), .A2(n9834), .ZN(n9836) );
  NAND2_X1 U12440 ( .A1(n14782), .A2(n6445), .ZN(n9841) );
  INV_X1 U12441 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n15794) );
  NAND2_X1 U12442 ( .A1(n9920), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9838) );
  NAND2_X1 U12443 ( .A1(n9927), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9837) );
  OAI211_X1 U12444 ( .C1(n15794), .C2(n9930), .A(n9838), .B(n9837), .ZN(n9839)
         );
  INV_X1 U12445 ( .A(n9839), .ZN(n9840) );
  NOR2_X1 U12446 ( .A1(n9842), .A2(P1_U3086), .ZN(n9975) );
  NAND2_X1 U12447 ( .A1(n9843), .A2(n9975), .ZN(n11046) );
  INV_X1 U12448 ( .A(n10406), .ZN(n9845) );
  NAND2_X1 U12449 ( .A1(n14491), .A2(n14903), .ZN(n14482) );
  INV_X1 U12450 ( .A(n14482), .ZN(n14473) );
  NAND2_X1 U12451 ( .A1(n14800), .A2(n14473), .ZN(n9847) );
  INV_X1 U12452 ( .A(n15167), .ZN(n10511) );
  AOI22_X1 U12453 ( .A1(n14830), .A2(n14478), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9846) );
  OAI211_X1 U12454 ( .C1(n14494), .C2(n14801), .A(n9847), .B(n9846), .ZN(n9848) );
  AOI21_X1 U12455 ( .B1(n14795), .B2(n14496), .A(n9848), .ZN(n9849) );
  MUX2_X1 U12456 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n10338), .Z(n9854) );
  INV_X1 U12457 ( .A(SI_31_), .ZN(n9853) );
  XNOR2_X1 U12458 ( .A(n9854), .B(n9853), .ZN(n9859) );
  MUX2_X1 U12459 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n10338), .Z(n9855) );
  NAND2_X1 U12460 ( .A1(n9855), .A2(SI_30_), .ZN(n9914) );
  NAND2_X1 U12461 ( .A1(n9859), .A2(n9914), .ZN(n9865) );
  INV_X1 U12462 ( .A(n9855), .ZN(n9856) );
  INV_X1 U12463 ( .A(SI_30_), .ZN(n12460) );
  NAND2_X1 U12464 ( .A1(n9856), .A2(n12460), .ZN(n9913) );
  INV_X1 U12465 ( .A(SI_29_), .ZN(n13240) );
  NAND2_X1 U12466 ( .A1(n9857), .A2(n13240), .ZN(n9911) );
  NAND2_X1 U12467 ( .A1(n9913), .A2(n9911), .ZN(n9861) );
  NOR2_X1 U12468 ( .A1(n9861), .A2(n9859), .ZN(n9858) );
  NAND2_X1 U12469 ( .A1(n9912), .A2(n9858), .ZN(n9864) );
  INV_X1 U12470 ( .A(n9859), .ZN(n9862) );
  XNOR2_X1 U12471 ( .A(n9859), .B(n9914), .ZN(n9860) );
  OAI21_X1 U12472 ( .B1(n9862), .B2(n9861), .A(n9860), .ZN(n9863) );
  NAND2_X1 U12473 ( .A1(n14355), .A2(n9461), .ZN(n9867) );
  NAND2_X1 U12474 ( .A1(n9924), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n9866) );
  NAND2_X1 U12475 ( .A1(n9919), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n9870) );
  NAND2_X1 U12476 ( .A1(n9920), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9869) );
  NAND2_X1 U12477 ( .A1(n9927), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9868) );
  NAND3_X1 U12478 ( .A1(n9870), .A2(n9869), .A3(n9868), .ZN(n14653) );
  XNOR2_X1 U12479 ( .A(n9939), .B(n14653), .ZN(n9963) );
  NAND2_X1 U12480 ( .A1(n9924), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9871) );
  INV_X1 U12481 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9873) );
  NAND2_X1 U12482 ( .A1(n9874), .A2(n9873), .ZN(n9875) );
  INV_X1 U12483 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9879) );
  NAND2_X1 U12484 ( .A1(n9444), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9878) );
  NAND2_X1 U12485 ( .A1(n9927), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9877) );
  OAI211_X1 U12486 ( .C1(n9879), .C2(n9930), .A(n9878), .B(n9877), .ZN(n9880)
         );
  INV_X1 U12487 ( .A(n9880), .ZN(n9881) );
  XNOR2_X2 U12488 ( .A(n15027), .B(n14741), .ZN(n14772) );
  NAND2_X1 U12489 ( .A1(n9924), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9882) );
  XNOR2_X1 U12490 ( .A(n14731), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n12433) );
  NAND2_X1 U12491 ( .A1(n12433), .A2(n6445), .ZN(n9889) );
  INV_X1 U12492 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n14743) );
  NAND2_X1 U12493 ( .A1(n9919), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n9885) );
  NAND2_X1 U12494 ( .A1(n9927), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n9884) );
  OAI211_X1 U12495 ( .C1(n9886), .C2(n14743), .A(n9885), .B(n9884), .ZN(n9887)
         );
  INV_X1 U12496 ( .A(n9887), .ZN(n9888) );
  XNOR2_X1 U12497 ( .A(n15046), .B(n14798), .ZN(n14818) );
  XNOR2_X1 U12498 ( .A(n15051), .B(n14856), .ZN(n14829) );
  INV_X1 U12499 ( .A(n14829), .ZN(n14842) );
  NAND2_X1 U12500 ( .A1(n14854), .A2(n14870), .ZN(n14681) );
  NAND2_X1 U12501 ( .A1(n15058), .A2(n14831), .ZN(n9890) );
  NAND2_X1 U12502 ( .A1(n14681), .A2(n9890), .ZN(n14849) );
  INV_X1 U12503 ( .A(n14849), .ZN(n14852) );
  XNOR2_X1 U12504 ( .A(n14702), .B(n14869), .ZN(n14884) );
  OR2_X1 U12505 ( .A1(n15076), .A2(n14922), .ZN(n10073) );
  NAND2_X1 U12506 ( .A1(n15076), .A2(n14922), .ZN(n14678) );
  NAND2_X1 U12507 ( .A1(n10073), .A2(n14678), .ZN(n14697) );
  INV_X1 U12508 ( .A(n14697), .ZN(n14901) );
  NOR2_X1 U12509 ( .A1(n15088), .A2(n14500), .ZN(n14694) );
  NAND2_X1 U12510 ( .A1(n15088), .A2(n14500), .ZN(n14695) );
  OR2_X1 U12511 ( .A1(n14694), .A2(n6926), .ZN(n14928) );
  NAND2_X1 U12512 ( .A1(n15107), .A2(n14981), .ZN(n14665) );
  INV_X1 U12513 ( .A(n12031), .ZN(n12034) );
  OR2_X1 U12514 ( .A1(n11073), .A2(n14994), .ZN(n9984) );
  NAND2_X1 U12515 ( .A1(n9984), .A2(n10992), .ZN(n14991) );
  NOR2_X1 U12516 ( .A1(n14991), .A2(n7190), .ZN(n9893) );
  NAND2_X1 U12517 ( .A1(n15356), .A2(n14510), .ZN(n10995) );
  NAND2_X1 U12518 ( .A1(n10996), .A2(n10995), .ZN(n10979) );
  INV_X1 U12519 ( .A(n10979), .ZN(n11308) );
  INV_X1 U12520 ( .A(n9892), .ZN(n14511) );
  NAND2_X1 U12521 ( .A1(n14511), .A2(n9891), .ZN(n9996) );
  NAND2_X1 U12522 ( .A1(n9892), .A2(n10657), .ZN(n10994) );
  NAND4_X1 U12523 ( .A1(n9893), .A2(n11308), .A3(n11362), .A4(n11102), .ZN(
        n9894) );
  XNOR2_X1 U12524 ( .A(n11250), .B(n14507), .ZN(n11248) );
  XNOR2_X1 U12525 ( .A(n15373), .B(n14508), .ZN(n15320) );
  NOR3_X1 U12526 ( .A1(n9894), .A2(n11248), .A3(n15320), .ZN(n9897) );
  XNOR2_X1 U12527 ( .A(n11987), .B(n11832), .ZN(n15289) );
  XNOR2_X1 U12528 ( .A(n15397), .B(n11983), .ZN(n11829) );
  NOR2_X1 U12529 ( .A1(n15289), .A2(n11829), .ZN(n9896) );
  AND2_X1 U12530 ( .A1(n15417), .A2(n11981), .ZN(n12009) );
  INV_X1 U12531 ( .A(n12009), .ZN(n9895) );
  NAND2_X1 U12532 ( .A1(n12046), .A2(n9895), .ZN(n12026) );
  INV_X1 U12533 ( .A(n12026), .ZN(n11833) );
  XNOR2_X1 U12534 ( .A(n15389), .B(n14506), .ZN(n15304) );
  NAND4_X1 U12535 ( .A1(n9897), .A2(n9896), .A3(n11833), .A4(n15304), .ZN(
        n9898) );
  XNOR2_X1 U12536 ( .A(n15126), .B(n12071), .ZN(n12045) );
  NOR2_X1 U12537 ( .A1(n9898), .A2(n12045), .ZN(n9899) );
  XNOR2_X1 U12538 ( .A(n15121), .B(n14983), .ZN(n12063) );
  XNOR2_X1 U12539 ( .A(n15116), .B(n14661), .ZN(n12030) );
  NAND4_X1 U12540 ( .A1(n12034), .A2(n9899), .A3(n12063), .A4(n7695), .ZN(
        n9901) );
  INV_X1 U12541 ( .A(n15103), .ZN(n14966) );
  INV_X1 U12542 ( .A(n14669), .ZN(n9900) );
  NAND2_X1 U12543 ( .A1(n14943), .A2(n9900), .ZN(n14959) );
  NOR2_X1 U12544 ( .A1(n9901), .A2(n14959), .ZN(n9902) );
  AND2_X1 U12545 ( .A1(n14928), .A2(n9902), .ZN(n9903) );
  XNOR2_X1 U12546 ( .A(n14692), .B(n14932), .ZN(n14944) );
  XNOR2_X1 U12547 ( .A(n15083), .B(n14902), .ZN(n14919) );
  NAND4_X1 U12548 ( .A1(n14901), .A2(n9903), .A3(n6927), .A4(n14919), .ZN(
        n9904) );
  NOR2_X1 U12549 ( .A1(n14884), .A2(n9904), .ZN(n9905) );
  XNOR2_X1 U12550 ( .A(n15066), .B(n14855), .ZN(n14867) );
  NAND3_X1 U12551 ( .A1(n14852), .A2(n9905), .A3(n14867), .ZN(n9906) );
  NOR3_X1 U12552 ( .A1(n14818), .A2(n14842), .A3(n9906), .ZN(n9910) );
  XNOR2_X1 U12553 ( .A(n14795), .B(n14812), .ZN(n14793) );
  INV_X1 U12554 ( .A(n14793), .ZN(n14790) );
  NAND2_X1 U12555 ( .A1(n9924), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9908) );
  NAND2_X4 U12556 ( .A1(n9909), .A2(n9908), .ZN(n15033) );
  AND2_X1 U12557 ( .A1(n9914), .A2(n9913), .ZN(n9915) );
  NAND2_X1 U12558 ( .A1(n12454), .A2(n9461), .ZN(n9918) );
  NAND2_X1 U12559 ( .A1(n9924), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9917) );
  NAND2_X1 U12560 ( .A1(n9919), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n9923) );
  NAND2_X1 U12561 ( .A1(n9920), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9922) );
  NAND2_X1 U12562 ( .A1(n9927), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9921) );
  NAND3_X1 U12563 ( .A1(n9923), .A2(n9922), .A3(n9921), .ZN(n14727) );
  XNOR2_X1 U12564 ( .A(n14656), .B(n14727), .ZN(n9935) );
  NAND2_X1 U12565 ( .A1(n9924), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n9925) );
  NAND2_X1 U12566 ( .A1(n6445), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9926) );
  OR2_X1 U12567 ( .A1(n14731), .A2(n9926), .ZN(n9934) );
  INV_X1 U12568 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9931) );
  NAND2_X1 U12569 ( .A1(n9444), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9929) );
  NAND2_X1 U12570 ( .A1(n9927), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9928) );
  OAI211_X1 U12571 ( .C1(n9931), .C2(n9930), .A(n9929), .B(n9928), .ZN(n9932)
         );
  INV_X1 U12572 ( .A(n9932), .ZN(n9933) );
  NAND3_X1 U12573 ( .A1(n9936), .A2(n9935), .A3(n14717), .ZN(n9937) );
  XNOR2_X1 U12574 ( .A(n9937), .B(n14817), .ZN(n9938) );
  INV_X1 U12575 ( .A(n11513), .ZN(n10986) );
  NAND2_X1 U12576 ( .A1(n11710), .A2(n10986), .ZN(n9947) );
  NOR2_X1 U12577 ( .A1(n9938), .A2(n9947), .ZN(n9954) );
  NAND2_X1 U12578 ( .A1(n9940), .A2(n11050), .ZN(n9941) );
  OR2_X1 U12579 ( .A1(n9939), .A2(n10124), .ZN(n9970) );
  INV_X1 U12580 ( .A(n9970), .ZN(n9945) );
  INV_X1 U12581 ( .A(n9942), .ZN(n11049) );
  NAND2_X1 U12582 ( .A1(n11049), .A2(n10406), .ZN(n9944) );
  NAND2_X1 U12583 ( .A1(n9943), .A2(n9940), .ZN(n11067) );
  AND2_X1 U12584 ( .A1(n9944), .A2(n11067), .ZN(n9962) );
  INV_X1 U12585 ( .A(n9962), .ZN(n9948) );
  INV_X1 U12586 ( .A(n14653), .ZN(n9969) );
  INV_X1 U12587 ( .A(n9947), .ZN(n11000) );
  NOR4_X1 U12588 ( .A1(n9946), .A2(n9969), .A3(n11000), .A4(n9939), .ZN(n9953)
         );
  NAND2_X1 U12589 ( .A1(n9939), .A2(n9955), .ZN(n9966) );
  NOR3_X1 U12590 ( .A1(n9966), .A2(n14653), .A3(n9948), .ZN(n9952) );
  INV_X1 U12591 ( .A(n9966), .ZN(n9950) );
  AND2_X1 U12592 ( .A1(n9948), .A2(n9947), .ZN(n9968) );
  INV_X1 U12593 ( .A(n9968), .ZN(n9949) );
  NOR4_X1 U12594 ( .A1(n9950), .A2(n15004), .A3(n14653), .A4(n9949), .ZN(n9951) );
  OR2_X1 U12595 ( .A1(n10404), .A2(P1_U3086), .ZN(n10133) );
  OAI21_X1 U12596 ( .B1(n14653), .B2(n11513), .A(n14727), .ZN(n9956) );
  MUX2_X1 U12597 ( .A(n9956), .B(n15009), .S(n10124), .Z(n9965) );
  INV_X1 U12598 ( .A(n9965), .ZN(n9961) );
  NAND2_X1 U12599 ( .A1(n14656), .A2(n10082), .ZN(n9959) );
  OAI22_X1 U12600 ( .A1(n10082), .A2(n9969), .B1(n10987), .B2(n6667), .ZN(
        n9957) );
  NAND2_X1 U12601 ( .A1(n9957), .A2(n14727), .ZN(n9958) );
  NAND2_X1 U12602 ( .A1(n9959), .A2(n9958), .ZN(n9964) );
  INV_X1 U12603 ( .A(n9964), .ZN(n9960) );
  NOR2_X1 U12604 ( .A1(n9961), .A2(n9960), .ZN(n10135) );
  INV_X1 U12605 ( .A(n10135), .ZN(n9972) );
  NAND2_X1 U12606 ( .A1(n9963), .A2(n9962), .ZN(n10131) );
  NOR2_X1 U12607 ( .A1(n9965), .A2(n9964), .ZN(n10132) );
  INV_X1 U12608 ( .A(n10132), .ZN(n9971) );
  OR2_X1 U12609 ( .A1(n9966), .A2(n14653), .ZN(n9967) );
  OAI211_X1 U12610 ( .C1(n9970), .C2(n9969), .A(n9968), .B(n9967), .ZN(n10134)
         );
  OAI22_X1 U12611 ( .A1(n9972), .A2(n10131), .B1(n9971), .B2(n10134), .ZN(
        n9973) );
  INV_X1 U12612 ( .A(n10133), .ZN(n11837) );
  NAND2_X1 U12613 ( .A1(n9973), .A2(n11837), .ZN(n9978) );
  INV_X1 U12614 ( .A(n14651), .ZN(n9974) );
  NAND3_X1 U12615 ( .A1(n9975), .A2(n9974), .A3(n14982), .ZN(n9976) );
  OAI211_X1 U12616 ( .C1(n15176), .C2(n10133), .A(n9976), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9977) );
  OAI211_X1 U12617 ( .C1(n9979), .C2(n10133), .A(n9978), .B(n9977), .ZN(n9980)
         );
  INV_X1 U12618 ( .A(n9980), .ZN(n10137) );
  MUX2_X1 U12619 ( .A(n14726), .B(n14740), .S(n10124), .Z(n10130) );
  MUX2_X1 U12620 ( .A(n11104), .B(n14509), .S(n10002), .Z(n10003) );
  OR2_X1 U12621 ( .A1(n10996), .A2(n9955), .ZN(n10000) );
  INV_X1 U12622 ( .A(n10995), .ZN(n9981) );
  NAND2_X1 U12623 ( .A1(n9981), .A2(n9955), .ZN(n9999) );
  AND4_X1 U12624 ( .A1(n10000), .A2(n10657), .A3(n14511), .A4(n9999), .ZN(
        n9995) );
  NAND3_X1 U12625 ( .A1(n10996), .A2(n10085), .A3(n9891), .ZN(n9983) );
  NAND3_X1 U12626 ( .A1(n10995), .A2(n9892), .A3(n9955), .ZN(n9982) );
  NAND2_X1 U12627 ( .A1(n9983), .A2(n9982), .ZN(n9994) );
  NAND2_X1 U12628 ( .A1(n10992), .A2(n10973), .ZN(n9985) );
  NAND2_X1 U12629 ( .A1(n9985), .A2(n9984), .ZN(n9987) );
  INV_X1 U12630 ( .A(n10992), .ZN(n9986) );
  MUX2_X1 U12631 ( .A(n9987), .B(n9986), .S(n9955), .Z(n9988) );
  INV_X1 U12632 ( .A(n7190), .ZN(n11072) );
  NAND2_X1 U12633 ( .A1(n9988), .A2(n11072), .ZN(n9992) );
  NAND2_X1 U12634 ( .A1(n10085), .A2(n6441), .ZN(n9990) );
  NAND2_X1 U12635 ( .A1(n9955), .A2(n15341), .ZN(n9989) );
  NAND2_X1 U12636 ( .A1(n9992), .A2(n9991), .ZN(n9993) );
  NAND2_X1 U12637 ( .A1(n9996), .A2(n10085), .ZN(n9997) );
  OR2_X1 U12638 ( .A1(n10979), .A2(n9997), .ZN(n10001) );
  NAND3_X1 U12639 ( .A1(n10996), .A2(n10994), .A3(n9955), .ZN(n9998) );
  INV_X1 U12640 ( .A(n15373), .ZN(n11153) );
  MUX2_X1 U12641 ( .A(n11153), .B(n14508), .S(n10124), .Z(n10007) );
  MUX2_X1 U12642 ( .A(n11153), .B(n14508), .S(n10085), .Z(n10004) );
  NAND2_X1 U12643 ( .A1(n10005), .A2(n10004), .ZN(n10011) );
  INV_X1 U12644 ( .A(n10006), .ZN(n10009) );
  NAND2_X1 U12645 ( .A1(n10009), .A2(n10008), .ZN(n10010) );
  MUX2_X1 U12646 ( .A(n14507), .B(n15380), .S(n9955), .Z(n10014) );
  NAND2_X1 U12647 ( .A1(n10015), .A2(n10014), .ZN(n10013) );
  MUX2_X1 U12648 ( .A(n15380), .B(n14507), .S(n10124), .Z(n10012) );
  NAND2_X1 U12649 ( .A1(n10013), .A2(n10012), .ZN(n10017) );
  MUX2_X1 U12650 ( .A(n14506), .B(n15389), .S(n10085), .Z(n10019) );
  MUX2_X1 U12651 ( .A(n15389), .B(n14506), .S(n10085), .Z(n10018) );
  INV_X1 U12652 ( .A(n10019), .ZN(n10020) );
  INV_X1 U12653 ( .A(n11983), .ZN(n14505) );
  MUX2_X1 U12654 ( .A(n15397), .B(n14505), .S(n10002), .Z(n10022) );
  INV_X1 U12655 ( .A(n15397), .ZN(n11242) );
  MUX2_X1 U12656 ( .A(n11983), .B(n11242), .S(n10002), .Z(n10021) );
  MUX2_X1 U12657 ( .A(n11981), .B(n11824), .S(n10002), .Z(n10040) );
  MUX2_X1 U12658 ( .A(n14503), .B(n15417), .S(n10124), .Z(n10033) );
  INV_X1 U12659 ( .A(n11987), .ZN(n15407) );
  MUX2_X1 U12660 ( .A(n11832), .B(n15407), .S(n10085), .Z(n10030) );
  INV_X1 U12661 ( .A(n11832), .ZN(n14504) );
  MUX2_X1 U12662 ( .A(n11987), .B(n14504), .S(n10002), .Z(n10029) );
  AOI22_X1 U12663 ( .A1(n10040), .A2(n10033), .B1(n10030), .B2(n10029), .ZN(
        n10023) );
  MUX2_X1 U12664 ( .A(n14661), .B(n14977), .S(n10002), .Z(n10044) );
  INV_X1 U12665 ( .A(n10044), .ZN(n10026) );
  NOR2_X1 U12666 ( .A1(n14661), .A2(n10124), .ZN(n10024) );
  AOI21_X1 U12667 ( .B1(n15116), .B2(n9955), .A(n10024), .ZN(n10025) );
  AND2_X1 U12668 ( .A1(n10026), .A2(n10025), .ZN(n10027) );
  MUX2_X1 U12669 ( .A(n12013), .B(n7770), .S(n10124), .Z(n10052) );
  MUX2_X1 U12670 ( .A(n14983), .B(n15121), .S(n10085), .Z(n10051) );
  NAND2_X1 U12671 ( .A1(n10052), .A2(n10051), .ZN(n10028) );
  NAND2_X1 U12672 ( .A1(n10055), .A2(n10028), .ZN(n10050) );
  INV_X1 U12673 ( .A(n10029), .ZN(n10032) );
  INV_X1 U12674 ( .A(n10030), .ZN(n10031) );
  AND2_X1 U12675 ( .A1(n10032), .A2(n10031), .ZN(n10036) );
  INV_X1 U12676 ( .A(n10036), .ZN(n10039) );
  MUX2_X1 U12677 ( .A(n12071), .B(n7772), .S(n10124), .Z(n10049) );
  MUX2_X1 U12678 ( .A(n14502), .B(n15126), .S(n10085), .Z(n10048) );
  NAND2_X1 U12679 ( .A1(n10049), .A2(n10048), .ZN(n10038) );
  INV_X1 U12680 ( .A(n10040), .ZN(n10035) );
  INV_X1 U12681 ( .A(n10033), .ZN(n10034) );
  OAI21_X1 U12682 ( .B1(n10036), .B2(n10035), .A(n10034), .ZN(n10037) );
  OAI211_X1 U12683 ( .C1(n10040), .C2(n10039), .A(n10038), .B(n10037), .ZN(
        n10041) );
  NOR2_X1 U12684 ( .A1(n10050), .A2(n10041), .ZN(n10061) );
  INV_X1 U12685 ( .A(n14666), .ZN(n10042) );
  OR2_X1 U12686 ( .A1(n14671), .A2(n10042), .ZN(n10047) );
  INV_X1 U12687 ( .A(n14661), .ZN(n14501) );
  MUX2_X1 U12688 ( .A(n14501), .B(n15116), .S(n10124), .Z(n10043) );
  NAND2_X1 U12689 ( .A1(n10044), .A2(n10043), .ZN(n10045) );
  NOR2_X1 U12690 ( .A1(n10045), .A2(n12031), .ZN(n10046) );
  AOI21_X1 U12691 ( .B1(n10047), .B2(n10082), .A(n10046), .ZN(n10060) );
  OR3_X1 U12692 ( .A1(n10050), .A2(n10049), .A3(n10048), .ZN(n10059) );
  INV_X1 U12693 ( .A(n10051), .ZN(n10054) );
  INV_X1 U12694 ( .A(n10052), .ZN(n10053) );
  NAND3_X1 U12695 ( .A1(n10055), .A2(n10054), .A3(n10053), .ZN(n10058) );
  INV_X1 U12696 ( .A(n14665), .ZN(n10056) );
  OAI21_X1 U12697 ( .B1(n14669), .B2(n10056), .A(n10124), .ZN(n10057) );
  MUX2_X1 U12698 ( .A(n14669), .B(n14671), .S(n10124), .Z(n10062) );
  MUX2_X1 U12699 ( .A(n14691), .B(n14692), .S(n10082), .Z(n10064) );
  MUX2_X1 U12700 ( .A(n14932), .B(n15095), .S(n10124), .Z(n10063) );
  AOI21_X1 U12701 ( .B1(n10065), .B2(n10064), .A(n10063), .ZN(n10072) );
  NOR2_X1 U12702 ( .A1(n10065), .A2(n10064), .ZN(n10071) );
  NAND2_X1 U12703 ( .A1(n15088), .A2(n9955), .ZN(n10066) );
  OAI21_X1 U12704 ( .B1(n14921), .B2(n9955), .A(n10066), .ZN(n10067) );
  NOR2_X1 U12705 ( .A1(n14694), .A2(n10067), .ZN(n10068) );
  NOR2_X1 U12706 ( .A1(n14697), .A2(n10068), .ZN(n10069) );
  MUX2_X1 U12707 ( .A(n14678), .B(n10073), .S(n10082), .Z(n10080) );
  MUX2_X1 U12708 ( .A(n14500), .B(n15088), .S(n10124), .Z(n10074) );
  NAND3_X1 U12709 ( .A1(n14919), .A2(n10074), .A3(n14695), .ZN(n10077) );
  INV_X1 U12710 ( .A(n14902), .ZN(n14933) );
  NAND3_X1 U12711 ( .A1(n15083), .A2(n14933), .A3(n9955), .ZN(n10076) );
  OR3_X1 U12712 ( .A1(n15083), .A2(n14933), .A3(n9955), .ZN(n10075) );
  NAND3_X1 U12713 ( .A1(n10077), .A2(n10076), .A3(n10075), .ZN(n10078) );
  NAND2_X1 U12714 ( .A1(n10078), .A2(n14901), .ZN(n10079) );
  NAND3_X1 U12715 ( .A1(n10081), .A2(n10080), .A3(n10079), .ZN(n10088) );
  NAND2_X1 U12716 ( .A1(n10088), .A2(n10087), .ZN(n10090) );
  MUX2_X1 U12717 ( .A(n14702), .B(n14904), .S(n10082), .Z(n10086) );
  OAI21_X1 U12718 ( .B1(n10088), .B2(n10087), .A(n10086), .ZN(n10089) );
  MUX2_X1 U12719 ( .A(n14855), .B(n15066), .S(n10124), .Z(n10093) );
  MUX2_X1 U12720 ( .A(n14855), .B(n15066), .S(n10082), .Z(n10091) );
  MUX2_X1 U12721 ( .A(n14854), .B(n14831), .S(n10124), .Z(n10095) );
  MUX2_X1 U12722 ( .A(n14854), .B(n14831), .S(n10082), .Z(n10094) );
  MUX2_X1 U12723 ( .A(n15051), .B(n14856), .S(n10082), .Z(n10099) );
  MUX2_X1 U12724 ( .A(n15051), .B(n14856), .S(n10124), .Z(n10096) );
  NAND2_X1 U12725 ( .A1(n10097), .A2(n10096), .ZN(n10103) );
  INV_X1 U12726 ( .A(n10098), .ZN(n10101) );
  INV_X1 U12727 ( .A(n10099), .ZN(n10100) );
  NAND2_X1 U12728 ( .A1(n10101), .A2(n10100), .ZN(n10102) );
  MUX2_X1 U12729 ( .A(n14830), .B(n15046), .S(n10082), .Z(n10105) );
  MUX2_X1 U12730 ( .A(n15046), .B(n14830), .S(n10082), .Z(n10104) );
  INV_X1 U12731 ( .A(n10105), .ZN(n10106) );
  MUX2_X1 U12732 ( .A(n14711), .B(n14795), .S(n10124), .Z(n10109) );
  MUX2_X1 U12733 ( .A(n14711), .B(n14795), .S(n10082), .Z(n10107) );
  MUX2_X1 U12734 ( .A(n14800), .B(n15033), .S(n10082), .Z(n10111) );
  MUX2_X1 U12735 ( .A(n15033), .B(n14800), .S(n10082), .Z(n10110) );
  INV_X1 U12736 ( .A(n10111), .ZN(n10112) );
  MUX2_X1 U12737 ( .A(n14741), .B(n15027), .S(n10124), .Z(n10116) );
  NAND2_X1 U12738 ( .A1(n10115), .A2(n10116), .ZN(n10114) );
  MUX2_X1 U12739 ( .A(n14741), .B(n15027), .S(n10082), .Z(n10113) );
  NAND2_X1 U12740 ( .A1(n10114), .A2(n10113), .ZN(n10120) );
  INV_X1 U12741 ( .A(n10115), .ZN(n10118) );
  INV_X1 U12742 ( .A(n10116), .ZN(n10117) );
  NAND2_X1 U12743 ( .A1(n10118), .A2(n10117), .ZN(n10119) );
  MUX2_X1 U12744 ( .A(n14758), .B(n14748), .S(n10082), .Z(n10122) );
  MUX2_X1 U12745 ( .A(n14758), .B(n14748), .S(n10124), .Z(n10121) );
  INV_X1 U12746 ( .A(n10122), .ZN(n10123) );
  MUX2_X1 U12747 ( .A(n14740), .B(n14726), .S(n10124), .Z(n10126) );
  NAND2_X1 U12748 ( .A1(n10125), .A2(n10126), .ZN(n10129) );
  INV_X1 U12749 ( .A(n10125), .ZN(n10128) );
  INV_X1 U12750 ( .A(n10126), .ZN(n10127) );
  INV_X1 U12751 ( .A(n10230), .ZN(n11854) );
  NAND2_X1 U12752 ( .A1(n7438), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10138) );
  NAND2_X1 U12753 ( .A1(n10440), .A2(n10138), .ZN(n10140) );
  NAND2_X1 U12754 ( .A1(n10139), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10141) );
  NAND2_X1 U12755 ( .A1(n10140), .A2(n10141), .ZN(n10948) );
  XNOR2_X1 U12756 ( .A(n10947), .B(n10203), .ZN(n10938) );
  NAND2_X1 U12757 ( .A1(n10937), .A2(n10938), .ZN(n10936) );
  NAND2_X1 U12758 ( .A1(n10947), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10142) );
  NAND2_X1 U12759 ( .A1(n10936), .A2(n10142), .ZN(n10143) );
  NAND2_X1 U12760 ( .A1(n10143), .A2(n10423), .ZN(n10815) );
  XNOR2_X1 U12761 ( .A(n10436), .B(n11529), .ZN(n10814) );
  NAND2_X1 U12762 ( .A1(n10436), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n10145) );
  NAND2_X1 U12763 ( .A1(n10818), .A2(n10145), .ZN(n10146) );
  OR2_X1 U12764 ( .A1(n10218), .A2(n11518), .ZN(n10149) );
  NAND2_X1 U12765 ( .A1(n10218), .A2(n11518), .ZN(n10148) );
  AND2_X1 U12766 ( .A1(n10149), .A2(n10148), .ZN(n11084) );
  AOI22_X1 U12767 ( .A1(n11035), .A2(P3_REG2_REG_7__SCAN_IN), .B1(n10433), 
        .B2(n7437), .ZN(n11195) );
  XNOR2_X1 U12768 ( .A(n10428), .B(P3_REG2_REG_8__SCAN_IN), .ZN(n11196) );
  INV_X1 U12769 ( .A(n11466), .ZN(n10222) );
  INV_X1 U12770 ( .A(n10150), .ZN(n11609) );
  XNOR2_X1 U12771 ( .A(n11607), .B(P3_REG2_REG_10__SCAN_IN), .ZN(n11610) );
  INV_X1 U12772 ( .A(n10354), .ZN(n11783) );
  INV_X1 U12773 ( .A(n10152), .ZN(n11840) );
  XNOR2_X1 U12774 ( .A(n10230), .B(n10153), .ZN(n11841) );
  OR2_X1 U12775 ( .A1(n10560), .A2(n12970), .ZN(n10236) );
  NAND2_X1 U12776 ( .A1(n10560), .A2(n12970), .ZN(n10155) );
  AND2_X1 U12777 ( .A1(n10236), .A2(n10155), .ZN(n12665) );
  NAND2_X1 U12778 ( .A1(n12663), .A2(n10236), .ZN(n10156) );
  INV_X1 U12779 ( .A(n10156), .ZN(n10158) );
  INV_X1 U12780 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12688) );
  INV_X1 U12781 ( .A(n10159), .ZN(n12710) );
  XNOR2_X1 U12782 ( .A(n12722), .B(P3_REG2_REG_16__SCAN_IN), .ZN(n12709) );
  INV_X1 U12783 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n10240) );
  NAND2_X1 U12784 ( .A1(n12726), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n12743) );
  INV_X1 U12785 ( .A(n12752), .ZN(n10637) );
  NAND2_X1 U12786 ( .A1(n10637), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n10163) );
  INV_X1 U12787 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12919) );
  NAND2_X1 U12788 ( .A1(n12752), .A2(n12919), .ZN(n10162) );
  NAND2_X1 U12789 ( .A1(n10163), .A2(n10162), .ZN(n12742) );
  INV_X1 U12790 ( .A(n10163), .ZN(n10164) );
  XNOR2_X1 U12791 ( .A(n12357), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n10199) );
  INV_X1 U12792 ( .A(n10828), .ZN(n10165) );
  OR2_X1 U12793 ( .A1(n12267), .A2(n10165), .ZN(n10167) );
  NAND2_X1 U12794 ( .A1(n10167), .A2(n10166), .ZN(n10196) );
  NOR2_X1 U12795 ( .A1(n10828), .A2(P3_U3151), .ZN(n12363) );
  INV_X1 U12796 ( .A(n12363), .ZN(n12367) );
  NAND2_X1 U12797 ( .A1(n10840), .A2(n12367), .ZN(n10195) );
  INV_X1 U12798 ( .A(n10195), .ZN(n10168) );
  NOR2_X1 U12799 ( .A1(n10196), .A2(n10168), .ZN(n10171) );
  INV_X1 U12800 ( .A(n10171), .ZN(n10170) );
  NOR2_X2 U12801 ( .A1(n10170), .A2(n10169), .ZN(n12744) );
  MUX2_X1 U12802 ( .A(P3_U3897), .B(n10171), .S(n13243), .Z(n12751) );
  NAND2_X1 U12803 ( .A1(n10171), .A2(n13246), .ZN(n12750) );
  INV_X1 U12804 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13095) );
  XNOR2_X1 U12805 ( .A(n12722), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n12705) );
  INV_X1 U12806 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13103) );
  OR2_X1 U12807 ( .A1(n10560), .A2(n13103), .ZN(n10235) );
  INV_X1 U12808 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n13112) );
  AOI22_X1 U12809 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n11854), .B1(n10230), 
        .B2(n13112), .ZN(n11847) );
  INV_X1 U12810 ( .A(n10218), .ZN(n11086) );
  NAND2_X1 U12811 ( .A1(n10440), .A2(n10174), .ZN(n10175) );
  NAND2_X1 U12812 ( .A1(n10175), .A2(n6486), .ZN(n10956) );
  INV_X1 U12813 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10955) );
  NAND2_X1 U12814 ( .A1(n10931), .A2(n10930), .ZN(n10929) );
  NAND2_X1 U12815 ( .A1(n10947), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10176) );
  NAND2_X1 U12816 ( .A1(n10929), .A2(n10176), .ZN(n10177) );
  INV_X1 U12817 ( .A(n10423), .ZN(n10801) );
  XNOR2_X1 U12818 ( .A(n10801), .B(n10177), .ZN(n10794) );
  NAND2_X1 U12819 ( .A1(n10794), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n10179) );
  NAND2_X1 U12820 ( .A1(n10177), .A2(n10423), .ZN(n10178) );
  INV_X1 U12821 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10180) );
  MUX2_X1 U12822 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n10180), .S(n10436), .Z(
        n10810) );
  INV_X1 U12823 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15672) );
  MUX2_X1 U12824 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n15672), .S(n10218), .Z(
        n11088) );
  INV_X1 U12825 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n10181) );
  INV_X1 U12826 ( .A(n10428), .ZN(n11198) );
  XNOR2_X1 U12827 ( .A(n11198), .B(P3_REG1_REG_8__SCAN_IN), .ZN(n11191) );
  INV_X1 U12828 ( .A(n10182), .ZN(n10183) );
  XOR2_X1 U12829 ( .A(P3_REG1_REG_10__SCAN_IN), .B(n11607), .Z(n11599) );
  INV_X1 U12830 ( .A(n11599), .ZN(n10186) );
  INV_X1 U12831 ( .A(n11607), .ZN(n10185) );
  INV_X1 U12832 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n10184) );
  NAND2_X1 U12833 ( .A1(n10354), .A2(n10187), .ZN(n10188) );
  NAND2_X1 U12834 ( .A1(n6841), .A2(n10189), .ZN(n10190) );
  NAND2_X1 U12835 ( .A1(n10560), .A2(n13103), .ZN(n10191) );
  AND2_X1 U12836 ( .A1(n10235), .A2(n10191), .ZN(n12671) );
  NAND2_X1 U12837 ( .A1(n10501), .A2(n10192), .ZN(n10193) );
  INV_X1 U12838 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13089) );
  XNOR2_X1 U12839 ( .A(n12752), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n12748) );
  AOI22_X1 U12840 ( .A1(n12747), .A2(n12748), .B1(P3_REG1_REG_18__SCAN_IN), 
        .B2(n10637), .ZN(n10194) );
  XNOR2_X1 U12841 ( .A(n12357), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n10200) );
  NAND2_X1 U12842 ( .A1(n15581), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n10197) );
  NAND2_X1 U12843 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12526)
         );
  MUX2_X1 U12844 ( .A(n10200), .B(n10199), .S(n10198), .Z(n10245) );
  MUX2_X1 U12845 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13246), .Z(n10242) );
  INV_X1 U12846 ( .A(n10436), .ZN(n10825) );
  MUX2_X1 U12847 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n13246), .Z(n10212) );
  INV_X1 U12848 ( .A(n10212), .ZN(n10213) );
  NAND2_X1 U12849 ( .A1(n10201), .A2(n10440), .ZN(n10202) );
  OAI21_X1 U12850 ( .B1(n10201), .B2(n10440), .A(n10202), .ZN(n10952) );
  MUX2_X1 U12851 ( .A(n8822), .B(n15725), .S(n13246), .Z(n11143) );
  NAND2_X1 U12852 ( .A1(n11143), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11148) );
  NOR2_X1 U12853 ( .A1(n10952), .A2(n11148), .ZN(n10951) );
  INV_X1 U12854 ( .A(n10202), .ZN(n10932) );
  MUX2_X1 U12855 ( .A(n10203), .B(n10173), .S(n13246), .Z(n10205) );
  INV_X1 U12856 ( .A(n10947), .ZN(n10204) );
  NAND2_X1 U12857 ( .A1(n10205), .A2(n10204), .ZN(n10803) );
  INV_X1 U12858 ( .A(n10205), .ZN(n10206) );
  NAND2_X1 U12859 ( .A1(n10206), .A2(n10947), .ZN(n10207) );
  AND2_X1 U12860 ( .A1(n10803), .A2(n10207), .ZN(n10933) );
  INV_X1 U12861 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10793) );
  MUX2_X1 U12862 ( .A(n11453), .B(n10793), .S(n13246), .Z(n10208) );
  NAND2_X1 U12863 ( .A1(n10208), .A2(n10801), .ZN(n10211) );
  INV_X1 U12864 ( .A(n10208), .ZN(n10209) );
  NAND2_X1 U12865 ( .A1(n10209), .A2(n10423), .ZN(n10210) );
  NAND2_X1 U12866 ( .A1(n10211), .A2(n10210), .ZN(n10802) );
  XNOR2_X1 U12867 ( .A(n10212), .B(n10436), .ZN(n10808) );
  INV_X1 U12868 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10214) );
  MUX2_X1 U12869 ( .A(n11539), .B(n10214), .S(n13246), .Z(n10215) );
  NOR2_X1 U12870 ( .A1(n10215), .A2(n6979), .ZN(n11121) );
  NAND2_X1 U12871 ( .A1(n10215), .A2(n6979), .ZN(n11119) );
  OAI21_X1 U12872 ( .B1(n11123), .B2(n11121), .A(n11119), .ZN(n11081) );
  MUX2_X1 U12873 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n13246), .Z(n10216) );
  XNOR2_X1 U12874 ( .A(n10216), .B(n10218), .ZN(n11082) );
  INV_X1 U12875 ( .A(n10216), .ZN(n10217) );
  MUX2_X1 U12876 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n13246), .Z(n10219) );
  XNOR2_X1 U12877 ( .A(n10219), .B(n10433), .ZN(n11033) );
  MUX2_X1 U12878 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n13246), .Z(n10220) );
  XOR2_X1 U12879 ( .A(n10428), .B(n10220), .Z(n11192) );
  INV_X1 U12880 ( .A(n10220), .ZN(n10221) );
  MUX2_X1 U12881 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n13246), .Z(n10224) );
  INV_X1 U12882 ( .A(n10224), .ZN(n10223) );
  NAND2_X1 U12883 ( .A1(n10223), .A2(n10222), .ZN(n11459) );
  MUX2_X1 U12884 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n13246), .Z(n10225) );
  NOR2_X1 U12885 ( .A1(n10225), .A2(n11607), .ZN(n10226) );
  AOI21_X1 U12886 ( .B1(n10225), .B2(n11607), .A(n10226), .ZN(n11603) );
  INV_X1 U12887 ( .A(n10226), .ZN(n10227) );
  NAND2_X1 U12888 ( .A1(n11601), .A2(n10227), .ZN(n11782) );
  MUX2_X1 U12889 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13246), .Z(n10228) );
  XNOR2_X1 U12890 ( .A(n10228), .B(n11783), .ZN(n11781) );
  INV_X1 U12891 ( .A(n10228), .ZN(n10229) );
  NAND2_X1 U12892 ( .A1(n10229), .A2(n11783), .ZN(n11848) );
  MUX2_X1 U12893 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n13246), .Z(n10231) );
  XNOR2_X1 U12894 ( .A(n10231), .B(n10230), .ZN(n11850) );
  NAND2_X1 U12895 ( .A1(n10231), .A2(n11854), .ZN(n12652) );
  MUX2_X1 U12896 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13246), .Z(n10232) );
  XNOR2_X1 U12897 ( .A(n10232), .B(n10233), .ZN(n12651) );
  INV_X1 U12898 ( .A(n10232), .ZN(n10234) );
  NAND2_X1 U12899 ( .A1(n10234), .A2(n10233), .ZN(n12672) );
  MUX2_X1 U12900 ( .A(n12665), .B(n12671), .S(n13246), .Z(n12676) );
  MUX2_X1 U12901 ( .A(n10236), .B(n10235), .S(n13246), .Z(n10237) );
  INV_X1 U12902 ( .A(n10238), .ZN(n10239) );
  XNOR2_X1 U12903 ( .A(n10238), .B(n10501), .ZN(n12697) );
  MUX2_X1 U12904 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n13246), .Z(n12696) );
  MUX2_X1 U12905 ( .A(n10240), .B(n13095), .S(n13246), .Z(n10241) );
  NOR2_X1 U12906 ( .A1(n10241), .A2(n12722), .ZN(n12716) );
  XNOR2_X1 U12907 ( .A(n10242), .B(n10565), .ZN(n12733) );
  XNOR2_X1 U12908 ( .A(n10243), .B(n12752), .ZN(n12740) );
  MUX2_X1 U12909 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n13246), .Z(n12741) );
  NOR2_X1 U12910 ( .A1(n12740), .A2(n12741), .ZN(n12739) );
  AOI21_X1 U12911 ( .B1(n10243), .B2(n12752), .A(n12739), .ZN(n10244) );
  XOR2_X1 U12912 ( .A(n10245), .B(n10244), .Z(n10246) );
  NAND2_X1 U12913 ( .A1(n12647), .A2(n13243), .ZN(n12755) );
  NOR2_X1 U12914 ( .A1(n10246), .A2(n12755), .ZN(n10247) );
  INV_X1 U12915 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12455) );
  INV_X1 U12916 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n10249) );
  OR2_X1 U12917 ( .A1(n7177), .A2(n10249), .ZN(n10251) );
  INV_X1 U12918 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n10261) );
  NAND2_X1 U12919 ( .A1(n8111), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n10256) );
  INV_X1 U12920 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n10253) );
  OR2_X1 U12921 ( .A1(n10254), .A2(n10253), .ZN(n10255) );
  OAI211_X1 U12922 ( .C1(n8131), .C2(n10261), .A(n10256), .B(n10255), .ZN(
        n13807) );
  AND2_X1 U12923 ( .A1(n13807), .A2(n10257), .ZN(n14204) );
  NOR2_X1 U12924 ( .A1(n13939), .A2(n14204), .ZN(n10260) );
  NAND2_X1 U12925 ( .A1(n15571), .A2(n15525), .ZN(n14350) );
  NAND2_X1 U12926 ( .A1(n13718), .A2(n10258), .ZN(n10259) );
  MUX2_X1 U12927 ( .A(n10261), .B(n10260), .S(n15580), .Z(n10263) );
  NAND2_X1 U12928 ( .A1(n15580), .A2(n15525), .ZN(n14294) );
  NAND2_X1 U12929 ( .A1(n10263), .A2(n10262), .ZN(P2_U3530) );
  OAI21_X1 U12930 ( .B1(n10265), .B2(n10264), .A(n13786), .ZN(n10266) );
  NOR2_X1 U12931 ( .A1(n10268), .A2(n15493), .ZN(n10269) );
  NOR2_X1 U12932 ( .A1(n10269), .A2(n7943), .ZN(n10270) );
  INV_X1 U12933 ( .A(n10292), .ZN(n10273) );
  INV_X1 U12934 ( .A(n10271), .ZN(n10272) );
  AND2_X1 U12935 ( .A1(n13969), .A2(n14271), .ZN(n10276) );
  INV_X1 U12936 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n10280) );
  XNOR2_X1 U12937 ( .A(n10281), .B(n10283), .ZN(n13981) );
  INV_X1 U12938 ( .A(n10282), .ZN(n10284) );
  NAND2_X1 U12939 ( .A1(n14004), .A2(n14188), .ZN(n10286) );
  NAND2_X1 U12940 ( .A1(n13974), .A2(n13988), .ZN(n10290) );
  NAND2_X1 U12941 ( .A1(n10290), .A2(n14181), .ZN(n10291) );
  OR2_X1 U12942 ( .A1(n10292), .A2(n10291), .ZN(n13977) );
  INV_X1 U12943 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n10293) );
  INV_X1 U12944 ( .A(n10397), .ZN(n10297) );
  OR2_X2 U12945 ( .A1(n10297), .A2(n10296), .ZN(n14525) );
  INV_X1 U12946 ( .A(n10298), .ZN(n10299) );
  OR2_X2 U12947 ( .A1(n10578), .A2(n10299), .ZN(n13830) );
  INV_X1 U12948 ( .A(n13830), .ZN(P2_U3947) );
  NOR2_X1 U12949 ( .A1(n10902), .A2(n10301), .ZN(n10305) );
  XNOR2_X1 U12950 ( .A(n10303), .B(n10302), .ZN(n10304) );
  XNOR2_X1 U12951 ( .A(n10305), .B(n10304), .ZN(n10306) );
  NOR2_X1 U12952 ( .A1(n10306), .A2(n14498), .ZN(n10311) );
  NOR2_X1 U12953 ( .A1(n14494), .A2(n11002), .ZN(n10310) );
  AND2_X1 U12954 ( .A1(n14496), .A2(n11104), .ZN(n10309) );
  INV_X1 U12955 ( .A(n14508), .ZN(n11099) );
  NAND2_X1 U12956 ( .A1(n14478), .A2(n14510), .ZN(n10307) );
  NAND2_X1 U12957 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n15284) );
  OAI211_X1 U12958 ( .C1(n11099), .C2(n14482), .A(n10307), .B(n15284), .ZN(
        n10308) );
  OR4_X1 U12959 ( .A1(n10311), .A2(n10310), .A3(n10309), .A4(n10308), .ZN(
        P1_U3230) );
  NAND2_X1 U12960 ( .A1(n10338), .A2(P2_U3088), .ZN(n14367) );
  AND2_X1 U12961 ( .A1(n10339), .A2(P2_U3088), .ZN(n14359) );
  OAI222_X1 U12962 ( .A1(n13851), .A2(P2_U3088), .B1(n14367), .B2(n10320), 
        .C1(n10313), .C2(n14372), .ZN(P2_U3325) );
  OAI222_X1 U12963 ( .A1(n13838), .A2(P2_U3088), .B1(n14367), .B2(n10343), 
        .C1(n10314), .C2(n14372), .ZN(P2_U3326) );
  OAI222_X1 U12964 ( .A1(n15452), .A2(P2_U3088), .B1(n14367), .B2(n10323), 
        .C1(n10315), .C2(n14372), .ZN(P2_U3324) );
  OAI222_X1 U12965 ( .A1(n13861), .A2(P2_U3088), .B1(n14367), .B2(n10318), 
        .C1(n10316), .C2(n14372), .ZN(P2_U3323) );
  AND2_X1 U12966 ( .A1(n10338), .A2(P1_U3086), .ZN(n15155) );
  INV_X2 U12967 ( .A(n15155), .ZN(n15164) );
  OAI222_X1 U12968 ( .A1(n15271), .A2(P1_U3086), .B1(n15169), .B2(n10318), 
        .C1(n10317), .C2(n15164), .ZN(P1_U3351) );
  INV_X1 U12969 ( .A(n14537), .ZN(n10321) );
  OAI222_X1 U12970 ( .A1(n10321), .A2(P1_U3086), .B1(n15169), .B2(n10320), 
        .C1(n10319), .C2(n15164), .ZN(P1_U3353) );
  OAI222_X1 U12971 ( .A1(n14553), .A2(P1_U3086), .B1(n15169), .B2(n10323), 
        .C1(n10322), .C2(n15164), .ZN(P1_U3352) );
  NAND2_X1 U12972 ( .A1(n12154), .A2(P3_D_REG_0__SCAN_IN), .ZN(n10324) );
  OAI21_X1 U12973 ( .B1(n10848), .B2(n12154), .A(n10324), .ZN(P3_U3376) );
  INV_X1 U12974 ( .A(n10325), .ZN(n10328) );
  OAI222_X1 U12975 ( .A1(n10471), .A2(P1_U3086), .B1(n15169), .B2(n10328), 
        .C1(n10326), .C2(n15164), .ZN(P1_U3350) );
  OAI222_X1 U12976 ( .A1(n10680), .A2(P2_U3088), .B1(n14367), .B2(n10328), 
        .C1(n10327), .C2(n14372), .ZN(P2_U3322) );
  INV_X1 U12977 ( .A(n10329), .ZN(n10332) );
  OAI222_X1 U12978 ( .A1(n10495), .A2(P1_U3086), .B1(n15169), .B2(n10332), 
        .C1(n10330), .C2(n15164), .ZN(P1_U3349) );
  OAI222_X1 U12979 ( .A1(n15464), .A2(P2_U3088), .B1(n14367), .B2(n10332), 
        .C1(n10331), .C2(n14372), .ZN(P2_U3321) );
  INV_X1 U12980 ( .A(n10627), .ZN(n10573) );
  INV_X1 U12981 ( .A(n10333), .ZN(n10336) );
  INV_X2 U12982 ( .A(n14359), .ZN(n14372) );
  OAI222_X1 U12983 ( .A1(n10573), .A2(P2_U3088), .B1(n14367), .B2(n10336), 
        .C1(n10334), .C2(n14372), .ZN(P2_U3319) );
  INV_X1 U12984 ( .A(n10524), .ZN(n10337) );
  OAI222_X1 U12985 ( .A1(n10337), .A2(P1_U3086), .B1(n15169), .B2(n10336), 
        .C1(n10335), .C2(n15164), .ZN(P1_U3347) );
  NAND2_X1 U12986 ( .A1(n10338), .A2(P3_U3151), .ZN(n13256) );
  NAND2_X1 U12987 ( .A1(n10339), .A2(P3_U3151), .ZN(n13248) );
  OAI222_X1 U12988 ( .A1(n13256), .A2(n10341), .B1(n13248), .B2(n10340), .C1(
        P3_U3151), .C2(n11466), .ZN(P3_U3286) );
  INV_X1 U12989 ( .A(n14517), .ZN(n10344) );
  OAI222_X1 U12990 ( .A1(n10344), .A2(P1_U3086), .B1(n15169), .B2(n10343), 
        .C1(n10342), .C2(n15164), .ZN(P1_U3354) );
  INV_X1 U12991 ( .A(n10345), .ZN(n10348) );
  OAI222_X1 U12992 ( .A1(n10540), .A2(P1_U3086), .B1(n15169), .B2(n10348), 
        .C1(n10346), .C2(n15164), .ZN(P1_U3348) );
  INV_X1 U12993 ( .A(n10612), .ZN(n10623) );
  OAI222_X1 U12994 ( .A1(n10623), .A2(P2_U3088), .B1(n14367), .B2(n10348), 
        .C1(n10347), .C2(n14372), .ZN(P2_U3320) );
  INV_X1 U12995 ( .A(n10720), .ZN(n10607) );
  INV_X1 U12996 ( .A(n10349), .ZN(n10352) );
  OAI222_X1 U12997 ( .A1(n10607), .A2(P2_U3088), .B1(n14367), .B2(n10352), 
        .C1(n10350), .C2(n14372), .ZN(P2_U3318) );
  INV_X1 U12998 ( .A(n10644), .ZN(n10353) );
  OAI222_X1 U12999 ( .A1(n10353), .A2(P1_U3086), .B1(n15169), .B2(n10352), 
        .C1(n10351), .C2(n15164), .ZN(P1_U3346) );
  OAI222_X1 U13000 ( .A1(n13256), .A2(n10356), .B1(n13248), .B2(n10355), .C1(
        P3_U3151), .C2(n10354), .ZN(P3_U3284) );
  NAND2_X1 U13001 ( .A1(n10365), .A2(n10366), .ZN(n10358) );
  NAND2_X1 U13002 ( .A1(n14513), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n10357) );
  NAND2_X1 U13003 ( .A1(n14531), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n10359) );
  NAND2_X1 U13004 ( .A1(n10361), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n10362) );
  INV_X1 U13005 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n10364) );
  XNOR2_X1 U13006 ( .A(n10382), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n10381) );
  INV_X1 U13007 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n13858) );
  XNOR2_X1 U13008 ( .A(n10381), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15840) );
  INV_X1 U13009 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n11140) );
  AOI21_X1 U13010 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n11140), .A(n10365), .ZN(
        n15842) );
  INV_X1 U13011 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15841) );
  NOR2_X1 U13012 ( .A1(n15842), .A2(n15841), .ZN(n15848) );
  XNOR2_X1 U13013 ( .A(n10366), .B(n10365), .ZN(n10367) );
  NAND2_X1 U13014 ( .A1(n15848), .A2(n15847), .ZN(n10369) );
  NAND2_X1 U13015 ( .A1(n10367), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n10368) );
  NAND2_X1 U13016 ( .A1(n10369), .A2(n10368), .ZN(n10372) );
  XNOR2_X1 U13017 ( .A(n10370), .B(n10371), .ZN(n10373) );
  NAND2_X1 U13018 ( .A1(n10372), .A2(n10373), .ZN(n15261) );
  INV_X1 U13019 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n15731) );
  NAND2_X1 U13020 ( .A1(n15261), .A2(n15731), .ZN(n10376) );
  INV_X1 U13021 ( .A(n10372), .ZN(n10375) );
  INV_X1 U13022 ( .A(n10373), .ZN(n10374) );
  NAND2_X1 U13023 ( .A1(n10375), .A2(n10374), .ZN(n15262) );
  NAND2_X1 U13024 ( .A1(n10376), .A2(n15262), .ZN(n15843) );
  INV_X1 U13025 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15845) );
  NAND2_X1 U13026 ( .A1(n15843), .A2(n15845), .ZN(n10378) );
  XNOR2_X1 U13027 ( .A(n10377), .B(n14546), .ZN(n15844) );
  NAND2_X1 U13028 ( .A1(n10378), .A2(n15844), .ZN(n10380) );
  OR2_X1 U13029 ( .A1(n15843), .A2(n15845), .ZN(n10379) );
  NAND2_X1 U13030 ( .A1(n10380), .A2(n10379), .ZN(n15839) );
  INV_X1 U13031 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n15286) );
  NAND2_X1 U13032 ( .A1(n10382), .A2(n15286), .ZN(n10385) );
  NAND2_X1 U13033 ( .A1(n10383), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n10384) );
  INV_X1 U13034 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n10386) );
  INV_X1 U13035 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10387) );
  XNOR2_X1 U13036 ( .A(n10755), .B(n10387), .ZN(n10388) );
  NAND2_X1 U13037 ( .A1(n10389), .A2(n10388), .ZN(n10390) );
  OAI21_X1 U13038 ( .B1(n6675), .B2(n7457), .A(n10754), .ZN(SUB_1596_U58) );
  INV_X1 U13039 ( .A(n10391), .ZN(n10392) );
  INV_X1 U13040 ( .A(n10393), .ZN(n10394) );
  AOI22_X1 U13041 ( .A1(n15338), .A2(n10395), .B1(n10394), .B2(n10397), .ZN(
        P1_U3445) );
  INV_X1 U13042 ( .A(n10396), .ZN(n10398) );
  AOI22_X1 U13043 ( .A1(n15338), .A2(n10399), .B1(n10398), .B2(n10397), .ZN(
        P1_U3446) );
  INV_X1 U13044 ( .A(n10703), .ZN(n10653) );
  INV_X1 U13045 ( .A(n10400), .ZN(n10403) );
  OAI222_X1 U13046 ( .A1(n10653), .A2(P1_U3086), .B1(n15169), .B2(n10403), 
        .C1(n10401), .C2(n15164), .ZN(P1_U3345) );
  INV_X1 U13047 ( .A(n10723), .ZN(n10792) );
  OAI222_X1 U13048 ( .A1(n10792), .A2(P2_U3088), .B1(n14367), .B2(n10403), 
        .C1(n10402), .C2(n14372), .ZN(P2_U3317) );
  INV_X1 U13049 ( .A(n10404), .ZN(n10405) );
  OR2_X1 U13050 ( .A1(n10406), .A2(n10405), .ZN(n10408) );
  NAND2_X1 U13051 ( .A1(n10408), .A2(n7215), .ZN(n10455) );
  NAND2_X1 U13052 ( .A1(n10457), .A2(n10455), .ZN(n15287) );
  INV_X1 U13053 ( .A(n15287), .ZN(n14631) );
  NOR2_X1 U13054 ( .A1(n14631), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U13055 ( .A(n10409), .ZN(n10413) );
  INV_X1 U13056 ( .A(n11317), .ZN(n10410) );
  OAI222_X1 U13057 ( .A1(n15164), .A2(n10411), .B1(n15169), .B2(n10413), .C1(
        P1_U3086), .C2(n10410), .ZN(P1_U3344) );
  INV_X1 U13058 ( .A(n10917), .ZN(n10911) );
  OAI222_X1 U13059 ( .A1(n10911), .A2(P2_U3088), .B1(n14367), .B2(n10413), 
        .C1(n10412), .C2(n14372), .ZN(P2_U3316) );
  INV_X1 U13060 ( .A(n10414), .ZN(n10415) );
  OAI222_X1 U13061 ( .A1(n13256), .A2(n10416), .B1(n13248), .B2(n10415), .C1(
        P3_U3151), .C2(n11854), .ZN(P3_U3283) );
  INV_X1 U13062 ( .A(n13256), .ZN(n13234) );
  INV_X1 U13063 ( .A(n13234), .ZN(n13250) );
  INV_X1 U13064 ( .A(SI_6_), .ZN(n10418) );
  OAI222_X1 U13065 ( .A1(n13250), .A2(n10418), .B1(n13248), .B2(n10417), .C1(
        P3_U3151), .C2(n11086), .ZN(P3_U3289) );
  INV_X1 U13066 ( .A(n13248), .ZN(n11556) );
  AOI22_X1 U13067 ( .A1(n11556), .A2(n10419), .B1(P3_STATE_REG_SCAN_IN), .B2(
        P3_IR_REG_0__SCAN_IN), .ZN(n10420) );
  OAI21_X1 U13068 ( .B1(n10421), .B2(n13250), .A(n10420), .ZN(P3_U3295) );
  INV_X1 U13069 ( .A(n11556), .ZN(n13260) );
  OAI222_X1 U13070 ( .A1(n13260), .A2(n10424), .B1(n10423), .B2(P3_U3151), 
        .C1(n10422), .C2(n13256), .ZN(P3_U3292) );
  OAI222_X1 U13071 ( .A1(n13260), .A2(n10426), .B1(n11130), .B2(P3_U3151), 
        .C1(n10425), .C2(n13256), .ZN(P3_U3290) );
  OAI222_X1 U13072 ( .A1(n13260), .A2(n10429), .B1(n10428), .B2(P3_U3151), 
        .C1(n10427), .C2(n13256), .ZN(P3_U3287) );
  OAI222_X1 U13073 ( .A1(n13260), .A2(n10431), .B1(n10947), .B2(P3_U3151), 
        .C1(n10430), .C2(n13256), .ZN(P3_U3293) );
  INV_X1 U13074 ( .A(SI_7_), .ZN(n10432) );
  OAI222_X1 U13075 ( .A1(n13260), .A2(n10434), .B1(n10433), .B2(P3_U3151), 
        .C1(n10432), .C2(n13256), .ZN(P3_U3288) );
  OAI222_X1 U13076 ( .A1(n13260), .A2(n10437), .B1(n10436), .B2(P3_U3151), 
        .C1(n10435), .C2(n13256), .ZN(P3_U3291) );
  OAI222_X1 U13077 ( .A1(n13260), .A2(n10439), .B1(n11607), .B2(P3_U3151), 
        .C1(n10438), .C2(n13256), .ZN(P3_U3285) );
  INV_X1 U13078 ( .A(n10440), .ZN(n10963) );
  OAI222_X1 U13079 ( .A1(n13250), .A2(n8837), .B1(n10963), .B2(P3_U3151), .C1(
        n13260), .C2(n10441), .ZN(P3_U3294) );
  INV_X1 U13080 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n10443) );
  NAND2_X1 U13081 ( .A1(n13507), .A2(P2_U3947), .ZN(n10442) );
  OAI21_X1 U13082 ( .B1(P2_U3947), .B2(n10443), .A(n10442), .ZN(P2_U3531) );
  INV_X1 U13083 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10444) );
  MUX2_X1 U13084 ( .A(n10444), .B(P1_REG1_REG_8__SCAN_IN), .S(n10524), .Z(
        n10454) );
  INV_X1 U13085 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n15435) );
  INV_X1 U13086 ( .A(n10471), .ZN(n14563) );
  INV_X1 U13087 ( .A(n15271), .ZN(n15278) );
  INV_X1 U13088 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10445) );
  MUX2_X1 U13089 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10445), .S(n14537), .Z(
        n10448) );
  INV_X1 U13090 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10446) );
  AND2_X1 U13091 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14516) );
  NAND2_X1 U13092 ( .A1(n14517), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n14533) );
  NAND2_X1 U13093 ( .A1(n14534), .A2(n14533), .ZN(n10447) );
  NAND2_X1 U13094 ( .A1(n14537), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n14549) );
  NAND2_X1 U13095 ( .A1(n14551), .A2(n14549), .ZN(n10451) );
  INV_X1 U13096 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10449) );
  MUX2_X1 U13097 ( .A(n10449), .B(P1_REG1_REG_3__SCAN_IN), .S(n14553), .Z(
        n10450) );
  OR2_X1 U13098 ( .A1(n14553), .A2(n10449), .ZN(n15266) );
  INV_X1 U13099 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n15429) );
  MUX2_X1 U13100 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n15429), .S(n15271), .Z(
        n15265) );
  INV_X1 U13101 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n15431) );
  MUX2_X1 U13102 ( .A(n15431), .B(P1_REG1_REG_5__SCAN_IN), .S(n10471), .Z(
        n14566) );
  OAI21_X1 U13103 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n14563), .A(n14564), .ZN(
        n10497) );
  INV_X1 U13104 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n15433) );
  MUX2_X1 U13105 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n15433), .S(n10495), .Z(
        n10496) );
  NOR2_X1 U13106 ( .A1(n10495), .A2(n15433), .ZN(n10541) );
  MUX2_X1 U13107 ( .A(n15435), .B(P1_REG1_REG_7__SCAN_IN), .S(n10540), .Z(
        n10452) );
  AOI21_X1 U13108 ( .B1(n10454), .B2(n10453), .A(n10527), .ZN(n10483) );
  INV_X1 U13109 ( .A(n10455), .ZN(n10456) );
  AND2_X1 U13110 ( .A1(n10457), .A2(n10456), .ZN(n10515) );
  NAND2_X1 U13111 ( .A1(n10515), .A2(n14651), .ZN(n14645) );
  NAND2_X1 U13112 ( .A1(n10515), .A2(n15167), .ZN(n14644) );
  INV_X1 U13113 ( .A(n14644), .ZN(n15279) );
  INV_X1 U13114 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10458) );
  NAND2_X1 U13115 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11593) );
  OAI21_X1 U13116 ( .B1(n15287), .B2(n10458), .A(n11593), .ZN(n10459) );
  AOI21_X1 U13117 ( .B1(n15279), .B2(n10524), .A(n10459), .ZN(n10482) );
  INV_X1 U13118 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n14538) );
  MUX2_X1 U13119 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n14538), .S(n14537), .Z(
        n10464) );
  INV_X1 U13120 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10460) );
  MUX2_X1 U13121 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n10460), .S(n14517), .Z(
        n10462) );
  AND2_X1 U13122 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10461) );
  NAND2_X1 U13123 ( .A1(n10462), .A2(n10461), .ZN(n14540) );
  NAND2_X1 U13124 ( .A1(n14517), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n14539) );
  NAND2_X1 U13125 ( .A1(n14540), .A2(n14539), .ZN(n10463) );
  NAND2_X1 U13126 ( .A1(n10464), .A2(n10463), .ZN(n14556) );
  NAND2_X1 U13127 ( .A1(n14537), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14554) );
  NAND2_X1 U13128 ( .A1(n14556), .A2(n14554), .ZN(n10466) );
  INV_X1 U13129 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n11311) );
  MUX2_X1 U13130 ( .A(n11311), .B(P1_REG2_REG_3__SCAN_IN), .S(n14553), .Z(
        n10465) );
  OR2_X1 U13131 ( .A1(n14553), .A2(n11311), .ZN(n15273) );
  NAND2_X1 U13132 ( .A1(n15274), .A2(n15273), .ZN(n10469) );
  INV_X1 U13133 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10467) );
  MUX2_X1 U13134 ( .A(n10467), .B(P1_REG2_REG_4__SCAN_IN), .S(n15271), .Z(
        n10468) );
  NAND2_X1 U13135 ( .A1(n10469), .A2(n10468), .ZN(n15276) );
  NAND2_X1 U13136 ( .A1(n15278), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n14569) );
  INV_X1 U13137 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10470) );
  MUX2_X1 U13138 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10470), .S(n10471), .Z(
        n14570) );
  AOI21_X1 U13139 ( .B1(n15276), .B2(n14569), .A(n14570), .ZN(n14568) );
  NOR2_X1 U13140 ( .A1(n10471), .A2(n10470), .ZN(n10489) );
  INV_X1 U13141 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11112) );
  MUX2_X1 U13142 ( .A(n11112), .B(P1_REG2_REG_6__SCAN_IN), .S(n10495), .Z(
        n10472) );
  INV_X1 U13143 ( .A(n10495), .ZN(n10473) );
  NAND2_X1 U13144 ( .A1(n10473), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10535) );
  INV_X1 U13145 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10474) );
  MUX2_X1 U13146 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10474), .S(n10540), .Z(
        n10534) );
  AOI21_X1 U13147 ( .B1(n10536), .B2(n10535), .A(n10534), .ZN(n10550) );
  INV_X1 U13148 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11241) );
  MUX2_X1 U13149 ( .A(n11241), .B(P1_REG2_REG_8__SCAN_IN), .S(n10524), .Z(
        n10476) );
  NOR2_X1 U13150 ( .A1(n10540), .A2(n10474), .ZN(n10478) );
  INV_X1 U13151 ( .A(n10478), .ZN(n10475) );
  NAND2_X1 U13152 ( .A1(n10476), .A2(n10475), .ZN(n10480) );
  MUX2_X1 U13153 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n11241), .S(n10524), .Z(
        n10477) );
  NOR2_X1 U13154 ( .A1(n14651), .A2(n15167), .ZN(n10479) );
  OAI211_X1 U13155 ( .C1(n10550), .C2(n10480), .A(n10522), .B(n15277), .ZN(
        n10481) );
  OAI211_X1 U13156 ( .C1(n10483), .C2(n14645), .A(n10482), .B(n10481), .ZN(
        P1_U3251) );
  INV_X1 U13157 ( .A(n11258), .ZN(n11265) );
  INV_X1 U13158 ( .A(n14367), .ZN(n11859) );
  INV_X1 U13159 ( .A(n11859), .ZN(n14374) );
  INV_X1 U13160 ( .A(n10484), .ZN(n10486) );
  OAI222_X1 U13161 ( .A1(P2_U3088), .A2(n11265), .B1(n14372), .B2(n10485), 
        .C1(n14374), .C2(n10486), .ZN(P2_U3315) );
  INV_X1 U13162 ( .A(n14585), .ZN(n10488) );
  OAI222_X1 U13163 ( .A1(P1_U3086), .A2(n10488), .B1(n15164), .B2(n10487), 
        .C1(n15169), .C2(n10486), .ZN(P1_U3343) );
  MUX2_X1 U13164 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n11112), .S(n10495), .Z(
        n10491) );
  INV_X1 U13165 ( .A(n10489), .ZN(n10490) );
  NAND2_X1 U13166 ( .A1(n10491), .A2(n10490), .ZN(n10492) );
  OAI211_X1 U13167 ( .C1(n14568), .C2(n10492), .A(n15277), .B(n10536), .ZN(
        n10494) );
  NOR2_X1 U13168 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9392), .ZN(n11440) );
  AOI21_X1 U13169 ( .B1(n14631), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n11440), .ZN(
        n10493) );
  OAI211_X1 U13170 ( .C1(n14644), .C2(n10495), .A(n10494), .B(n10493), .ZN(
        n10499) );
  AOI211_X1 U13171 ( .C1(n10497), .C2(n10496), .A(n10546), .B(n14645), .ZN(
        n10498) );
  OR2_X1 U13172 ( .A1(n10499), .A2(n10498), .ZN(P1_U3249) );
  INV_X1 U13173 ( .A(n10500), .ZN(n10502) );
  OAI222_X1 U13174 ( .A1(n13250), .A2(n10503), .B1(n13248), .B2(n10502), .C1(
        P3_U3151), .C2(n10501), .ZN(P3_U3280) );
  INV_X1 U13175 ( .A(n10504), .ZN(n10506) );
  OAI222_X1 U13176 ( .A1(P2_U3088), .A2(n11268), .B1(n14372), .B2(n10505), 
        .C1(n14374), .C2(n10506), .ZN(P2_U3314) );
  INV_X1 U13177 ( .A(n11340), .ZN(n11333) );
  OAI222_X1 U13178 ( .A1(P1_U3086), .A2(n11333), .B1(n15164), .B2(n10507), 
        .C1(n15169), .C2(n10506), .ZN(P1_U3342) );
  INV_X1 U13179 ( .A(n10508), .ZN(n10509) );
  OAI222_X1 U13180 ( .A1(n13250), .A2(n10510), .B1(n6841), .B2(P3_U3151), .C1(
        n13260), .C2(n10509), .ZN(P3_U3282) );
  INV_X1 U13181 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10512) );
  NAND3_X1 U13182 ( .A1(n15270), .A2(P1_IR_REG_0__SCAN_IN), .A3(n10512), .ZN(
        n10517) );
  OAI21_X1 U13183 ( .B1(n14651), .B2(P1_REG2_REG_0__SCAN_IN), .A(n10511), .ZN(
        n14526) );
  AOI21_X1 U13184 ( .B1(n14651), .B2(n10512), .A(n14526), .ZN(n10513) );
  INV_X1 U13185 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14527) );
  MUX2_X1 U13186 ( .A(n14526), .B(n10513), .S(n14527), .Z(n10514) );
  AOI22_X1 U13187 ( .A1(n10515), .A2(n10514), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10516) );
  OAI211_X1 U13188 ( .C1(n15287), .C2(n10518), .A(n10517), .B(n10516), .ZN(
        P1_U3243) );
  NAND2_X1 U13189 ( .A1(n10524), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10521) );
  INV_X1 U13190 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10519) );
  MUX2_X1 U13191 ( .A(n10519), .B(P1_REG2_REG_9__SCAN_IN), .S(n10644), .Z(
        n10520) );
  AOI21_X1 U13192 ( .B1(n10522), .B2(n10521), .A(n10520), .ZN(n10643) );
  NAND3_X1 U13193 ( .A1(n10522), .A2(n10521), .A3(n10520), .ZN(n10523) );
  NAND2_X1 U13194 ( .A1(n10523), .A2(n15277), .ZN(n10533) );
  NOR2_X1 U13195 ( .A1(n10524), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10525) );
  INV_X1 U13196 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n15438) );
  MUX2_X1 U13197 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n15438), .S(n10644), .Z(
        n10526) );
  INV_X1 U13198 ( .A(n10639), .ZN(n10529) );
  NOR3_X1 U13199 ( .A1(n10527), .A2(n10526), .A3(n10525), .ZN(n10528) );
  OAI21_X1 U13200 ( .B1(n10529), .B2(n10528), .A(n15270), .ZN(n10532) );
  INV_X1 U13201 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n11281) );
  NAND2_X1 U13202 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n11984) );
  OAI21_X1 U13203 ( .B1(n15287), .B2(n11281), .A(n11984), .ZN(n10530) );
  AOI21_X1 U13204 ( .B1(n15279), .B2(n10644), .A(n10530), .ZN(n10531) );
  OAI211_X1 U13205 ( .C1(n10643), .C2(n10533), .A(n10532), .B(n10531), .ZN(
        P1_U3252) );
  NAND3_X1 U13206 ( .A1(n10536), .A2(n10535), .A3(n10534), .ZN(n10537) );
  NAND2_X1 U13207 ( .A1(n15277), .A2(n10537), .ZN(n10549) );
  NAND2_X1 U13208 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n11507) );
  INV_X1 U13209 ( .A(n11507), .ZN(n10539) );
  NOR2_X1 U13210 ( .A1(n14644), .A2(n10540), .ZN(n10538) );
  AOI211_X1 U13211 ( .C1(n14631), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n10539), .B(
        n10538), .ZN(n10548) );
  MUX2_X1 U13212 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n15435), .S(n10540), .Z(
        n10543) );
  INV_X1 U13213 ( .A(n10541), .ZN(n10542) );
  NAND2_X1 U13214 ( .A1(n10543), .A2(n10542), .ZN(n10545) );
  OAI211_X1 U13215 ( .C1(n10546), .C2(n10545), .A(n10544), .B(n15270), .ZN(
        n10547) );
  OAI211_X1 U13216 ( .C1(n10550), .C2(n10549), .A(n10548), .B(n10547), .ZN(
        P1_U3250) );
  INV_X1 U13217 ( .A(n10551), .ZN(n10552) );
  OAI222_X1 U13218 ( .A1(n13250), .A2(n10553), .B1(n13248), .B2(n10552), .C1(
        P3_U3151), .C2(n7639), .ZN(P3_U3279) );
  INV_X1 U13219 ( .A(n11721), .ZN(n10556) );
  INV_X1 U13220 ( .A(n10554), .ZN(n10557) );
  OAI222_X1 U13221 ( .A1(P1_U3086), .A2(n10556), .B1(n15164), .B2(n10555), 
        .C1(n15169), .C2(n10557), .ZN(P1_U3341) );
  INV_X1 U13222 ( .A(n11378), .ZN(n11672) );
  OAI222_X1 U13223 ( .A1(P2_U3088), .A2(n11672), .B1(n14372), .B2(n10558), 
        .C1(n14374), .C2(n10557), .ZN(P2_U3313) );
  INV_X1 U13224 ( .A(SI_14_), .ZN(n10562) );
  INV_X1 U13225 ( .A(n10559), .ZN(n10561) );
  INV_X1 U13226 ( .A(n10560), .ZN(n12681) );
  OAI222_X1 U13227 ( .A1(n13256), .A2(n10562), .B1(n13248), .B2(n10561), .C1(
        P3_U3151), .C2(n12681), .ZN(P3_U3281) );
  INV_X1 U13228 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n15705) );
  NAND2_X1 U13229 ( .A1(n15639), .A2(n12647), .ZN(n10563) );
  OAI21_X1 U13230 ( .B1(P3_U3897), .B2(n15705), .A(n10563), .ZN(P3_U3496) );
  OAI222_X1 U13231 ( .A1(n13250), .A2(n10566), .B1(n10565), .B2(P3_U3151), 
        .C1(n13260), .C2(n10564), .ZN(P3_U3278) );
  XNOR2_X1 U13232 ( .A(n10720), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n10718) );
  NOR2_X1 U13233 ( .A1(n10680), .A2(n10672), .ZN(n10571) );
  OAI21_X1 U13234 ( .B1(n10567), .B2(n13838), .A(n13835), .ZN(n13849) );
  MUX2_X1 U13235 ( .A(n10568), .B(P2_REG1_REG_2__SCAN_IN), .S(n13851), .Z(
        n13850) );
  NAND2_X1 U13236 ( .A1(n13849), .A2(n13850), .ZN(n13848) );
  INV_X1 U13237 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10569) );
  MUX2_X1 U13238 ( .A(n10569), .B(P2_REG1_REG_3__SCAN_IN), .S(n15452), .Z(
        n15459) );
  INV_X1 U13239 ( .A(n15452), .ZN(n10570) );
  NAND2_X1 U13240 ( .A1(n10570), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n13868) );
  INV_X1 U13241 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n15576) );
  MUX2_X1 U13242 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n15576), .S(n13861), .Z(
        n13867) );
  NOR2_X1 U13243 ( .A1(n13861), .A2(n15576), .ZN(n10674) );
  NOR2_X1 U13244 ( .A1(n10676), .A2(n10571), .ZN(n15473) );
  XNOR2_X1 U13245 ( .A(n15464), .B(n8179), .ZN(n15474) );
  OAI22_X1 U13246 ( .A1(n15473), .A2(n15474), .B1(n8179), .B2(n15464), .ZN(
        n10616) );
  INV_X1 U13247 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10572) );
  XNOR2_X1 U13248 ( .A(n10612), .B(n10572), .ZN(n10617) );
  XNOR2_X1 U13249 ( .A(n10627), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n10624) );
  INV_X1 U13250 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10574) );
  OAI22_X1 U13251 ( .A1(n10625), .A2(n10624), .B1(n10574), .B2(n10573), .ZN(
        n10719) );
  XOR2_X1 U13252 ( .A(n10718), .B(n10719), .Z(n10611) );
  AND2_X1 U13253 ( .A1(n10578), .A2(n11861), .ZN(n10744) );
  INV_X1 U13254 ( .A(n10575), .ZN(n10736) );
  NAND2_X1 U13255 ( .A1(n10744), .A2(n10736), .ZN(n10580) );
  INV_X1 U13256 ( .A(n11861), .ZN(n10577) );
  OAI21_X1 U13257 ( .B1(n10578), .B2(n10577), .A(n10576), .ZN(n10579) );
  NAND2_X1 U13258 ( .A1(n10580), .A2(n10579), .ZN(n10605) );
  NOR2_X1 U13259 ( .A1(n10604), .A2(n8615), .ZN(n10581) );
  INV_X1 U13260 ( .A(n14366), .ZN(n13793) );
  NAND2_X1 U13261 ( .A1(n10581), .A2(n13793), .ZN(n15444) );
  AND2_X1 U13262 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10582) );
  OR2_X1 U13263 ( .A1(n13838), .A2(n6966), .ZN(n10583) );
  INV_X1 U13264 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10584) );
  MUX2_X1 U13265 ( .A(n10584), .B(P2_REG2_REG_2__SCAN_IN), .S(n13851), .Z(
        n10585) );
  OR2_X1 U13266 ( .A1(n13851), .A2(n10584), .ZN(n10586) );
  NAND2_X1 U13267 ( .A1(n13845), .A2(n10586), .ZN(n15455) );
  MUX2_X1 U13268 ( .A(n11216), .B(P2_REG2_REG_3__SCAN_IN), .S(n15452), .Z(
        n15456) );
  OR2_X1 U13269 ( .A1(n15452), .A2(n11216), .ZN(n13863) );
  NAND2_X1 U13270 ( .A1(n15454), .A2(n13863), .ZN(n10588) );
  MUX2_X1 U13271 ( .A(n10589), .B(P2_REG2_REG_4__SCAN_IN), .S(n13861), .Z(
        n10587) );
  NAND2_X1 U13272 ( .A1(n10588), .A2(n10587), .ZN(n13865) );
  OR2_X1 U13273 ( .A1(n13861), .A2(n10589), .ZN(n10682) );
  NAND2_X1 U13274 ( .A1(n13865), .A2(n10682), .ZN(n10592) );
  INV_X1 U13275 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10590) );
  MUX2_X1 U13276 ( .A(n10590), .B(P2_REG2_REG_5__SCAN_IN), .S(n10680), .Z(
        n10591) );
  INV_X1 U13277 ( .A(n10680), .ZN(n10679) );
  NAND2_X1 U13278 ( .A1(n10679), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10593) );
  MUX2_X1 U13279 ( .A(n11357), .B(P2_REG2_REG_6__SCAN_IN), .S(n15464), .Z(
        n15472) );
  OR2_X1 U13280 ( .A1(n15464), .A2(n11357), .ZN(n10614) );
  MUX2_X1 U13281 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n11412), .S(n10612), .Z(
        n10594) );
  NAND2_X1 U13282 ( .A1(n10595), .A2(n10594), .ZN(n10630) );
  NAND2_X1 U13283 ( .A1(n10612), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10629) );
  NAND2_X1 U13284 ( .A1(n10630), .A2(n10629), .ZN(n10598) );
  INV_X1 U13285 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10596) );
  MUX2_X1 U13286 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10596), .S(n10627), .Z(
        n10597) );
  NAND2_X1 U13287 ( .A1(n10598), .A2(n10597), .ZN(n10632) );
  NAND2_X1 U13288 ( .A1(n10627), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10599) );
  INV_X1 U13289 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10600) );
  MUX2_X1 U13290 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n10600), .S(n10720), .Z(
        n10602) );
  MUX2_X1 U13291 ( .A(n10600), .B(P2_REG2_REG_9__SCAN_IN), .S(n10720), .Z(
        n10601) );
  OAI21_X1 U13292 ( .B1(n6662), .B2(n10602), .A(n10722), .ZN(n10609) );
  NAND2_X1 U13293 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n11630) );
  NAND2_X1 U13294 ( .A1(n15468), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n10606) );
  OAI211_X1 U13295 ( .C1(n15465), .C2(n10607), .A(n11630), .B(n10606), .ZN(
        n10608) );
  AOI21_X1 U13296 ( .B1(n15470), .B2(n10609), .A(n10608), .ZN(n10610) );
  OAI21_X1 U13297 ( .B1(n10611), .B2(n15445), .A(n10610), .ZN(P2_U3223) );
  MUX2_X1 U13298 ( .A(n11412), .B(P2_REG2_REG_7__SCAN_IN), .S(n10612), .Z(
        n10613) );
  NAND3_X1 U13299 ( .A1(n15469), .A2(n10614), .A3(n10613), .ZN(n10615) );
  NAND3_X1 U13300 ( .A1(n15470), .A2(n10630), .A3(n10615), .ZN(n10622) );
  NAND2_X1 U13301 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n11581) );
  XOR2_X1 U13302 ( .A(n10617), .B(n10616), .Z(n10618) );
  NAND2_X1 U13303 ( .A1(n15475), .A2(n10618), .ZN(n10619) );
  NAND2_X1 U13304 ( .A1(n11581), .A2(n10619), .ZN(n10620) );
  AOI21_X1 U13305 ( .B1(n15468), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n10620), .ZN(
        n10621) );
  OAI211_X1 U13306 ( .C1(n15465), .C2(n10623), .A(n10622), .B(n10621), .ZN(
        P2_U3221) );
  XNOR2_X1 U13307 ( .A(n10625), .B(n10624), .ZN(n10635) );
  INV_X1 U13308 ( .A(n15468), .ZN(n13938) );
  NAND2_X1 U13309 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n11688) );
  OAI21_X1 U13310 ( .B1(n13938), .B2(n7206), .A(n11688), .ZN(n10626) );
  AOI21_X1 U13311 ( .B1(n10627), .B2(n15447), .A(n10626), .ZN(n10634) );
  MUX2_X1 U13312 ( .A(n10596), .B(P2_REG2_REG_8__SCAN_IN), .S(n10627), .Z(
        n10628) );
  NAND3_X1 U13313 ( .A1(n10630), .A2(n10629), .A3(n10628), .ZN(n10631) );
  NAND3_X1 U13314 ( .A1(n15470), .A2(n10632), .A3(n10631), .ZN(n10633) );
  OAI211_X1 U13315 ( .C1(n10635), .C2(n15445), .A(n10634), .B(n10633), .ZN(
        P2_U3222) );
  OAI222_X1 U13316 ( .A1(n13250), .A2(n10638), .B1(n10637), .B2(P3_U3151), 
        .C1(n13248), .C2(n10636), .ZN(P3_U3277) );
  OAI21_X1 U13317 ( .B1(n10644), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10639), .ZN(
        n10641) );
  INV_X1 U13318 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n15441) );
  MUX2_X1 U13319 ( .A(n15441), .B(P1_REG1_REG_10__SCAN_IN), .S(n10703), .Z(
        n10640) );
  NOR2_X1 U13320 ( .A1(n10641), .A2(n10640), .ZN(n10702) );
  AOI211_X1 U13321 ( .C1(n10641), .C2(n10640), .A(n14645), .B(n10702), .ZN(
        n10642) );
  INV_X1 U13322 ( .A(n10642), .ZN(n10652) );
  NAND2_X1 U13323 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11948)
         );
  INV_X1 U13324 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10645) );
  MUX2_X1 U13325 ( .A(n10645), .B(P1_REG2_REG_10__SCAN_IN), .S(n10703), .Z(
        n10646) );
  INV_X1 U13326 ( .A(n15277), .ZN(n11724) );
  AOI21_X1 U13327 ( .B1(n10647), .B2(n10646), .A(n11724), .ZN(n10648) );
  NAND2_X1 U13328 ( .A1(n10648), .A2(n10700), .ZN(n10649) );
  NAND2_X1 U13329 ( .A1(n11948), .A2(n10649), .ZN(n10650) );
  AOI21_X1 U13330 ( .B1(n14631), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n10650), 
        .ZN(n10651) );
  OAI211_X1 U13331 ( .C1(n14644), .C2(n10653), .A(n10652), .B(n10651), .ZN(
        P1_U3253) );
  XOR2_X1 U13332 ( .A(n10655), .B(n10654), .Z(n10661) );
  NAND2_X1 U13333 ( .A1(n14510), .A2(n14903), .ZN(n10656) );
  OAI21_X1 U13334 ( .B1(n10991), .B2(n14931), .A(n10656), .ZN(n11364) );
  AOI22_X1 U13335 ( .A1(n14496), .A2(n10657), .B1(n14491), .B2(n11364), .ZN(
        n10660) );
  OR2_X1 U13336 ( .A1(n10658), .A2(P1_U3086), .ZN(n10691) );
  NAND2_X1 U13337 ( .A1(n10691), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n10659) );
  OAI211_X1 U13338 ( .C1(n10661), .C2(n14498), .A(n10660), .B(n10659), .ZN(
        P1_U3237) );
  XOR2_X1 U13339 ( .A(n10663), .B(n10662), .Z(n10667) );
  INV_X1 U13340 ( .A(n14496), .ZN(n14468) );
  AOI22_X1 U13341 ( .A1(n14473), .A2(n14511), .B1(n14478), .B2(n9435), .ZN(
        n10664) );
  OAI21_X1 U13342 ( .B1(n14468), .B2(n7698), .A(n10664), .ZN(n10665) );
  AOI21_X1 U13343 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n10691), .A(n10665), .ZN(
        n10666) );
  OAI21_X1 U13344 ( .B1(n14498), .B2(n10667), .A(n10666), .ZN(P1_U3222) );
  INV_X1 U13345 ( .A(n10668), .ZN(n10671) );
  OAI222_X1 U13346 ( .A1(n7307), .A2(P2_U3088), .B1(n14367), .B2(n10671), .C1(
        n10669), .C2(n14372), .ZN(P2_U3312) );
  OAI222_X1 U13347 ( .A1(n14598), .A2(P1_U3086), .B1(n15169), .B2(n10671), 
        .C1(n10670), .C2(n15164), .ZN(P1_U3340) );
  NAND2_X1 U13348 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n13419) );
  OAI21_X1 U13349 ( .B1(n13938), .B2(n7457), .A(n13419), .ZN(n10678) );
  MUX2_X1 U13350 ( .A(n10672), .B(P2_REG1_REG_5__SCAN_IN), .S(n10680), .Z(
        n10673) );
  NOR3_X1 U13351 ( .A1(n13866), .A2(n10674), .A3(n10673), .ZN(n10675) );
  NOR3_X1 U13352 ( .A1(n15445), .A2(n10676), .A3(n10675), .ZN(n10677) );
  AOI211_X1 U13353 ( .C1(n15447), .C2(n10679), .A(n10678), .B(n10677), .ZN(
        n10686) );
  MUX2_X1 U13354 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10590), .S(n10680), .Z(
        n10681) );
  NAND3_X1 U13355 ( .A1(n13865), .A2(n10682), .A3(n10681), .ZN(n10683) );
  NAND3_X1 U13356 ( .A1(n15470), .A2(n10684), .A3(n10683), .ZN(n10685) );
  NAND2_X1 U13357 ( .A1(n10686), .A2(n10685), .ZN(P2_U3219) );
  INV_X1 U13358 ( .A(n14994), .ZN(n10696) );
  NAND2_X1 U13359 ( .A1(n7192), .A2(n10688), .ZN(n10689) );
  NAND2_X1 U13360 ( .A1(n10690), .A2(n10689), .ZN(n14523) );
  INV_X1 U13361 ( .A(n14523), .ZN(n10693) );
  NAND2_X1 U13362 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n10691), .ZN(n10692) );
  OAI21_X1 U13363 ( .B1(n14498), .B2(n10693), .A(n10692), .ZN(n10694) );
  AOI21_X1 U13364 ( .B1(n14473), .B2(n14512), .A(n10694), .ZN(n10695) );
  OAI21_X1 U13365 ( .B1(n10696), .B2(n14468), .A(n10695), .ZN(P1_U3232) );
  NAND2_X1 U13366 ( .A1(n10703), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10699) );
  INV_X1 U13367 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10697) );
  MUX2_X1 U13368 ( .A(n10697), .B(P1_REG2_REG_11__SCAN_IN), .S(n11317), .Z(
        n10698) );
  NAND3_X1 U13369 ( .A1(n10700), .A2(n10699), .A3(n10698), .ZN(n10701) );
  NAND2_X1 U13370 ( .A1(n10701), .A2(n15277), .ZN(n10711) );
  NOR2_X1 U13371 ( .A1(n11317), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n11323) );
  AOI21_X1 U13372 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n11317), .A(n11323), 
        .ZN(n10704) );
  OAI21_X1 U13373 ( .B1(n10705), .B2(n10704), .A(n11325), .ZN(n10706) );
  NAND2_X1 U13374 ( .A1(n10706), .A2(n15270), .ZN(n10710) );
  INV_X1 U13375 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10707) );
  NAND2_X1 U13376 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n11936)
         );
  OAI21_X1 U13377 ( .B1(n15287), .B2(n10707), .A(n11936), .ZN(n10708) );
  AOI21_X1 U13378 ( .B1(n15279), .B2(n11317), .A(n10708), .ZN(n10709) );
  OAI211_X1 U13379 ( .C1(n11316), .C2(n10711), .A(n10710), .B(n10709), .ZN(
        P1_U3254) );
  INV_X1 U13380 ( .A(n13885), .ZN(n13893) );
  INV_X1 U13381 ( .A(n10712), .ZN(n10714) );
  OAI222_X1 U13382 ( .A1(P2_U3088), .A2(n13893), .B1(n14372), .B2(n10713), 
        .C1(n14374), .C2(n10714), .ZN(P2_U3311) );
  OAI222_X1 U13383 ( .A1(P1_U3086), .A2(n14612), .B1(n15164), .B2(n10715), 
        .C1(n15169), .C2(n10714), .ZN(P1_U3339) );
  OAI222_X1 U13384 ( .A1(n13260), .A2(n10717), .B1(n12357), .B2(P3_U3151), 
        .C1(n10716), .C2(n13250), .ZN(P3_U3276) );
  XNOR2_X1 U13385 ( .A(n10723), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n10786) );
  NOR2_X1 U13386 ( .A1(n10785), .A2(n10786), .ZN(n10784) );
  XNOR2_X1 U13387 ( .A(n10917), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n10912) );
  XNOR2_X1 U13388 ( .A(n10913), .B(n10912), .ZN(n10733) );
  OR2_X1 U13389 ( .A1(n10720), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10721) );
  MUX2_X1 U13390 ( .A(n11872), .B(P2_REG2_REG_10__SCAN_IN), .S(n10723), .Z(
        n10780) );
  NAND2_X1 U13391 ( .A1(n10723), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10724) );
  NAND2_X1 U13392 ( .A1(n10782), .A2(n10724), .ZN(n10726) );
  INV_X1 U13393 ( .A(n10726), .ZN(n10728) );
  INV_X1 U13394 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11810) );
  MUX2_X1 U13395 ( .A(n11810), .B(P2_REG2_REG_11__SCAN_IN), .S(n10917), .Z(
        n10725) );
  INV_X1 U13396 ( .A(n10725), .ZN(n10727) );
  OAI21_X1 U13397 ( .B1(n10728), .B2(n10727), .A(n10921), .ZN(n10731) );
  NAND2_X1 U13398 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n11888)
         );
  NAND2_X1 U13399 ( .A1(n15468), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n10729) );
  OAI211_X1 U13400 ( .C1(n15465), .C2(n10911), .A(n11888), .B(n10729), .ZN(
        n10730) );
  AOI21_X1 U13401 ( .B1(n10731), .B2(n15470), .A(n10730), .ZN(n10732) );
  OAI21_X1 U13402 ( .B1(n10733), .B2(n15445), .A(n10732), .ZN(P2_U3225) );
  INV_X1 U13403 ( .A(n15516), .ZN(n11019) );
  NAND2_X1 U13404 ( .A1(n10734), .A2(n11019), .ZN(n10743) );
  INV_X1 U13405 ( .A(n10743), .ZN(n10735) );
  NAND2_X1 U13406 ( .A1(n10735), .A2(n15517), .ZN(n10749) );
  AND2_X1 U13407 ( .A1(n12371), .A2(n13300), .ZN(n12375) );
  AOI21_X1 U13408 ( .B1(n13314), .B2(n7237), .A(n12375), .ZN(n10739) );
  XNOR2_X1 U13409 ( .A(n10875), .B(n10876), .ZN(n10738) );
  NAND2_X1 U13410 ( .A1(n10738), .A2(n10739), .ZN(n10879) );
  OAI21_X1 U13411 ( .B1(n10739), .B2(n10738), .A(n10879), .ZN(n10752) );
  OR2_X1 U13412 ( .A1(n15518), .A2(n8558), .ZN(n11021) );
  OR2_X1 U13413 ( .A1(n10749), .A2(n11021), .ZN(n10741) );
  NAND2_X1 U13414 ( .A1(n10743), .A2(n10742), .ZN(n10746) );
  AND2_X1 U13415 ( .A1(n10744), .A2(n10747), .ZN(n10745) );
  NAND2_X1 U13416 ( .A1(n10746), .A2(n10745), .ZN(n11232) );
  NOR2_X1 U13417 ( .A1(n11232), .A2(P2_U3088), .ZN(n12370) );
  INV_X1 U13418 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n11302) );
  OAI22_X1 U13419 ( .A1(n13498), .A2(n13512), .B1(n12370), .B2(n11302), .ZN(
        n10751) );
  INV_X1 U13420 ( .A(n10747), .ZN(n10748) );
  OR3_X1 U13421 ( .A1(n10749), .A2(n10748), .A3(n15495), .ZN(n13492) );
  INV_X1 U13422 ( .A(n13507), .ZN(n12372) );
  OAI22_X1 U13423 ( .A1(n13492), .A2(n12372), .B1(n11298), .B2(n13491), .ZN(
        n10750) );
  AOI211_X1 U13424 ( .C1(n13487), .C2(n10752), .A(n10751), .B(n10750), .ZN(
        n10753) );
  INV_X1 U13425 ( .A(n10753), .ZN(P2_U3194) );
  NAND2_X1 U13426 ( .A1(n10755), .A2(n10387), .ZN(n10758) );
  NAND2_X1 U13427 ( .A1(n10756), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n10757) );
  XNOR2_X1 U13428 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n10759) );
  XNOR2_X1 U13429 ( .A(n10768), .B(n10759), .ZN(n15180) );
  NAND2_X1 U13430 ( .A1(n15179), .A2(n15180), .ZN(n10763) );
  INV_X1 U13431 ( .A(n10760), .ZN(n10761) );
  NAND2_X1 U13432 ( .A1(n10761), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n10762) );
  INV_X1 U13433 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10764) );
  INV_X1 U13434 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10765) );
  OR2_X1 U13435 ( .A1(n10765), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n10767) );
  AND2_X1 U13436 ( .A1(n10765), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n10766) );
  XNOR2_X1 U13437 ( .A(n10773), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n10772) );
  INV_X1 U13438 ( .A(n10772), .ZN(n10769) );
  XNOR2_X1 U13439 ( .A(n10769), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15182) );
  NAND2_X1 U13440 ( .A1(n10770), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n10771) );
  NAND2_X1 U13441 ( .A1(n10772), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n10775) );
  INV_X1 U13442 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n11036) );
  NAND2_X1 U13443 ( .A1(n10773), .A2(n11036), .ZN(n10774) );
  XNOR2_X1 U13444 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(P3_ADDR_REG_8__SCAN_IN), 
        .ZN(n11276) );
  INV_X1 U13445 ( .A(n11276), .ZN(n10776) );
  NAND2_X1 U13446 ( .A1(n11275), .A2(n10779), .ZN(SUB_1596_U55) );
  AOI21_X1 U13447 ( .B1(n10781), .B2(n10780), .A(n15444), .ZN(n10783) );
  NAND2_X1 U13448 ( .A1(n10783), .A2(n10782), .ZN(n10791) );
  NAND2_X1 U13449 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n11775)
         );
  AOI211_X1 U13450 ( .C1(n10786), .C2(n10785), .A(n10784), .B(n15445), .ZN(
        n10787) );
  INV_X1 U13451 ( .A(n10787), .ZN(n10788) );
  NAND2_X1 U13452 ( .A1(n11775), .A2(n10788), .ZN(n10789) );
  AOI21_X1 U13453 ( .B1(n15468), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n10789), 
        .ZN(n10790) );
  OAI211_X1 U13454 ( .C1(n15465), .C2(n10792), .A(n10791), .B(n10790), .ZN(
        P2_U3224) );
  XNOR2_X1 U13455 ( .A(n10794), .B(n10793), .ZN(n10799) );
  OAI21_X1 U13456 ( .B1(P3_REG2_REG_3__SCAN_IN), .B2(n6676), .A(n10795), .ZN(
        n10796) );
  NAND2_X1 U13457 ( .A1(n12744), .A2(n10796), .ZN(n10798) );
  AOI22_X1 U13458 ( .A1(n15581), .A2(P3_ADDR_REG_3__SCAN_IN), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(P3_U3151), .ZN(n10797) );
  OAI211_X1 U13459 ( .C1(n12750), .C2(n10799), .A(n10798), .B(n10797), .ZN(
        n10800) );
  AOI21_X1 U13460 ( .B1(n10801), .B2(n12751), .A(n10800), .ZN(n10807) );
  AND3_X1 U13461 ( .A1(n10935), .A2(n10803), .A3(n10802), .ZN(n10804) );
  OAI21_X1 U13462 ( .B1(n10805), .B2(n10804), .A(n12675), .ZN(n10806) );
  NAND2_X1 U13463 ( .A1(n10807), .A2(n10806), .ZN(P3_U3185) );
  AOI21_X1 U13464 ( .B1(n10809), .B2(n10808), .A(n6670), .ZN(n10827) );
  NOR2_X1 U13465 ( .A1(n10811), .A2(n10810), .ZN(n10812) );
  NOR2_X1 U13466 ( .A1(n10813), .A2(n10812), .ZN(n10823) );
  INV_X1 U13467 ( .A(n10814), .ZN(n10816) );
  NAND3_X1 U13468 ( .A1(n10795), .A2(n10816), .A3(n10815), .ZN(n10817) );
  NAND2_X1 U13469 ( .A1(n10818), .A2(n10817), .ZN(n10819) );
  NAND2_X1 U13470 ( .A1(n12744), .A2(n10819), .ZN(n10822) );
  NAND2_X1 U13471 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n11168) );
  INV_X1 U13472 ( .A(n11168), .ZN(n10820) );
  AOI21_X1 U13473 ( .B1(n15581), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n10820), .ZN(
        n10821) );
  OAI211_X1 U13474 ( .C1(n12750), .C2(n10823), .A(n10822), .B(n10821), .ZN(
        n10824) );
  AOI21_X1 U13475 ( .B1(n10825), .B2(n12751), .A(n10824), .ZN(n10826) );
  OAI21_X1 U13476 ( .B1(n10827), .B2(n12755), .A(n10826), .ZN(P3_U3186) );
  INV_X1 U13477 ( .A(n10858), .ZN(n10833) );
  OR2_X1 U13478 ( .A1(n10862), .A2(n10860), .ZN(n10832) );
  AND3_X1 U13479 ( .A1(n10830), .A2(n10829), .A3(n10828), .ZN(n10831) );
  OAI211_X1 U13480 ( .C1(n10859), .C2(n10833), .A(n10832), .B(n10831), .ZN(
        n10834) );
  NAND2_X1 U13481 ( .A1(n10834), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10838) );
  INV_X1 U13482 ( .A(n10862), .ZN(n10836) );
  NAND2_X1 U13483 ( .A1(n10836), .A2(n12365), .ZN(n10837) );
  NAND2_X2 U13484 ( .A1(n10838), .A2(n10837), .ZN(n12630) );
  NOR2_X1 U13485 ( .A1(n12630), .A2(P3_U3151), .ZN(n10901) );
  INV_X1 U13486 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10870) );
  NAND2_X1 U13487 ( .A1(n10844), .A2(n10839), .ZN(n12593) );
  NOR2_X1 U13488 ( .A1(n10840), .A2(n15651), .ZN(n10841) );
  NAND2_X1 U13489 ( .A1(n10859), .A2(n10841), .ZN(n10842) );
  INV_X1 U13490 ( .A(n15586), .ZN(n11394) );
  NAND2_X2 U13491 ( .A1(n10844), .A2(n10843), .ZN(n12628) );
  OAI22_X1 U13492 ( .A1(n10845), .A2(n12610), .B1(n12628), .B2(n15608), .ZN(
        n10846) );
  AOI21_X1 U13493 ( .B1(n12626), .B2(n15605), .A(n10846), .ZN(n10869) );
  NAND2_X1 U13494 ( .A1(n10850), .A2(n12316), .ZN(n10851) );
  NAND3_X1 U13495 ( .A1(n12646), .A2(n12494), .A3(n13014), .ZN(n10852) );
  INV_X1 U13496 ( .A(n10853), .ZN(n12168) );
  NAND2_X1 U13497 ( .A1(n13017), .A2(n12494), .ZN(n10854) );
  OAI21_X1 U13498 ( .B1(n12168), .B2(n13008), .A(n10854), .ZN(n10855) );
  NAND3_X1 U13499 ( .A1(n13018), .A2(n13008), .A3(n12463), .ZN(n10856) );
  OAI211_X1 U13500 ( .C1(n10857), .C2(n13017), .A(n10892), .B(n10856), .ZN(
        n10867) );
  NAND3_X1 U13501 ( .A1(n10859), .A2(n10858), .A3(n15651), .ZN(n10864) );
  INV_X1 U13502 ( .A(n10860), .ZN(n10861) );
  NAND2_X1 U13503 ( .A1(n10862), .A2(n10861), .ZN(n10863) );
  NAND2_X1 U13504 ( .A1(n10864), .A2(n10863), .ZN(n10866) );
  NAND2_X1 U13505 ( .A1(n10867), .A2(n12589), .ZN(n10868) );
  OAI211_X1 U13506 ( .C1(n10901), .C2(n10870), .A(n10869), .B(n10868), .ZN(
        P3_U3162) );
  INV_X1 U13507 ( .A(n10871), .ZN(n10873) );
  OAI222_X1 U13508 ( .A1(P1_U3086), .A2(n14625), .B1(n15164), .B2(n10872), 
        .C1(n15169), .C2(n10873), .ZN(P1_U3338) );
  INV_X1 U13509 ( .A(n13915), .ZN(n13908) );
  OAI222_X1 U13510 ( .A1(P2_U3088), .A2(n13908), .B1(n14372), .B2(n10874), 
        .C1(n14374), .C2(n10873), .ZN(P2_U3310) );
  XNOR2_X1 U13511 ( .A(n13515), .B(n13379), .ZN(n11225) );
  NAND2_X1 U13512 ( .A1(n13829), .A2(n13300), .ZN(n11223) );
  XNOR2_X1 U13513 ( .A(n11225), .B(n11223), .ZN(n10881) );
  INV_X1 U13514 ( .A(n10875), .ZN(n10877) );
  NAND2_X1 U13515 ( .A1(n10879), .A2(n10878), .ZN(n10880) );
  NAND2_X1 U13516 ( .A1(n10880), .A2(n10881), .ZN(n11224) );
  OAI21_X1 U13517 ( .B1(n10881), .B2(n10880), .A(n11224), .ZN(n10885) );
  OAI22_X1 U13518 ( .A1(n13498), .A2(n15533), .B1(n12370), .B2(n11185), .ZN(
        n10884) );
  OAI22_X1 U13519 ( .A1(n13492), .A2(n10882), .B1(n15496), .B2(n13491), .ZN(
        n10883) );
  AOI211_X1 U13520 ( .C1(n13487), .C2(n10885), .A(n10884), .B(n10883), .ZN(
        n10886) );
  INV_X1 U13521 ( .A(n10886), .ZN(P2_U3209) );
  INV_X1 U13522 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10889) );
  INV_X1 U13523 ( .A(n11397), .ZN(n11059) );
  NAND2_X1 U13524 ( .A1(n15605), .A2(n11059), .ZN(n12164) );
  NAND2_X1 U13525 ( .A1(n13008), .A2(n12164), .ZN(n12319) );
  OAI22_X1 U13526 ( .A1(n11059), .A2(n12610), .B1(n12628), .B2(n15592), .ZN(
        n10887) );
  AOI21_X1 U13527 ( .B1(n12589), .B2(n12319), .A(n10887), .ZN(n10888) );
  OAI21_X1 U13528 ( .B1(n10901), .B2(n10889), .A(n10888), .ZN(P3_U3172) );
  INV_X1 U13529 ( .A(P3_DATAO_REG_21__SCAN_IN), .ZN(n15704) );
  NAND2_X1 U13530 ( .A1(n12860), .A2(n12647), .ZN(n10890) );
  OAI21_X1 U13531 ( .B1(P3_U3897), .B2(n15704), .A(n10890), .ZN(P3_U3512) );
  INV_X1 U13532 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10900) );
  XNOR2_X1 U13533 ( .A(n11007), .B(n13012), .ZN(n10894) );
  NAND2_X1 U13534 ( .A1(n10892), .A2(n10891), .ZN(n10893) );
  OAI21_X1 U13535 ( .B1(n10894), .B2(n10893), .A(n11010), .ZN(n10895) );
  NAND2_X1 U13536 ( .A1(n10895), .A2(n12589), .ZN(n10899) );
  OAI22_X1 U13537 ( .A1(n12610), .A2(n10896), .B1(n12628), .B2(n15591), .ZN(
        n10897) );
  AOI21_X1 U13538 ( .B1(n12626), .B2(n12646), .A(n10897), .ZN(n10898) );
  OAI211_X1 U13539 ( .C1(n10901), .C2(n10900), .A(n10899), .B(n10898), .ZN(
        P3_U3177) );
  AOI211_X1 U13540 ( .C1(n10904), .C2(n10903), .A(n14498), .B(n10902), .ZN(
        n10909) );
  MUX2_X1 U13541 ( .A(n14479), .B(P1_U3086), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n10908) );
  OR2_X1 U13542 ( .A1(n9892), .A2(n14931), .ZN(n10906) );
  NAND2_X1 U13543 ( .A1(n14509), .A2(n14903), .ZN(n10905) );
  AND2_X1 U13544 ( .A1(n10906), .A2(n10905), .ZN(n15355) );
  INV_X1 U13545 ( .A(n14491), .ZN(n14433) );
  OAI22_X1 U13546 ( .A1(n14468), .A2(n15356), .B1(n15355), .B2(n14433), .ZN(
        n10907) );
  OR3_X1 U13547 ( .A1(n10909), .A2(n10908), .A3(n10907), .ZN(P1_U3218) );
  XNOR2_X1 U13548 ( .A(n11258), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n10915) );
  OAI22_X1 U13549 ( .A1(n10913), .A2(n10912), .B1(n10911), .B2(n10910), .ZN(
        n10914) );
  AOI21_X1 U13550 ( .B1(n10915), .B2(n10914), .A(n11260), .ZN(n10928) );
  AND2_X1 U13551 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n12136) );
  INV_X1 U13552 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n11965) );
  NOR2_X1 U13553 ( .A1(n13938), .A2(n11965), .ZN(n10916) );
  AOI211_X1 U13554 ( .C1(n15447), .C2(n11258), .A(n12136), .B(n10916), .ZN(
        n10927) );
  INV_X1 U13555 ( .A(n10921), .ZN(n10919) );
  MUX2_X1 U13556 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n11899), .S(n11258), .Z(
        n10922) );
  OR2_X1 U13557 ( .A1(n10917), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10920) );
  INV_X1 U13558 ( .A(n10920), .ZN(n10918) );
  NOR3_X1 U13559 ( .A1(n10919), .A2(n10922), .A3(n10918), .ZN(n10925) );
  NAND2_X1 U13560 ( .A1(n10921), .A2(n10920), .ZN(n10923) );
  NAND2_X1 U13561 ( .A1(n10923), .A2(n10922), .ZN(n11267) );
  INV_X1 U13562 ( .A(n11267), .ZN(n10924) );
  OAI21_X1 U13563 ( .B1(n10925), .B2(n10924), .A(n15470), .ZN(n10926) );
  OAI211_X1 U13564 ( .C1(n10928), .C2(n15445), .A(n10927), .B(n10926), .ZN(
        P2_U3226) );
  INV_X1 U13565 ( .A(n12751), .ZN(n12682) );
  OAI21_X1 U13566 ( .B1(n10931), .B2(n10930), .A(n10929), .ZN(n10945) );
  OR3_X1 U13567 ( .A1(n10933), .A2(n10951), .A3(n10932), .ZN(n10934) );
  AOI21_X1 U13568 ( .B1(n10935), .B2(n10934), .A(n12755), .ZN(n10944) );
  OAI21_X1 U13569 ( .B1(n10938), .B2(n10937), .A(n10936), .ZN(n10939) );
  NAND2_X1 U13570 ( .A1(n12744), .A2(n10939), .ZN(n10942) );
  NOR2_X1 U13571 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10900), .ZN(n10940) );
  AOI21_X1 U13572 ( .B1(n15581), .B2(P3_ADDR_REG_2__SCAN_IN), .A(n10940), .ZN(
        n10941) );
  NAND2_X1 U13573 ( .A1(n10942), .A2(n10941), .ZN(n10943) );
  AOI211_X1 U13574 ( .C1(n12692), .C2(n10945), .A(n10944), .B(n10943), .ZN(
        n10946) );
  OAI21_X1 U13575 ( .B1(n10947), .B2(n12682), .A(n10946), .ZN(P3_U3184) );
  INV_X1 U13576 ( .A(n10948), .ZN(n10950) );
  OAI21_X1 U13577 ( .B1(n10950), .B2(P3_REG2_REG_1__SCAN_IN), .A(n10949), .ZN(
        n10961) );
  AOI21_X1 U13578 ( .B1(n10952), .B2(n11148), .A(n10951), .ZN(n10954) );
  AOI22_X1 U13579 ( .A1(n15581), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10953) );
  OAI21_X1 U13580 ( .B1(n10954), .B2(n12755), .A(n10953), .ZN(n10960) );
  NAND2_X1 U13581 ( .A1(n10956), .A2(n10955), .ZN(n10957) );
  AOI21_X1 U13582 ( .B1(n10958), .B2(n10957), .A(n12750), .ZN(n10959) );
  AOI211_X1 U13583 ( .C1(n12744), .C2(n10961), .A(n10960), .B(n10959), .ZN(
        n10962) );
  OAI21_X1 U13584 ( .B1(n10963), .B2(n12682), .A(n10962), .ZN(P3_U3183) );
  OAI222_X1 U13585 ( .A1(n13260), .A2(n10965), .B1(n12316), .B2(P3_U3151), 
        .C1(n10964), .C2(n13250), .ZN(P3_U3275) );
  NAND3_X1 U13586 ( .A1(n12319), .A2(n10966), .A3(n15651), .ZN(n10967) );
  OAI21_X1 U13587 ( .B1(n15592), .B2(n15642), .A(n10967), .ZN(n11057) );
  INV_X1 U13588 ( .A(n11057), .ZN(n11393) );
  MUX2_X1 U13589 ( .A(n15725), .B(n11393), .S(n15676), .Z(n10968) );
  OAI21_X1 U13590 ( .B1(n11059), .B2(n9283), .A(n10968), .ZN(P3_U3459) );
  INV_X1 U13591 ( .A(n11046), .ZN(n10970) );
  INV_X1 U13592 ( .A(n11045), .ZN(n10969) );
  NAND3_X1 U13593 ( .A1(n10970), .A2(n10969), .A3(n15005), .ZN(n14729) );
  INV_X1 U13594 ( .A(n11044), .ZN(n10972) );
  INV_X4 U13595 ( .A(n14935), .ZN(n15336) );
  OAI21_X1 U13596 ( .B1(n10974), .B2(n10973), .A(n12425), .ZN(n14910) );
  INV_X1 U13597 ( .A(n11102), .ZN(n11095) );
  NAND2_X1 U13598 ( .A1(n11066), .A2(n11064), .ZN(n10976) );
  NAND2_X1 U13599 ( .A1(n10991), .A2(n7698), .ZN(n10975) );
  NAND2_X1 U13600 ( .A1(n9892), .A2(n9891), .ZN(n10977) );
  NAND2_X1 U13601 ( .A1(n11306), .A2(n10979), .ZN(n10982) );
  NAND2_X1 U13602 ( .A1(n10980), .A2(n15356), .ZN(n10981) );
  NAND2_X1 U13603 ( .A1(n10982), .A2(n10981), .ZN(n11096) );
  XNOR2_X1 U13604 ( .A(n11095), .B(n11096), .ZN(n15370) );
  INV_X1 U13605 ( .A(n15370), .ZN(n11006) );
  INV_X1 U13606 ( .A(n11104), .ZN(n15368) );
  NAND2_X1 U13608 ( .A1(n11368), .A2(n9891), .ZN(n11367) );
  INV_X1 U13609 ( .A(n10984), .ZN(n11309) );
  NOR2_X2 U13610 ( .A1(n10984), .A2(n11104), .ZN(n15330) );
  INV_X1 U13611 ( .A(n15330), .ZN(n10985) );
  OAI211_X1 U13612 ( .C1(n15368), .C2(n11309), .A(n10985), .B(n15328), .ZN(
        n15366) );
  NAND2_X1 U13613 ( .A1(n15176), .A2(n9940), .ZN(n10989) );
  NAND2_X1 U13614 ( .A1(n10987), .A2(n10986), .ZN(n10988) );
  NAND2_X1 U13615 ( .A1(n14512), .A2(n7698), .ZN(n10993) );
  NAND2_X1 U13616 ( .A1(n11361), .A2(n10994), .ZN(n11307) );
  NAND2_X1 U13617 ( .A1(n11307), .A2(n10995), .ZN(n10997) );
  NAND2_X1 U13618 ( .A1(n10997), .A2(n10996), .ZN(n11103) );
  XNOR2_X1 U13619 ( .A(n11103), .B(n11102), .ZN(n10998) );
  AOI222_X1 U13620 ( .A1(n15359), .A2(n10998), .B1(n14510), .B2(n14982), .C1(
        n14508), .C2(n14903), .ZN(n15367) );
  OAI21_X1 U13621 ( .B1(n9940), .B2(n15366), .A(n15367), .ZN(n10999) );
  NAND2_X1 U13622 ( .A1(n10999), .A2(n14935), .ZN(n11005) );
  NAND2_X1 U13623 ( .A1(n11000), .A2(n11050), .ZN(n11001) );
  OR2_X2 U13624 ( .A1(n15336), .A2(n11001), .ZN(n15311) );
  OAI22_X1 U13625 ( .A1(n14935), .A2(n10467), .B1(n11002), .B2(n14997), .ZN(
        n11003) );
  AOI21_X1 U13626 ( .B1(n14995), .B2(n11104), .A(n11003), .ZN(n11004) );
  OAI211_X1 U13627 ( .C1(n14990), .C2(n11006), .A(n11005), .B(n11004), .ZN(
        P1_U3289) );
  NAND2_X1 U13628 ( .A1(n11007), .A2(n15608), .ZN(n11008) );
  XNOR2_X1 U13629 ( .A(n11160), .B(n15620), .ZN(n11009) );
  AOI21_X1 U13630 ( .B1(n11010), .B2(n11008), .A(n11009), .ZN(n11016) );
  NAND2_X1 U13631 ( .A1(n11163), .A2(n12589), .ZN(n11015) );
  OAI22_X1 U13632 ( .A1(n12610), .A2(n11011), .B1(n12628), .B2(n15628), .ZN(
        n11013) );
  MUX2_X1 U13633 ( .A(P3_U3151), .B(n12630), .S(n15680), .Z(n11012) );
  AOI211_X1 U13634 ( .C1(n12626), .C2(n13012), .A(n11013), .B(n11012), .ZN(
        n11014) );
  OAI21_X1 U13635 ( .B1(n11016), .B2(n11015), .A(n11014), .ZN(P3_U3158) );
  NAND4_X1 U13636 ( .A1(n11019), .A2(n11018), .A3(n11017), .A4(n15513), .ZN(
        n11020) );
  INV_X1 U13637 ( .A(n11021), .ZN(n11022) );
  AOI21_X1 U13638 ( .B1(n15484), .B2(n11023), .A(n15827), .ZN(n11031) );
  NAND2_X1 U13639 ( .A1(n12372), .A2(n7237), .ZN(n11024) );
  NAND2_X1 U13640 ( .A1(n11025), .A2(n11024), .ZN(n15519) );
  INV_X1 U13641 ( .A(n15556), .ZN(n14274) );
  AND2_X1 U13642 ( .A1(n14274), .A2(n15501), .ZN(n11026) );
  OAI22_X1 U13643 ( .A1(n15519), .A2(n11026), .B1(n10882), .B2(n15493), .ZN(
        n15521) );
  OAI22_X1 U13644 ( .A1(n15831), .A2(n8127), .B1(n11027), .B2(n15503), .ZN(
        n11029) );
  NAND2_X1 U13645 ( .A1(n15831), .A2(n13499), .ZN(n14172) );
  NOR2_X1 U13646 ( .A1(n15519), .A2(n14172), .ZN(n11028) );
  AOI211_X1 U13647 ( .C1(n15831), .C2(n15521), .A(n11029), .B(n11028), .ZN(
        n11030) );
  OAI21_X1 U13648 ( .B1(n11031), .B2(n7237), .A(n11030), .ZN(P2_U3265) );
  XNOR2_X1 U13649 ( .A(n11032), .B(P3_REG1_REG_7__SCAN_IN), .ZN(n11043) );
  XNOR2_X1 U13650 ( .A(n11034), .B(n11033), .ZN(n11041) );
  INV_X1 U13651 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11571) );
  XNOR2_X1 U13652 ( .A(n11035), .B(n11571), .ZN(n11039) );
  INV_X1 U13653 ( .A(n12744), .ZN(n12702) );
  NOR2_X1 U13654 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8912), .ZN(n11665) );
  INV_X1 U13655 ( .A(n15581), .ZN(n12715) );
  NOR2_X1 U13656 ( .A1(n12715), .A2(n11036), .ZN(n11037) );
  AOI211_X1 U13657 ( .C1(n12751), .C2(n7436), .A(n11665), .B(n11037), .ZN(
        n11038) );
  OAI21_X1 U13658 ( .B1(n11039), .B2(n12702), .A(n11038), .ZN(n11040) );
  AOI21_X1 U13659 ( .B1(n11041), .B2(n12675), .A(n11040), .ZN(n11042) );
  OAI21_X1 U13660 ( .B1(n11043), .B2(n12750), .A(n11042), .ZN(P3_U3189) );
  NAND2_X1 U13661 ( .A1(n11045), .A2(n11044), .ZN(n11047) );
  OR2_X1 U13662 ( .A1(n11047), .A2(n11046), .ZN(n15006) );
  INV_X1 U13663 ( .A(n15005), .ZN(n11048) );
  INV_X1 U13664 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n11054) );
  OR2_X1 U13665 ( .A1(n14910), .A2(n9940), .ZN(n15305) );
  OR2_X1 U13666 ( .A1(n11049), .A2(n14817), .ZN(n15393) );
  OAI21_X1 U13667 ( .B1(n15359), .B2(n15402), .A(n14991), .ZN(n11052) );
  OR2_X1 U13668 ( .A1(n10991), .A2(n14980), .ZN(n14998) );
  NAND3_X1 U13669 ( .A1(n14994), .A2(n11710), .A3(n11050), .ZN(n11051) );
  NAND3_X1 U13670 ( .A1(n11052), .A2(n14998), .A3(n11051), .ZN(n15130) );
  NAND2_X1 U13671 ( .A1(n15425), .A2(n15130), .ZN(n11053) );
  OAI21_X1 U13672 ( .B1(n15425), .B2(n11054), .A(n11053), .ZN(P1_U3459) );
  INV_X1 U13673 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11055) );
  NOR2_X1 U13674 ( .A1(n15666), .A2(n11055), .ZN(n11056) );
  AOI21_X1 U13675 ( .B1(n15666), .B2(n11057), .A(n11056), .ZN(n11058) );
  OAI21_X1 U13676 ( .B1(n11059), .B2(n9296), .A(n11058), .ZN(P3_U3390) );
  INV_X1 U13677 ( .A(n14640), .ZN(n14634) );
  INV_X1 U13678 ( .A(n11060), .ZN(n11062) );
  OAI222_X1 U13679 ( .A1(P1_U3086), .A2(n14634), .B1(n15164), .B2(n11061), 
        .C1(n15169), .C2(n11062), .ZN(P1_U3337) );
  INV_X1 U13680 ( .A(n13927), .ZN(n13920) );
  OAI222_X1 U13681 ( .A1(P2_U3088), .A2(n13920), .B1(n14372), .B2(n11063), 
        .C1(n14374), .C2(n11062), .ZN(P2_U3309) );
  INV_X1 U13682 ( .A(n11064), .ZN(n11065) );
  XNOR2_X1 U13683 ( .A(n7190), .B(n11065), .ZN(n15339) );
  NOR2_X1 U13684 ( .A1(n15336), .A2(n11067), .ZN(n15333) );
  INV_X1 U13685 ( .A(n15333), .ZN(n11080) );
  OAI22_X1 U13686 ( .A1(n14935), .A2(n10460), .B1(n7003), .B2(n14997), .ZN(
        n11071) );
  NAND2_X1 U13687 ( .A1(n15332), .A2(n15328), .ZN(n14840) );
  INV_X1 U13688 ( .A(n11368), .ZN(n11069) );
  NAND2_X1 U13689 ( .A1(n14994), .A2(n15341), .ZN(n11068) );
  NAND2_X1 U13690 ( .A1(n11069), .A2(n11068), .ZN(n15343) );
  NOR2_X1 U13691 ( .A1(n14840), .A2(n15343), .ZN(n11070) );
  AOI211_X1 U13692 ( .C1(n14995), .C2(n15341), .A(n11071), .B(n11070), .ZN(
        n11079) );
  AOI21_X1 U13693 ( .B1(n11072), .B2(n9435), .A(n15400), .ZN(n11076) );
  XNOR2_X1 U13694 ( .A(n15343), .B(n10991), .ZN(n11074) );
  OAI21_X1 U13695 ( .B1(n11074), .B2(n15400), .A(n11073), .ZN(n11075) );
  OAI21_X1 U13696 ( .B1(n14982), .B2(n11076), .A(n11075), .ZN(n11077) );
  OAI21_X1 U13697 ( .B1(n15305), .B2(n15339), .A(n11077), .ZN(n15345) );
  NOR2_X1 U13698 ( .A1(n9892), .A2(n14980), .ZN(n15340) );
  OAI21_X1 U13699 ( .B1(n15345), .B2(n15340), .A(n14935), .ZN(n11078) );
  OAI211_X1 U13700 ( .C1(n15339), .C2(n11080), .A(n11079), .B(n11078), .ZN(
        P1_U3292) );
  XOR2_X1 U13701 ( .A(n11082), .B(n11081), .Z(n11094) );
  OAI21_X1 U13702 ( .B1(n11084), .B2(n11083), .A(n6664), .ZN(n11092) );
  AND2_X1 U13703 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n11551) );
  AOI21_X1 U13704 ( .B1(n15581), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n11551), .ZN(
        n11085) );
  OAI21_X1 U13705 ( .B1(n12682), .B2(n11086), .A(n11085), .ZN(n11091) );
  AOI21_X1 U13706 ( .B1(n11088), .B2(n11087), .A(n6665), .ZN(n11089) );
  NOR2_X1 U13707 ( .A1(n11089), .A2(n12750), .ZN(n11090) );
  AOI211_X1 U13708 ( .C1(n12744), .C2(n11092), .A(n11091), .B(n11090), .ZN(
        n11093) );
  OAI21_X1 U13709 ( .B1(n11094), .B2(n12755), .A(n11093), .ZN(P3_U3188) );
  NAND2_X1 U13710 ( .A1(n11096), .A2(n11095), .ZN(n11098) );
  INV_X1 U13711 ( .A(n14509), .ZN(n11105) );
  NAND2_X1 U13712 ( .A1(n11105), .A2(n15368), .ZN(n11097) );
  NAND2_X1 U13713 ( .A1(n11098), .A2(n11097), .ZN(n15318) );
  NAND2_X1 U13714 ( .A1(n15318), .A2(n15320), .ZN(n11101) );
  NAND2_X1 U13715 ( .A1(n11099), .A2(n15373), .ZN(n11100) );
  NAND2_X1 U13716 ( .A1(n11101), .A2(n11100), .ZN(n11249) );
  XOR2_X1 U13717 ( .A(n11249), .B(n11248), .Z(n15383) );
  NAND2_X1 U13718 ( .A1(n11105), .A2(n11104), .ZN(n11106) );
  NAND2_X1 U13719 ( .A1(n15373), .A2(n14508), .ZN(n11108) );
  XNOR2_X1 U13720 ( .A(n11238), .B(n11248), .ZN(n11111) );
  NAND2_X1 U13721 ( .A1(n14508), .A2(n14982), .ZN(n11110) );
  NAND2_X1 U13722 ( .A1(n14506), .A2(n14903), .ZN(n11109) );
  NAND2_X1 U13723 ( .A1(n11110), .A2(n11109), .ZN(n11441) );
  AOI21_X1 U13724 ( .B1(n11111), .B2(n15359), .A(n11441), .ZN(n15381) );
  MUX2_X1 U13725 ( .A(n15381), .B(n11112), .S(n15336), .Z(n11118) );
  NAND2_X1 U13726 ( .A1(n15330), .A2(n15373), .ZN(n15329) );
  INV_X1 U13727 ( .A(n15314), .ZN(n11114) );
  AOI211_X1 U13728 ( .C1(n15380), .C2(n15329), .A(n15344), .B(n11114), .ZN(
        n15379) );
  INV_X1 U13729 ( .A(n11115), .ZN(n11444) );
  OAI22_X1 U13730 ( .A1(n15311), .A2(n11250), .B1(n14997), .B2(n11444), .ZN(
        n11116) );
  AOI21_X1 U13731 ( .B1(n15379), .B2(n15332), .A(n11116), .ZN(n11117) );
  OAI211_X1 U13732 ( .C1(n14990), .C2(n15383), .A(n11118), .B(n11117), .ZN(
        P1_U3287) );
  INV_X1 U13733 ( .A(n11119), .ZN(n11120) );
  NOR2_X1 U13734 ( .A1(n11121), .A2(n11120), .ZN(n11122) );
  XNOR2_X1 U13735 ( .A(n11123), .B(n11122), .ZN(n11134) );
  XNOR2_X1 U13736 ( .A(n11124), .B(P3_REG1_REG_5__SCAN_IN), .ZN(n11132) );
  AND2_X1 U13737 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n11426) );
  AOI21_X1 U13738 ( .B1(n15581), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11426), .ZN(
        n11129) );
  OAI21_X1 U13739 ( .B1(P3_REG2_REG_5__SCAN_IN), .B2(n11126), .A(n11125), .ZN(
        n11127) );
  NAND2_X1 U13740 ( .A1(n12744), .A2(n11127), .ZN(n11128) );
  OAI211_X1 U13741 ( .C1(n12682), .C2(n11130), .A(n11129), .B(n11128), .ZN(
        n11131) );
  AOI21_X1 U13742 ( .B1(n12692), .B2(n11132), .A(n11131), .ZN(n11133) );
  OAI21_X1 U13743 ( .B1(n11134), .B2(n12755), .A(n11133), .ZN(P3_U3187) );
  INV_X1 U13744 ( .A(n11135), .ZN(n11139) );
  OAI222_X1 U13745 ( .A1(P2_U3088), .A2(n11137), .B1(n14374), .B2(n11139), 
        .C1(n11136), .C2(n14372), .ZN(P2_U3308) );
  OAI222_X1 U13746 ( .A1(n14817), .A2(P1_U3086), .B1(n15169), .B2(n11139), 
        .C1(n11138), .C2(n15164), .ZN(P1_U3336) );
  NOR3_X1 U13747 ( .A1(n12692), .A2(n12744), .A3(n12675), .ZN(n11149) );
  OAI22_X1 U13748 ( .A1(n12715), .A2(n11140), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10889), .ZN(n11141) );
  AOI21_X1 U13749 ( .B1(n12692), .B2(n11142), .A(n11141), .ZN(n11147) );
  NOR2_X1 U13750 ( .A1(n12755), .A2(n11143), .ZN(n11144) );
  AOI21_X1 U13751 ( .B1(n12744), .B2(P3_REG2_REG_0__SCAN_IN), .A(n11144), .ZN(
        n11145) );
  MUX2_X1 U13752 ( .A(n11145), .B(n12682), .S(P3_IR_REG_0__SCAN_IN), .Z(n11146) );
  OAI211_X1 U13753 ( .C1(n11149), .C2(n11148), .A(n11147), .B(n11146), .ZN(
        P3_U3182) );
  XNOR2_X1 U13754 ( .A(n11431), .B(n11432), .ZN(n11150) );
  XNOR2_X1 U13755 ( .A(n11433), .B(n11150), .ZN(n11158) );
  INV_X1 U13756 ( .A(n15325), .ZN(n11156) );
  NAND2_X1 U13757 ( .A1(n14509), .A2(n14982), .ZN(n11152) );
  NAND2_X1 U13758 ( .A1(n14507), .A2(n14903), .ZN(n11151) );
  NAND2_X1 U13759 ( .A1(n11152), .A2(n11151), .ZN(n15323) );
  AOI22_X1 U13760 ( .A1(n14491), .A2(n15323), .B1(P1_REG3_REG_5__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11155) );
  NAND2_X1 U13761 ( .A1(n14496), .A2(n11153), .ZN(n11154) );
  OAI211_X1 U13762 ( .C1(n14494), .C2(n11156), .A(n11155), .B(n11154), .ZN(
        n11157) );
  AOI21_X1 U13763 ( .B1(n11158), .B2(n14462), .A(n11157), .ZN(n11159) );
  INV_X1 U13764 ( .A(n11159), .ZN(P1_U3227) );
  INV_X1 U13765 ( .A(n11160), .ZN(n11161) );
  NAND2_X1 U13766 ( .A1(n11161), .A2(n15620), .ZN(n11162) );
  XNOR2_X1 U13767 ( .A(n12463), .B(n15619), .ZN(n11164) );
  NAND2_X1 U13768 ( .A1(n11164), .A2(n15628), .ZN(n11420) );
  INV_X1 U13769 ( .A(n11421), .ZN(n11165) );
  AOI21_X1 U13770 ( .B1(n11167), .B2(n11166), .A(n11165), .ZN(n11173) );
  INV_X1 U13771 ( .A(n12628), .ZN(n12511) );
  AOI22_X1 U13772 ( .A1(n12511), .A2(n15639), .B1(n12626), .B2(n15620), .ZN(
        n11169) );
  OAI211_X1 U13773 ( .C1(n12610), .C2(n11170), .A(n11169), .B(n11168), .ZN(
        n11171) );
  AOI21_X1 U13774 ( .B1(n11530), .B2(n12630), .A(n11171), .ZN(n11172) );
  OAI21_X1 U13775 ( .B1(n11173), .B2(n12634), .A(n11172), .ZN(P3_U3170) );
  INV_X1 U13776 ( .A(n15501), .ZN(n15550) );
  NAND2_X1 U13777 ( .A1(n11295), .A2(n11174), .ZN(n11175) );
  NAND2_X1 U13778 ( .A1(n11175), .A2(n11179), .ZN(n11207) );
  OAI21_X1 U13779 ( .B1(n11175), .B2(n11179), .A(n11207), .ZN(n15537) );
  OAI22_X1 U13780 ( .A1(n15496), .A2(n15493), .B1(n10882), .B2(n15495), .ZN(
        n11182) );
  INV_X1 U13781 ( .A(n11179), .ZN(n13760) );
  NAND2_X1 U13782 ( .A1(n11176), .A2(n13760), .ZN(n11211) );
  NAND3_X1 U13783 ( .A1(n11177), .A2(n11179), .A3(n11178), .ZN(n11180) );
  AOI21_X1 U13784 ( .B1(n11211), .B2(n11180), .A(n14274), .ZN(n11181) );
  AOI211_X1 U13785 ( .C1(n15550), .C2(n15537), .A(n11182), .B(n11181), .ZN(
        n15534) );
  INV_X1 U13786 ( .A(n14172), .ZN(n15835) );
  NAND2_X1 U13787 ( .A1(n11183), .A2(n14181), .ZN(n11184) );
  OR2_X1 U13788 ( .A1(n11184), .A2(n11217), .ZN(n15532) );
  OAI22_X1 U13789 ( .A1(n15831), .A2(n10584), .B1(n11185), .B2(n15503), .ZN(
        n11186) );
  AOI21_X1 U13790 ( .B1(n15827), .B2(n13515), .A(n11186), .ZN(n11187) );
  OAI21_X1 U13791 ( .B1(n15829), .B2(n15532), .A(n11187), .ZN(n11188) );
  AOI21_X1 U13792 ( .B1(n15835), .B2(n15537), .A(n11188), .ZN(n11189) );
  OAI21_X1 U13793 ( .B1(n15534), .B2(n14180), .A(n11189), .ZN(P2_U3263) );
  XOR2_X1 U13794 ( .A(n11190), .B(n11191), .Z(n11204) );
  XNOR2_X1 U13795 ( .A(n11193), .B(n11192), .ZN(n11202) );
  AOI21_X1 U13796 ( .B1(n11196), .B2(n11195), .A(n11194), .ZN(n11200) );
  NOR2_X1 U13797 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n6704), .ZN(n11799) );
  INV_X1 U13798 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n11278) );
  NOR2_X1 U13799 ( .A1(n12715), .A2(n11278), .ZN(n11197) );
  AOI211_X1 U13800 ( .C1(n12751), .C2(n11198), .A(n11799), .B(n11197), .ZN(
        n11199) );
  OAI21_X1 U13801 ( .B1(n11200), .B2(n12702), .A(n11199), .ZN(n11201) );
  AOI21_X1 U13802 ( .B1(n11202), .B2(n12675), .A(n11201), .ZN(n11203) );
  OAI21_X1 U13803 ( .B1(n11204), .B2(n12750), .A(n11203), .ZN(P3_U3190) );
  INV_X1 U13804 ( .A(n13763), .ZN(n11206) );
  NAND3_X1 U13805 ( .A1(n11207), .A2(n11206), .A3(n11205), .ZN(n11209) );
  NAND2_X1 U13806 ( .A1(n11209), .A2(n11208), .ZN(n11404) );
  OAI22_X1 U13807 ( .A1(n11298), .A2(n15495), .B1(n15544), .B2(n15493), .ZN(
        n11215) );
  AOI21_X1 U13808 ( .B1(n11211), .B2(n11210), .A(n13763), .ZN(n15492) );
  INV_X1 U13809 ( .A(n15492), .ZN(n11213) );
  NAND3_X1 U13810 ( .A1(n11211), .A2(n13763), .A3(n11210), .ZN(n11212) );
  AOI21_X1 U13811 ( .B1(n11213), .B2(n11212), .A(n14274), .ZN(n11214) );
  AOI211_X1 U13812 ( .C1(n15550), .C2(n11404), .A(n11215), .B(n11214), .ZN(
        n11401) );
  MUX2_X1 U13813 ( .A(n11216), .B(n11401), .S(n15831), .Z(n11221) );
  OAI211_X1 U13814 ( .C1(n11217), .C2(n13535), .A(n14181), .B(n15481), .ZN(
        n11400) );
  NOR2_X1 U13815 ( .A1(n15829), .A2(n11400), .ZN(n11219) );
  OAI22_X1 U13816 ( .A1(n15504), .A2(n13535), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n15503), .ZN(n11218) );
  AOI211_X1 U13817 ( .C1(n11404), .C2(n15835), .A(n11219), .B(n11218), .ZN(
        n11220) );
  NAND2_X1 U13818 ( .A1(n11221), .A2(n11220), .ZN(P2_U3262) );
  XNOR2_X1 U13819 ( .A(n13762), .B(n13379), .ZN(n11471) );
  INV_X1 U13820 ( .A(n11472), .ZN(n11222) );
  XNOR2_X1 U13821 ( .A(n11471), .B(n11222), .ZN(n11474) );
  INV_X1 U13822 ( .A(n11474), .ZN(n11231) );
  INV_X1 U13823 ( .A(n11223), .ZN(n11226) );
  AND2_X1 U13824 ( .A1(n13828), .A2(n13300), .ZN(n11228) );
  XNOR2_X1 U13825 ( .A(n13531), .B(n13379), .ZN(n11227) );
  NOR2_X1 U13826 ( .A1(n11228), .A2(n11227), .ZN(n11473) );
  NAND2_X1 U13827 ( .A1(n11228), .A2(n11227), .ZN(n11475) );
  INV_X1 U13828 ( .A(n11475), .ZN(n11229) );
  NOR2_X1 U13829 ( .A1(n11473), .A2(n11229), .ZN(n13351) );
  NAND2_X1 U13830 ( .A1(n6458), .A2(n13351), .ZN(n13350) );
  NAND2_X1 U13831 ( .A1(n13350), .A2(n11475), .ZN(n11230) );
  NOR2_X1 U13832 ( .A1(n11230), .A2(n11231), .ZN(n13413) );
  AOI21_X1 U13833 ( .B1(n11231), .B2(n11230), .A(n13413), .ZN(n11236) );
  NAND2_X1 U13834 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n13857) );
  OAI21_X1 U13835 ( .B1(n13492), .B2(n15496), .A(n13857), .ZN(n11234) );
  OAI22_X1 U13836 ( .A1(n15545), .A2(n13498), .B1(n13459), .B2(n15502), .ZN(
        n11233) );
  AOI211_X1 U13837 ( .C1(n13474), .C2(n13826), .A(n11234), .B(n11233), .ZN(
        n11235) );
  OAI21_X1 U13838 ( .B1(n11236), .B2(n13481), .A(n11235), .ZN(P2_U3202) );
  AND2_X1 U13839 ( .A1(n11250), .A2(n14507), .ZN(n11237) );
  INV_X1 U13840 ( .A(n14506), .ZN(n11239) );
  NAND2_X1 U13841 ( .A1(n15389), .A2(n11239), .ZN(n11240) );
  XNOR2_X1 U13842 ( .A(n11828), .B(n11829), .ZN(n15399) );
  OAI22_X1 U13843 ( .A1(n14935), .A2(n11241), .B1(n11598), .B2(n14997), .ZN(
        n11247) );
  AOI211_X1 U13844 ( .C1(n15397), .C2(n7758), .A(n15344), .B(n6478), .ZN(
        n15395) );
  OR2_X1 U13845 ( .A1(n11832), .A2(n14980), .ZN(n11244) );
  NAND2_X1 U13846 ( .A1(n14506), .A2(n14982), .ZN(n11243) );
  NAND2_X1 U13847 ( .A1(n11244), .A2(n11243), .ZN(n15396) );
  AOI21_X1 U13848 ( .B1(n15395), .B2(n14817), .A(n15396), .ZN(n11245) );
  NOR2_X1 U13849 ( .A1(n11245), .A2(n15336), .ZN(n11246) );
  AOI211_X1 U13850 ( .C1(n14995), .C2(n15397), .A(n11247), .B(n11246), .ZN(
        n11257) );
  NAND2_X1 U13851 ( .A1(n11249), .A2(n11248), .ZN(n11253) );
  NAND2_X1 U13852 ( .A1(n11251), .A2(n11250), .ZN(n11252) );
  INV_X1 U13853 ( .A(n15304), .ZN(n11254) );
  OR2_X1 U13854 ( .A1(n14506), .A2(n15389), .ZN(n11255) );
  XNOR2_X1 U13855 ( .A(n11821), .B(n11829), .ZN(n15403) );
  NAND2_X1 U13856 ( .A1(n15403), .A2(n14992), .ZN(n11256) );
  OAI211_X1 U13857 ( .C1(n15399), .C2(n14970), .A(n11257), .B(n11256), .ZN(
        P1_U3285) );
  INV_X1 U13858 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n15184) );
  NAND2_X1 U13859 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n12147)
         );
  OAI21_X1 U13860 ( .B1(n13938), .B2(n15184), .A(n12147), .ZN(n11264) );
  XNOR2_X1 U13861 ( .A(n11375), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n11262) );
  NOR2_X1 U13862 ( .A1(n11258), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n11259) );
  OR2_X1 U13863 ( .A1(n11260), .A2(n11259), .ZN(n11261) );
  AOI211_X1 U13864 ( .C1(n11262), .C2(n11261), .A(n15445), .B(n11373), .ZN(
        n11263) );
  AOI211_X1 U13865 ( .C1(n15447), .C2(n11375), .A(n11264), .B(n11263), .ZN(
        n11273) );
  NAND2_X1 U13866 ( .A1(n11265), .A2(n11899), .ZN(n11266) );
  INV_X1 U13867 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11269) );
  MUX2_X1 U13868 ( .A(n11269), .B(P2_REG2_REG_13__SCAN_IN), .S(n11268), .Z(
        n11270) );
  NAND2_X1 U13869 ( .A1(n11271), .A2(n11270), .ZN(n11377) );
  OAI211_X1 U13870 ( .C1(n11271), .C2(n11270), .A(n11377), .B(n15470), .ZN(
        n11272) );
  NAND2_X1 U13871 ( .A1(n11273), .A2(n11272), .ZN(P2_U3227) );
  NAND2_X1 U13872 ( .A1(n11277), .A2(n11276), .ZN(n11280) );
  NAND2_X1 U13873 ( .A1(n11278), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n11279) );
  XNOR2_X1 U13874 ( .A(n11281), .B(P3_ADDR_REG_9__SCAN_IN), .ZN(n11287) );
  XNOR2_X1 U13875 ( .A(n11286), .B(n11287), .ZN(n11283) );
  INV_X1 U13876 ( .A(n11282), .ZN(n11284) );
  NAND2_X1 U13877 ( .A1(n11284), .A2(n11283), .ZN(n11285) );
  XNOR2_X1 U13878 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(P3_ADDR_REG_10__SCAN_IN), 
        .ZN(n11288) );
  XNOR2_X1 U13879 ( .A(n11499), .B(n11288), .ZN(n11496) );
  INV_X1 U13880 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n11493) );
  XNOR2_X1 U13881 ( .A(n11496), .B(n11493), .ZN(n11289) );
  XNOR2_X1 U13882 ( .A(n11495), .B(n11289), .ZN(SUB_1596_U70) );
  NOR2_X1 U13883 ( .A1(n13256), .A2(SI_22_), .ZN(n11290) );
  AOI21_X1 U13884 ( .B1(n11291), .B2(P3_STATE_REG_SCAN_IN), .A(n11290), .ZN(
        n11292) );
  OAI21_X1 U13885 ( .B1(n11293), .B2(n13248), .A(n11292), .ZN(n11294) );
  INV_X1 U13886 ( .A(n11294), .ZN(P3_U3273) );
  INV_X1 U13887 ( .A(n11295), .ZN(n11296) );
  AOI21_X1 U13888 ( .B1(n12371), .B2(n8563), .A(n11296), .ZN(n15529) );
  OAI21_X1 U13889 ( .B1(n11297), .B2(n8563), .A(n11177), .ZN(n11301) );
  OAI22_X1 U13890 ( .A1(n12372), .A2(n15495), .B1(n11298), .B2(n15493), .ZN(
        n11300) );
  NOR2_X1 U13891 ( .A1(n15529), .A2(n15501), .ZN(n11299) );
  AOI211_X1 U13892 ( .C1(n15556), .C2(n11301), .A(n11300), .B(n11299), .ZN(
        n15527) );
  MUX2_X1 U13893 ( .A(n6966), .B(n15527), .S(n15831), .Z(n11305) );
  AOI211_X1 U13894 ( .C1(n13503), .C2(n15524), .A(n15561), .B(n6661), .ZN(
        n15523) );
  OAI22_X1 U13895 ( .A1(n15504), .A2(n13512), .B1(n11302), .B2(n15503), .ZN(
        n11303) );
  AOI21_X1 U13896 ( .B1(n15484), .B2(n15523), .A(n11303), .ZN(n11304) );
  OAI211_X1 U13897 ( .C1(n15529), .C2(n14172), .A(n11305), .B(n11304), .ZN(
        P2_U3264) );
  XNOR2_X1 U13898 ( .A(n11306), .B(n11308), .ZN(n15362) );
  INV_X1 U13899 ( .A(n14970), .ZN(n14993) );
  XNOR2_X1 U13900 ( .A(n11307), .B(n11308), .ZN(n15360) );
  AOI211_X1 U13901 ( .C1(n11310), .C2(n11367), .A(n15344), .B(n11309), .ZN(
        n15357) );
  INV_X1 U13902 ( .A(n14997), .ZN(n15324) );
  AOI22_X1 U13903 ( .A1(n15357), .A2(n15332), .B1(n15324), .B2(n9457), .ZN(
        n11313) );
  MUX2_X1 U13904 ( .A(n15355), .B(n11311), .S(n15336), .Z(n11312) );
  OAI211_X1 U13905 ( .C1(n15356), .C2(n15311), .A(n11313), .B(n11312), .ZN(
        n11314) );
  AOI21_X1 U13906 ( .B1(n14993), .B2(n15360), .A(n11314), .ZN(n11315) );
  OAI21_X1 U13907 ( .B1(n14990), .B2(n15362), .A(n11315), .ZN(P1_U3290) );
  INV_X1 U13908 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11318) );
  MUX2_X1 U13909 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n11318), .S(n14585), .Z(
        n14583) );
  NAND2_X1 U13910 ( .A1(n14582), .A2(n14583), .ZN(n14581) );
  OAI21_X1 U13911 ( .B1(n14585), .B2(P1_REG2_REG_12__SCAN_IN), .A(n14581), 
        .ZN(n11321) );
  INV_X1 U13912 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11319) );
  MUX2_X1 U13913 ( .A(n11319), .B(P1_REG2_REG_13__SCAN_IN), .S(n11340), .Z(
        n11320) );
  AOI21_X1 U13914 ( .B1(n11321), .B2(n11320), .A(n11724), .ZN(n11322) );
  NAND2_X1 U13915 ( .A1(n11322), .A2(n11337), .ZN(n11332) );
  NAND2_X1 U13916 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n14454)
         );
  XNOR2_X1 U13917 ( .A(n11340), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n11327) );
  INV_X1 U13918 ( .A(n11323), .ZN(n11324) );
  XOR2_X1 U13919 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n14585), .Z(n14578) );
  NOR2_X1 U13920 ( .A1(n11326), .A2(n11327), .ZN(n11339) );
  AOI211_X1 U13921 ( .C1(n11327), .C2(n11326), .A(n11339), .B(n14645), .ZN(
        n11328) );
  INV_X1 U13922 ( .A(n11328), .ZN(n11329) );
  NAND2_X1 U13923 ( .A1(n14454), .A2(n11329), .ZN(n11330) );
  AOI21_X1 U13924 ( .B1(n14631), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n11330), 
        .ZN(n11331) );
  OAI211_X1 U13925 ( .C1(n14644), .C2(n11333), .A(n11332), .B(n11331), .ZN(
        P1_U3256) );
  NAND2_X1 U13926 ( .A1(n11340), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11336) );
  INV_X1 U13927 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11334) );
  MUX2_X1 U13928 ( .A(n11334), .B(P1_REG2_REG_14__SCAN_IN), .S(n11721), .Z(
        n11335) );
  NAND3_X1 U13929 ( .A1(n11337), .A2(n11336), .A3(n11335), .ZN(n11338) );
  NAND2_X1 U13930 ( .A1(n11338), .A2(n15277), .ZN(n11349) );
  XOR2_X1 U13931 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n11721), .Z(n11342) );
  OAI21_X1 U13932 ( .B1(n11342), .B2(n11341), .A(n11718), .ZN(n11343) );
  NAND2_X1 U13933 ( .A1(n11343), .A2(n15270), .ZN(n11348) );
  NOR2_X1 U13934 ( .A1(n11344), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14382) );
  INV_X1 U13935 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n11345) );
  NOR2_X1 U13936 ( .A1(n15287), .A2(n11345), .ZN(n11346) );
  AOI211_X1 U13937 ( .C1(n15279), .C2(n11721), .A(n14382), .B(n11346), .ZN(
        n11347) );
  OAI211_X1 U13938 ( .C1(n11720), .C2(n11349), .A(n11348), .B(n11347), .ZN(
        P1_U3257) );
  INV_X1 U13939 ( .A(n13499), .ZN(n11350) );
  NAND2_X1 U13940 ( .A1(n15501), .A2(n11350), .ZN(n11351) );
  XNOR2_X1 U13941 ( .A(n11352), .B(n13765), .ZN(n14309) );
  XNOR2_X1 U13942 ( .A(n11353), .B(n11354), .ZN(n11355) );
  OAI222_X1 U13943 ( .A1(n15495), .A2(n15494), .B1(n15493), .B2(n11487), .C1(
        n14274), .C2(n11355), .ZN(n14305) );
  INV_X1 U13944 ( .A(n14305), .ZN(n11356) );
  MUX2_X1 U13945 ( .A(n11357), .B(n11356), .S(n15831), .Z(n11360) );
  AOI211_X1 U13946 ( .C1(n14307), .C2(n15563), .A(n15561), .B(n11415), .ZN(
        n14306) );
  OAI22_X1 U13947 ( .A1(n15504), .A2(n13554), .B1(n11486), .B2(n15503), .ZN(
        n11358) );
  AOI21_X1 U13948 ( .B1(n14306), .B2(n15484), .A(n11358), .ZN(n11359) );
  OAI211_X1 U13949 ( .C1(n14200), .C2(n14309), .A(n11360), .B(n11359), .ZN(
        P2_U3259) );
  OAI21_X1 U13950 ( .B1(n11363), .B2(n11362), .A(n11361), .ZN(n11365) );
  AOI21_X1 U13951 ( .B1(n11365), .B2(n15359), .A(n11364), .ZN(n15350) );
  NAND2_X1 U13952 ( .A1(n14992), .A2(n15353), .ZN(n11372) );
  OAI211_X1 U13953 ( .C1(n11368), .C2(n9891), .A(n15328), .B(n11367), .ZN(
        n15349) );
  INV_X1 U13954 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n14530) );
  OAI22_X1 U13955 ( .A1(n14952), .A2(n15349), .B1(n14530), .B2(n14997), .ZN(
        n11370) );
  NOR2_X1 U13956 ( .A1(n15311), .A2(n9891), .ZN(n11369) );
  AOI211_X1 U13957 ( .C1(n15336), .C2(P1_REG2_REG_2__SCAN_IN), .A(n11370), .B(
        n11369), .ZN(n11371) );
  OAI211_X1 U13958 ( .C1(n15336), .C2(n15350), .A(n11372), .B(n11371), .ZN(
        P1_U3291) );
  AOI21_X1 U13959 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n11375), .A(n11373), 
        .ZN(n11674) );
  XNOR2_X1 U13960 ( .A(n11378), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n11673) );
  XNOR2_X1 U13961 ( .A(n11674), .B(n11673), .ZN(n11386) );
  INV_X1 U13962 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n15197) );
  NAND2_X1 U13963 ( .A1(P2_U3088), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n13334)
         );
  OAI21_X1 U13964 ( .B1(n13938), .B2(n15197), .A(n13334), .ZN(n11374) );
  AOI21_X1 U13965 ( .B1(n11378), .B2(n15447), .A(n11374), .ZN(n11385) );
  NAND2_X1 U13966 ( .A1(n11375), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11376) );
  NAND2_X1 U13967 ( .A1(n11379), .A2(n11378), .ZN(n11380) );
  INV_X1 U13968 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n11381) );
  NAND2_X1 U13969 ( .A1(n11382), .A2(n11381), .ZN(n11671) );
  OAI21_X1 U13970 ( .B1(n11382), .B2(n11381), .A(n11671), .ZN(n11383) );
  NAND2_X1 U13971 ( .A1(n11383), .A2(n15470), .ZN(n11384) );
  OAI211_X1 U13972 ( .C1(n11386), .C2(n15445), .A(n11385), .B(n11384), .ZN(
        P2_U3228) );
  INV_X1 U13973 ( .A(n11387), .ZN(n11392) );
  NAND2_X1 U13974 ( .A1(n11388), .A2(n11391), .ZN(n11389) );
  OAI211_X1 U13975 ( .C1(n11392), .C2(n11391), .A(n11390), .B(n11389), .ZN(
        n11396) );
  MUX2_X1 U13976 ( .A(n11393), .B(n8822), .S(n15601), .Z(n11399) );
  OR2_X1 U13977 ( .A1(n15651), .A2(n11394), .ZN(n11395) );
  INV_X1 U13978 ( .A(n12991), .ZN(n12804) );
  INV_X2 U13979 ( .A(n15588), .ZN(n13011) );
  AOI22_X1 U13980 ( .A1(n13004), .A2(n11397), .B1(P3_REG3_REG_0__SCAN_IN), 
        .B2(n13011), .ZN(n11398) );
  NAND2_X1 U13981 ( .A1(n11399), .A2(n11398), .ZN(P3_U3233) );
  INV_X1 U13982 ( .A(n15528), .ZN(n15560) );
  INV_X1 U13983 ( .A(n11400), .ZN(n11403) );
  INV_X1 U13984 ( .A(n11401), .ZN(n11402) );
  AOI211_X1 U13985 ( .C1(n15560), .C2(n11404), .A(n11403), .B(n11402), .ZN(
        n11409) );
  INV_X1 U13986 ( .A(n14294), .ZN(n14280) );
  AOI22_X1 U13987 ( .A1(n14280), .A2(n13531), .B1(n15578), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n11405) );
  OAI21_X1 U13988 ( .B1(n11409), .B2(n15578), .A(n11405), .ZN(P2_U3502) );
  INV_X1 U13989 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n11406) );
  OAI22_X1 U13990 ( .A1(n14350), .A2(n13535), .B1(n15571), .B2(n11406), .ZN(
        n11407) );
  INV_X1 U13991 ( .A(n11407), .ZN(n11408) );
  OAI21_X1 U13992 ( .B1(n11409), .B2(n15569), .A(n11408), .ZN(P2_U3439) );
  XNOR2_X1 U13993 ( .A(n11410), .B(n8571), .ZN(n11411) );
  AOI222_X1 U13994 ( .A1(n15556), .A2(n11411), .B1(n13825), .B2(n14188), .C1(
        n13823), .C2(n14190), .ZN(n11561) );
  MUX2_X1 U13995 ( .A(n11412), .B(n11561), .S(n15831), .Z(n11419) );
  XNOR2_X1 U13996 ( .A(n11413), .B(n11414), .ZN(n11563) );
  INV_X1 U13997 ( .A(n14200), .ZN(n14134) );
  OAI22_X1 U13998 ( .A1(n15504), .A2(n11588), .B1(n11583), .B2(n15503), .ZN(
        n11417) );
  OAI211_X1 U13999 ( .C1(n11415), .C2(n11588), .A(n11695), .B(n14181), .ZN(
        n11560) );
  NOR2_X1 U14000 ( .A1(n11560), .A2(n15829), .ZN(n11416) );
  AOI211_X1 U14001 ( .C1(n11563), .C2(n14134), .A(n11417), .B(n11416), .ZN(
        n11418) );
  NAND2_X1 U14002 ( .A1(n11419), .A2(n11418), .ZN(P2_U3258) );
  INV_X1 U14003 ( .A(n11540), .ZN(n11429) );
  INV_X1 U14004 ( .A(n12630), .ZN(n11554) );
  XNOR2_X1 U14005 ( .A(n12463), .B(n11541), .ZN(n11547) );
  XNOR2_X1 U14006 ( .A(n11547), .B(n15639), .ZN(n11423) );
  OAI21_X1 U14007 ( .B1(n11423), .B2(n11422), .A(n11640), .ZN(n11424) );
  NAND2_X1 U14008 ( .A1(n11424), .A2(n12589), .ZN(n11428) );
  OAI22_X1 U14009 ( .A1(n15653), .A2(n12628), .B1(n12593), .B2(n15628), .ZN(
        n11425) );
  AOI211_X1 U14010 ( .C1(n11541), .C2(n12631), .A(n11426), .B(n11425), .ZN(
        n11427) );
  OAI211_X1 U14011 ( .C1(n11429), .C2(n11554), .A(n11428), .B(n11427), .ZN(
        P3_U3167) );
  INV_X1 U14012 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n15762) );
  NAND2_X1 U14013 ( .A1(n12861), .A2(n12647), .ZN(n11430) );
  OAI21_X1 U14014 ( .B1(P3_U3897), .B2(n15762), .A(n11430), .ZN(P3_U3514) );
  INV_X1 U14015 ( .A(n11433), .ZN(n11435) );
  OAI21_X1 U14016 ( .B1(n11433), .B2(n11432), .A(n11431), .ZN(n11434) );
  OAI21_X1 U14017 ( .B1(n11435), .B2(n7896), .A(n11434), .ZN(n11439) );
  XNOR2_X1 U14018 ( .A(n11437), .B(n11436), .ZN(n11438) );
  XNOR2_X1 U14019 ( .A(n11439), .B(n11438), .ZN(n11446) );
  AOI21_X1 U14020 ( .B1(n14491), .B2(n11441), .A(n11440), .ZN(n11443) );
  NAND2_X1 U14021 ( .A1(n14496), .A2(n15380), .ZN(n11442) );
  OAI211_X1 U14022 ( .C1(n14494), .C2(n11444), .A(n11443), .B(n11442), .ZN(
        n11445) );
  AOI21_X1 U14023 ( .B1(n11446), .B2(n14462), .A(n11445), .ZN(n11447) );
  INV_X1 U14024 ( .A(n11447), .ZN(P1_U3239) );
  OAI21_X1 U14025 ( .B1(n11449), .B2(n12323), .A(n11448), .ZN(n15616) );
  INV_X1 U14026 ( .A(n15616), .ZN(n11457) );
  OR2_X1 U14027 ( .A1(n15586), .A2(n10849), .ZN(n15582) );
  NOR2_X1 U14028 ( .A1(n15601), .A2(n15582), .ZN(n12806) );
  INV_X1 U14029 ( .A(n12806), .ZN(n11456) );
  INV_X1 U14030 ( .A(n15644), .ZN(n15662) );
  OAI22_X1 U14031 ( .A1(n15628), .A2(n15642), .B1(n15608), .B2(n15652), .ZN(
        n11452) );
  NOR2_X1 U14032 ( .A1(n11450), .A2(n12323), .ZN(n11525) );
  AOI211_X1 U14033 ( .C1(n12323), .C2(n11450), .A(n13052), .B(n11525), .ZN(
        n11451) );
  AOI211_X1 U14034 ( .C1(n15662), .C2(n15616), .A(n11452), .B(n11451), .ZN(
        n15618) );
  MUX2_X1 U14035 ( .A(n11453), .B(n15618), .S(n15599), .Z(n11455) );
  AOI22_X1 U14036 ( .A1(n13004), .A2(n15615), .B1(n13011), .B2(n15680), .ZN(
        n11454) );
  OAI211_X1 U14037 ( .C1(n11457), .C2(n11456), .A(n11455), .B(n11454), .ZN(
        P3_U3230) );
  XOR2_X1 U14038 ( .A(n11458), .B(P3_REG1_REG_9__SCAN_IN), .Z(n11470) );
  NAND2_X1 U14039 ( .A1(n6668), .A2(n11459), .ZN(n11460) );
  XNOR2_X1 U14040 ( .A(n11461), .B(n11460), .ZN(n11468) );
  OAI21_X1 U14041 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n11462), .A(n11611), .ZN(
        n11463) );
  NAND2_X1 U14042 ( .A1(n11463), .A2(n12744), .ZN(n11465) );
  AND2_X1 U14043 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n11656) );
  AOI21_X1 U14044 ( .B1(n15581), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n11656), .ZN(
        n11464) );
  OAI211_X1 U14045 ( .C1(n12682), .C2(n11466), .A(n11465), .B(n11464), .ZN(
        n11467) );
  AOI21_X1 U14046 ( .B1(n12675), .B2(n11468), .A(n11467), .ZN(n11469) );
  OAI21_X1 U14047 ( .B1(n11470), .B2(n12750), .A(n11469), .ZN(P3_U3191) );
  NAND2_X1 U14048 ( .A1(n13826), .A2(n13300), .ZN(n11478) );
  XNOR2_X1 U14049 ( .A(n15826), .B(n13379), .ZN(n11477) );
  INV_X1 U14050 ( .A(n11477), .ZN(n11479) );
  AND2_X1 U14051 ( .A1(n11479), .A2(n11478), .ZN(n11480) );
  NAND2_X1 U14052 ( .A1(n13825), .A2(n13300), .ZN(n11483) );
  INV_X1 U14053 ( .A(n11483), .ZN(n11482) );
  XNOR2_X1 U14054 ( .A(n14307), .B(n13314), .ZN(n11484) );
  INV_X1 U14055 ( .A(n11484), .ZN(n11481) );
  NAND2_X1 U14056 ( .A1(n11482), .A2(n11481), .ZN(n11627) );
  NAND2_X1 U14057 ( .A1(n11484), .A2(n11483), .ZN(n11618) );
  AND2_X1 U14058 ( .A1(n11627), .A2(n11618), .ZN(n11485) );
  NAND2_X1 U14059 ( .A1(n11620), .A2(n11485), .ZN(n11576) );
  OAI211_X1 U14060 ( .C1(n11620), .C2(n11485), .A(n11576), .B(n13487), .ZN(
        n11492) );
  INV_X1 U14061 ( .A(n11486), .ZN(n11490) );
  NAND2_X1 U14062 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n15463) );
  OAI21_X1 U14063 ( .B1(n13492), .B2(n15494), .A(n15463), .ZN(n11489) );
  OAI22_X1 U14064 ( .A1(n13498), .A2(n13554), .B1(n13491), .B2(n11487), .ZN(
        n11488) );
  AOI211_X1 U14065 ( .C1(n11490), .C2(n13495), .A(n11489), .B(n11488), .ZN(
        n11491) );
  NAND2_X1 U14066 ( .A1(n11492), .A2(n11491), .ZN(P2_U3211) );
  NAND2_X1 U14067 ( .A1(n11496), .A2(n11493), .ZN(n11494) );
  INV_X1 U14068 ( .A(n11496), .ZN(n11497) );
  NOR2_X1 U14069 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n11499), .ZN(n11501) );
  NAND2_X1 U14070 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n11499), .ZN(n11500) );
  XNOR2_X1 U14071 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n11733) );
  XNOR2_X1 U14072 ( .A(n11730), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(n11502) );
  XNOR2_X1 U14073 ( .A(n11731), .B(n11502), .ZN(SUB_1596_U69) );
  INV_X1 U14074 ( .A(n15309), .ZN(n11512) );
  XOR2_X1 U14075 ( .A(n11504), .B(n11503), .Z(n11505) );
  NAND2_X1 U14076 ( .A1(n11505), .A2(n14462), .ZN(n11511) );
  NAND2_X1 U14077 ( .A1(n14507), .A2(n14982), .ZN(n11506) );
  OAI21_X1 U14078 ( .B1(n11983), .B2(n14980), .A(n11506), .ZN(n15307) );
  NAND2_X1 U14079 ( .A1(n14491), .A2(n15307), .ZN(n11508) );
  NAND2_X1 U14080 ( .A1(n11508), .A2(n11507), .ZN(n11509) );
  AOI21_X1 U14081 ( .B1(n14496), .B2(n15389), .A(n11509), .ZN(n11510) );
  OAI211_X1 U14082 ( .C1(n14494), .C2(n11512), .A(n11511), .B(n11510), .ZN(
        P1_U3213) );
  OAI222_X1 U14083 ( .A1(P1_U3086), .A2(n11513), .B1(n15164), .B2(n7230), .C1(
        n15169), .C2(n12447), .ZN(P1_U3335) );
  AND2_X1 U14084 ( .A1(n15644), .A2(n15582), .ZN(n11514) );
  NAND2_X1 U14085 ( .A1(n11515), .A2(n12180), .ZN(n11516) );
  XNOR2_X1 U14086 ( .A(n11516), .B(n12321), .ZN(n15645) );
  OAI211_X1 U14087 ( .C1(n6653), .C2(n12321), .A(n11517), .B(n15611), .ZN(
        n15641) );
  MUX2_X1 U14088 ( .A(n15641), .B(n11518), .S(n15601), .Z(n11522) );
  NOR2_X1 U14089 ( .A1(n15601), .A2(n15642), .ZN(n13013) );
  AOI22_X1 U14090 ( .A1(n13004), .A2(n15636), .B1(n13011), .B2(n11546), .ZN(
        n11519) );
  OAI21_X1 U14091 ( .B1(n15623), .B2(n12989), .A(n11519), .ZN(n11520) );
  AOI21_X1 U14092 ( .B1(n13013), .B2(n12644), .A(n11520), .ZN(n11521) );
  OAI211_X1 U14093 ( .C1(n13007), .C2(n15645), .A(n11522), .B(n11521), .ZN(
        P3_U3227) );
  XNOR2_X1 U14094 ( .A(n11523), .B(n11526), .ZN(n15624) );
  NOR2_X1 U14095 ( .A1(n11525), .A2(n11524), .ZN(n11527) );
  XNOR2_X1 U14096 ( .A(n11527), .B(n11526), .ZN(n11528) );
  NAND2_X1 U14097 ( .A1(n11528), .A2(n15611), .ZN(n15622) );
  MUX2_X1 U14098 ( .A(n11529), .B(n15622), .S(n15599), .Z(n11534) );
  AOI22_X1 U14099 ( .A1(n13004), .A2(n15619), .B1(n13011), .B2(n11530), .ZN(
        n11531) );
  OAI21_X1 U14100 ( .B1(n15591), .B2(n12989), .A(n11531), .ZN(n11532) );
  AOI21_X1 U14101 ( .B1(n13013), .B2(n15639), .A(n11532), .ZN(n11533) );
  OAI211_X1 U14102 ( .C1(n13007), .C2(n15624), .A(n11534), .B(n11533), .ZN(
        P3_U3229) );
  XNOR2_X1 U14103 ( .A(n11535), .B(n7845), .ZN(n15633) );
  OAI21_X1 U14104 ( .B1(n11537), .B2(n12320), .A(n11536), .ZN(n11538) );
  NAND2_X1 U14105 ( .A1(n11538), .A2(n15611), .ZN(n15631) );
  MUX2_X1 U14106 ( .A(n15631), .B(n11539), .S(n15601), .Z(n11545) );
  AOI22_X1 U14107 ( .A1(n13004), .A2(n11541), .B1(n13011), .B2(n11540), .ZN(
        n11542) );
  OAI21_X1 U14108 ( .B1(n15628), .B2(n12989), .A(n11542), .ZN(n11543) );
  AOI21_X1 U14109 ( .B1(n13013), .B2(n15630), .A(n11543), .ZN(n11544) );
  OAI211_X1 U14110 ( .C1(n13007), .C2(n15633), .A(n11545), .B(n11544), .ZN(
        P3_U3228) );
  INV_X1 U14111 ( .A(n11546), .ZN(n11555) );
  NAND2_X1 U14112 ( .A1(n11547), .A2(n15623), .ZN(n11638) );
  AND2_X1 U14113 ( .A1(n11640), .A2(n11638), .ZN(n11549) );
  XNOR2_X1 U14114 ( .A(n12463), .B(n15636), .ZN(n11642) );
  XNOR2_X1 U14115 ( .A(n11642), .B(n15630), .ZN(n11548) );
  NAND2_X1 U14116 ( .A1(n11549), .A2(n11548), .ZN(n11662) );
  OAI211_X1 U14117 ( .C1(n11549), .C2(n11548), .A(n11662), .B(n12589), .ZN(
        n11553) );
  OAI22_X1 U14118 ( .A1(n15643), .A2(n12628), .B1(n12593), .B2(n15623), .ZN(
        n11550) );
  AOI211_X1 U14119 ( .C1(n15636), .C2(n12631), .A(n11551), .B(n11550), .ZN(
        n11552) );
  OAI211_X1 U14120 ( .C1(n11555), .C2(n11554), .A(n11553), .B(n11552), .ZN(
        P3_U3179) );
  NAND2_X1 U14121 ( .A1(n11557), .A2(n11556), .ZN(n11558) );
  OAI211_X1 U14122 ( .C1(n11559), .C2(n13250), .A(n11558), .B(n12367), .ZN(
        P3_U3272) );
  OAI211_X1 U14123 ( .C1(n11588), .C2(n15565), .A(n11561), .B(n11560), .ZN(
        n11562) );
  AOI21_X1 U14124 ( .B1(n11563), .B2(n14271), .A(n11562), .ZN(n11566) );
  NAND2_X1 U14125 ( .A1(n15569), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n11564) );
  OAI21_X1 U14126 ( .B1(n11566), .B2(n15569), .A(n11564), .ZN(P2_U3451) );
  NAND2_X1 U14127 ( .A1(n15578), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n11565) );
  OAI21_X1 U14128 ( .B1(n11566), .B2(n15578), .A(n11565), .ZN(P2_U3506) );
  AND2_X1 U14129 ( .A1(n11567), .A2(n12182), .ZN(n11568) );
  XNOR2_X1 U14130 ( .A(n11568), .B(n11636), .ZN(n15660) );
  OAI211_X1 U14131 ( .C1(n11570), .C2(n11636), .A(n11569), .B(n15611), .ZN(
        n15657) );
  MUX2_X1 U14132 ( .A(n15657), .B(n11571), .S(n15601), .Z(n11575) );
  AOI22_X1 U14133 ( .A1(n13004), .A2(n12188), .B1(n13011), .B2(n11666), .ZN(
        n11572) );
  OAI21_X1 U14134 ( .B1(n15653), .B2(n12989), .A(n11572), .ZN(n11573) );
  AOI21_X1 U14135 ( .B1(n13013), .B2(n15655), .A(n11573), .ZN(n11574) );
  OAI211_X1 U14136 ( .C1(n13007), .C2(n15660), .A(n11575), .B(n11574), .ZN(
        P3_U3226) );
  NAND2_X1 U14137 ( .A1(n11576), .A2(n11627), .ZN(n11580) );
  XNOR2_X1 U14138 ( .A(n6752), .B(n13379), .ZN(n11578) );
  AND2_X1 U14139 ( .A1(n13824), .A2(n13300), .ZN(n11577) );
  NOR2_X1 U14140 ( .A1(n11578), .A2(n11577), .ZN(n11617) );
  NAND2_X1 U14141 ( .A1(n11578), .A2(n11577), .ZN(n11680) );
  INV_X1 U14142 ( .A(n11680), .ZN(n11622) );
  NOR2_X1 U14143 ( .A1(n11617), .A2(n11622), .ZN(n11579) );
  NAND2_X1 U14144 ( .A1(n11580), .A2(n11579), .ZN(n11681) );
  OAI211_X1 U14145 ( .C1(n11580), .C2(n11579), .A(n11681), .B(n13487), .ZN(
        n11587) );
  OAI21_X1 U14146 ( .B1(n13492), .B2(n11582), .A(n11581), .ZN(n11585) );
  NOR2_X1 U14147 ( .A1(n13459), .A2(n11583), .ZN(n11584) );
  AOI211_X1 U14148 ( .C1(n13474), .C2(n13823), .A(n11585), .B(n11584), .ZN(
        n11586) );
  OAI211_X1 U14149 ( .C1(n11588), .C2(n13498), .A(n11587), .B(n11586), .ZN(
        P2_U3185) );
  OAI21_X1 U14150 ( .B1(n11591), .B2(n11590), .A(n11589), .ZN(n11592) );
  NAND2_X1 U14151 ( .A1(n11592), .A2(n14462), .ZN(n11597) );
  INV_X1 U14152 ( .A(n15396), .ZN(n11594) );
  OAI21_X1 U14153 ( .B1(n14433), .B2(n11594), .A(n11593), .ZN(n11595) );
  AOI21_X1 U14154 ( .B1(n14496), .B2(n15397), .A(n11595), .ZN(n11596) );
  OAI211_X1 U14155 ( .C1(n14494), .C2(n11598), .A(n11597), .B(n11596), .ZN(
        P1_U3221) );
  XNOR2_X1 U14156 ( .A(n11600), .B(n11599), .ZN(n11616) );
  OAI21_X1 U14157 ( .B1(n11603), .B2(n11602), .A(n11601), .ZN(n11604) );
  NAND2_X1 U14158 ( .A1(n11604), .A2(n12675), .ZN(n11606) );
  NOR2_X1 U14159 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n6702), .ZN(n11751) );
  AOI21_X1 U14160 ( .B1(n15581), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n11751), 
        .ZN(n11605) );
  OAI211_X1 U14161 ( .C1(n12682), .C2(n11607), .A(n11606), .B(n11605), .ZN(
        n11608) );
  INV_X1 U14162 ( .A(n11608), .ZN(n11615) );
  AND3_X1 U14163 ( .A1(n11611), .A2(n11610), .A3(n11609), .ZN(n11612) );
  OAI21_X1 U14164 ( .B1(n11613), .B2(n11612), .A(n12744), .ZN(n11614) );
  OAI211_X1 U14165 ( .C1(n11616), .C2(n12750), .A(n11615), .B(n11614), .ZN(
        P3_U3192) );
  XNOR2_X1 U14166 ( .A(n13567), .B(n13314), .ZN(n11683) );
  NAND2_X1 U14167 ( .A1(n13823), .A2(n13300), .ZN(n11621) );
  INV_X1 U14168 ( .A(n11619), .ZN(n11628) );
  INV_X1 U14169 ( .A(n11683), .ZN(n11624) );
  NAND2_X1 U14170 ( .A1(n11680), .A2(n11621), .ZN(n11623) );
  INV_X1 U14171 ( .A(n11621), .ZN(n11682) );
  AOI22_X1 U14172 ( .A1(n11624), .A2(n11623), .B1(n11622), .B2(n11682), .ZN(
        n11625) );
  NAND2_X1 U14173 ( .A1(n13822), .A2(n13300), .ZN(n11771) );
  XNOR2_X1 U14174 ( .A(n14301), .B(n13379), .ZN(n11770) );
  XOR2_X1 U14175 ( .A(n11771), .B(n11770), .Z(n11769) );
  XNOR2_X1 U14176 ( .A(n11768), .B(n11769), .ZN(n11629) );
  NAND2_X1 U14177 ( .A1(n11629), .A2(n13487), .ZN(n11635) );
  INV_X1 U14178 ( .A(n13823), .ZN(n11631) );
  OAI21_X1 U14179 ( .B1(n13492), .B2(n11631), .A(n11630), .ZN(n11633) );
  NOR2_X1 U14180 ( .A1(n13459), .A2(n11764), .ZN(n11632) );
  AOI211_X1 U14181 ( .C1(n13474), .C2(n13821), .A(n11633), .B(n11632), .ZN(
        n11634) );
  OAI211_X1 U14182 ( .C1(n7920), .C2(n13498), .A(n11635), .B(n11634), .ZN(
        P2_U3203) );
  XNOR2_X1 U14183 ( .A(n12057), .B(n12463), .ZN(n11745) );
  XNOR2_X1 U14184 ( .A(n11745), .B(n12643), .ZN(n11654) );
  XNOR2_X1 U14185 ( .A(n12463), .B(n13127), .ZN(n11645) );
  XNOR2_X1 U14186 ( .A(n11645), .B(n15655), .ZN(n11796) );
  NAND2_X1 U14187 ( .A1(n11642), .A2(n15653), .ZN(n11637) );
  NAND2_X1 U14188 ( .A1(n11640), .A2(n11639), .ZN(n11650) );
  INV_X1 U14189 ( .A(n11796), .ZN(n11644) );
  INV_X1 U14190 ( .A(n11794), .ZN(n11641) );
  OAI21_X1 U14191 ( .B1(n11644), .B2(n15643), .A(n11641), .ZN(n11648) );
  INV_X1 U14192 ( .A(n11642), .ZN(n11643) );
  NAND2_X1 U14193 ( .A1(n11643), .A2(n15630), .ZN(n11661) );
  OAI21_X1 U14194 ( .B1(n11644), .B2(n11661), .A(n11794), .ZN(n11647) );
  INV_X1 U14195 ( .A(n11645), .ZN(n11646) );
  AOI22_X1 U14196 ( .A1(n11648), .A2(n11647), .B1(n11646), .B2(n15655), .ZN(
        n11649) );
  INV_X1 U14197 ( .A(n11749), .ZN(n11652) );
  AOI21_X1 U14198 ( .B1(n11654), .B2(n11653), .A(n11652), .ZN(n11660) );
  NOR2_X1 U14199 ( .A1(n12593), .A2(n11663), .ZN(n11655) );
  AOI211_X1 U14200 ( .C1(n12511), .C2(n12998), .A(n11656), .B(n11655), .ZN(
        n11657) );
  OAI21_X1 U14201 ( .B1(n12610), .B2(n12057), .A(n11657), .ZN(n11658) );
  AOI21_X1 U14202 ( .B1(n11922), .B2(n12630), .A(n11658), .ZN(n11659) );
  OAI21_X1 U14203 ( .B1(n11660), .B2(n12634), .A(n11659), .ZN(P3_U3171) );
  NAND2_X1 U14204 ( .A1(n11662), .A2(n11661), .ZN(n11795) );
  XNOR2_X1 U14205 ( .A(n11795), .B(n11794), .ZN(n11669) );
  OAI22_X1 U14206 ( .A1(n11663), .A2(n12628), .B1(n12593), .B2(n15653), .ZN(
        n11664) );
  AOI211_X1 U14207 ( .C1(n12188), .C2(n12631), .A(n11665), .B(n11664), .ZN(
        n11668) );
  NAND2_X1 U14208 ( .A1(n12630), .A2(n11666), .ZN(n11667) );
  OAI211_X1 U14209 ( .C1(n11669), .C2(n12634), .A(n11668), .B(n11667), .ZN(
        P3_U3153) );
  NAND2_X1 U14210 ( .A1(n11671), .A2(n11670), .ZN(n13877) );
  XNOR2_X1 U14211 ( .A(n13877), .B(n13884), .ZN(n13876) );
  XNOR2_X1 U14212 ( .A(n13876), .B(P2_REG2_REG_15__SCAN_IN), .ZN(n11679) );
  INV_X1 U14213 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n14292) );
  INV_X1 U14214 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14285) );
  XNOR2_X1 U14215 ( .A(n13883), .B(n14285), .ZN(n11677) );
  AND2_X1 U14216 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n13494) );
  AOI21_X1 U14217 ( .B1(n15468), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n13494), 
        .ZN(n11675) );
  OAI21_X1 U14218 ( .B1(n15465), .B2(n7307), .A(n11675), .ZN(n11676) );
  AOI21_X1 U14219 ( .B1(n11677), .B2(n15475), .A(n11676), .ZN(n11678) );
  OAI21_X1 U14220 ( .B1(n15444), .B2(n11679), .A(n11678), .ZN(P2_U3229) );
  NAND2_X1 U14221 ( .A1(n11681), .A2(n11680), .ZN(n11685) );
  XNOR2_X1 U14222 ( .A(n11683), .B(n11682), .ZN(n11684) );
  XNOR2_X1 U14223 ( .A(n11685), .B(n11684), .ZN(n11692) );
  NAND2_X1 U14224 ( .A1(n13822), .A2(n14190), .ZN(n11687) );
  NAND2_X1 U14225 ( .A1(n13824), .A2(n14188), .ZN(n11686) );
  AND2_X1 U14226 ( .A1(n11687), .A2(n11686), .ZN(n11702) );
  OAI21_X1 U14227 ( .B1(n13461), .B2(n11702), .A(n11688), .ZN(n11690) );
  NOR2_X1 U14228 ( .A1(n13459), .A2(n11697), .ZN(n11689) );
  AOI211_X1 U14229 ( .C1(n13567), .C2(n13479), .A(n11690), .B(n11689), .ZN(
        n11691) );
  OAI21_X1 U14230 ( .B1(n11692), .B2(n13481), .A(n11691), .ZN(P2_U3193) );
  OR2_X1 U14231 ( .A1(n11693), .A2(n13766), .ZN(n11759) );
  INV_X1 U14232 ( .A(n11759), .ZN(n11694) );
  AOI21_X1 U14233 ( .B1(n13766), .B2(n11693), .A(n11694), .ZN(n11714) );
  AOI21_X1 U14234 ( .B1(n11695), .B2(n13567), .A(n15561), .ZN(n11696) );
  NAND2_X1 U14235 ( .A1(n11696), .A2(n11763), .ZN(n11711) );
  INV_X1 U14236 ( .A(n11697), .ZN(n11698) );
  INV_X1 U14237 ( .A(n15503), .ZN(n15825) );
  AOI22_X1 U14238 ( .A1(n15827), .A2(n13567), .B1(n11698), .B2(n15825), .ZN(
        n11699) );
  OAI21_X1 U14239 ( .B1(n11711), .B2(n15829), .A(n11699), .ZN(n11705) );
  OAI211_X1 U14240 ( .C1(n11701), .C2(n13766), .A(n11700), .B(n15556), .ZN(
        n11703) );
  NAND2_X1 U14241 ( .A1(n11703), .A2(n11702), .ZN(n11713) );
  MUX2_X1 U14242 ( .A(n11713), .B(P2_REG2_REG_8__SCAN_IN), .S(n14180), .Z(
        n11704) );
  AOI211_X1 U14243 ( .C1(n11714), .C2(n14134), .A(n11705), .B(n11704), .ZN(
        n11706) );
  INV_X1 U14244 ( .A(n11706), .ZN(P2_U3257) );
  INV_X1 U14245 ( .A(n11707), .ZN(n11709) );
  OAI222_X1 U14246 ( .A1(P2_U3088), .A2(n13744), .B1(n14374), .B2(n11709), 
        .C1(n15733), .C2(n14372), .ZN(P2_U3306) );
  OAI222_X1 U14247 ( .A1(n11710), .A2(P1_U3086), .B1(n15169), .B2(n11709), 
        .C1(n11708), .C2(n15164), .ZN(P1_U3334) );
  OAI21_X1 U14248 ( .B1(n7921), .B2(n15565), .A(n11711), .ZN(n11712) );
  AOI211_X1 U14249 ( .C1(n11714), .C2(n14271), .A(n11713), .B(n11712), .ZN(
        n11717) );
  NAND2_X1 U14250 ( .A1(n15578), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n11715) );
  OAI21_X1 U14251 ( .B1(n11717), .B2(n15578), .A(n11715), .ZN(P2_U3507) );
  NAND2_X1 U14252 ( .A1(n15569), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n11716) );
  OAI21_X1 U14253 ( .B1(n11717), .B2(n15569), .A(n11716), .ZN(P2_U3454) );
  XNOR2_X1 U14254 ( .A(n14600), .B(P1_REG1_REG_15__SCAN_IN), .ZN(n11729) );
  INV_X1 U14255 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n11719) );
  NAND2_X1 U14256 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14493)
         );
  OAI21_X1 U14257 ( .B1(n15287), .B2(n11719), .A(n14493), .ZN(n11727) );
  OAI21_X1 U14258 ( .B1(n11722), .B2(n14598), .A(n14590), .ZN(n11723) );
  NOR2_X1 U14259 ( .A1(n11723), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n14592) );
  AOI21_X1 U14260 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n11723), .A(n14592), 
        .ZN(n11725) );
  NOR2_X1 U14261 ( .A1(n11725), .A2(n11724), .ZN(n11726) );
  AOI211_X1 U14262 ( .C1(n15279), .C2(n7339), .A(n11727), .B(n11726), .ZN(
        n11728) );
  OAI21_X1 U14263 ( .B1(n14645), .B2(n11729), .A(n11728), .ZN(P1_U3258) );
  NAND2_X1 U14264 ( .A1(n11733), .A2(n11732), .ZN(n11735) );
  INV_X1 U14265 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n11785) );
  NAND2_X1 U14266 ( .A1(n11785), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n11734) );
  INV_X1 U14267 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n11736) );
  NAND2_X1 U14268 ( .A1(n11736), .A2(P3_ADDR_REG_12__SCAN_IN), .ZN(n11972) );
  INV_X1 U14269 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n11737) );
  NAND2_X1 U14270 ( .A1(n11737), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n11738) );
  AND2_X1 U14271 ( .A1(n11972), .A2(n11738), .ZN(n11740) );
  INV_X1 U14272 ( .A(n11739), .ZN(n11742) );
  INV_X1 U14273 ( .A(n11740), .ZN(n11741) );
  NAND2_X1 U14274 ( .A1(n11742), .A2(n11741), .ZN(n11743) );
  AND2_X1 U14275 ( .A1(n11973), .A2(n11743), .ZN(n11967) );
  XNOR2_X1 U14276 ( .A(n11969), .B(n11967), .ZN(n11966) );
  XNOR2_X1 U14277 ( .A(n11966), .B(n11965), .ZN(SUB_1596_U68) );
  XNOR2_X1 U14278 ( .A(n11744), .B(n12494), .ZN(n11910) );
  XNOR2_X1 U14279 ( .A(n11910), .B(n12998), .ZN(n11747) );
  OR2_X1 U14280 ( .A1(n11745), .A2(n12643), .ZN(n11748) );
  AND2_X1 U14281 ( .A1(n11747), .A2(n11748), .ZN(n11746) );
  AOI21_X1 U14282 ( .B1(n11749), .B2(n11748), .A(n11747), .ZN(n11750) );
  NOR3_X1 U14283 ( .A1(n6640), .A2(n11750), .A3(n12634), .ZN(n11757) );
  AOI21_X1 U14284 ( .B1(n12626), .B2(n12643), .A(n11751), .ZN(n11755) );
  NAND2_X1 U14285 ( .A1(n12630), .A2(n12120), .ZN(n11754) );
  NAND2_X1 U14286 ( .A1(n12631), .A2(n13122), .ZN(n11753) );
  NAND2_X1 U14287 ( .A1(n12511), .A2(n12642), .ZN(n11752) );
  NAND4_X1 U14288 ( .A1(n11755), .A2(n11754), .A3(n11753), .A4(n11752), .ZN(
        n11756) );
  OR2_X1 U14289 ( .A1(n11757), .A2(n11756), .ZN(P3_U3157) );
  XNOR2_X1 U14290 ( .A(n13822), .B(n14301), .ZN(n13768) );
  NAND2_X1 U14291 ( .A1(n11759), .A2(n11758), .ZN(n11760) );
  XOR2_X1 U14292 ( .A(n13768), .B(n11760), .Z(n14304) );
  XOR2_X1 U14293 ( .A(n11761), .B(n13768), .Z(n11762) );
  AOI222_X1 U14294 ( .A1(n15556), .A2(n11762), .B1(n13821), .B2(n14190), .C1(
        n13823), .C2(n14188), .ZN(n14303) );
  MUX2_X1 U14295 ( .A(n10600), .B(n14303), .S(n15831), .Z(n11767) );
  AOI211_X1 U14296 ( .C1(n14301), .C2(n11763), .A(n15561), .B(n11873), .ZN(
        n14300) );
  OAI22_X1 U14297 ( .A1(n15504), .A2(n7920), .B1(n15503), .B2(n11764), .ZN(
        n11765) );
  AOI21_X1 U14298 ( .B1(n14300), .B2(n15484), .A(n11765), .ZN(n11766) );
  OAI211_X1 U14299 ( .C1(n14200), .C2(n14304), .A(n11767), .B(n11766), .ZN(
        P2_U3256) );
  INV_X1 U14300 ( .A(n11770), .ZN(n11772) );
  XNOR2_X1 U14301 ( .A(n13581), .B(n7172), .ZN(n11880) );
  NAND2_X1 U14302 ( .A1(n13821), .A2(n13300), .ZN(n11878) );
  XNOR2_X1 U14303 ( .A(n11880), .B(n11878), .ZN(n11773) );
  OAI211_X1 U14304 ( .C1(n11774), .C2(n11773), .A(n11882), .B(n13487), .ZN(
        n11779) );
  OAI21_X1 U14305 ( .B1(n13492), .B2(n11867), .A(n11775), .ZN(n11777) );
  NOR2_X1 U14306 ( .A1(n13459), .A2(n11871), .ZN(n11776) );
  AOI211_X1 U14307 ( .C1(n13474), .C2(n13820), .A(n11777), .B(n11776), .ZN(
        n11778) );
  OAI211_X1 U14308 ( .C1(n12099), .C2(n13498), .A(n11779), .B(n11778), .ZN(
        P2_U3189) );
  INV_X1 U14309 ( .A(n11842), .ZN(n11780) );
  AOI21_X1 U14310 ( .B1(n13001), .B2(n6644), .A(n11780), .ZN(n11793) );
  OAI21_X1 U14311 ( .B1(n11782), .B2(n11781), .A(n11849), .ZN(n11787) );
  NAND2_X1 U14312 ( .A1(n12751), .A2(n11783), .ZN(n11784) );
  NAND2_X1 U14313 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n11912)
         );
  OAI211_X1 U14314 ( .C1(n12715), .C2(n11785), .A(n11784), .B(n11912), .ZN(
        n11786) );
  AOI21_X1 U14315 ( .B1(n11787), .B2(n12675), .A(n11786), .ZN(n11792) );
  OAI21_X1 U14316 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n11789), .A(n11788), 
        .ZN(n11790) );
  NAND2_X1 U14317 ( .A1(n11790), .A2(n12692), .ZN(n11791) );
  OAI211_X1 U14318 ( .C1(n11793), .C2(n12702), .A(n11792), .B(n11791), .ZN(
        P3_U3193) );
  MUX2_X1 U14319 ( .A(n12644), .B(n11795), .S(n11794), .Z(n11797) );
  XNOR2_X1 U14320 ( .A(n11797), .B(n11796), .ZN(n11802) );
  INV_X1 U14321 ( .A(n12643), .ZN(n13120) );
  OAI22_X1 U14322 ( .A1(n13120), .A2(n12628), .B1(n12593), .B2(n15643), .ZN(
        n11798) );
  AOI211_X1 U14323 ( .C1(n13127), .C2(n12631), .A(n11799), .B(n11798), .ZN(
        n11801) );
  NAND2_X1 U14324 ( .A1(n12630), .A2(n11962), .ZN(n11800) );
  OAI211_X1 U14325 ( .C1(n11802), .C2(n12634), .A(n11801), .B(n11800), .ZN(
        P3_U3161) );
  XOR2_X1 U14326 ( .A(n11803), .B(n13772), .Z(n11806) );
  NAND2_X1 U14327 ( .A1(n13821), .A2(n14188), .ZN(n11805) );
  NAND2_X1 U14328 ( .A1(n14189), .A2(n14190), .ZN(n11804) );
  AND2_X1 U14329 ( .A1(n11805), .A2(n11804), .ZN(n11890) );
  OAI21_X1 U14330 ( .B1(n11806), .B2(n14274), .A(n11890), .ZN(n12091) );
  INV_X1 U14331 ( .A(n12091), .ZN(n11816) );
  INV_X1 U14332 ( .A(n11807), .ZN(n11808) );
  AOI211_X1 U14333 ( .C1(n13585), .C2(n6636), .A(n15561), .B(n11808), .ZN(
        n12092) );
  NOR2_X1 U14334 ( .A1(n15504), .A2(n11809), .ZN(n11812) );
  OAI22_X1 U14335 ( .A1(n15831), .A2(n11810), .B1(n11886), .B2(n15503), .ZN(
        n11811) );
  AOI211_X1 U14336 ( .C1(n12092), .C2(n15484), .A(n11812), .B(n11811), .ZN(
        n11815) );
  XNOR2_X1 U14337 ( .A(n11813), .B(n13772), .ZN(n12093) );
  NAND2_X1 U14338 ( .A1(n12093), .A2(n14134), .ZN(n11814) );
  OAI211_X1 U14339 ( .C1(n11816), .C2(n14180), .A(n11815), .B(n11814), .ZN(
        P2_U3254) );
  INV_X1 U14340 ( .A(n11817), .ZN(n11819) );
  OAI222_X1 U14341 ( .A1(n13250), .A2(n11820), .B1(n13248), .B2(n11819), .C1(
        n11818), .C2(P3_U3151), .ZN(P3_U3271) );
  OR2_X1 U14342 ( .A1(n14504), .A2(n11987), .ZN(n11822) );
  XNOR2_X1 U14343 ( .A(n12027), .B(n11833), .ZN(n15421) );
  INV_X2 U14344 ( .A(n15298), .ZN(n11825) );
  OAI211_X1 U14345 ( .C1(n11825), .C2(n11824), .A(n15328), .B(n12039), .ZN(
        n11826) );
  OAI21_X1 U14346 ( .B1(n12071), .B2(n14980), .A(n11826), .ZN(n15415) );
  AOI22_X1 U14347 ( .A1(n15336), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n11952), 
        .B2(n15324), .ZN(n11827) );
  OAI21_X1 U14348 ( .B1(n15311), .B2(n11824), .A(n11827), .ZN(n11835) );
  OR2_X1 U14349 ( .A1(n11983), .A2(n15397), .ZN(n11830) );
  NAND2_X1 U14350 ( .A1(n6652), .A2(n11833), .ZN(n12048) );
  OAI211_X1 U14351 ( .C1(n6652), .C2(n11833), .A(n12048), .B(n15359), .ZN(
        n15420) );
  NAND2_X1 U14352 ( .A1(n14504), .A2(n14982), .ZN(n15414) );
  AOI21_X1 U14353 ( .B1(n15420), .B2(n15414), .A(n15336), .ZN(n11834) );
  AOI211_X1 U14354 ( .C1(n15332), .C2(n15415), .A(n11835), .B(n11834), .ZN(
        n11836) );
  OAI21_X1 U14355 ( .B1(n15421), .B2(n14990), .A(n11836), .ZN(P1_U3283) );
  INV_X1 U14356 ( .A(n11860), .ZN(n11839) );
  AOI21_X1 U14357 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n15155), .A(n11837), 
        .ZN(n11838) );
  OAI21_X1 U14358 ( .B1(n11839), .B2(n15169), .A(n11838), .ZN(P1_U3332) );
  AND3_X1 U14359 ( .A1(n11842), .A2(n11841), .A3(n11840), .ZN(n11843) );
  OAI21_X1 U14360 ( .B1(n11844), .B2(n11843), .A(n12744), .ZN(n11858) );
  OAI21_X1 U14361 ( .B1(n11847), .B2(n11846), .A(n11845), .ZN(n11856) );
  AND2_X1 U14362 ( .A1(n11849), .A2(n11848), .ZN(n11851) );
  OAI211_X1 U14363 ( .C1(n11851), .C2(n11850), .A(n12675), .B(n12653), .ZN(
        n11853) );
  AND2_X1 U14364 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n12085) );
  AOI21_X1 U14365 ( .B1(n15581), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n12085), 
        .ZN(n11852) );
  OAI211_X1 U14366 ( .C1(n12682), .C2(n11854), .A(n11853), .B(n11852), .ZN(
        n11855) );
  AOI21_X1 U14367 ( .B1(n12692), .B2(n11856), .A(n11855), .ZN(n11857) );
  NAND2_X1 U14368 ( .A1(n11858), .A2(n11857), .ZN(P3_U3194) );
  NAND2_X1 U14369 ( .A1(n11860), .A2(n11859), .ZN(n11862) );
  OR2_X1 U14370 ( .A1(n11861), .A2(P2_U3088), .ZN(n13805) );
  OAI211_X1 U14371 ( .C1(n11863), .C2(n14372), .A(n11862), .B(n13805), .ZN(
        P2_U3304) );
  XNOR2_X1 U14372 ( .A(n13581), .B(n13821), .ZN(n13771) );
  XOR2_X1 U14373 ( .A(n11864), .B(n13771), .Z(n12097) );
  XOR2_X1 U14374 ( .A(n11865), .B(n13771), .Z(n11869) );
  OAI22_X1 U14375 ( .A1(n11867), .A2(n15495), .B1(n11866), .B2(n15493), .ZN(
        n11868) );
  AOI21_X1 U14376 ( .B1(n11869), .B2(n15556), .A(n11868), .ZN(n11870) );
  OAI21_X1 U14377 ( .B1(n12097), .B2(n15501), .A(n11870), .ZN(n12100) );
  NAND2_X1 U14378 ( .A1(n12100), .A2(n15831), .ZN(n11877) );
  OAI22_X1 U14379 ( .A1(n15831), .A2(n11872), .B1(n11871), .B2(n15503), .ZN(
        n11875) );
  OAI211_X1 U14380 ( .C1(n12099), .C2(n11873), .A(n6636), .B(n14181), .ZN(
        n12098) );
  NOR2_X1 U14381 ( .A1(n12098), .A2(n15829), .ZN(n11874) );
  AOI211_X1 U14382 ( .C1(n15827), .C2(n13581), .A(n11875), .B(n11874), .ZN(
        n11876) );
  OAI211_X1 U14383 ( .C1(n12097), .C2(n14172), .A(n11877), .B(n11876), .ZN(
        P2_U3255) );
  INV_X1 U14384 ( .A(n11878), .ZN(n11879) );
  NAND2_X1 U14385 ( .A1(n11880), .A2(n11879), .ZN(n11881) );
  XNOR2_X1 U14386 ( .A(n13585), .B(n13314), .ZN(n11884) );
  NAND2_X1 U14387 ( .A1(n13820), .A2(n15561), .ZN(n11883) );
  NOR2_X1 U14388 ( .A1(n11884), .A2(n11883), .ZN(n12132) );
  NAND2_X1 U14389 ( .A1(n11884), .A2(n11883), .ZN(n12131) );
  NOR2_X1 U14390 ( .A1(n12132), .A2(n7062), .ZN(n11885) );
  XNOR2_X1 U14391 ( .A(n12133), .B(n11885), .ZN(n11893) );
  INV_X1 U14392 ( .A(n11886), .ZN(n11887) );
  NAND2_X1 U14393 ( .A1(n13495), .A2(n11887), .ZN(n11889) );
  OAI211_X1 U14394 ( .C1(n11890), .C2(n13461), .A(n11889), .B(n11888), .ZN(
        n11891) );
  AOI21_X1 U14395 ( .B1(n13585), .B2(n13479), .A(n11891), .ZN(n11892) );
  OAI21_X1 U14396 ( .B1(n11893), .B2(n13481), .A(n11892), .ZN(P2_U3208) );
  XNOR2_X1 U14397 ( .A(n13590), .B(n14189), .ZN(n13773) );
  XNOR2_X1 U14398 ( .A(n11894), .B(n13773), .ZN(n12108) );
  XNOR2_X1 U14399 ( .A(n11895), .B(n13773), .ZN(n12110) );
  NOR2_X1 U14400 ( .A1(n14180), .A2(n14274), .ZN(n14177) );
  NAND2_X1 U14401 ( .A1(n12110), .A2(n14177), .ZN(n11906) );
  AOI21_X1 U14402 ( .B1(n11807), .B2(n13590), .A(n15561), .ZN(n11896) );
  NAND2_X1 U14403 ( .A1(n11896), .A2(n14194), .ZN(n12106) );
  INV_X1 U14404 ( .A(n12106), .ZN(n11904) );
  NAND2_X1 U14405 ( .A1(n13820), .A2(n14188), .ZN(n11898) );
  NAND2_X1 U14406 ( .A1(n13819), .A2(n14190), .ZN(n11897) );
  NAND2_X1 U14407 ( .A1(n11898), .A2(n11897), .ZN(n12137) );
  OAI22_X1 U14408 ( .A1(n15831), .A2(n11899), .B1(n12140), .B2(n15503), .ZN(
        n11900) );
  AOI21_X1 U14409 ( .B1(n15831), .B2(n12137), .A(n11900), .ZN(n11901) );
  OAI21_X1 U14410 ( .B1(n11902), .B2(n15504), .A(n11901), .ZN(n11903) );
  AOI21_X1 U14411 ( .B1(n11904), .B2(n15484), .A(n11903), .ZN(n11905) );
  OAI211_X1 U14412 ( .C1(n12108), .C2(n14200), .A(n11906), .B(n11905), .ZN(
        P2_U3253) );
  INV_X1 U14413 ( .A(n11907), .ZN(n11908) );
  OAI222_X1 U14414 ( .A1(n14372), .A2(n11909), .B1(P2_U3088), .B2(n8559), .C1(
        n14374), .C2(n11908), .ZN(P2_U3305) );
  INV_X1 U14415 ( .A(n11910), .ZN(n11911) );
  XNOR2_X1 U14416 ( .A(n13002), .B(n12494), .ZN(n12078) );
  XNOR2_X1 U14417 ( .A(n11991), .B(n12078), .ZN(n12080) );
  XNOR2_X1 U14418 ( .A(n12080), .B(n12642), .ZN(n11917) );
  NOR2_X1 U14419 ( .A1(n12610), .A2(n13002), .ZN(n11915) );
  NAND2_X1 U14420 ( .A1(n12626), .A2(n12998), .ZN(n11913) );
  OAI211_X1 U14421 ( .C1(n11996), .C2(n12628), .A(n11913), .B(n11912), .ZN(
        n11914) );
  AOI211_X1 U14422 ( .C1(n13003), .C2(n12630), .A(n11915), .B(n11914), .ZN(
        n11916) );
  OAI21_X1 U14423 ( .B1(n11917), .B2(n12634), .A(n11916), .ZN(P3_U3176) );
  INV_X1 U14424 ( .A(n11920), .ZN(n12332) );
  XNOR2_X1 U14425 ( .A(n11918), .B(n12332), .ZN(n12059) );
  INV_X1 U14426 ( .A(n12059), .ZN(n11929) );
  OAI211_X1 U14427 ( .C1(n11921), .C2(n11920), .A(n11919), .B(n15611), .ZN(
        n12056) );
  OR2_X1 U14428 ( .A1(n12056), .A2(n15601), .ZN(n11927) );
  AOI22_X1 U14429 ( .A1(n15601), .A2(P3_REG2_REG_9__SCAN_IN), .B1(n13011), 
        .B2(n11922), .ZN(n11926) );
  INV_X1 U14430 ( .A(n12989), .ZN(n13009) );
  AOI22_X1 U14431 ( .A1(n13013), .A2(n12998), .B1(n13009), .B2(n15655), .ZN(
        n11925) );
  NAND2_X1 U14432 ( .A1(n13004), .A2(n11923), .ZN(n11924) );
  AND4_X1 U14433 ( .A1(n11927), .A2(n11926), .A3(n11925), .A4(n11924), .ZN(
        n11928) );
  OAI21_X1 U14434 ( .B1(n13007), .B2(n11929), .A(n11928), .ZN(P3_U3224) );
  INV_X1 U14435 ( .A(n11930), .ZN(n11931) );
  AOI21_X1 U14436 ( .B1(n11933), .B2(n11932), .A(n11931), .ZN(n11940) );
  INV_X1 U14437 ( .A(n12041), .ZN(n11937) );
  NAND2_X1 U14438 ( .A1(n14983), .A2(n14903), .ZN(n11934) );
  OAI21_X1 U14439 ( .B1(n11981), .B2(n14931), .A(n11934), .ZN(n12050) );
  NAND2_X1 U14440 ( .A1(n14491), .A2(n12050), .ZN(n11935) );
  OAI211_X1 U14441 ( .C1(n14494), .C2(n11937), .A(n11936), .B(n11935), .ZN(
        n11938) );
  AOI21_X1 U14442 ( .B1(n14496), .B2(n15126), .A(n11938), .ZN(n11939) );
  OAI21_X1 U14443 ( .B1(n11940), .B2(n14498), .A(n11939), .ZN(P1_U3236) );
  XOR2_X1 U14444 ( .A(n11942), .B(n11941), .Z(n11978) );
  AOI22_X1 U14445 ( .A1(n11978), .A2(n11979), .B1(n11942), .B2(n11941), .ZN(
        n11947) );
  OAI21_X1 U14446 ( .B1(n11945), .B2(n11944), .A(n11943), .ZN(n11946) );
  XNOR2_X1 U14447 ( .A(n11947), .B(n11946), .ZN(n11954) );
  NAND2_X1 U14448 ( .A1(n14478), .A2(n14504), .ZN(n11949) );
  OAI211_X1 U14449 ( .C1(n12071), .C2(n14482), .A(n11949), .B(n11948), .ZN(
        n11951) );
  NOR2_X1 U14450 ( .A1(n14468), .A2(n11824), .ZN(n11950) );
  AOI211_X1 U14451 ( .C1(n14479), .C2(n11952), .A(n11951), .B(n11950), .ZN(
        n11953) );
  OAI21_X1 U14452 ( .B1(n11954), .B2(n14498), .A(n11953), .ZN(P1_U3217) );
  XOR2_X1 U14453 ( .A(n11955), .B(n12326), .Z(n13129) );
  INV_X1 U14454 ( .A(n11956), .ZN(n11957) );
  AOI21_X1 U14455 ( .B1(n12326), .B2(n11958), .A(n11957), .ZN(n11959) );
  OAI222_X1 U14456 ( .A1(n15652), .A2(n15643), .B1(n15642), .B2(n13120), .C1(
        n13052), .C2(n11959), .ZN(n13126) );
  INV_X1 U14457 ( .A(n13126), .ZN(n11960) );
  MUX2_X1 U14458 ( .A(n11961), .B(n11960), .S(n15599), .Z(n11964) );
  AOI22_X1 U14459 ( .A1(n13004), .A2(n13127), .B1(n13011), .B2(n11962), .ZN(
        n11963) );
  OAI211_X1 U14460 ( .C1(n13007), .C2(n13129), .A(n11964), .B(n11963), .ZN(
        P3_U3225) );
  NAND2_X1 U14461 ( .A1(n11966), .A2(n11965), .ZN(n11971) );
  INV_X1 U14462 ( .A(n11967), .ZN(n11968) );
  OR2_X1 U14463 ( .A1(n11969), .A2(n11968), .ZN(n11970) );
  NAND2_X1 U14464 ( .A1(n11971), .A2(n11970), .ZN(n11976) );
  INV_X1 U14465 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15187) );
  XNOR2_X1 U14466 ( .A(n15187), .B(P1_ADDR_REG_13__SCAN_IN), .ZN(n11974) );
  XNOR2_X1 U14467 ( .A(n15189), .B(n11974), .ZN(n11975) );
  OR2_X2 U14468 ( .A1(n11976), .A2(n11975), .ZN(n15185) );
  NAND2_X1 U14469 ( .A1(n11976), .A2(n11975), .ZN(n15186) );
  NAND2_X1 U14470 ( .A1(n15185), .A2(n15186), .ZN(n11977) );
  XNOR2_X1 U14471 ( .A(n11977), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  INV_X1 U14472 ( .A(n15295), .ZN(n11990) );
  XOR2_X1 U14473 ( .A(n11979), .B(n11978), .Z(n11980) );
  NAND2_X1 U14474 ( .A1(n11980), .A2(n14462), .ZN(n11989) );
  OR2_X1 U14475 ( .A1(n11981), .A2(n14980), .ZN(n11982) );
  OAI21_X1 U14476 ( .B1(n11983), .B2(n14931), .A(n11982), .ZN(n15294) );
  NAND2_X1 U14477 ( .A1(n14491), .A2(n15294), .ZN(n11985) );
  NAND2_X1 U14478 ( .A1(n11985), .A2(n11984), .ZN(n11986) );
  AOI21_X1 U14479 ( .B1(n14496), .B2(n11987), .A(n11986), .ZN(n11988) );
  OAI211_X1 U14480 ( .C1(n14494), .C2(n11990), .A(n11989), .B(n11988), .ZN(
        P1_U3231) );
  XNOR2_X1 U14481 ( .A(n13111), .B(n12494), .ZN(n11995) );
  NAND2_X1 U14482 ( .A1(n11995), .A2(n12999), .ZN(n12082) );
  OAI21_X1 U14483 ( .B1(n13119), .B2(n12078), .A(n12082), .ZN(n11992) );
  INV_X1 U14484 ( .A(n11992), .ZN(n11993) );
  NAND3_X1 U14485 ( .A1(n12082), .A2(n13119), .A3(n12078), .ZN(n11998) );
  INV_X1 U14486 ( .A(n11995), .ZN(n11997) );
  NAND2_X1 U14487 ( .A1(n11997), .A2(n11996), .ZN(n12081) );
  AND2_X1 U14488 ( .A1(n11998), .A2(n12081), .ZN(n11999) );
  XNOR2_X1 U14489 ( .A(n13206), .B(n12463), .ZN(n12000) );
  AND2_X1 U14490 ( .A1(n12000), .A2(n12985), .ZN(n12465) );
  INV_X1 U14491 ( .A(n12465), .ZN(n12002) );
  INV_X1 U14492 ( .A(n12000), .ZN(n12001) );
  NAND2_X1 U14493 ( .A1(n12001), .A2(n12967), .ZN(n12464) );
  NAND2_X1 U14494 ( .A1(n12002), .A2(n12464), .ZN(n12003) );
  XNOR2_X1 U14495 ( .A(n12466), .B(n12003), .ZN(n12008) );
  AND2_X1 U14496 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n12656) );
  AOI21_X1 U14497 ( .B1(n12626), .B2(n12999), .A(n12656), .ZN(n12005) );
  NAND2_X1 U14498 ( .A1(n12630), .A2(n12979), .ZN(n12004) );
  OAI211_X1 U14499 ( .C1(n12953), .C2(n12628), .A(n12005), .B(n12004), .ZN(
        n12006) );
  AOI21_X1 U14500 ( .B1(n13206), .B2(n12631), .A(n12006), .ZN(n12007) );
  OAI21_X1 U14501 ( .B1(n12008), .B2(n12634), .A(n12007), .ZN(P3_U3174) );
  AOI21_X1 U14502 ( .B1(n12071), .B2(n15126), .A(n12009), .ZN(n12010) );
  NAND2_X1 U14503 ( .A1(n12046), .A2(n12071), .ZN(n12011) );
  AOI22_X1 U14504 ( .A1(n7772), .A2(n12011), .B1(n12043), .B2(n14502), .ZN(
        n12012) );
  OR2_X1 U14505 ( .A1(n15121), .A2(n12013), .ZN(n12014) );
  INV_X1 U14506 ( .A(n14979), .ZN(n12015) );
  NOR2_X1 U14507 ( .A1(n12015), .A2(n12030), .ZN(n12016) );
  NOR2_X1 U14508 ( .A1(n15116), .A2(n14661), .ZN(n14664) );
  OAI21_X1 U14509 ( .B1(n12016), .B2(n14664), .A(n12034), .ZN(n12020) );
  INV_X1 U14510 ( .A(n12016), .ZN(n14978) );
  NOR2_X1 U14511 ( .A1(n12034), .A2(n14664), .ZN(n12017) );
  AOI21_X1 U14512 ( .B1(n14978), .B2(n12017), .A(n15400), .ZN(n12019) );
  OAI22_X1 U14513 ( .A1(n12018), .A2(n14980), .B1(n14661), .B2(n14931), .ZN(
        n14383) );
  AOI21_X1 U14514 ( .B1(n12020), .B2(n12019), .A(n14383), .ZN(n15113) );
  NOR2_X2 U14515 ( .A1(n14973), .A2(n15107), .ZN(n12021) );
  INV_X1 U14516 ( .A(n12021), .ZN(n14961) );
  NAND2_X1 U14517 ( .A1(n14973), .A2(n15107), .ZN(n12022) );
  AND2_X1 U14518 ( .A1(n14961), .A2(n12022), .ZN(n15108) );
  INV_X1 U14519 ( .A(n14840), .ZN(n14996) );
  NAND2_X1 U14520 ( .A1(n15107), .A2(n14995), .ZN(n12024) );
  AOI22_X1 U14521 ( .A1(n15336), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n14381), 
        .B2(n15324), .ZN(n12023) );
  NAND2_X1 U14522 ( .A1(n12024), .A2(n12023), .ZN(n12025) );
  AOI21_X1 U14523 ( .B1(n15108), .B2(n14996), .A(n12025), .ZN(n12037) );
  OR2_X1 U14524 ( .A1(n15417), .A2(n14503), .ZN(n12028) );
  OR2_X1 U14525 ( .A1(n15121), .A2(n14983), .ZN(n12029) );
  OR2_X1 U14526 ( .A1(n15116), .A2(n14501), .ZN(n12032) );
  NAND2_X1 U14527 ( .A1(n12033), .A2(n12032), .ZN(n12035) );
  NAND2_X1 U14528 ( .A1(n12035), .A2(n12034), .ZN(n15109) );
  NAND3_X1 U14529 ( .A1(n15110), .A2(n15109), .A3(n14992), .ZN(n12036) );
  OAI211_X1 U14530 ( .C1(n15113), .C2(n15336), .A(n12037), .B(n12036), .ZN(
        P1_U3279) );
  XOR2_X1 U14531 ( .A(n12038), .B(n12045), .Z(n15129) );
  AOI21_X1 U14532 ( .B1(n12039), .B2(n15126), .A(n15344), .ZN(n12040) );
  AND2_X1 U14533 ( .A1(n12065), .A2(n12040), .ZN(n15125) );
  AOI22_X1 U14534 ( .A1(n15336), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n12041), 
        .B2(n15324), .ZN(n12042) );
  OAI21_X1 U14535 ( .B1(n15311), .B2(n7772), .A(n12042), .ZN(n12053) );
  INV_X1 U14536 ( .A(n12045), .ZN(n12044) );
  NOR2_X1 U14537 ( .A1(n12044), .A2(n12043), .ZN(n12049) );
  AOI21_X1 U14538 ( .B1(n12048), .B2(n12046), .A(n12045), .ZN(n12047) );
  AOI211_X1 U14539 ( .C1(n12049), .C2(n12048), .A(n15400), .B(n12047), .ZN(
        n12051) );
  NOR2_X1 U14540 ( .A1(n12051), .A2(n12050), .ZN(n15128) );
  NOR2_X1 U14541 ( .A1(n15128), .A2(n15336), .ZN(n12052) );
  AOI211_X1 U14542 ( .C1(n15125), .C2(n15332), .A(n12053), .B(n12052), .ZN(
        n12054) );
  OAI21_X1 U14543 ( .B1(n14990), .B2(n15129), .A(n12054), .ZN(P1_U3282) );
  INV_X1 U14544 ( .A(n13138), .ZN(n15602) );
  AOI22_X1 U14545 ( .A1(n15655), .A2(n15638), .B1(n15656), .B2(n12998), .ZN(
        n12055) );
  OAI211_X1 U14546 ( .C1(n15651), .C2(n12057), .A(n12056), .B(n12055), .ZN(
        n12058) );
  AOI21_X1 U14547 ( .B1(n12059), .B2(n15602), .A(n12058), .ZN(n12062) );
  NAND2_X1 U14548 ( .A1(n15674), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n12060) );
  OAI21_X1 U14549 ( .B1(n12062), .B2(n15674), .A(n12060), .ZN(P3_U3468) );
  NAND2_X1 U14550 ( .A1(n15664), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n12061) );
  OAI21_X1 U14551 ( .B1(n12062), .B2(n15664), .A(n12061), .ZN(P3_U3417) );
  XNOR2_X1 U14552 ( .A(n12064), .B(n12063), .ZN(n15124) );
  NAND2_X1 U14553 ( .A1(n12065), .A2(n15121), .ZN(n12066) );
  NAND2_X1 U14554 ( .A1(n12066), .A2(n15328), .ZN(n12067) );
  NOR2_X1 U14555 ( .A1(n14972), .A2(n12067), .ZN(n15120) );
  AOI22_X1 U14556 ( .A1(n15336), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n14418), 
        .B2(n15324), .ZN(n12068) );
  OAI21_X1 U14557 ( .B1(n15311), .B2(n7770), .A(n12068), .ZN(n12076) );
  INV_X1 U14558 ( .A(n12069), .ZN(n12070) );
  AOI21_X1 U14559 ( .B1(n12070), .B2(n7134), .A(n15400), .ZN(n12074) );
  OR2_X1 U14560 ( .A1(n12071), .A2(n14931), .ZN(n12072) );
  OAI21_X1 U14561 ( .B1(n14661), .B2(n14980), .A(n12072), .ZN(n14421) );
  AOI21_X1 U14562 ( .B1(n12074), .B2(n12073), .A(n14421), .ZN(n15123) );
  NOR2_X1 U14563 ( .A1(n15123), .A2(n15336), .ZN(n12075) );
  AOI211_X1 U14564 ( .C1(n15120), .C2(n15332), .A(n12076), .B(n12075), .ZN(
        n12077) );
  OAI21_X1 U14565 ( .B1(n14990), .B2(n15124), .A(n12077), .ZN(P1_U3281) );
  INV_X1 U14566 ( .A(n12078), .ZN(n12079) );
  AOI22_X1 U14567 ( .A1(n12080), .A2(n12642), .B1(n11991), .B2(n12079), .ZN(
        n12084) );
  NAND2_X1 U14568 ( .A1(n12082), .A2(n12081), .ZN(n12083) );
  XNOR2_X1 U14569 ( .A(n12084), .B(n12083), .ZN(n12090) );
  AOI21_X1 U14570 ( .B1(n12626), .B2(n12642), .A(n12085), .ZN(n12087) );
  NAND2_X1 U14571 ( .A1(n12630), .A2(n12987), .ZN(n12086) );
  OAI211_X1 U14572 ( .C1(n12985), .C2(n12628), .A(n12087), .B(n12086), .ZN(
        n12088) );
  AOI21_X1 U14573 ( .B1(n13111), .B2(n12631), .A(n12088), .ZN(n12089) );
  OAI21_X1 U14574 ( .B1(n12090), .B2(n12634), .A(n12089), .ZN(P3_U3164) );
  AOI211_X1 U14575 ( .C1(n14271), .C2(n12093), .A(n12092), .B(n12091), .ZN(
        n12096) );
  AOI22_X1 U14576 ( .A1(n14280), .A2(n13585), .B1(P2_REG1_REG_11__SCAN_IN), 
        .B2(n15578), .ZN(n12094) );
  OAI21_X1 U14577 ( .B1(n12096), .B2(n15578), .A(n12094), .ZN(P2_U3510) );
  AOI22_X1 U14578 ( .A1(n10258), .A2(n13585), .B1(P2_REG0_REG_11__SCAN_IN), 
        .B2(n15569), .ZN(n12095) );
  OAI21_X1 U14579 ( .B1(n12096), .B2(n15569), .A(n12095), .ZN(P2_U3463) );
  INV_X1 U14580 ( .A(n12097), .ZN(n12102) );
  OAI21_X1 U14581 ( .B1(n12099), .B2(n15565), .A(n12098), .ZN(n12101) );
  AOI211_X1 U14582 ( .C1(n15560), .C2(n12102), .A(n12101), .B(n12100), .ZN(
        n12105) );
  NAND2_X1 U14583 ( .A1(n15569), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n12103) );
  OAI21_X1 U14584 ( .B1(n12105), .B2(n15569), .A(n12103), .ZN(P2_U3460) );
  NAND2_X1 U14585 ( .A1(n15578), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n12104) );
  OAI21_X1 U14586 ( .B1(n12105), .B2(n15578), .A(n12104), .ZN(P2_U3509) );
  AOI21_X1 U14587 ( .B1(n13590), .B2(n15525), .A(n12137), .ZN(n12107) );
  OAI211_X1 U14588 ( .C1(n12108), .C2(n14310), .A(n12107), .B(n12106), .ZN(
        n12109) );
  AOI21_X1 U14589 ( .B1(n15556), .B2(n12110), .A(n12109), .ZN(n12113) );
  NAND2_X1 U14590 ( .A1(n15578), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n12111) );
  OAI21_X1 U14591 ( .B1(n12113), .B2(n15578), .A(n12111), .ZN(P2_U3511) );
  NAND2_X1 U14592 ( .A1(n15569), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n12112) );
  OAI21_X1 U14593 ( .B1(n12113), .B2(n15569), .A(n12112), .ZN(P2_U3466) );
  INV_X1 U14594 ( .A(n12114), .ZN(n12126) );
  OAI222_X1 U14595 ( .A1(n12116), .A2(P1_U3086), .B1(n15169), .B2(n12126), 
        .C1(n12115), .C2(n15164), .ZN(P1_U3331) );
  INV_X1 U14596 ( .A(n12201), .ZN(n12331) );
  XNOR2_X1 U14597 ( .A(n12117), .B(n12331), .ZN(n13125) );
  OAI211_X1 U14598 ( .C1(n12119), .C2(n12201), .A(n12118), .B(n15611), .ZN(
        n13124) );
  OR2_X1 U14599 ( .A1(n13124), .A2(n15601), .ZN(n12124) );
  AOI22_X1 U14600 ( .A1(n15601), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n13011), 
        .B2(n12120), .ZN(n12123) );
  AOI22_X1 U14601 ( .A1(n13013), .A2(n12642), .B1(n13009), .B2(n12643), .ZN(
        n12122) );
  NAND2_X1 U14602 ( .A1(n13004), .A2(n13122), .ZN(n12121) );
  AND4_X1 U14603 ( .A1(n12124), .A2(n12123), .A3(n12122), .A4(n12121), .ZN(
        n12125) );
  OAI21_X1 U14604 ( .B1(n13007), .B2(n13125), .A(n12125), .ZN(P3_U3223) );
  OAI222_X1 U14605 ( .A1(P2_U3088), .A2(n12128), .B1(n14372), .B2(n12127), 
        .C1(n14374), .C2(n12126), .ZN(P2_U3303) );
  AND2_X1 U14606 ( .A1(n14189), .A2(n13300), .ZN(n12130) );
  XNOR2_X1 U14607 ( .A(n13590), .B(n7172), .ZN(n12129) );
  NOR2_X1 U14608 ( .A1(n12129), .A2(n12130), .ZN(n12144) );
  AOI21_X1 U14609 ( .B1(n12130), .B2(n12129), .A(n12144), .ZN(n12135) );
  OAI21_X1 U14610 ( .B1(n12135), .B2(n12134), .A(n12145), .ZN(n12142) );
  INV_X1 U14611 ( .A(n13461), .ZN(n13448) );
  AOI21_X1 U14612 ( .B1(n13448), .B2(n12137), .A(n12136), .ZN(n12139) );
  NAND2_X1 U14613 ( .A1(n13479), .A2(n13590), .ZN(n12138) );
  OAI211_X1 U14614 ( .C1(n13459), .C2(n12140), .A(n12139), .B(n12138), .ZN(
        n12141) );
  AOI21_X1 U14615 ( .B1(n12142), .B2(n13487), .A(n12141), .ZN(n12143) );
  INV_X1 U14616 ( .A(n12143), .ZN(P2_U3196) );
  NAND2_X1 U14617 ( .A1(n13819), .A2(n15561), .ZN(n13265) );
  XNOR2_X1 U14618 ( .A(n14296), .B(n7172), .ZN(n13267) );
  XOR2_X1 U14619 ( .A(n13265), .B(n13267), .Z(n13262) );
  XNOR2_X1 U14620 ( .A(n13261), .B(n13262), .ZN(n12153) );
  INV_X1 U14621 ( .A(n12146), .ZN(n14195) );
  OAI21_X1 U14622 ( .B1(n13492), .B2(n12148), .A(n12147), .ZN(n12149) );
  AOI21_X1 U14623 ( .B1(n14195), .B2(n13495), .A(n12149), .ZN(n12150) );
  OAI21_X1 U14624 ( .B1(n14160), .B2(n13491), .A(n12150), .ZN(n12151) );
  AOI21_X1 U14625 ( .B1(n14296), .B2(n13479), .A(n12151), .ZN(n12152) );
  OAI21_X1 U14626 ( .B1(n12153), .B2(n13481), .A(n12152), .ZN(P2_U3206) );
  AND2_X1 U14627 ( .A1(n12156), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U14628 ( .A1(n12156), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U14629 ( .A1(n12156), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U14630 ( .A1(n12156), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U14631 ( .A1(n12156), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U14632 ( .A1(n12156), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U14633 ( .A1(n12156), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U14634 ( .A1(n12156), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U14635 ( .A1(n12156), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U14636 ( .A1(n12156), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U14637 ( .A1(n12156), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U14638 ( .A1(n12156), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U14639 ( .A1(n12156), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U14640 ( .A1(n12156), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U14641 ( .A1(n12156), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U14642 ( .A1(n12156), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U14643 ( .A1(n12156), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U14644 ( .A1(n12156), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U14645 ( .A1(n12156), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U14646 ( .A1(n12156), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U14647 ( .A1(n12156), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U14648 ( .A1(n12156), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U14649 ( .A1(n12156), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U14650 ( .A1(n12156), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U14651 ( .A1(n12156), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U14652 ( .A1(n12156), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U14653 ( .A1(n12156), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U14654 ( .A1(n12156), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U14655 ( .A1(n12156), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U14656 ( .A1(n12156), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U14657 ( .A1(n12158), .A2(n12157), .ZN(n12782) );
  INV_X1 U14658 ( .A(n12782), .ZN(n12266) );
  INV_X1 U14659 ( .A(n12159), .ZN(n12896) );
  AND2_X1 U14660 ( .A1(n12898), .A2(n12269), .ZN(n12160) );
  NAND2_X1 U14661 ( .A1(n12238), .A2(n12160), .ZN(n12231) );
  INV_X1 U14662 ( .A(n12222), .ZN(n12227) );
  AOI211_X1 U14663 ( .C1(n12163), .C2(n12164), .A(n12269), .B(n12162), .ZN(
        n12170) );
  INV_X1 U14664 ( .A(n12164), .ZN(n12166) );
  OAI21_X1 U14665 ( .B1(n12168), .B2(n12166), .A(n12165), .ZN(n12167) );
  MUX2_X1 U14666 ( .A(n12168), .B(n12167), .S(n12269), .Z(n12169) );
  AOI21_X1 U14667 ( .B1(n12174), .B2(n12171), .A(n12269), .ZN(n12173) );
  NAND3_X1 U14668 ( .A1(n12182), .A2(n12175), .A3(n12269), .ZN(n12178) );
  NAND2_X1 U14669 ( .A1(n12176), .A2(n12267), .ZN(n12177) );
  AOI21_X1 U14670 ( .B1(n12178), .B2(n12177), .A(n12320), .ZN(n12185) );
  INV_X1 U14671 ( .A(n12182), .ZN(n12179) );
  AOI211_X1 U14672 ( .C1(n12180), .C2(n12187), .A(n12267), .B(n12179), .ZN(
        n12184) );
  AOI21_X1 U14673 ( .B1(n12182), .B2(n12181), .A(n12269), .ZN(n12183) );
  OAI21_X1 U14674 ( .B1(n12269), .B2(n12187), .A(n12324), .ZN(n12192) );
  NAND2_X1 U14675 ( .A1(n12188), .A2(n12269), .ZN(n12190) );
  NAND2_X1 U14676 ( .A1(n15650), .A2(n12267), .ZN(n12189) );
  MUX2_X1 U14677 ( .A(n12190), .B(n12189), .S(n12644), .Z(n12191) );
  OAI211_X1 U14678 ( .C1(n12193), .C2(n12192), .A(n12326), .B(n12191), .ZN(
        n12197) );
  MUX2_X1 U14679 ( .A(n12195), .B(n12194), .S(n12267), .Z(n12196) );
  NAND3_X1 U14680 ( .A1(n12197), .A2(n12332), .A3(n12196), .ZN(n12203) );
  INV_X1 U14681 ( .A(n12198), .ZN(n12199) );
  MUX2_X1 U14682 ( .A(n12200), .B(n12199), .S(n12269), .Z(n12202) );
  AOI21_X1 U14683 ( .B1(n12203), .B2(n12202), .A(n12201), .ZN(n12207) );
  MUX2_X1 U14684 ( .A(n12205), .B(n7870), .S(n12269), .Z(n12206) );
  INV_X1 U14685 ( .A(n12997), .ZN(n12994) );
  NAND2_X1 U14686 ( .A1(n12213), .A2(n12208), .ZN(n12211) );
  NAND2_X1 U14687 ( .A1(n12212), .A2(n12209), .ZN(n12210) );
  MUX2_X1 U14688 ( .A(n12211), .B(n12210), .S(n12269), .Z(n12215) );
  MUX2_X1 U14689 ( .A(n12213), .B(n12212), .S(n12267), .Z(n12214) );
  MUX2_X1 U14690 ( .A(n12217), .B(n12216), .S(n12267), .Z(n12218) );
  MUX2_X1 U14691 ( .A(n12220), .B(n12219), .S(n12269), .Z(n12224) );
  AOI21_X1 U14692 ( .B1(n12222), .B2(n12221), .A(n12269), .ZN(n12223) );
  AOI21_X1 U14693 ( .B1(n12225), .B2(n12224), .A(n12223), .ZN(n12226) );
  AOI211_X1 U14694 ( .C1(n12229), .C2(n12228), .A(n12267), .B(n12227), .ZN(
        n12230) );
  INV_X1 U14695 ( .A(n12231), .ZN(n12236) );
  INV_X1 U14696 ( .A(n12232), .ZN(n12233) );
  NOR2_X1 U14697 ( .A1(n12233), .A2(n12269), .ZN(n12234) );
  AOI22_X1 U14698 ( .A1(n12236), .A2(n12235), .B1(n12234), .B2(n12237), .ZN(
        n12240) );
  MUX2_X1 U14699 ( .A(n12238), .B(n12237), .S(n12269), .Z(n12239) );
  MUX2_X1 U14700 ( .A(n12242), .B(n12241), .S(n12269), .Z(n12246) );
  INV_X1 U14701 ( .A(n12243), .ZN(n12245) );
  MUX2_X1 U14702 ( .A(n12248), .B(n12247), .S(n12267), .Z(n12249) );
  NAND2_X1 U14703 ( .A1(n12250), .A2(n12251), .ZN(n12859) );
  INV_X1 U14704 ( .A(n12847), .ZN(n12842) );
  MUX2_X1 U14705 ( .A(n12251), .B(n12250), .S(n12269), .Z(n12252) );
  NAND2_X1 U14706 ( .A1(n12253), .A2(n12255), .ZN(n12835) );
  NAND2_X1 U14707 ( .A1(n12254), .A2(n12267), .ZN(n12256) );
  MUX2_X1 U14708 ( .A(n12267), .B(n12256), .S(n12255), .Z(n12257) );
  OAI211_X1 U14709 ( .C1(n12258), .C2(n12835), .A(n12821), .B(n12257), .ZN(
        n12262) );
  NAND2_X1 U14710 ( .A1(n12264), .A2(n12536), .ZN(n12265) );
  AND2_X1 U14711 ( .A1(n15165), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12271) );
  XNOR2_X1 U14712 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n12276) );
  XNOR2_X1 U14713 ( .A(n12279), .B(n12276), .ZN(n13237) );
  NAND2_X1 U14714 ( .A1(n13237), .A2(n12294), .ZN(n12274) );
  NAND2_X1 U14715 ( .A1(n12297), .A2(SI_29_), .ZN(n12273) );
  INV_X1 U14716 ( .A(n12636), .ZN(n12539) );
  INV_X1 U14717 ( .A(n12345), .ZN(n12275) );
  INV_X1 U14718 ( .A(n12276), .ZN(n12278) );
  NAND2_X1 U14719 ( .A1(n15163), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12277) );
  XNOR2_X1 U14720 ( .A(n12455), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n12280) );
  XNOR2_X1 U14721 ( .A(n13229), .B(n12280), .ZN(n12459) );
  NAND2_X1 U14722 ( .A1(n12459), .A2(n12294), .ZN(n12282) );
  NAND2_X1 U14723 ( .A1(n12297), .A2(SI_30_), .ZN(n12281) );
  NAND2_X1 U14724 ( .A1(n12282), .A2(n12281), .ZN(n12309) );
  INV_X1 U14725 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n12285) );
  NAND2_X1 U14726 ( .A1(n8851), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n12284) );
  INV_X1 U14727 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n12767) );
  OR2_X1 U14728 ( .A1(n12300), .A2(n12767), .ZN(n12283) );
  OAI211_X1 U14729 ( .C1(n8880), .C2(n12285), .A(n12284), .B(n12283), .ZN(
        n12286) );
  INV_X1 U14730 ( .A(n12286), .ZN(n12287) );
  NAND2_X1 U14731 ( .A1(n12306), .A2(n12287), .ZN(n12773) );
  INV_X1 U14732 ( .A(n12773), .ZN(n12347) );
  OR2_X1 U14733 ( .A1(n12309), .A2(n12347), .ZN(n12351) );
  XNOR2_X1 U14734 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12289) );
  INV_X1 U14735 ( .A(n12289), .ZN(n13230) );
  INV_X1 U14736 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n15159) );
  NAND2_X1 U14737 ( .A1(n15159), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13226) );
  NAND2_X1 U14738 ( .A1(n13230), .A2(n13226), .ZN(n12288) );
  OR2_X1 U14739 ( .A1(n13229), .A2(n12288), .ZN(n12296) );
  NAND2_X1 U14740 ( .A1(n12455), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13227) );
  NAND3_X1 U14741 ( .A1(n13229), .A2(n12289), .A3(n13227), .ZN(n12295) );
  OAI21_X1 U14742 ( .B1(n12289), .B2(n15159), .A(n12455), .ZN(n12292) );
  NAND2_X1 U14743 ( .A1(n12289), .A2(n15159), .ZN(n12290) );
  NAND2_X1 U14744 ( .A1(n12290), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12291) );
  NAND2_X1 U14745 ( .A1(n12292), .A2(n12291), .ZN(n12293) );
  NAND4_X1 U14746 ( .A1(n12296), .A2(n12295), .A3(n12294), .A4(n12293), .ZN(
        n12299) );
  NAND2_X1 U14747 ( .A1(n12297), .A2(SI_31_), .ZN(n12298) );
  INV_X1 U14748 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12303) );
  NAND2_X1 U14749 ( .A1(n8851), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12302) );
  INV_X1 U14750 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12764) );
  OR2_X1 U14751 ( .A1(n12300), .A2(n12764), .ZN(n12301) );
  OAI211_X1 U14752 ( .C1(n8880), .C2(n12303), .A(n12302), .B(n12301), .ZN(
        n12304) );
  INV_X1 U14753 ( .A(n12304), .ZN(n12305) );
  NAND2_X1 U14754 ( .A1(n12757), .A2(n12352), .ZN(n12307) );
  INV_X1 U14755 ( .A(n12757), .ZN(n13132) );
  NOR2_X1 U14756 ( .A1(n12315), .A2(n12343), .ZN(n12312) );
  NAND2_X1 U14757 ( .A1(n12309), .A2(n12347), .ZN(n12341) );
  NAND2_X1 U14758 ( .A1(n13139), .A2(n12539), .ZN(n12349) );
  OAI21_X1 U14759 ( .B1(n12348), .B2(n12357), .A(n12316), .ZN(n12317) );
  INV_X1 U14760 ( .A(n12821), .ZN(n12818) );
  INV_X1 U14761 ( .A(n12873), .ZN(n12338) );
  INV_X1 U14762 ( .A(n12932), .ZN(n12897) );
  NOR2_X1 U14763 ( .A1(n12320), .A2(n12319), .ZN(n12325) );
  NAND4_X1 U14764 ( .A1(n12325), .A2(n12324), .A3(n12323), .A4(n12322), .ZN(
        n12330) );
  INV_X1 U14765 ( .A(n15590), .ZN(n15583) );
  INV_X1 U14766 ( .A(n13018), .ZN(n12328) );
  NOR2_X1 U14767 ( .A1(n12330), .A2(n12329), .ZN(n12333) );
  NOR2_X1 U14768 ( .A1(n12966), .A2(n12334), .ZN(n12335) );
  NAND3_X1 U14769 ( .A1(n12897), .A2(n12336), .A3(n12335), .ZN(n12337) );
  OR4_X1 U14770 ( .A1(n12847), .A2(n12338), .A3(n12859), .A4(n6634), .ZN(
        n12339) );
  NAND2_X1 U14771 ( .A1(n12345), .A2(n12783), .ZN(n12346) );
  OAI21_X1 U14772 ( .B1(n12347), .B2(n12352), .A(n12309), .ZN(n12350) );
  NAND3_X1 U14773 ( .A1(n12350), .A2(n12349), .A3(n12348), .ZN(n12355) );
  INV_X1 U14774 ( .A(n12351), .ZN(n12353) );
  OAI21_X1 U14775 ( .B1(n12353), .B2(n12352), .A(n12757), .ZN(n12354) );
  OAI21_X1 U14776 ( .B1(n12356), .B2(n12355), .A(n12354), .ZN(n12358) );
  XNOR2_X1 U14777 ( .A(n12358), .B(n12357), .ZN(n12360) );
  OAI22_X1 U14778 ( .A1(n12362), .A2(n12361), .B1(n12360), .B2(n12359), .ZN(
        n12364) );
  NAND3_X1 U14779 ( .A1(n12365), .A2(n12758), .A3(n13246), .ZN(n12366) );
  OAI211_X1 U14780 ( .C1(n12368), .C2(n12367), .A(n12366), .B(P3_B_REG_SCAN_IN), .ZN(n12369) );
  INV_X1 U14781 ( .A(n12370), .ZN(n12374) );
  NOR4_X1 U14782 ( .A1(n13481), .A2(n14181), .A3(n12372), .A4(n12371), .ZN(
        n12373) );
  AOI21_X1 U14783 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n12374), .A(n12373), .ZN(
        n12378) );
  OAI21_X1 U14784 ( .B1(n12375), .B2(n13481), .A(n13498), .ZN(n12376) );
  NAND2_X1 U14785 ( .A1(n12376), .A2(n13503), .ZN(n12377) );
  OAI211_X1 U14786 ( .C1(n10882), .C2(n13491), .A(n12378), .B(n12377), .ZN(
        P2_U3204) );
  OAI222_X1 U14787 ( .A1(n13260), .A2(n12380), .B1(n10849), .B2(P3_U3151), 
        .C1(n12379), .C2(n13250), .ZN(P3_U3274) );
  OAI211_X1 U14788 ( .C1(n12383), .C2(n12382), .A(n12381), .B(n14462), .ZN(
        n12387) );
  INV_X1 U14789 ( .A(n14922), .ZN(n14698) );
  AOI22_X1 U14790 ( .A1(n14855), .A2(n14903), .B1(n14698), .B2(n14982), .ZN(
        n15069) );
  OAI22_X1 U14791 ( .A1(n15069), .A2(n14433), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12384), .ZN(n12385) );
  AOI21_X1 U14792 ( .B1(n14886), .B2(n14479), .A(n12385), .ZN(n12386) );
  OAI211_X1 U14793 ( .C1(n15071), .C2(n14468), .A(n12387), .B(n12386), .ZN(
        P1_U3233) );
  INV_X1 U14794 ( .A(n12388), .ZN(n12391) );
  INV_X1 U14795 ( .A(n12389), .ZN(n12390) );
  NAND2_X1 U14796 ( .A1(n12391), .A2(n12390), .ZN(n12398) );
  AND2_X1 U14797 ( .A1(n14390), .A2(n12394), .ZN(n12393) );
  AND2_X1 U14798 ( .A1(n12396), .A2(n12395), .ZN(n12397) );
  INV_X1 U14799 ( .A(n12398), .ZN(n12400) );
  NAND2_X1 U14800 ( .A1(n15033), .A2(n12427), .ZN(n12402) );
  NAND2_X1 U14801 ( .A1(n14800), .A2(n12422), .ZN(n12401) );
  NAND2_X1 U14802 ( .A1(n12402), .A2(n12401), .ZN(n12403) );
  XNOR2_X1 U14803 ( .A(n12403), .B(n12425), .ZN(n12404) );
  AOI22_X1 U14804 ( .A1(n15033), .A2(n12422), .B1(n9434), .B2(n14800), .ZN(
        n12405) );
  INV_X1 U14805 ( .A(n12404), .ZN(n12406) );
  NAND2_X1 U14806 ( .A1(n12406), .A2(n12405), .ZN(n12407) );
  NAND2_X1 U14807 ( .A1(n12408), .A2(n12407), .ZN(n12421) );
  NAND2_X1 U14808 ( .A1(n15027), .A2(n12427), .ZN(n12410) );
  NAND2_X1 U14809 ( .A1(n14741), .A2(n12422), .ZN(n12409) );
  NAND2_X1 U14810 ( .A1(n12410), .A2(n12409), .ZN(n12412) );
  XNOR2_X1 U14811 ( .A(n12412), .B(n12411), .ZN(n12431) );
  AND2_X1 U14812 ( .A1(n14741), .A2(n9434), .ZN(n12413) );
  AOI21_X1 U14813 ( .B1(n15027), .B2(n12422), .A(n12413), .ZN(n12430) );
  XNOR2_X1 U14814 ( .A(n12431), .B(n12430), .ZN(n12419) );
  XNOR2_X1 U14815 ( .A(n12421), .B(n12419), .ZN(n12418) );
  INV_X1 U14816 ( .A(n14758), .ZN(n14686) );
  NOR2_X1 U14817 ( .A1(n14686), .A2(n14482), .ZN(n12416) );
  AOI22_X1 U14818 ( .A1(n14800), .A2(n14478), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12414) );
  OAI21_X1 U14819 ( .B1(n14766), .B2(n14494), .A(n12414), .ZN(n12415) );
  AOI211_X1 U14820 ( .C1(n15027), .C2(n14496), .A(n12416), .B(n12415), .ZN(
        n12417) );
  OAI21_X1 U14821 ( .B1(n12418), .B2(n14498), .A(n12417), .ZN(P1_U3214) );
  INV_X1 U14822 ( .A(n12419), .ZN(n12420) );
  NAND2_X1 U14823 ( .A1(n12421), .A2(n12420), .ZN(n12445) );
  NAND2_X1 U14824 ( .A1(n14748), .A2(n12422), .ZN(n12424) );
  NAND2_X1 U14825 ( .A1(n14758), .A2(n9434), .ZN(n12423) );
  NAND2_X1 U14826 ( .A1(n12424), .A2(n12423), .ZN(n12426) );
  XNOR2_X1 U14827 ( .A(n12426), .B(n12425), .ZN(n12429) );
  AOI22_X1 U14828 ( .A1(n14748), .A2(n12427), .B1(n12422), .B2(n14758), .ZN(
        n12428) );
  XNOR2_X1 U14829 ( .A(n12429), .B(n12428), .ZN(n12436) );
  NAND2_X1 U14830 ( .A1(n12436), .A2(n14462), .ZN(n12444) );
  AND2_X1 U14831 ( .A1(n12431), .A2(n12430), .ZN(n12437) );
  NOR3_X1 U14832 ( .A1(n12436), .A2(n12437), .A3(n14498), .ZN(n12432) );
  NAND2_X1 U14833 ( .A1(n12445), .A2(n12432), .ZN(n12443) );
  INV_X1 U14834 ( .A(n12433), .ZN(n14744) );
  AOI22_X1 U14835 ( .A1(n14740), .A2(n14473), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12435) );
  NAND2_X1 U14836 ( .A1(n14741), .A2(n14478), .ZN(n12434) );
  OAI211_X1 U14837 ( .C1(n14744), .C2(n14494), .A(n12435), .B(n12434), .ZN(
        n12441) );
  INV_X1 U14838 ( .A(n12436), .ZN(n12439) );
  INV_X1 U14839 ( .A(n12437), .ZN(n12438) );
  NOR3_X1 U14840 ( .A1(n12439), .A2(n14498), .A3(n12438), .ZN(n12440) );
  AOI211_X1 U14841 ( .C1(n14496), .C2(n14748), .A(n12441), .B(n12440), .ZN(
        n12442) );
  OAI211_X1 U14842 ( .C1(n12445), .C2(n12444), .A(n12443), .B(n12442), .ZN(
        P1_U3220) );
  OAI222_X1 U14843 ( .A1(n14374), .A2(n12447), .B1(n14372), .B2(n12446), .C1(
        P2_U3088), .C2(n8558), .ZN(P2_U3307) );
  INV_X1 U14844 ( .A(n12448), .ZN(n14365) );
  OAI222_X1 U14845 ( .A1(n14651), .A2(P1_U3086), .B1(n15169), .B2(n14365), 
        .C1(n12449), .C2(n15164), .ZN(P1_U3328) );
  AOI22_X1 U14846 ( .A1(n12540), .A2(n13011), .B1(n15601), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12450) );
  OAI21_X1 U14847 ( .B1(n12618), .B2(n12989), .A(n12450), .ZN(n12451) );
  OAI21_X1 U14848 ( .B1(n12453), .B2(n13007), .A(n12452), .ZN(P3_U3205) );
  INV_X1 U14849 ( .A(n12454), .ZN(n15160) );
  OAI222_X1 U14850 ( .A1(n12456), .A2(P2_U3088), .B1(n14372), .B2(n12455), 
        .C1(n14367), .C2(n15160), .ZN(P2_U3297) );
  INV_X1 U14851 ( .A(n12457), .ZN(n15166) );
  OAI222_X1 U14852 ( .A1(P2_U3088), .A2(n8615), .B1(n14374), .B2(n15166), .C1(
        n12458), .C2(n14372), .ZN(P2_U3299) );
  INV_X1 U14853 ( .A(n12459), .ZN(n12462) );
  OAI222_X1 U14854 ( .A1(n13248), .A2(n12462), .B1(n12461), .B2(P3_U3151), 
        .C1(n12460), .C2(n13256), .ZN(P3_U3265) );
  XNOR2_X1 U14855 ( .A(n12801), .B(n12463), .ZN(n12533) );
  XNOR2_X1 U14856 ( .A(n12533), .B(n13036), .ZN(n12534) );
  XNOR2_X1 U14857 ( .A(n13200), .B(n12463), .ZN(n12467) );
  XNOR2_X1 U14858 ( .A(n12467), .B(n12976), .ZN(n12509) );
  INV_X1 U14859 ( .A(n12467), .ZN(n12468) );
  NAND2_X1 U14860 ( .A1(n12468), .A2(n12976), .ZN(n12469) );
  INV_X1 U14861 ( .A(n12624), .ZN(n12471) );
  XNOR2_X1 U14862 ( .A(n13100), .B(n12463), .ZN(n12472) );
  XNOR2_X1 U14863 ( .A(n12472), .B(n12943), .ZN(n12625) );
  NAND2_X1 U14864 ( .A1(n12472), .A2(n12943), .ZN(n12473) );
  XNOR2_X1 U14865 ( .A(n13094), .B(n12463), .ZN(n12474) );
  XNOR2_X1 U14866 ( .A(n12474), .B(n13097), .ZN(n12562) );
  INV_X1 U14867 ( .A(n12474), .ZN(n12475) );
  XNOR2_X1 U14868 ( .A(n13088), .B(n12463), .ZN(n12476) );
  XNOR2_X1 U14869 ( .A(n12476), .B(n12640), .ZN(n12572) );
  INV_X1 U14870 ( .A(n12476), .ZN(n12477) );
  NAND2_X1 U14871 ( .A1(n12477), .A2(n12640), .ZN(n12478) );
  NAND2_X1 U14872 ( .A1(n12571), .A2(n12478), .ZN(n12607) );
  XNOR2_X1 U14873 ( .A(n12924), .B(n12463), .ZN(n12480) );
  XNOR2_X1 U14874 ( .A(n12480), .B(n13085), .ZN(n12608) );
  INV_X1 U14875 ( .A(n12608), .ZN(n12479) );
  NAND2_X1 U14876 ( .A1(n12480), .A2(n13085), .ZN(n12481) );
  XNOR2_X1 U14877 ( .A(n12910), .B(n12463), .ZN(n12482) );
  XNOR2_X1 U14878 ( .A(n12482), .B(n13070), .ZN(n12524) );
  INV_X1 U14879 ( .A(n12482), .ZN(n12483) );
  XNOR2_X1 U14880 ( .A(n13073), .B(n12463), .ZN(n12484) );
  XNOR2_X1 U14881 ( .A(n12484), .B(n12908), .ZN(n12591) );
  INV_X1 U14882 ( .A(n12484), .ZN(n12485) );
  XNOR2_X1 U14883 ( .A(n13168), .B(n12463), .ZN(n12487) );
  XNOR2_X1 U14884 ( .A(n12487), .B(n12889), .ZN(n12549) );
  INV_X1 U14885 ( .A(n12549), .ZN(n12486) );
  NAND2_X1 U14886 ( .A1(n12487), .A2(n12889), .ZN(n12488) );
  XNOR2_X1 U14887 ( .A(n12489), .B(n12463), .ZN(n12490) );
  INV_X1 U14888 ( .A(n12490), .ZN(n12491) );
  AND2_X1 U14889 ( .A1(n12492), .A2(n12491), .ZN(n12493) );
  AOI21_X2 U14890 ( .B1(n12599), .B2(n12848), .A(n12493), .ZN(n12517) );
  XNOR2_X1 U14891 ( .A(n13056), .B(n12463), .ZN(n12581) );
  XNOR2_X1 U14892 ( .A(n13061), .B(n12494), .ZN(n12579) );
  INV_X1 U14893 ( .A(n12579), .ZN(n12495) );
  OAI22_X1 U14894 ( .A1(n12581), .A2(n13058), .B1(n13050), .B2(n12495), .ZN(
        n12499) );
  OAI21_X1 U14895 ( .B1(n12579), .B2(n12861), .A(n12637), .ZN(n12497) );
  NOR2_X1 U14896 ( .A1(n12637), .A2(n12861), .ZN(n12496) );
  AOI22_X1 U14897 ( .A1(n12581), .A2(n12497), .B1(n12496), .B2(n12495), .ZN(
        n12498) );
  XNOR2_X1 U14898 ( .A(n13046), .B(n12463), .ZN(n12500) );
  XNOR2_X1 U14899 ( .A(n12500), .B(n13035), .ZN(n12556) );
  XNOR2_X1 U14900 ( .A(n13034), .B(n12463), .ZN(n12501) );
  XNOR2_X1 U14901 ( .A(n12501), .B(n13043), .ZN(n12615) );
  INV_X1 U14902 ( .A(n12501), .ZN(n12502) );
  XOR2_X1 U14903 ( .A(n12534), .B(n12535), .Z(n12507) );
  NOR2_X1 U14904 ( .A1(n12796), .A2(n12628), .ZN(n12505) );
  AOI22_X1 U14905 ( .A1(n12802), .A2(n12630), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12503) );
  OAI21_X1 U14906 ( .B1(n13043), .B2(n12593), .A(n12503), .ZN(n12504) );
  AOI211_X1 U14907 ( .C1(n12801), .C2(n12631), .A(n12505), .B(n12504), .ZN(
        n12506) );
  OAI21_X1 U14908 ( .B1(n12507), .B2(n12634), .A(n12506), .ZN(P3_U3154) );
  INV_X1 U14909 ( .A(n13200), .ZN(n12516) );
  OAI211_X1 U14910 ( .C1(n12510), .C2(n12509), .A(n12508), .B(n12589), .ZN(
        n12515) );
  AND2_X1 U14911 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12678) );
  AOI21_X1 U14912 ( .B1(n12511), .B2(n12968), .A(n12678), .ZN(n12512) );
  OAI21_X1 U14913 ( .B1(n12985), .B2(n12593), .A(n12512), .ZN(n12513) );
  AOI21_X1 U14914 ( .B1(n12971), .B2(n12630), .A(n12513), .ZN(n12514) );
  OAI211_X1 U14915 ( .C1(n12516), .C2(n12610), .A(n12515), .B(n12514), .ZN(
        P3_U3155) );
  XNOR2_X1 U14916 ( .A(n12517), .B(n12579), .ZN(n12580) );
  XNOR2_X1 U14917 ( .A(n12580), .B(n13050), .ZN(n12523) );
  INV_X1 U14918 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n12518) );
  OAI22_X1 U14919 ( .A1(n12848), .A2(n12593), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12518), .ZN(n12520) );
  NOR2_X1 U14920 ( .A1(n13058), .A2(n12628), .ZN(n12519) );
  AOI211_X1 U14921 ( .C1(n12843), .C2(n12630), .A(n12520), .B(n12519), .ZN(
        n12522) );
  NAND2_X1 U14922 ( .A1(n13061), .A2(n12631), .ZN(n12521) );
  OAI211_X1 U14923 ( .C1(n12523), .C2(n12634), .A(n12522), .B(n12521), .ZN(
        P3_U3156) );
  XOR2_X1 U14924 ( .A(n12525), .B(n12524), .Z(n12532) );
  NAND2_X1 U14925 ( .A1(n12639), .A2(n12626), .ZN(n12527) );
  OAI211_X1 U14926 ( .C1(n12528), .C2(n12628), .A(n12527), .B(n12526), .ZN(
        n12530) );
  NOR2_X1 U14927 ( .A1(n12910), .A2(n12610), .ZN(n12529) );
  AOI211_X1 U14928 ( .C1(n12911), .C2(n12630), .A(n12530), .B(n12529), .ZN(
        n12531) );
  OAI21_X1 U14929 ( .B1(n12532), .B2(n12634), .A(n12531), .ZN(P3_U3159) );
  XNOR2_X1 U14930 ( .A(n12536), .B(n12463), .ZN(n12537) );
  XNOR2_X1 U14931 ( .A(n12538), .B(n12537), .ZN(n12545) );
  NOR2_X1 U14932 ( .A1(n12539), .A2(n12628), .ZN(n12543) );
  AOI22_X1 U14933 ( .A1(n12540), .A2(n12630), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12541) );
  OAI21_X1 U14934 ( .B1(n12618), .B2(n12593), .A(n12541), .ZN(n12542) );
  AOI211_X1 U14935 ( .C1(n12772), .C2(n12631), .A(n12543), .B(n12542), .ZN(
        n12544) );
  OAI21_X1 U14936 ( .B1(n12545), .B2(n12634), .A(n12544), .ZN(P3_U3160) );
  INV_X1 U14937 ( .A(n12546), .ZN(n12547) );
  AOI21_X1 U14938 ( .B1(n12549), .B2(n12548), .A(n12547), .ZN(n12554) );
  AOI22_X1 U14939 ( .A1(n12908), .A2(n12626), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12551) );
  NAND2_X1 U14940 ( .A1(n12878), .A2(n12630), .ZN(n12550) );
  OAI211_X1 U14941 ( .C1(n12848), .C2(n12628), .A(n12551), .B(n12550), .ZN(
        n12552) );
  AOI21_X1 U14942 ( .B1(n13168), .B2(n12631), .A(n12552), .ZN(n12553) );
  OAI21_X1 U14943 ( .B1(n12554), .B2(n12634), .A(n12553), .ZN(P3_U3163) );
  XOR2_X1 U14944 ( .A(n12556), .B(n12555), .Z(n12561) );
  AOI22_X1 U14945 ( .A1(n12637), .A2(n12626), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12558) );
  NAND2_X1 U14946 ( .A1(n12823), .A2(n12630), .ZN(n12557) );
  OAI211_X1 U14947 ( .C1(n13043), .C2(n12628), .A(n12558), .B(n12557), .ZN(
        n12559) );
  AOI21_X1 U14948 ( .B1(n13046), .B2(n12631), .A(n12559), .ZN(n12560) );
  OAI21_X1 U14949 ( .B1(n12561), .B2(n12634), .A(n12560), .ZN(P3_U3165) );
  INV_X1 U14950 ( .A(n13094), .ZN(n12570) );
  AOI21_X1 U14951 ( .B1(n12563), .B2(n12562), .A(n12634), .ZN(n12565) );
  NAND2_X1 U14952 ( .A1(n12565), .A2(n12564), .ZN(n12569) );
  NAND2_X1 U14953 ( .A1(n12626), .A2(n12968), .ZN(n12566) );
  NAND2_X1 U14954 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12714)
         );
  OAI211_X1 U14955 ( .C1(n13091), .C2(n12628), .A(n12566), .B(n12714), .ZN(
        n12567) );
  AOI21_X1 U14956 ( .B1(n12945), .B2(n12630), .A(n12567), .ZN(n12568) );
  OAI211_X1 U14957 ( .C1(n12570), .C2(n12610), .A(n12569), .B(n12568), .ZN(
        P3_U3166) );
  INV_X1 U14958 ( .A(n13088), .ZN(n12578) );
  OAI211_X1 U14959 ( .C1(n12573), .C2(n12572), .A(n12571), .B(n12589), .ZN(
        n12577) );
  NAND2_X1 U14960 ( .A1(n12626), .A2(n12641), .ZN(n12574) );
  NAND2_X1 U14961 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12730)
         );
  OAI211_X1 U14962 ( .C1(n13085), .C2(n12628), .A(n12574), .B(n12730), .ZN(
        n12575) );
  AOI21_X1 U14963 ( .B1(n12935), .B2(n12630), .A(n12575), .ZN(n12576) );
  OAI211_X1 U14964 ( .C1(n12578), .C2(n12610), .A(n12577), .B(n12576), .ZN(
        P3_U3168) );
  OAI22_X1 U14965 ( .A1(n12580), .A2(n12861), .B1(n12517), .B2(n12579), .ZN(
        n12583) );
  XNOR2_X1 U14966 ( .A(n12581), .B(n13058), .ZN(n12582) );
  XNOR2_X1 U14967 ( .A(n12583), .B(n12582), .ZN(n12588) );
  AOI22_X1 U14968 ( .A1(n12861), .A2(n12626), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12585) );
  NAND2_X1 U14969 ( .A1(n12832), .A2(n12630), .ZN(n12584) );
  OAI211_X1 U14970 ( .C1(n13051), .C2(n12628), .A(n12585), .B(n12584), .ZN(
        n12586) );
  AOI21_X1 U14971 ( .B1(n13056), .B2(n12631), .A(n12586), .ZN(n12587) );
  OAI21_X1 U14972 ( .B1(n12588), .B2(n12634), .A(n12587), .ZN(P3_U3169) );
  INV_X1 U14973 ( .A(n13073), .ZN(n12598) );
  OAI211_X1 U14974 ( .C1(n12592), .C2(n12591), .A(n12590), .B(n12589), .ZN(
        n12597) );
  NOR2_X1 U14975 ( .A1(n13070), .A2(n12593), .ZN(n12595) );
  OAI22_X1 U14976 ( .A1(n12889), .A2(n12628), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15793), .ZN(n12594) );
  AOI211_X1 U14977 ( .C1(n12891), .C2(n12630), .A(n12595), .B(n12594), .ZN(
        n12596) );
  OAI211_X1 U14978 ( .C1(n12598), .C2(n12610), .A(n12597), .B(n12596), .ZN(
        P3_U3173) );
  XNOR2_X1 U14979 ( .A(n12599), .B(n12875), .ZN(n12604) );
  AOI22_X1 U14980 ( .A1(n12860), .A2(n12626), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12601) );
  NAND2_X1 U14981 ( .A1(n12864), .A2(n12630), .ZN(n12600) );
  OAI211_X1 U14982 ( .C1(n13050), .C2(n12628), .A(n12601), .B(n12600), .ZN(
        n12602) );
  AOI21_X1 U14983 ( .B1(n13162), .B2(n12631), .A(n12602), .ZN(n12603) );
  OAI21_X1 U14984 ( .B1(n12604), .B2(n12634), .A(n12603), .ZN(P3_U3175) );
  INV_X1 U14985 ( .A(n12605), .ZN(n12606) );
  AOI21_X1 U14986 ( .B1(n12608), .B2(n12607), .A(n12606), .ZN(n12614) );
  NAND2_X1 U14987 ( .A1(n12626), .A2(n12640), .ZN(n12609) );
  NAND2_X1 U14988 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12749)
         );
  OAI211_X1 U14989 ( .C1(n13070), .C2(n12628), .A(n12609), .B(n12749), .ZN(
        n12612) );
  INV_X1 U14990 ( .A(n12924), .ZN(n13185) );
  NOR2_X1 U14991 ( .A1(n13185), .A2(n12610), .ZN(n12611) );
  AOI211_X1 U14992 ( .C1(n12917), .C2(n12630), .A(n12612), .B(n12611), .ZN(
        n12613) );
  OAI21_X1 U14993 ( .B1(n12614), .B2(n12634), .A(n12613), .ZN(P3_U3178) );
  AOI22_X1 U14994 ( .A1(n12810), .A2(n12630), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12617) );
  NAND2_X1 U14995 ( .A1(n13035), .A2(n12626), .ZN(n12616) );
  OAI211_X1 U14996 ( .C1(n12618), .C2(n12628), .A(n12617), .B(n12616), .ZN(
        n12619) );
  AOI21_X1 U14997 ( .B1(n13034), .B2(n12631), .A(n12619), .ZN(n12620) );
  OAI21_X1 U14998 ( .B1(n12621), .B2(n12634), .A(n12620), .ZN(P3_U3180) );
  INV_X1 U14999 ( .A(n12622), .ZN(n12623) );
  AOI21_X1 U15000 ( .B1(n12625), .B2(n12624), .A(n12623), .ZN(n12635) );
  NAND2_X1 U15001 ( .A1(n12626), .A2(n12976), .ZN(n12627) );
  NAND2_X1 U15002 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12693)
         );
  OAI211_X1 U15003 ( .C1(n13097), .C2(n12628), .A(n12627), .B(n12693), .ZN(
        n12629) );
  AOI21_X1 U15004 ( .B1(n12955), .B2(n12630), .A(n12629), .ZN(n12633) );
  NAND2_X1 U15005 ( .A1(n13100), .A2(n12631), .ZN(n12632) );
  OAI211_X1 U15006 ( .C1(n12635), .C2(n12634), .A(n12633), .B(n12632), .ZN(
        P3_U3181) );
  MUX2_X1 U15007 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12760), .S(n12647), .Z(
        P3_U3522) );
  MUX2_X1 U15008 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n12773), .S(P3_U3897), .Z(
        P3_U3521) );
  MUX2_X1 U15009 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n12636), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U15010 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12775), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U15011 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n13036), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U15012 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12822), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U15013 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n13035), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U15014 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12637), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U15015 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12875), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15016 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12908), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15017 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12638), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U15018 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12639), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15019 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12640), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U15020 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12641), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U15021 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12968), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U15022 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12976), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U15023 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12967), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U15024 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12999), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U15025 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12642), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U15026 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12998), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15027 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12643), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U15028 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n15655), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U15029 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12644), .S(n12647), .Z(
        P3_U3498) );
  MUX2_X1 U15030 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n15630), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U15031 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12645), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U15032 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n15620), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15033 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n13012), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15034 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12646), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15035 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n15605), .S(n12647), .Z(
        P3_U3491) );
  AOI21_X1 U15036 ( .B1(n12978), .B2(n12648), .A(n12664), .ZN(n12662) );
  OAI21_X1 U15037 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n12650), .A(n12649), 
        .ZN(n12660) );
  INV_X1 U15038 ( .A(n12673), .ZN(n12655) );
  AOI21_X1 U15039 ( .B1(n12653), .B2(n12652), .A(n12651), .ZN(n12654) );
  OAI21_X1 U15040 ( .B1(n12655), .B2(n12654), .A(n12675), .ZN(n12658) );
  AOI21_X1 U15041 ( .B1(n15581), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12656), 
        .ZN(n12657) );
  OAI211_X1 U15042 ( .C1(n12682), .C2(n6841), .A(n12658), .B(n12657), .ZN(
        n12659) );
  AOI21_X1 U15043 ( .B1(n12692), .B2(n12660), .A(n12659), .ZN(n12661) );
  OAI21_X1 U15044 ( .B1(n12662), .B2(n12702), .A(n12661), .ZN(P3_U3195) );
  INV_X1 U15045 ( .A(n12663), .ZN(n12668) );
  NOR3_X1 U15046 ( .A1(n12666), .A2(n12665), .A3(n12664), .ZN(n12667) );
  OAI21_X1 U15047 ( .B1(n12668), .B2(n12667), .A(n12744), .ZN(n12686) );
  OAI21_X1 U15048 ( .B1(n12671), .B2(n12670), .A(n12669), .ZN(n12684) );
  AND2_X1 U15049 ( .A1(n12673), .A2(n12672), .ZN(n12677) );
  OAI211_X1 U15050 ( .C1(n12677), .C2(n12676), .A(n12675), .B(n12674), .ZN(
        n12680) );
  AOI21_X1 U15051 ( .B1(n15581), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12678), 
        .ZN(n12679) );
  OAI211_X1 U15052 ( .C1(n12682), .C2(n12681), .A(n12680), .B(n12679), .ZN(
        n12683) );
  AOI21_X1 U15053 ( .B1(n12692), .B2(n12684), .A(n12683), .ZN(n12685) );
  NAND2_X1 U15054 ( .A1(n12686), .A2(n12685), .ZN(P3_U3196) );
  AOI21_X1 U15055 ( .B1(n12688), .B2(n12687), .A(n12711), .ZN(n12703) );
  INV_X1 U15056 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n15213) );
  OAI21_X1 U15057 ( .B1(n12690), .B2(P3_REG1_REG_15__SCAN_IN), .A(n12689), 
        .ZN(n12691) );
  NAND2_X1 U15058 ( .A1(n12692), .A2(n12691), .ZN(n12694) );
  OAI211_X1 U15059 ( .C1(n12715), .C2(n15213), .A(n12694), .B(n12693), .ZN(
        n12700) );
  AOI21_X1 U15060 ( .B1(n12697), .B2(n12696), .A(n12695), .ZN(n12698) );
  NOR2_X1 U15061 ( .A1(n12698), .A2(n12755), .ZN(n12699) );
  AOI211_X1 U15062 ( .C1(n12751), .C2(n10157), .A(n12700), .B(n12699), .ZN(
        n12701) );
  OAI21_X1 U15063 ( .B1(n12703), .B2(n12702), .A(n12701), .ZN(P3_U3197) );
  OAI21_X1 U15064 ( .B1(n12706), .B2(n12705), .A(n12704), .ZN(n12707) );
  INV_X1 U15065 ( .A(n12707), .ZN(n12725) );
  INV_X1 U15066 ( .A(n12708), .ZN(n12713) );
  NOR3_X1 U15067 ( .A1(n12711), .A2(n12710), .A3(n12709), .ZN(n12712) );
  OAI21_X1 U15068 ( .B1(n12713), .B2(n12712), .A(n12744), .ZN(n12724) );
  INV_X1 U15069 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n15226) );
  OAI21_X1 U15070 ( .B1(n12715), .B2(n15226), .A(n12714), .ZN(n12721) );
  NOR2_X1 U15071 ( .A1(n12716), .A2(n6660), .ZN(n12717) );
  XNOR2_X1 U15072 ( .A(n12718), .B(n12717), .ZN(n12719) );
  NOR2_X1 U15073 ( .A1(n12719), .A2(n12755), .ZN(n12720) );
  AOI211_X1 U15074 ( .C1(n12751), .C2(n12722), .A(n12721), .B(n12720), .ZN(
        n12723) );
  OAI211_X1 U15075 ( .C1(n12725), .C2(n12750), .A(n12724), .B(n12723), .ZN(
        P3_U3198) );
  OAI21_X1 U15076 ( .B1(P3_REG2_REG_17__SCAN_IN), .B2(n12726), .A(n12743), 
        .ZN(n12727) );
  NAND2_X1 U15077 ( .A1(n12727), .A2(n12744), .ZN(n12738) );
  XNOR2_X1 U15078 ( .A(n12728), .B(P3_REG1_REG_17__SCAN_IN), .ZN(n12731) );
  NAND2_X1 U15079 ( .A1(n15581), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n12729) );
  OAI211_X1 U15080 ( .C1(n12750), .C2(n12731), .A(n12730), .B(n12729), .ZN(
        n12735) );
  AOI211_X1 U15081 ( .C1(n12733), .C2(n12732), .A(n12755), .B(n6546), .ZN(
        n12734) );
  AOI211_X1 U15082 ( .C1(n12751), .C2(n12736), .A(n12735), .B(n12734), .ZN(
        n12737) );
  NAND2_X1 U15083 ( .A1(n12738), .A2(n12737), .ZN(P3_U3199) );
  AOI21_X1 U15084 ( .B1(n12741), .B2(n12740), .A(n12739), .ZN(n12756) );
  AND3_X1 U15085 ( .A1(n12743), .A2(n7265), .A3(n12742), .ZN(n12745) );
  OAI21_X1 U15086 ( .B1(n12746), .B2(n12745), .A(n12744), .ZN(n12754) );
  OAI211_X1 U15087 ( .C1(n12756), .C2(n12755), .A(n12754), .B(n12753), .ZN(
        P3_U3200) );
  NAND2_X1 U15088 ( .A1(n12757), .A2(n13004), .ZN(n12763) );
  NAND2_X1 U15089 ( .A1(n12758), .A2(P3_B_REG_SCAN_IN), .ZN(n12759) );
  AND2_X1 U15090 ( .A1(n15656), .A2(n12759), .ZN(n12774) );
  NAND2_X1 U15091 ( .A1(n12760), .A2(n12774), .ZN(n13130) );
  INV_X1 U15092 ( .A(n13130), .ZN(n12762) );
  NOR2_X1 U15093 ( .A1(n12761), .A2(n15588), .ZN(n12781) );
  OAI21_X1 U15094 ( .B1(n12762), .B2(n12781), .A(n15599), .ZN(n12765) );
  OAI211_X1 U15095 ( .C1(n15599), .C2(n12764), .A(n12763), .B(n12765), .ZN(
        P3_U3202) );
  NAND2_X1 U15096 ( .A1(n12309), .A2(n13004), .ZN(n12766) );
  OAI211_X1 U15097 ( .C1(n15599), .C2(n12767), .A(n12766), .B(n12765), .ZN(
        P3_U3203) );
  AOI21_X1 U15098 ( .B1(n12772), .B2(n12775), .A(n13052), .ZN(n12769) );
  NAND2_X1 U15099 ( .A1(n12785), .A2(n12769), .ZN(n12770) );
  NAND3_X1 U15100 ( .A1(n12768), .A2(n12771), .A3(n15611), .ZN(n12779) );
  NAND3_X1 U15101 ( .A1(n12772), .A2(n12775), .A3(n15611), .ZN(n12777) );
  AOI22_X1 U15102 ( .A1(n12775), .A2(n15638), .B1(n12774), .B2(n12773), .ZN(
        n12776) );
  OAI21_X1 U15103 ( .B1(n12785), .B2(n12777), .A(n12776), .ZN(n12778) );
  INV_X1 U15104 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n12780) );
  AOI21_X1 U15105 ( .B1(n13139), .B2(n12991), .A(n12781), .ZN(n12788) );
  NAND2_X1 U15106 ( .A1(n12792), .A2(n12782), .ZN(n12784) );
  NAND2_X1 U15107 ( .A1(n12784), .A2(n12783), .ZN(n12786) );
  NAND2_X1 U15108 ( .A1(n13140), .A2(n13010), .ZN(n12787) );
  NAND3_X1 U15109 ( .A1(n12789), .A2(n12788), .A3(n12787), .ZN(P3_U3204) );
  INV_X1 U15110 ( .A(n12790), .ZN(n12793) );
  OAI21_X1 U15111 ( .B1(n12795), .B2(n9269), .A(n12794), .ZN(n12798) );
  OAI22_X1 U15112 ( .A1(n12796), .A2(n15642), .B1(n13043), .B2(n15652), .ZN(
        n12797) );
  AOI21_X1 U15113 ( .B1(n12798), .B2(n15611), .A(n12797), .ZN(n12799) );
  INV_X1 U15114 ( .A(n13030), .ZN(n12808) );
  INV_X1 U15115 ( .A(n12800), .ZN(n13031) );
  INV_X1 U15116 ( .A(n12801), .ZN(n13145) );
  AOI22_X1 U15117 ( .A1(n12802), .A2(n13011), .B1(n15601), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12803) );
  OAI21_X1 U15118 ( .B1(n13145), .B2(n12804), .A(n12803), .ZN(n12805) );
  AOI21_X1 U15119 ( .B1(n13031), .B2(n12806), .A(n12805), .ZN(n12807) );
  OAI21_X1 U15120 ( .B1(n12808), .B2(n15601), .A(n12807), .ZN(P3_U3206) );
  XNOR2_X1 U15121 ( .A(n6596), .B(n12809), .ZN(n13038) );
  NAND2_X1 U15122 ( .A1(n13036), .A2(n13013), .ZN(n12812) );
  AOI22_X1 U15123 ( .A1(n12810), .A2(n13011), .B1(n15601), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12811) );
  OAI211_X1 U15124 ( .C1(n13051), .C2(n12989), .A(n12812), .B(n12811), .ZN(
        n12813) );
  AOI21_X1 U15125 ( .B1(n13034), .B2(n12991), .A(n12813), .ZN(n12817) );
  XNOR2_X1 U15126 ( .A(n12814), .B(n12815), .ZN(n13040) );
  NOR2_X1 U15127 ( .A1(n15601), .A2(n13052), .ZN(n13019) );
  NAND2_X1 U15128 ( .A1(n13040), .A2(n13019), .ZN(n12816) );
  OAI211_X1 U15129 ( .C1(n13038), .C2(n13007), .A(n12817), .B(n12816), .ZN(
        P3_U3207) );
  XNOR2_X1 U15130 ( .A(n12819), .B(n12818), .ZN(n13048) );
  AOI211_X1 U15131 ( .C1(n12821), .C2(n12820), .A(n13052), .B(n6530), .ZN(
        n13044) );
  NAND2_X1 U15132 ( .A1(n13044), .A2(n15599), .ZN(n12828) );
  NAND2_X1 U15133 ( .A1(n12822), .A2(n13013), .ZN(n12825) );
  AOI22_X1 U15134 ( .A1(n12823), .A2(n13011), .B1(n15601), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12824) );
  OAI211_X1 U15135 ( .C1(n13058), .C2(n12989), .A(n12825), .B(n12824), .ZN(
        n12826) );
  AOI21_X1 U15136 ( .B1(n13046), .B2(n13004), .A(n12826), .ZN(n12827) );
  OAI211_X1 U15137 ( .C1(n13007), .C2(n13048), .A(n12828), .B(n12827), .ZN(
        P3_U3208) );
  NAND2_X1 U15138 ( .A1(n12829), .A2(n12842), .ZN(n12841) );
  NAND2_X1 U15139 ( .A1(n12841), .A2(n12830), .ZN(n12831) );
  XOR2_X1 U15140 ( .A(n12835), .B(n12831), .Z(n13155) );
  NAND2_X1 U15141 ( .A1(n13035), .A2(n13013), .ZN(n12834) );
  AOI22_X1 U15142 ( .A1(n12832), .A2(n13011), .B1(n15601), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n12833) );
  OAI211_X1 U15143 ( .C1(n13050), .C2(n12989), .A(n12834), .B(n12833), .ZN(
        n12839) );
  XNOR2_X1 U15144 ( .A(n12836), .B(n12835), .ZN(n13053) );
  INV_X1 U15145 ( .A(n13019), .ZN(n12837) );
  NOR2_X1 U15146 ( .A1(n13053), .A2(n12837), .ZN(n12838) );
  AOI211_X1 U15147 ( .C1(n12991), .C2(n13056), .A(n12839), .B(n12838), .ZN(
        n12840) );
  OAI21_X1 U15148 ( .B1(n13155), .B2(n13007), .A(n12840), .ZN(P3_U3209) );
  OAI21_X1 U15149 ( .B1(n12829), .B2(n12842), .A(n12841), .ZN(n13159) );
  INV_X1 U15150 ( .A(n13013), .ZN(n12957) );
  AOI22_X1 U15151 ( .A1(n12843), .A2(n13011), .B1(n15601), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n12844) );
  OAI21_X1 U15152 ( .B1(n13058), .B2(n12957), .A(n12844), .ZN(n12845) );
  AOI21_X1 U15153 ( .B1(n13061), .B2(n12991), .A(n12845), .ZN(n12851) );
  XNOR2_X1 U15154 ( .A(n12846), .B(n12847), .ZN(n12849) );
  OAI22_X1 U15155 ( .A1(n12849), .A2(n13052), .B1(n12848), .B2(n15652), .ZN(
        n13059) );
  NAND2_X1 U15156 ( .A1(n13059), .A2(n15599), .ZN(n12850) );
  OAI211_X1 U15157 ( .C1(n13159), .C2(n13007), .A(n12851), .B(n12850), .ZN(
        P3_U3210) );
  XOR2_X1 U15158 ( .A(n12852), .B(n12859), .Z(n13165) );
  INV_X1 U15159 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12863) );
  NOR2_X1 U15160 ( .A1(n12915), .A2(n12854), .ZN(n12857) );
  OAI21_X1 U15161 ( .B1(n12857), .B2(n12856), .A(n12855), .ZN(n12858) );
  XOR2_X1 U15162 ( .A(n12859), .B(n12858), .Z(n12862) );
  AOI222_X1 U15163 ( .A1(n15611), .A2(n12862), .B1(n12861), .B2(n15656), .C1(
        n12860), .C2(n15638), .ZN(n13160) );
  MUX2_X1 U15164 ( .A(n12863), .B(n13160), .S(n15599), .Z(n12866) );
  AOI22_X1 U15165 ( .A1(n13162), .A2(n12991), .B1(n13011), .B2(n12864), .ZN(
        n12865) );
  OAI211_X1 U15166 ( .C1(n13165), .C2(n13007), .A(n12866), .B(n12865), .ZN(
        P3_U3211) );
  XNOR2_X1 U15167 ( .A(n12867), .B(n12873), .ZN(n13171) );
  INV_X1 U15168 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12877) );
  INV_X1 U15169 ( .A(n12868), .ZN(n12869) );
  NOR2_X1 U15170 ( .A1(n12915), .A2(n12869), .ZN(n12872) );
  OAI21_X1 U15171 ( .B1(n12872), .B2(n12871), .A(n12870), .ZN(n12874) );
  XNOR2_X1 U15172 ( .A(n12874), .B(n12873), .ZN(n12876) );
  AOI222_X1 U15173 ( .A1(n15611), .A2(n12876), .B1(n12875), .B2(n15656), .C1(
        n12908), .C2(n15638), .ZN(n13166) );
  MUX2_X1 U15174 ( .A(n12877), .B(n13166), .S(n15599), .Z(n12880) );
  AOI22_X1 U15175 ( .A1(n13168), .A2(n12991), .B1(n13011), .B2(n12878), .ZN(
        n12879) );
  OAI211_X1 U15176 ( .C1(n13171), .C2(n13007), .A(n12880), .B(n12879), .ZN(
        P3_U3212) );
  NAND2_X1 U15177 ( .A1(n12881), .A2(n12887), .ZN(n12882) );
  NAND2_X1 U15178 ( .A1(n12883), .A2(n12882), .ZN(n13175) );
  NAND2_X1 U15179 ( .A1(n12903), .A2(n12886), .ZN(n12888) );
  XNOR2_X1 U15180 ( .A(n12888), .B(n12887), .ZN(n12890) );
  OAI22_X1 U15181 ( .A1(n12890), .A2(n13052), .B1(n12889), .B2(n15642), .ZN(
        n13071) );
  NAND2_X1 U15182 ( .A1(n13071), .A2(n15599), .ZN(n12895) );
  AOI22_X1 U15183 ( .A1(n12891), .A2(n13011), .B1(n15601), .B2(
        P3_REG2_REG_20__SCAN_IN), .ZN(n12892) );
  OAI21_X1 U15184 ( .B1(n13070), .B2(n12989), .A(n12892), .ZN(n12893) );
  AOI21_X1 U15185 ( .B1(n13073), .B2(n12991), .A(n12893), .ZN(n12894) );
  OAI211_X1 U15186 ( .C1(n13175), .C2(n13007), .A(n12895), .B(n12894), .ZN(
        P3_U3213) );
  AOI21_X1 U15187 ( .B1(n12927), .B2(n12897), .A(n12896), .ZN(n12920) );
  NAND2_X1 U15188 ( .A1(n12920), .A2(n6867), .ZN(n13081) );
  NAND2_X1 U15189 ( .A1(n13081), .A2(n12898), .ZN(n12899) );
  XOR2_X1 U15190 ( .A(n12900), .B(n12899), .Z(n13181) );
  INV_X1 U15191 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12909) );
  NOR2_X1 U15192 ( .A1(n13085), .A2(n15652), .ZN(n12907) );
  INV_X1 U15193 ( .A(n12914), .ZN(n12902) );
  AOI21_X1 U15194 ( .B1(n12902), .B2(n12901), .A(n12900), .ZN(n12905) );
  INV_X1 U15195 ( .A(n12903), .ZN(n12904) );
  NOR3_X1 U15196 ( .A1(n12905), .A2(n12904), .A3(n13052), .ZN(n12906) );
  AOI211_X1 U15197 ( .C1(n15656), .C2(n12908), .A(n12907), .B(n12906), .ZN(
        n13176) );
  MUX2_X1 U15198 ( .A(n12909), .B(n13176), .S(n15599), .Z(n12913) );
  INV_X1 U15199 ( .A(n12910), .ZN(n13178) );
  AOI22_X1 U15200 ( .A1(n13178), .A2(n13004), .B1(n13011), .B2(n12911), .ZN(
        n12912) );
  OAI211_X1 U15201 ( .C1(n13181), .C2(n13007), .A(n12913), .B(n12912), .ZN(
        P3_U3214) );
  AOI21_X1 U15202 ( .B1(n6867), .B2(n12915), .A(n12914), .ZN(n12916) );
  OAI222_X1 U15203 ( .A1(n15642), .A2(n13070), .B1(n15652), .B2(n13091), .C1(
        n13052), .C2(n12916), .ZN(n13080) );
  INV_X1 U15204 ( .A(n13080), .ZN(n12926) );
  INV_X1 U15205 ( .A(n12917), .ZN(n12918) );
  OAI22_X1 U15206 ( .A1(n15599), .A2(n12919), .B1(n12918), .B2(n15588), .ZN(
        n12923) );
  NOR2_X1 U15207 ( .A1(n12920), .A2(n6867), .ZN(n13079) );
  INV_X1 U15208 ( .A(n13081), .ZN(n12921) );
  NOR3_X1 U15209 ( .A1(n13079), .A2(n12921), .A3(n13007), .ZN(n12922) );
  AOI211_X1 U15210 ( .C1(n12991), .C2(n12924), .A(n12923), .B(n12922), .ZN(
        n12925) );
  OAI21_X1 U15211 ( .B1(n12926), .B2(n15601), .A(n12925), .ZN(P3_U3215) );
  XNOR2_X1 U15212 ( .A(n12927), .B(n12932), .ZN(n13189) );
  NAND2_X1 U15213 ( .A1(n12929), .A2(n12928), .ZN(n12942) );
  NAND2_X1 U15214 ( .A1(n12942), .A2(n12941), .ZN(n12931) );
  NAND2_X1 U15215 ( .A1(n12931), .A2(n12930), .ZN(n12933) );
  XNOR2_X1 U15216 ( .A(n12933), .B(n12932), .ZN(n12934) );
  OAI22_X1 U15217 ( .A1(n12934), .A2(n13052), .B1(n13097), .B2(n15652), .ZN(
        n13086) );
  NAND2_X1 U15218 ( .A1(n13086), .A2(n15599), .ZN(n12939) );
  AOI22_X1 U15219 ( .A1(n15601), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n13011), 
        .B2(n12935), .ZN(n12936) );
  OAI21_X1 U15220 ( .B1(n12957), .B2(n13085), .A(n12936), .ZN(n12937) );
  AOI21_X1 U15221 ( .B1(n13088), .B2(n13004), .A(n12937), .ZN(n12938) );
  OAI211_X1 U15222 ( .C1(n13189), .C2(n13007), .A(n12939), .B(n12938), .ZN(
        P3_U3216) );
  XNOR2_X1 U15223 ( .A(n12940), .B(n12941), .ZN(n13193) );
  XNOR2_X1 U15224 ( .A(n12942), .B(n12941), .ZN(n12944) );
  OAI22_X1 U15225 ( .A1(n12944), .A2(n13052), .B1(n12943), .B2(n15652), .ZN(
        n13092) );
  NAND2_X1 U15226 ( .A1(n13092), .A2(n15599), .ZN(n12949) );
  AOI22_X1 U15227 ( .A1(n15601), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n13011), 
        .B2(n12945), .ZN(n12946) );
  OAI21_X1 U15228 ( .B1(n12957), .B2(n13091), .A(n12946), .ZN(n12947) );
  AOI21_X1 U15229 ( .B1(n13094), .B2(n13004), .A(n12947), .ZN(n12948) );
  OAI211_X1 U15230 ( .C1(n13193), .C2(n13007), .A(n12949), .B(n12948), .ZN(
        P3_U3217) );
  XNOR2_X1 U15231 ( .A(n12950), .B(n12952), .ZN(n13197) );
  XNOR2_X1 U15232 ( .A(n12951), .B(n12952), .ZN(n12954) );
  OAI22_X1 U15233 ( .A1(n12954), .A2(n13052), .B1(n12953), .B2(n15652), .ZN(
        n13098) );
  NAND2_X1 U15234 ( .A1(n13098), .A2(n15599), .ZN(n12960) );
  AOI22_X1 U15235 ( .A1(n15601), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n13011), 
        .B2(n12955), .ZN(n12956) );
  OAI21_X1 U15236 ( .B1(n12957), .B2(n13097), .A(n12956), .ZN(n12958) );
  AOI21_X1 U15237 ( .B1(n13100), .B2(n13004), .A(n12958), .ZN(n12959) );
  OAI211_X1 U15238 ( .C1(n13197), .C2(n13007), .A(n12960), .B(n12959), .ZN(
        P3_U3218) );
  XOR2_X1 U15239 ( .A(n12961), .B(n12966), .Z(n13203) );
  NAND2_X1 U15240 ( .A1(n12962), .A2(n12974), .ZN(n12964) );
  NAND2_X1 U15241 ( .A1(n12964), .A2(n12963), .ZN(n12965) );
  XOR2_X1 U15242 ( .A(n12966), .B(n12965), .Z(n12969) );
  AOI222_X1 U15243 ( .A1(n15611), .A2(n12969), .B1(n12968), .B2(n15656), .C1(
        n12967), .C2(n15638), .ZN(n13198) );
  MUX2_X1 U15244 ( .A(n12970), .B(n13198), .S(n15599), .Z(n12973) );
  AOI22_X1 U15245 ( .A1(n13200), .A2(n13004), .B1(n13011), .B2(n12971), .ZN(
        n12972) );
  OAI211_X1 U15246 ( .C1(n13203), .C2(n13007), .A(n12973), .B(n12972), .ZN(
        P3_U3219) );
  XNOR2_X1 U15247 ( .A(n12974), .B(n12975), .ZN(n13209) );
  XNOR2_X1 U15248 ( .A(n12962), .B(n6695), .ZN(n12977) );
  AOI222_X1 U15249 ( .A1(n15611), .A2(n12977), .B1(n12976), .B2(n15656), .C1(
        n12999), .C2(n15638), .ZN(n13204) );
  MUX2_X1 U15250 ( .A(n12978), .B(n13204), .S(n15599), .Z(n12981) );
  AOI22_X1 U15251 ( .A1(n13206), .A2(n13004), .B1(n13011), .B2(n12979), .ZN(
        n12980) );
  OAI211_X1 U15252 ( .C1(n13209), .C2(n13007), .A(n12981), .B(n12980), .ZN(
        P3_U3220) );
  XNOR2_X1 U15253 ( .A(n12982), .B(n12984), .ZN(n13213) );
  XNOR2_X1 U15254 ( .A(n12983), .B(n12984), .ZN(n12986) );
  OAI22_X1 U15255 ( .A1(n12986), .A2(n13052), .B1(n12985), .B2(n15642), .ZN(
        n13109) );
  NAND2_X1 U15256 ( .A1(n13109), .A2(n15599), .ZN(n12993) );
  AOI22_X1 U15257 ( .A1(n15601), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n13011), 
        .B2(n12987), .ZN(n12988) );
  OAI21_X1 U15258 ( .B1(n12989), .B2(n13119), .A(n12988), .ZN(n12990) );
  AOI21_X1 U15259 ( .B1(n12991), .B2(n13111), .A(n12990), .ZN(n12992) );
  OAI211_X1 U15260 ( .C1(n13213), .C2(n13007), .A(n12993), .B(n12992), .ZN(
        P3_U3221) );
  XNOR2_X1 U15261 ( .A(n12995), .B(n12994), .ZN(n13221) );
  XNOR2_X1 U15262 ( .A(n12996), .B(n12997), .ZN(n13000) );
  AOI222_X1 U15263 ( .A1(n15611), .A2(n13000), .B1(n12999), .B2(n15656), .C1(
        n12998), .C2(n15638), .ZN(n13214) );
  MUX2_X1 U15264 ( .A(n13001), .B(n13214), .S(n15599), .Z(n13006) );
  INV_X1 U15265 ( .A(n13002), .ZN(n13216) );
  AOI22_X1 U15266 ( .A1(n13216), .A2(n13004), .B1(n13011), .B2(n13003), .ZN(
        n13005) );
  OAI211_X1 U15267 ( .C1(n13221), .C2(n13007), .A(n13006), .B(n13005), .ZN(
        P3_U3222) );
  XNOR2_X1 U15268 ( .A(n13018), .B(n13008), .ZN(n15603) );
  AOI22_X1 U15269 ( .A1(n13010), .A2(n15603), .B1(n13009), .B2(n15605), .ZN(
        n13023) );
  AOI22_X1 U15270 ( .A1(n13013), .A2(n13012), .B1(n13011), .B2(
        P3_REG3_REG_1__SCAN_IN), .ZN(n13022) );
  AND2_X1 U15271 ( .A1(n15637), .A2(n13014), .ZN(n15604) );
  NAND2_X1 U15272 ( .A1(n15604), .A2(n15586), .ZN(n13016) );
  MUX2_X1 U15273 ( .A(n13016), .B(n13015), .S(n15601), .Z(n13021) );
  XNOR2_X1 U15274 ( .A(n13018), .B(n13017), .ZN(n15610) );
  NAND2_X1 U15275 ( .A1(n13019), .A2(n15610), .ZN(n13020) );
  NAND4_X1 U15276 ( .A1(n13023), .A2(n13022), .A3(n13021), .A4(n13020), .ZN(
        P3_U3232) );
  NOR2_X1 U15277 ( .A1(n13130), .A2(n15674), .ZN(n13025) );
  AOI21_X1 U15278 ( .B1(P3_REG1_REG_31__SCAN_IN), .B2(n15674), .A(n13025), 
        .ZN(n13024) );
  OAI21_X1 U15279 ( .B1(n13132), .B2(n9283), .A(n13024), .ZN(P3_U3490) );
  INV_X1 U15280 ( .A(n12309), .ZN(n13135) );
  AOI21_X1 U15281 ( .B1(P3_REG1_REG_30__SCAN_IN), .B2(n15674), .A(n13025), 
        .ZN(n13026) );
  OAI21_X1 U15282 ( .B1(n13135), .B2(n9283), .A(n13026), .ZN(P3_U3489) );
  AOI22_X1 U15283 ( .A1(n13140), .A2(n13049), .B1(n13115), .B2(n13139), .ZN(
        n13028) );
  NAND2_X1 U15284 ( .A1(n13029), .A2(n13028), .ZN(P3_U3488) );
  INV_X1 U15285 ( .A(n15659), .ZN(n15648) );
  AOI21_X1 U15286 ( .B1(n15648), .B2(n13031), .A(n13030), .ZN(n13142) );
  MUX2_X1 U15287 ( .A(n13032), .B(n13142), .S(n15676), .Z(n13033) );
  INV_X1 U15288 ( .A(n13034), .ZN(n13149) );
  AOI22_X1 U15289 ( .A1(n13036), .A2(n15656), .B1(n15638), .B2(n13035), .ZN(
        n13037) );
  OAI21_X1 U15290 ( .B1(n13038), .B2(n13138), .A(n13037), .ZN(n13039) );
  AOI21_X1 U15291 ( .B1(n13040), .B2(n15611), .A(n13039), .ZN(n13146) );
  MUX2_X1 U15292 ( .A(n13041), .B(n13146), .S(n15676), .Z(n13042) );
  OAI21_X1 U15293 ( .B1(n13149), .B2(n9283), .A(n13042), .ZN(P3_U3485) );
  OAI22_X1 U15294 ( .A1(n13043), .A2(n15642), .B1(n13058), .B2(n15652), .ZN(
        n13045) );
  AOI211_X1 U15295 ( .C1(n15637), .C2(n13046), .A(n13045), .B(n13044), .ZN(
        n13047) );
  OAI21_X1 U15296 ( .B1(n13138), .B2(n13048), .A(n13047), .ZN(n13150) );
  MUX2_X1 U15297 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n13150), .S(n15676), .Z(
        P3_U3484) );
  OAI22_X1 U15298 ( .A1(n13051), .A2(n15642), .B1(n13050), .B2(n15652), .ZN(
        n13055) );
  NOR2_X1 U15299 ( .A1(n13053), .A2(n13052), .ZN(n13054) );
  AOI211_X1 U15300 ( .C1(n15637), .C2(n13056), .A(n13055), .B(n13054), .ZN(
        n13152) );
  MUX2_X1 U15301 ( .A(n15677), .B(n13152), .S(n15676), .Z(n13057) );
  OAI21_X1 U15302 ( .B1(n13155), .B2(n13118), .A(n13057), .ZN(P3_U3483) );
  NOR2_X1 U15303 ( .A1(n13058), .A2(n15642), .ZN(n13060) );
  AOI211_X1 U15304 ( .C1(n15637), .C2(n13061), .A(n13060), .B(n13059), .ZN(
        n13156) );
  MUX2_X1 U15305 ( .A(n13062), .B(n13156), .S(n15676), .Z(n13063) );
  OAI21_X1 U15306 ( .B1(n13118), .B2(n13159), .A(n13063), .ZN(P3_U3482) );
  MUX2_X1 U15307 ( .A(n13064), .B(n13160), .S(n15676), .Z(n13066) );
  NAND2_X1 U15308 ( .A1(n13162), .A2(n13115), .ZN(n13065) );
  OAI211_X1 U15309 ( .C1(n13165), .C2(n13118), .A(n13066), .B(n13065), .ZN(
        P3_U3481) );
  MUX2_X1 U15310 ( .A(n13067), .B(n13166), .S(n15676), .Z(n13069) );
  NAND2_X1 U15311 ( .A1(n13168), .A2(n13115), .ZN(n13068) );
  OAI211_X1 U15312 ( .C1(n13118), .C2(n13171), .A(n13069), .B(n13068), .ZN(
        P3_U3480) );
  NOR2_X1 U15313 ( .A1(n13070), .A2(n15652), .ZN(n13072) );
  AOI211_X1 U15314 ( .C1(n15637), .C2(n13073), .A(n13072), .B(n13071), .ZN(
        n13172) );
  MUX2_X1 U15315 ( .A(n13074), .B(n13172), .S(n15676), .Z(n13075) );
  OAI21_X1 U15316 ( .B1(n13118), .B2(n13175), .A(n13075), .ZN(P3_U3479) );
  MUX2_X1 U15317 ( .A(n13076), .B(n13176), .S(n15676), .Z(n13078) );
  NAND2_X1 U15318 ( .A1(n13178), .A2(n13115), .ZN(n13077) );
  OAI211_X1 U15319 ( .C1(n13181), .C2(n13118), .A(n13078), .B(n13077), .ZN(
        P3_U3478) );
  INV_X1 U15320 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13083) );
  NOR2_X1 U15321 ( .A1(n13079), .A2(n13138), .ZN(n13082) );
  AOI21_X1 U15322 ( .B1(n13082), .B2(n13081), .A(n13080), .ZN(n13182) );
  MUX2_X1 U15323 ( .A(n13083), .B(n13182), .S(n15676), .Z(n13084) );
  OAI21_X1 U15324 ( .B1(n13185), .B2(n9283), .A(n13084), .ZN(P3_U3477) );
  NOR2_X1 U15325 ( .A1(n13085), .A2(n15642), .ZN(n13087) );
  AOI211_X1 U15326 ( .C1(n15637), .C2(n13088), .A(n13087), .B(n13086), .ZN(
        n13186) );
  MUX2_X1 U15327 ( .A(n13089), .B(n13186), .S(n15676), .Z(n13090) );
  OAI21_X1 U15328 ( .B1(n13118), .B2(n13189), .A(n13090), .ZN(P3_U3476) );
  NOR2_X1 U15329 ( .A1(n13091), .A2(n15642), .ZN(n13093) );
  AOI211_X1 U15330 ( .C1(n15637), .C2(n13094), .A(n13093), .B(n13092), .ZN(
        n13190) );
  MUX2_X1 U15331 ( .A(n13095), .B(n13190), .S(n15676), .Z(n13096) );
  OAI21_X1 U15332 ( .B1(n13118), .B2(n13193), .A(n13096), .ZN(P3_U3475) );
  INV_X1 U15333 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13101) );
  NOR2_X1 U15334 ( .A1(n13097), .A2(n15642), .ZN(n13099) );
  AOI211_X1 U15335 ( .C1(n15637), .C2(n13100), .A(n13099), .B(n13098), .ZN(
        n13194) );
  MUX2_X1 U15336 ( .A(n13101), .B(n13194), .S(n15676), .Z(n13102) );
  OAI21_X1 U15337 ( .B1(n13118), .B2(n13197), .A(n13102), .ZN(P3_U3474) );
  MUX2_X1 U15338 ( .A(n13103), .B(n13198), .S(n15676), .Z(n13105) );
  NAND2_X1 U15339 ( .A1(n13200), .A2(n13115), .ZN(n13104) );
  OAI211_X1 U15340 ( .C1(n13203), .C2(n13118), .A(n13105), .B(n13104), .ZN(
        P3_U3473) );
  INV_X1 U15341 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n13106) );
  MUX2_X1 U15342 ( .A(n13106), .B(n13204), .S(n15676), .Z(n13108) );
  NAND2_X1 U15343 ( .A1(n13206), .A2(n13115), .ZN(n13107) );
  OAI211_X1 U15344 ( .C1(n13118), .C2(n13209), .A(n13108), .B(n13107), .ZN(
        P3_U3472) );
  NOR2_X1 U15345 ( .A1(n13119), .A2(n15652), .ZN(n13110) );
  AOI211_X1 U15346 ( .C1(n15637), .C2(n13111), .A(n13110), .B(n13109), .ZN(
        n13210) );
  MUX2_X1 U15347 ( .A(n13112), .B(n13210), .S(n15676), .Z(n13113) );
  OAI21_X1 U15348 ( .B1(n13118), .B2(n13213), .A(n13113), .ZN(P3_U3471) );
  INV_X1 U15349 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n13114) );
  MUX2_X1 U15350 ( .A(n13114), .B(n13214), .S(n15676), .Z(n13117) );
  NAND2_X1 U15351 ( .A1(n13115), .A2(n13216), .ZN(n13116) );
  OAI211_X1 U15352 ( .C1(n13118), .C2(n13221), .A(n13117), .B(n13116), .ZN(
        P3_U3470) );
  OAI22_X1 U15353 ( .A1(n13120), .A2(n15652), .B1(n13119), .B2(n15642), .ZN(
        n13121) );
  AOI21_X1 U15354 ( .B1(n13122), .B2(n15637), .A(n13121), .ZN(n13123) );
  OAI211_X1 U15355 ( .C1(n13138), .C2(n13125), .A(n13124), .B(n13123), .ZN(
        n13222) );
  MUX2_X1 U15356 ( .A(n13222), .B(P3_REG1_REG_10__SCAN_IN), .S(n15674), .Z(
        P3_U3469) );
  AOI21_X1 U15357 ( .B1(n15637), .B2(n13127), .A(n13126), .ZN(n13128) );
  OAI21_X1 U15358 ( .B1(n13138), .B2(n13129), .A(n13128), .ZN(n13223) );
  MUX2_X1 U15359 ( .A(P3_REG1_REG_8__SCAN_IN), .B(n13223), .S(n15676), .Z(
        P3_U3467) );
  NOR2_X1 U15360 ( .A1(n13130), .A2(n15664), .ZN(n13133) );
  AOI21_X1 U15361 ( .B1(n15664), .B2(P3_REG0_REG_31__SCAN_IN), .A(n13133), 
        .ZN(n13131) );
  OAI21_X1 U15362 ( .B1(n13132), .B2(n9296), .A(n13131), .ZN(P3_U3458) );
  AOI21_X1 U15363 ( .B1(n15664), .B2(P3_REG0_REG_30__SCAN_IN), .A(n13133), 
        .ZN(n13134) );
  OAI21_X1 U15364 ( .B1(n13135), .B2(n9296), .A(n13134), .ZN(P3_U3457) );
  INV_X1 U15365 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n13137) );
  NOR2_X1 U15366 ( .A1(n15664), .A2(n13138), .ZN(n13151) );
  AOI22_X1 U15367 ( .A1(n13140), .A2(n13151), .B1(n13217), .B2(n13139), .ZN(
        n13141) );
  INV_X1 U15368 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13143) );
  MUX2_X1 U15369 ( .A(n13143), .B(n13142), .S(n15666), .Z(n13144) );
  INV_X1 U15370 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13147) );
  MUX2_X1 U15371 ( .A(n13147), .B(n13146), .S(n15666), .Z(n13148) );
  OAI21_X1 U15372 ( .B1(n13149), .B2(n9296), .A(n13148), .ZN(P3_U3453) );
  MUX2_X1 U15373 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n13150), .S(n15666), .Z(
        P3_U3452) );
  INV_X1 U15374 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13153) );
  MUX2_X1 U15375 ( .A(n13153), .B(n13152), .S(n15666), .Z(n13154) );
  OAI21_X1 U15376 ( .B1(n13155), .B2(n13220), .A(n13154), .ZN(P3_U3451) );
  INV_X1 U15377 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13157) );
  MUX2_X1 U15378 ( .A(n13157), .B(n13156), .S(n15666), .Z(n13158) );
  OAI21_X1 U15379 ( .B1(n13159), .B2(n13220), .A(n13158), .ZN(P3_U3450) );
  INV_X1 U15380 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13161) );
  MUX2_X1 U15381 ( .A(n13161), .B(n13160), .S(n15666), .Z(n13164) );
  NAND2_X1 U15382 ( .A1(n13162), .A2(n13217), .ZN(n13163) );
  OAI211_X1 U15383 ( .C1(n13165), .C2(n13220), .A(n13164), .B(n13163), .ZN(
        P3_U3449) );
  INV_X1 U15384 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13167) );
  MUX2_X1 U15385 ( .A(n13167), .B(n13166), .S(n15666), .Z(n13170) );
  NAND2_X1 U15386 ( .A1(n13168), .A2(n13217), .ZN(n13169) );
  OAI211_X1 U15387 ( .C1(n13171), .C2(n13220), .A(n13170), .B(n13169), .ZN(
        P3_U3448) );
  INV_X1 U15388 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13173) );
  MUX2_X1 U15389 ( .A(n13173), .B(n13172), .S(n15666), .Z(n13174) );
  OAI21_X1 U15390 ( .B1(n13175), .B2(n13220), .A(n13174), .ZN(P3_U3447) );
  INV_X1 U15391 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13177) );
  MUX2_X1 U15392 ( .A(n13177), .B(n13176), .S(n15666), .Z(n13180) );
  NAND2_X1 U15393 ( .A1(n13178), .A2(n13217), .ZN(n13179) );
  OAI211_X1 U15394 ( .C1(n13181), .C2(n13220), .A(n13180), .B(n13179), .ZN(
        P3_U3446) );
  INV_X1 U15395 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13183) );
  MUX2_X1 U15396 ( .A(n13183), .B(n13182), .S(n15666), .Z(n13184) );
  OAI21_X1 U15397 ( .B1(n13185), .B2(n9296), .A(n13184), .ZN(P3_U3444) );
  INV_X1 U15398 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13187) );
  MUX2_X1 U15399 ( .A(n13187), .B(n13186), .S(n15666), .Z(n13188) );
  OAI21_X1 U15400 ( .B1(n13189), .B2(n13220), .A(n13188), .ZN(P3_U3441) );
  INV_X1 U15401 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13191) );
  MUX2_X1 U15402 ( .A(n13191), .B(n13190), .S(n15666), .Z(n13192) );
  OAI21_X1 U15403 ( .B1(n13193), .B2(n13220), .A(n13192), .ZN(P3_U3438) );
  INV_X1 U15404 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13195) );
  MUX2_X1 U15405 ( .A(n13195), .B(n13194), .S(n15666), .Z(n13196) );
  OAI21_X1 U15406 ( .B1(n13197), .B2(n13220), .A(n13196), .ZN(P3_U3435) );
  MUX2_X1 U15407 ( .A(n13199), .B(n13198), .S(n15666), .Z(n13202) );
  NAND2_X1 U15408 ( .A1(n13200), .A2(n13217), .ZN(n13201) );
  OAI211_X1 U15409 ( .C1(n13203), .C2(n13220), .A(n13202), .B(n13201), .ZN(
        P3_U3432) );
  MUX2_X1 U15410 ( .A(n13205), .B(n13204), .S(n15666), .Z(n13208) );
  NAND2_X1 U15411 ( .A1(n13206), .A2(n13217), .ZN(n13207) );
  OAI211_X1 U15412 ( .C1(n13209), .C2(n13220), .A(n13208), .B(n13207), .ZN(
        P3_U3429) );
  MUX2_X1 U15413 ( .A(n13211), .B(n13210), .S(n15666), .Z(n13212) );
  OAI21_X1 U15414 ( .B1(n13213), .B2(n13220), .A(n13212), .ZN(P3_U3426) );
  MUX2_X1 U15415 ( .A(n13215), .B(n13214), .S(n15666), .Z(n13219) );
  NAND2_X1 U15416 ( .A1(n13217), .A2(n13216), .ZN(n13218) );
  OAI211_X1 U15417 ( .C1(n13221), .C2(n13220), .A(n13219), .B(n13218), .ZN(
        P3_U3423) );
  MUX2_X1 U15418 ( .A(n13222), .B(P3_REG0_REG_10__SCAN_IN), .S(n15664), .Z(
        P3_U3420) );
  MUX2_X1 U15419 ( .A(P3_REG0_REG_8__SCAN_IN), .B(n13223), .S(n15666), .Z(
        P3_U3414) );
  MUX2_X1 U15420 ( .A(P3_D_REG_1__SCAN_IN), .B(n13225), .S(n13224), .Z(
        P3_U3377) );
  INV_X1 U15421 ( .A(n13226), .ZN(n13228) );
  OAI21_X1 U15422 ( .B1(n13229), .B2(n13228), .A(n13227), .ZN(n13231) );
  XNOR2_X1 U15423 ( .A(n13231), .B(n13230), .ZN(n13236) );
  NOR4_X1 U15424 ( .A1(n13232), .A2(P3_IR_REG_30__SCAN_IN), .A3(P3_U3151), 
        .A4(n7647), .ZN(n13233) );
  AOI21_X1 U15425 ( .B1(n13234), .B2(SI_31_), .A(n13233), .ZN(n13235) );
  OAI21_X1 U15426 ( .B1(n13236), .B2(n13248), .A(n13235), .ZN(P3_U3264) );
  INV_X1 U15427 ( .A(n13237), .ZN(n13239) );
  OAI222_X1 U15428 ( .A1(n13250), .A2(n13240), .B1(n13248), .B2(n13239), .C1(
        P3_U3151), .C2(n13238), .ZN(P3_U3266) );
  INV_X1 U15429 ( .A(n13241), .ZN(n13244) );
  OAI222_X1 U15430 ( .A1(n13260), .A2(n13244), .B1(n13243), .B2(P3_U3151), 
        .C1(n13242), .C2(n13256), .ZN(P3_U3267) );
  INV_X1 U15431 ( .A(n13245), .ZN(n13247) );
  OAI222_X1 U15432 ( .A1(n13250), .A2(n13249), .B1(n13248), .B2(n13247), .C1(
        P3_U3151), .C2(n13246), .ZN(P3_U3268) );
  INV_X1 U15433 ( .A(n13251), .ZN(n13254) );
  INV_X1 U15434 ( .A(SI_26_), .ZN(n13252) );
  OAI222_X1 U15435 ( .A1(n13260), .A2(n13254), .B1(P3_U3151), .B2(n13253), 
        .C1(n13252), .C2(n13256), .ZN(P3_U3269) );
  INV_X1 U15436 ( .A(n13255), .ZN(n13259) );
  INV_X1 U15437 ( .A(SI_25_), .ZN(n13257) );
  OAI222_X1 U15438 ( .A1(n13260), .A2(n13259), .B1(P3_U3151), .B2(n13258), 
        .C1(n13257), .C2(n13256), .ZN(P3_U3270) );
  XNOR2_X1 U15439 ( .A(n13974), .B(n7172), .ZN(n13374) );
  NAND2_X1 U15440 ( .A1(n13811), .A2(n13300), .ZN(n13370) );
  XNOR2_X1 U15441 ( .A(n13374), .B(n13370), .ZN(n13365) );
  INV_X1 U15442 ( .A(n13261), .ZN(n13264) );
  INV_X1 U15443 ( .A(n13262), .ZN(n13263) );
  INV_X1 U15444 ( .A(n13265), .ZN(n13266) );
  NAND2_X1 U15445 ( .A1(n13267), .A2(n13266), .ZN(n13268) );
  XNOR2_X1 U15446 ( .A(n14184), .B(n13314), .ZN(n13271) );
  NAND2_X1 U15447 ( .A1(n14191), .A2(n13300), .ZN(n13270) );
  NAND2_X1 U15448 ( .A1(n13271), .A2(n13270), .ZN(n13272) );
  OAI21_X1 U15449 ( .B1(n13271), .B2(n13270), .A(n13272), .ZN(n13332) );
  XNOR2_X1 U15450 ( .A(n14166), .B(n7172), .ZN(n13274) );
  AND2_X1 U15451 ( .A1(n13818), .A2(n13300), .ZN(n13273) );
  NOR2_X1 U15452 ( .A1(n13274), .A2(n13273), .ZN(n13485) );
  NAND2_X1 U15453 ( .A1(n13274), .A2(n13273), .ZN(n13483) );
  AND2_X1 U15454 ( .A1(n13817), .A2(n13300), .ZN(n13276) );
  XNOR2_X1 U15455 ( .A(n14341), .B(n7172), .ZN(n13275) );
  NOR2_X1 U15456 ( .A1(n13275), .A2(n13276), .ZN(n13282) );
  AOI21_X1 U15457 ( .B1(n13276), .B2(n13275), .A(n13282), .ZN(n13405) );
  XNOR2_X1 U15458 ( .A(n14127), .B(n7172), .ZN(n13278) );
  AND2_X1 U15459 ( .A1(n13816), .A2(n15561), .ZN(n13279) );
  NOR2_X1 U15460 ( .A1(n13278), .A2(n13279), .ZN(n13277) );
  INV_X1 U15461 ( .A(n13277), .ZN(n13283) );
  AOI21_X1 U15462 ( .B1(n13279), .B2(n13278), .A(n13277), .ZN(n13426) );
  OR2_X1 U15463 ( .A1(n13277), .A2(n13426), .ZN(n13281) );
  AND2_X1 U15464 ( .A1(n13405), .A2(n13281), .ZN(n13280) );
  INV_X1 U15465 ( .A(n13281), .ZN(n13285) );
  INV_X1 U15466 ( .A(n13282), .ZN(n13422) );
  AND2_X1 U15467 ( .A1(n13422), .A2(n13283), .ZN(n13284) );
  OR2_X1 U15468 ( .A1(n13285), .A2(n13284), .ZN(n13286) );
  NAND2_X1 U15469 ( .A1(n13287), .A2(n13286), .ZN(n13457) );
  NAND2_X1 U15470 ( .A1(n13815), .A2(n15561), .ZN(n13289) );
  XNOR2_X1 U15471 ( .A(n13648), .B(n7172), .ZN(n13288) );
  XOR2_X1 U15472 ( .A(n13289), .B(n13288), .Z(n13458) );
  XNOR2_X1 U15473 ( .A(n14105), .B(n13314), .ZN(n13291) );
  NAND2_X1 U15474 ( .A1(n13814), .A2(n15561), .ZN(n13290) );
  NAND2_X1 U15475 ( .A1(n13291), .A2(n13290), .ZN(n13292) );
  OAI21_X1 U15476 ( .B1(n13291), .B2(n13290), .A(n13292), .ZN(n13357) );
  AND2_X1 U15477 ( .A1(n13813), .A2(n13300), .ZN(n13294) );
  XNOR2_X1 U15478 ( .A(n14092), .B(n7172), .ZN(n13293) );
  NOR2_X1 U15479 ( .A1(n13293), .A2(n13294), .ZN(n13295) );
  AOI21_X1 U15480 ( .B1(n13294), .B2(n13293), .A(n13295), .ZN(n13442) );
  INV_X1 U15481 ( .A(n13295), .ZN(n13296) );
  NAND2_X1 U15482 ( .A1(n13812), .A2(n15561), .ZN(n13297) );
  XNOR2_X1 U15483 ( .A(n14073), .B(n7172), .ZN(n13299) );
  XOR2_X1 U15484 ( .A(n13297), .B(n13299), .Z(n13388) );
  INV_X1 U15485 ( .A(n13297), .ZN(n13298) );
  XNOR2_X1 U15486 ( .A(n14059), .B(n7172), .ZN(n13304) );
  INV_X1 U15487 ( .A(n13452), .ZN(n13303) );
  XNOR2_X1 U15488 ( .A(n14047), .B(n7172), .ZN(n13342) );
  AND2_X1 U15489 ( .A1(n14039), .A2(n13300), .ZN(n13339) );
  OAI21_X1 U15490 ( .B1(n13342), .B2(n14024), .A(n13339), .ZN(n13301) );
  NAND2_X1 U15491 ( .A1(n13305), .A2(n13304), .ZN(n13340) );
  AND2_X1 U15492 ( .A1(n14024), .A2(n15561), .ZN(n13306) );
  NOR2_X1 U15493 ( .A1(n13342), .A2(n13306), .ZN(n13308) );
  INV_X1 U15494 ( .A(n13342), .ZN(n13307) );
  INV_X1 U15495 ( .A(n13306), .ZN(n13341) );
  XNOR2_X1 U15496 ( .A(n14217), .B(n7172), .ZN(n13312) );
  NAND2_X1 U15497 ( .A1(n14041), .A2(n15561), .ZN(n13310) );
  XNOR2_X1 U15498 ( .A(n13312), .B(n13310), .ZN(n13432) );
  INV_X1 U15499 ( .A(n13310), .ZN(n13311) );
  NAND2_X1 U15500 ( .A1(n13312), .A2(n13311), .ZN(n13395) );
  XNOR2_X1 U15501 ( .A(n14008), .B(n7172), .ZN(n13319) );
  NAND2_X1 U15502 ( .A1(n14026), .A2(n15561), .ZN(n13318) );
  INV_X1 U15503 ( .A(n13318), .ZN(n13313) );
  NAND2_X1 U15504 ( .A1(n13319), .A2(n13313), .ZN(n13317) );
  AND2_X1 U15505 ( .A1(n13395), .A2(n13317), .ZN(n13466) );
  NAND2_X1 U15506 ( .A1(n14004), .A2(n15561), .ZN(n13315) );
  INV_X1 U15507 ( .A(n13317), .ZN(n13320) );
  XNOR2_X1 U15508 ( .A(n13319), .B(n13318), .ZN(n13396) );
  OR2_X1 U15509 ( .A1(n13473), .A2(n13468), .ZN(n13321) );
  NAND2_X1 U15510 ( .A1(n13470), .A2(n13368), .ZN(n13323) );
  XOR2_X1 U15511 ( .A(n13365), .B(n13323), .Z(n13328) );
  AOI22_X1 U15512 ( .A1(n13973), .A2(n13495), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13325) );
  INV_X1 U15513 ( .A(n13492), .ZN(n13352) );
  NAND2_X1 U15514 ( .A1(n14004), .A2(n13352), .ZN(n13324) );
  OAI211_X1 U15515 ( .C1(n13719), .C2(n13491), .A(n13325), .B(n13324), .ZN(
        n13326) );
  AOI21_X1 U15516 ( .B1(n13974), .B2(n13479), .A(n13326), .ZN(n13327) );
  OAI21_X1 U15517 ( .B1(n13328), .B2(n13481), .A(n13327), .ZN(P2_U3186) );
  INV_X1 U15518 ( .A(n13329), .ZN(n13330) );
  AOI21_X1 U15519 ( .B1(n13332), .B2(n13331), .A(n13330), .ZN(n13338) );
  AOI22_X1 U15520 ( .A1(n13818), .A2(n14190), .B1(n13819), .B2(n14188), .ZN(
        n14288) );
  INV_X1 U15521 ( .A(n13333), .ZN(n14178) );
  NAND2_X1 U15522 ( .A1(n13495), .A2(n14178), .ZN(n13335) );
  OAI211_X1 U15523 ( .C1(n14288), .C2(n13461), .A(n13335), .B(n13334), .ZN(
        n13336) );
  AOI21_X1 U15524 ( .B1(n14184), .B2(n13479), .A(n13336), .ZN(n13337) );
  OAI21_X1 U15525 ( .B1(n13338), .B2(n13481), .A(n13337), .ZN(P2_U3187) );
  INV_X1 U15526 ( .A(n13339), .ZN(n13451) );
  OAI21_X1 U15527 ( .B1(n13452), .B2(n13451), .A(n13340), .ZN(n13344) );
  XNOR2_X1 U15528 ( .A(n13342), .B(n13341), .ZN(n13343) );
  XNOR2_X1 U15529 ( .A(n13344), .B(n13343), .ZN(n13349) );
  OAI22_X1 U15530 ( .A1(n14043), .A2(n13459), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15749), .ZN(n13345) );
  AOI21_X1 U15531 ( .B1(n13352), .B2(n14039), .A(n13345), .ZN(n13346) );
  OAI21_X1 U15532 ( .B1(n13400), .B2(n13491), .A(n13346), .ZN(n13347) );
  AOI21_X1 U15533 ( .B1(n14047), .B2(n13479), .A(n13347), .ZN(n13348) );
  OAI21_X1 U15534 ( .B1(n13349), .B2(n13481), .A(n13348), .ZN(P2_U3188) );
  OAI211_X1 U15535 ( .C1(n6458), .C2(n13351), .A(n13350), .B(n13487), .ZN(
        n13356) );
  AOI22_X1 U15536 ( .A1(n13474), .A2(n13827), .B1(n13531), .B2(n13479), .ZN(
        n13355) );
  INV_X1 U15537 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n15451) );
  AOI22_X1 U15538 ( .A1(n13495), .A2(n15451), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13354) );
  NAND2_X1 U15539 ( .A1(n13352), .A2(n13829), .ZN(n13353) );
  NAND4_X1 U15540 ( .A1(n13356), .A2(n13355), .A3(n13354), .A4(n13353), .ZN(
        P2_U3190) );
  AOI21_X1 U15541 ( .B1(n13358), .B2(n13357), .A(n6529), .ZN(n13363) );
  AND2_X1 U15542 ( .A1(n13815), .A2(n14188), .ZN(n13359) );
  AOI21_X1 U15543 ( .B1(n13813), .B2(n14190), .A(n13359), .ZN(n14254) );
  NOR2_X1 U15544 ( .A1(n14254), .A2(n13461), .ZN(n13361) );
  NAND2_X1 U15545 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13937)
         );
  OAI21_X1 U15546 ( .B1(n13459), .B2(n14102), .A(n13937), .ZN(n13360) );
  AOI211_X1 U15547 ( .C1(n14105), .C2(n13479), .A(n13361), .B(n13360), .ZN(
        n13362) );
  OAI21_X1 U15548 ( .B1(n13363), .B2(n13481), .A(n13362), .ZN(P2_U3191) );
  INV_X1 U15549 ( .A(n13374), .ZN(n13364) );
  AND2_X1 U15550 ( .A1(n13810), .A2(n15561), .ZN(n13371) );
  INV_X1 U15551 ( .A(n13371), .ZN(n13369) );
  OAI21_X1 U15552 ( .B1(n13364), .B2(n13370), .A(n13369), .ZN(n13378) );
  INV_X1 U15553 ( .A(n13370), .ZN(n13367) );
  AOI21_X1 U15554 ( .B1(n13368), .B2(n13367), .A(n13371), .ZN(n13375) );
  MUX2_X1 U15555 ( .A(n13369), .B(n13368), .S(n13370), .Z(n13372) );
  AOI22_X1 U15556 ( .A1(n13372), .A2(n13374), .B1(n13371), .B2(n13370), .ZN(
        n13373) );
  OAI21_X1 U15557 ( .B1(n13375), .B2(n13374), .A(n13373), .ZN(n13376) );
  OAI211_X1 U15558 ( .C1(n13470), .C2(n13378), .A(n13377), .B(n13376), .ZN(
        n13381) );
  XOR2_X1 U15559 ( .A(n7172), .B(n13720), .Z(n13380) );
  XNOR2_X1 U15560 ( .A(n13381), .B(n13380), .ZN(n13387) );
  INV_X1 U15561 ( .A(n13382), .ZN(n13964) );
  AOI22_X1 U15562 ( .A1(n13964), .A2(n13495), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13384) );
  NAND2_X1 U15563 ( .A1(n13809), .A2(n13474), .ZN(n13383) );
  OAI211_X1 U15564 ( .C1(n13985), .C2(n13492), .A(n13384), .B(n13383), .ZN(
        n13385) );
  AOI21_X1 U15565 ( .B1(n13720), .B2(n13479), .A(n13385), .ZN(n13386) );
  OAI21_X1 U15566 ( .B1(n13387), .B2(n13481), .A(n13386), .ZN(P2_U3192) );
  XNOR2_X1 U15567 ( .A(n13389), .B(n13388), .ZN(n13394) );
  AND2_X1 U15568 ( .A1(n13813), .A2(n14188), .ZN(n13390) );
  AOI21_X1 U15569 ( .B1(n14039), .B2(n14190), .A(n13390), .ZN(n14239) );
  AOI22_X1 U15570 ( .A1(n14070), .A2(n13495), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13391) );
  OAI21_X1 U15571 ( .B1(n14239), .B2(n13461), .A(n13391), .ZN(n13392) );
  AOI21_X1 U15572 ( .B1(n14073), .B2(n13479), .A(n13392), .ZN(n13393) );
  OAI21_X1 U15573 ( .B1(n13394), .B2(n13481), .A(n13393), .ZN(P2_U3195) );
  NAND2_X1 U15574 ( .A1(n13467), .A2(n13395), .ZN(n13397) );
  XNOR2_X1 U15575 ( .A(n13397), .B(n13396), .ZN(n13403) );
  NAND2_X1 U15576 ( .A1(n14004), .A2(n13474), .ZN(n13399) );
  AOI22_X1 U15577 ( .A1(n14012), .A2(n13495), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13398) );
  OAI211_X1 U15578 ( .C1(n13400), .C2(n13492), .A(n13399), .B(n13398), .ZN(
        n13401) );
  AOI21_X1 U15579 ( .B1(n14008), .B2(n13479), .A(n13401), .ZN(n13402) );
  OAI21_X1 U15580 ( .B1(n13403), .B2(n13481), .A(n13402), .ZN(P2_U3197) );
  NAND2_X1 U15581 ( .A1(n13404), .A2(n13405), .ZN(n13423) );
  OAI21_X1 U15582 ( .B1(n13405), .B2(n13404), .A(n13423), .ZN(n13406) );
  NAND2_X1 U15583 ( .A1(n13406), .A2(n13487), .ZN(n13411) );
  INV_X1 U15584 ( .A(n14143), .ZN(n13409) );
  AND2_X1 U15585 ( .A1(n13818), .A2(n14188), .ZN(n13407) );
  AOI21_X1 U15586 ( .B1(n13816), .B2(n14190), .A(n13407), .ZN(n14141) );
  NAND2_X1 U15587 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n13874)
         );
  OAI21_X1 U15588 ( .B1(n14141), .B2(n13461), .A(n13874), .ZN(n13408) );
  AOI21_X1 U15589 ( .B1(n13409), .B2(n13495), .A(n13408), .ZN(n13410) );
  OAI211_X1 U15590 ( .C1(n7924), .C2(n13498), .A(n13411), .B(n13410), .ZN(
        P2_U3198) );
  NOR3_X1 U15591 ( .A1(n13413), .A2(n13412), .A3(n7930), .ZN(n13415) );
  OAI21_X1 U15592 ( .B1(n13415), .B2(n13414), .A(n13487), .ZN(n13421) );
  INV_X1 U15593 ( .A(n13416), .ZN(n15824) );
  AOI22_X1 U15594 ( .A1(n15826), .A2(n13479), .B1(n13495), .B2(n15824), .ZN(
        n13420) );
  NAND2_X1 U15595 ( .A1(n13825), .A2(n14190), .ZN(n13417) );
  OAI21_X1 U15596 ( .B1(n15544), .B2(n15495), .A(n13417), .ZN(n15555) );
  NAND2_X1 U15597 ( .A1(n13448), .A2(n15555), .ZN(n13418) );
  NAND4_X1 U15598 ( .A1(n13421), .A2(n13420), .A3(n13419), .A4(n13418), .ZN(
        P2_U3199) );
  NAND2_X1 U15599 ( .A1(n13423), .A2(n13422), .ZN(n13425) );
  NAND2_X1 U15600 ( .A1(n13425), .A2(n13426), .ZN(n13424) );
  OAI21_X1 U15601 ( .B1(n13426), .B2(n13425), .A(n13424), .ZN(n13427) );
  NAND2_X1 U15602 ( .A1(n13427), .A2(n13487), .ZN(n13431) );
  INV_X1 U15603 ( .A(n13428), .ZN(n14128) );
  AOI22_X1 U15604 ( .A1(n13815), .A2(n14190), .B1(n14188), .B2(n13817), .ZN(
        n14268) );
  NAND2_X1 U15605 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13904)
         );
  OAI21_X1 U15606 ( .B1(n14268), .B2(n13461), .A(n13904), .ZN(n13429) );
  AOI21_X1 U15607 ( .B1(n14128), .B2(n13495), .A(n13429), .ZN(n13430) );
  OAI211_X1 U15608 ( .C1(n7923), .C2(n13498), .A(n13431), .B(n13430), .ZN(
        P2_U3200) );
  XNOR2_X1 U15609 ( .A(n13433), .B(n13432), .ZN(n13439) );
  OAI22_X1 U15610 ( .A1(n14028), .A2(n13459), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13434), .ZN(n13436) );
  NOR2_X1 U15611 ( .A1(n13754), .A2(n13492), .ZN(n13435) );
  AOI211_X1 U15612 ( .C1(n13474), .C2(n14026), .A(n13436), .B(n13435), .ZN(
        n13438) );
  NAND2_X1 U15613 ( .A1(n14217), .A2(n13479), .ZN(n13437) );
  OAI211_X1 U15614 ( .C1(n13439), .C2(n13481), .A(n13438), .B(n13437), .ZN(
        P2_U3201) );
  OAI21_X1 U15615 ( .B1(n13442), .B2(n13441), .A(n13440), .ZN(n13443) );
  NAND2_X1 U15616 ( .A1(n13443), .A2(n13487), .ZN(n13450) );
  NAND2_X1 U15617 ( .A1(n13812), .A2(n14190), .ZN(n13445) );
  NAND2_X1 U15618 ( .A1(n13814), .A2(n14188), .ZN(n13444) );
  NAND2_X1 U15619 ( .A1(n13445), .A2(n13444), .ZN(n14087) );
  OAI22_X1 U15620 ( .A1(n13459), .A2(n14088), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13446), .ZN(n13447) );
  AOI21_X1 U15621 ( .B1(n14087), .B2(n13448), .A(n13447), .ZN(n13449) );
  OAI211_X1 U15622 ( .C1(n14335), .C2(n13498), .A(n13450), .B(n13449), .ZN(
        P2_U3205) );
  XNOR2_X1 U15623 ( .A(n13452), .B(n13451), .ZN(n13456) );
  AOI22_X1 U15624 ( .A1(n14024), .A2(n14190), .B1(n14188), .B2(n13812), .ZN(
        n14056) );
  AOI22_X1 U15625 ( .A1(n14060), .A2(n13495), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13453) );
  OAI21_X1 U15626 ( .B1(n14056), .B2(n13461), .A(n13453), .ZN(n13454) );
  AOI21_X1 U15627 ( .B1(n14059), .B2(n13479), .A(n13454), .ZN(n13455) );
  OAI21_X1 U15628 ( .B1(n13456), .B2(n13481), .A(n13455), .ZN(P2_U3207) );
  XNOR2_X1 U15629 ( .A(n13457), .B(n13458), .ZN(n13465) );
  NOR2_X1 U15630 ( .A1(n13459), .A2(n14115), .ZN(n13463) );
  AND2_X1 U15631 ( .A1(n13816), .A2(n14188), .ZN(n13460) );
  AOI21_X1 U15632 ( .B1(n13814), .B2(n14190), .A(n13460), .ZN(n14261) );
  NAND2_X1 U15633 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13919)
         );
  OAI21_X1 U15634 ( .B1(n14261), .B2(n13461), .A(n13919), .ZN(n13462) );
  AOI211_X1 U15635 ( .C1(n13648), .C2(n13479), .A(n13463), .B(n13462), .ZN(
        n13464) );
  OAI21_X1 U15636 ( .B1(n13465), .B2(n13481), .A(n13464), .ZN(P2_U3210) );
  NAND2_X1 U15637 ( .A1(n13467), .A2(n13466), .ZN(n13469) );
  AND2_X1 U15638 ( .A1(n13469), .A2(n13468), .ZN(n13472) );
  INV_X1 U15639 ( .A(n13470), .ZN(n13471) );
  AOI21_X1 U15640 ( .B1(n13473), .B2(n13472), .A(n13471), .ZN(n13482) );
  NAND2_X1 U15641 ( .A1(n13811), .A2(n13474), .ZN(n13477) );
  INV_X1 U15642 ( .A(n13475), .ZN(n13990) );
  AOI22_X1 U15643 ( .A1(n13990), .A2(n13495), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13476) );
  OAI211_X1 U15644 ( .C1(n13986), .C2(n13492), .A(n13477), .B(n13476), .ZN(
        n13478) );
  AOI21_X1 U15645 ( .B1(n14210), .B2(n13479), .A(n13478), .ZN(n13480) );
  OAI21_X1 U15646 ( .B1(n13482), .B2(n13481), .A(n13480), .ZN(P2_U3212) );
  INV_X1 U15647 ( .A(n13483), .ZN(n13488) );
  OAI21_X1 U15648 ( .B1(n13488), .B2(n13485), .A(n13484), .ZN(n13486) );
  OAI211_X1 U15649 ( .C1(n13489), .C2(n13488), .A(n13487), .B(n13486), .ZN(
        n13497) );
  INV_X1 U15650 ( .A(n13490), .ZN(n14167) );
  OAI22_X1 U15651 ( .A1(n13492), .A2(n14160), .B1(n14161), .B2(n13491), .ZN(
        n13493) );
  AOI211_X1 U15652 ( .C1(n13495), .C2(n14167), .A(n13494), .B(n13493), .ZN(
        n13496) );
  OAI211_X1 U15653 ( .C1(n14346), .C2(n13498), .A(n13497), .B(n13496), .ZN(
        P2_U3213) );
  NAND2_X1 U15654 ( .A1(n13499), .A2(n8559), .ZN(n13500) );
  INV_X2 U15655 ( .A(n13500), .ZN(n13530) );
  BUF_X4 U15656 ( .A(n13500), .Z(n13736) );
  OAI22_X1 U15657 ( .A1(n7918), .A2(n13738), .B1(n13501), .B2(n13736), .ZN(
        n13663) );
  INV_X1 U15658 ( .A(n13663), .ZN(n13666) );
  AOI22_X1 U15659 ( .A1(n14092), .A2(n13738), .B1(n13813), .B2(n13736), .ZN(
        n13661) );
  AOI21_X1 U15660 ( .B1(n13936), .B2(n8559), .A(n13742), .ZN(n13502) );
  AOI21_X1 U15661 ( .B1(n13503), .B2(n13736), .A(n13502), .ZN(n13506) );
  NAND2_X1 U15662 ( .A1(n13503), .A2(n13502), .ZN(n13505) );
  NAND3_X1 U15663 ( .A1(n13507), .A2(n13530), .A3(n7237), .ZN(n13504) );
  NAND2_X1 U15664 ( .A1(n13508), .A2(n13530), .ZN(n13510) );
  NAND2_X1 U15665 ( .A1(n13736), .A2(n15524), .ZN(n13509) );
  NAND2_X1 U15666 ( .A1(n13510), .A2(n13509), .ZN(n13519) );
  NAND2_X1 U15667 ( .A1(n13518), .A2(n13519), .ZN(n13514) );
  NAND2_X1 U15668 ( .A1(n13508), .A2(n13736), .ZN(n13511) );
  OAI21_X1 U15669 ( .B1(n13512), .B2(n13736), .A(n13511), .ZN(n13513) );
  NAND2_X1 U15670 ( .A1(n13514), .A2(n13513), .ZN(n13524) );
  AOI22_X1 U15671 ( .A1(n13829), .A2(n13738), .B1(n13515), .B2(n13736), .ZN(
        n13526) );
  NAND2_X1 U15672 ( .A1(n13829), .A2(n13736), .ZN(n13517) );
  NAND2_X1 U15673 ( .A1(n13526), .A2(n13525), .ZN(n13523) );
  NAND2_X1 U15674 ( .A1(n13521), .A2(n13520), .ZN(n13522) );
  INV_X1 U15675 ( .A(n13525), .ZN(n13528) );
  INV_X1 U15676 ( .A(n13526), .ZN(n13527) );
  NAND2_X1 U15677 ( .A1(n13528), .A2(n13527), .ZN(n13529) );
  NAND2_X1 U15678 ( .A1(n13828), .A2(n13738), .ZN(n13533) );
  NAND2_X1 U15679 ( .A1(n13736), .A2(n13531), .ZN(n13532) );
  NAND2_X1 U15680 ( .A1(n13533), .A2(n13532), .ZN(n13539) );
  NAND2_X1 U15681 ( .A1(n13538), .A2(n13539), .ZN(n13537) );
  NAND2_X1 U15682 ( .A1(n13828), .A2(n13736), .ZN(n13534) );
  OAI21_X1 U15683 ( .B1(n13535), .B2(n13736), .A(n13534), .ZN(n13536) );
  NAND2_X1 U15684 ( .A1(n13537), .A2(n13536), .ZN(n13543) );
  INV_X1 U15685 ( .A(n13538), .ZN(n13541) );
  INV_X1 U15686 ( .A(n13539), .ZN(n13540) );
  NAND2_X1 U15687 ( .A1(n13541), .A2(n13540), .ZN(n13542) );
  OAI22_X1 U15688 ( .A1(n15544), .A2(n13738), .B1(n15545), .B2(n13736), .ZN(
        n13545) );
  OAI22_X1 U15689 ( .A1(n15544), .A2(n13736), .B1(n15545), .B2(n13738), .ZN(
        n13544) );
  INV_X1 U15690 ( .A(n13545), .ZN(n13546) );
  NAND2_X1 U15691 ( .A1(n13826), .A2(n13738), .ZN(n13548) );
  NAND2_X1 U15692 ( .A1(n13736), .A2(n15826), .ZN(n13547) );
  NAND2_X1 U15693 ( .A1(n13826), .A2(n13736), .ZN(n13549) );
  OAI21_X1 U15694 ( .B1(n15566), .B2(n13736), .A(n13549), .ZN(n13550) );
  NAND2_X1 U15695 ( .A1(n13825), .A2(n13736), .ZN(n13552) );
  NAND2_X1 U15696 ( .A1(n14307), .A2(n13738), .ZN(n13551) );
  NAND2_X1 U15697 ( .A1(n13552), .A2(n13551), .ZN(n13556) );
  NAND2_X1 U15698 ( .A1(n13825), .A2(n13738), .ZN(n13553) );
  OAI21_X1 U15699 ( .B1(n13554), .B2(n13738), .A(n13553), .ZN(n13555) );
  INV_X1 U15700 ( .A(n13556), .ZN(n13557) );
  NAND2_X1 U15701 ( .A1(n13824), .A2(n13738), .ZN(n13559) );
  NAND2_X1 U15702 ( .A1(n6752), .A2(n13736), .ZN(n13558) );
  NAND2_X1 U15703 ( .A1(n13559), .A2(n13558), .ZN(n13561) );
  AOI22_X1 U15704 ( .A1(n13824), .A2(n13736), .B1(n6752), .B2(n13738), .ZN(
        n13560) );
  AOI21_X1 U15705 ( .B1(n13562), .B2(n13561), .A(n13560), .ZN(n13564) );
  NAND2_X1 U15706 ( .A1(n13823), .A2(n13736), .ZN(n13566) );
  NAND2_X1 U15707 ( .A1(n13567), .A2(n13738), .ZN(n13565) );
  NAND2_X1 U15708 ( .A1(n13566), .A2(n13565), .ZN(n13569) );
  AOI22_X1 U15709 ( .A1(n13823), .A2(n13738), .B1(n13567), .B2(n13736), .ZN(
        n13568) );
  NOR2_X1 U15710 ( .A1(n13570), .A2(n13569), .ZN(n13571) );
  NAND2_X1 U15711 ( .A1(n13822), .A2(n13738), .ZN(n13574) );
  NAND2_X1 U15712 ( .A1(n14301), .A2(n13736), .ZN(n13573) );
  NAND2_X1 U15713 ( .A1(n13574), .A2(n13573), .ZN(n13577) );
  NAND2_X1 U15714 ( .A1(n13822), .A2(n13736), .ZN(n13576) );
  NAND2_X1 U15715 ( .A1(n14301), .A2(n13738), .ZN(n13575) );
  NAND2_X1 U15716 ( .A1(n13581), .A2(n13738), .ZN(n13580) );
  NAND2_X1 U15717 ( .A1(n13821), .A2(n13736), .ZN(n13579) );
  AOI22_X1 U15718 ( .A1(n13581), .A2(n13736), .B1(n13738), .B2(n13821), .ZN(
        n13582) );
  NAND2_X1 U15719 ( .A1(n13585), .A2(n13736), .ZN(n13584) );
  NAND2_X1 U15720 ( .A1(n13820), .A2(n13738), .ZN(n13583) );
  NAND2_X1 U15721 ( .A1(n13584), .A2(n13583), .ZN(n13587) );
  AOI22_X1 U15722 ( .A1(n13585), .A2(n13738), .B1(n13820), .B2(n13736), .ZN(
        n13586) );
  NOR2_X1 U15723 ( .A1(n13588), .A2(n13587), .ZN(n13593) );
  AND2_X1 U15724 ( .A1(n14189), .A2(n13530), .ZN(n13589) );
  AOI21_X1 U15725 ( .B1(n13590), .B2(n13736), .A(n13589), .ZN(n13615) );
  NAND2_X1 U15726 ( .A1(n13590), .A2(n13738), .ZN(n13592) );
  NAND2_X1 U15727 ( .A1(n14189), .A2(n13736), .ZN(n13591) );
  NAND2_X1 U15728 ( .A1(n13592), .A2(n13591), .ZN(n13614) );
  AND2_X1 U15729 ( .A1(n13816), .A2(n13530), .ZN(n13595) );
  AOI21_X1 U15730 ( .B1(n14127), .B2(n13736), .A(n13595), .ZN(n13631) );
  NAND2_X1 U15731 ( .A1(n14127), .A2(n13738), .ZN(n13597) );
  NAND2_X1 U15732 ( .A1(n13816), .A2(n13736), .ZN(n13596) );
  NAND2_X1 U15733 ( .A1(n13597), .A2(n13596), .ZN(n13629) );
  NAND2_X1 U15734 ( .A1(n13631), .A2(n13629), .ZN(n13602) );
  AND2_X1 U15735 ( .A1(n13817), .A2(n13530), .ZN(n13598) );
  AOI21_X1 U15736 ( .B1(n14341), .B2(n13736), .A(n13598), .ZN(n13625) );
  NAND2_X1 U15737 ( .A1(n14341), .A2(n13738), .ZN(n13600) );
  NAND2_X1 U15738 ( .A1(n13817), .A2(n13736), .ZN(n13599) );
  NAND2_X1 U15739 ( .A1(n13600), .A2(n13599), .ZN(n13624) );
  NAND2_X1 U15740 ( .A1(n13625), .A2(n13624), .ZN(n13601) );
  NAND2_X1 U15741 ( .A1(n13602), .A2(n13601), .ZN(n13641) );
  AND2_X1 U15742 ( .A1(n13818), .A2(n13530), .ZN(n13603) );
  AOI21_X1 U15743 ( .B1(n14166), .B2(n13736), .A(n13603), .ZN(n13640) );
  NAND2_X1 U15744 ( .A1(n14166), .A2(n13738), .ZN(n13605) );
  NAND2_X1 U15745 ( .A1(n13818), .A2(n13736), .ZN(n13604) );
  NAND2_X1 U15746 ( .A1(n13605), .A2(n13604), .ZN(n13639) );
  AND2_X1 U15747 ( .A1(n13640), .A2(n13639), .ZN(n13606) );
  AND2_X1 U15748 ( .A1(n14191), .A2(n13530), .ZN(n13607) );
  AOI21_X1 U15749 ( .B1(n14184), .B2(n13736), .A(n13607), .ZN(n13637) );
  NAND2_X1 U15750 ( .A1(n14184), .A2(n13738), .ZN(n13609) );
  NAND2_X1 U15751 ( .A1(n14191), .A2(n13736), .ZN(n13608) );
  NAND2_X1 U15752 ( .A1(n13609), .A2(n13608), .ZN(n13636) );
  AND2_X1 U15753 ( .A1(n13637), .A2(n13636), .ZN(n13610) );
  NAND2_X1 U15754 ( .A1(n14296), .A2(n13738), .ZN(n13612) );
  NAND2_X1 U15755 ( .A1(n13819), .A2(n13736), .ZN(n13611) );
  NAND2_X1 U15756 ( .A1(n13612), .A2(n13611), .ZN(n13621) );
  INV_X1 U15757 ( .A(n13621), .ZN(n13619) );
  AND2_X1 U15758 ( .A1(n13819), .A2(n13530), .ZN(n13613) );
  AOI21_X1 U15759 ( .B1(n14296), .B2(n13736), .A(n13613), .ZN(n13622) );
  INV_X1 U15760 ( .A(n13622), .ZN(n13618) );
  INV_X1 U15761 ( .A(n13614), .ZN(n13617) );
  INV_X1 U15762 ( .A(n13615), .ZN(n13616) );
  OAI22_X1 U15763 ( .A1(n13619), .A2(n13618), .B1(n13617), .B2(n13616), .ZN(
        n13620) );
  INV_X1 U15764 ( .A(n13759), .ZN(n13628) );
  INV_X1 U15765 ( .A(n13624), .ZN(n13627) );
  INV_X1 U15766 ( .A(n13625), .ZN(n13626) );
  NAND2_X1 U15767 ( .A1(n13627), .A2(n13626), .ZN(n13630) );
  NAND2_X1 U15768 ( .A1(n13628), .A2(n13630), .ZN(n13635) );
  INV_X1 U15769 ( .A(n13629), .ZN(n13634) );
  INV_X1 U15770 ( .A(n13630), .ZN(n13633) );
  INV_X1 U15771 ( .A(n13631), .ZN(n13632) );
  AOI22_X1 U15772 ( .A1(n13635), .A2(n13634), .B1(n13633), .B2(n13632), .ZN(
        n13644) );
  OR3_X1 U15773 ( .A1(n13638), .A2(n13637), .A3(n13636), .ZN(n13643) );
  OR3_X1 U15774 ( .A1(n13641), .A2(n13640), .A3(n13639), .ZN(n13642) );
  NAND4_X1 U15775 ( .A1(n13645), .A2(n13644), .A3(n13643), .A4(n13642), .ZN(
        n13646) );
  NAND2_X1 U15776 ( .A1(n13648), .A2(n13738), .ZN(n13650) );
  NAND2_X1 U15777 ( .A1(n13815), .A2(n13736), .ZN(n13649) );
  OAI22_X1 U15778 ( .A1(n14262), .A2(n13738), .B1(n13651), .B2(n13736), .ZN(
        n13652) );
  OAI22_X1 U15779 ( .A1(n14256), .A2(n13738), .B1(n13653), .B2(n13736), .ZN(
        n13656) );
  INV_X1 U15780 ( .A(n13656), .ZN(n13655) );
  OAI22_X1 U15781 ( .A1(n14256), .A2(n13736), .B1(n13653), .B2(n13738), .ZN(
        n13654) );
  OAI22_X1 U15782 ( .A1(n14335), .A2(n13738), .B1(n13659), .B2(n13736), .ZN(
        n13660) );
  INV_X1 U15783 ( .A(n13664), .ZN(n13665) );
  AOI22_X1 U15784 ( .A1(n14073), .A2(n13738), .B1(n13812), .B2(n13736), .ZN(
        n13662) );
  AOI22_X1 U15785 ( .A1(n14059), .A2(n13738), .B1(n14039), .B2(n13736), .ZN(
        n13667) );
  AOI22_X1 U15786 ( .A1(n14059), .A2(n13736), .B1(n13530), .B2(n14039), .ZN(
        n13669) );
  OAI22_X1 U15787 ( .A1(n14227), .A2(n13738), .B1(n13754), .B2(n13736), .ZN(
        n13682) );
  AOI22_X1 U15788 ( .A1(n14047), .A2(n13738), .B1(n14024), .B2(n13736), .ZN(
        n13670) );
  AND2_X1 U15789 ( .A1(n14041), .A2(n13736), .ZN(n13671) );
  AOI21_X1 U15790 ( .B1(n14217), .B2(n13738), .A(n13671), .ZN(n13687) );
  NAND2_X1 U15791 ( .A1(n14217), .A2(n13736), .ZN(n13673) );
  NAND2_X1 U15792 ( .A1(n14041), .A2(n13738), .ZN(n13672) );
  NAND2_X1 U15793 ( .A1(n13673), .A2(n13672), .ZN(n13686) );
  AND2_X1 U15794 ( .A1(n14004), .A2(n13530), .ZN(n13674) );
  AOI21_X1 U15795 ( .B1(n14210), .B2(n13736), .A(n13674), .ZN(n13698) );
  NAND2_X1 U15796 ( .A1(n14210), .A2(n13738), .ZN(n13676) );
  NAND2_X1 U15797 ( .A1(n14004), .A2(n13736), .ZN(n13675) );
  NAND2_X1 U15798 ( .A1(n13676), .A2(n13675), .ZN(n13697) );
  NAND2_X1 U15799 ( .A1(n13698), .A2(n13697), .ZN(n13702) );
  AND2_X1 U15800 ( .A1(n14026), .A2(n13530), .ZN(n13677) );
  AOI21_X1 U15801 ( .B1(n14008), .B2(n13736), .A(n13677), .ZN(n13694) );
  NAND2_X1 U15802 ( .A1(n14008), .A2(n13738), .ZN(n13679) );
  NAND2_X1 U15803 ( .A1(n14026), .A2(n13736), .ZN(n13678) );
  NAND2_X1 U15804 ( .A1(n13679), .A2(n13678), .ZN(n13693) );
  NAND2_X1 U15805 ( .A1(n13694), .A2(n13693), .ZN(n13680) );
  AND2_X1 U15806 ( .A1(n13702), .A2(n13680), .ZN(n13685) );
  OAI21_X1 U15807 ( .B1(n13687), .B2(n13686), .A(n13685), .ZN(n13681) );
  INV_X1 U15808 ( .A(n13681), .ZN(n13684) );
  INV_X1 U15809 ( .A(n13682), .ZN(n13683) );
  INV_X1 U15810 ( .A(n13685), .ZN(n13706) );
  NAND2_X1 U15811 ( .A1(n13687), .A2(n13686), .ZN(n13705) );
  NAND2_X1 U15812 ( .A1(n13974), .A2(n13738), .ZN(n13689) );
  NAND2_X1 U15813 ( .A1(n13811), .A2(n13736), .ZN(n13688) );
  NAND2_X1 U15814 ( .A1(n13689), .A2(n13688), .ZN(n13721) );
  INV_X1 U15815 ( .A(n13721), .ZN(n13692) );
  AND2_X1 U15816 ( .A1(n13811), .A2(n13530), .ZN(n13690) );
  AOI21_X1 U15817 ( .B1(n13974), .B2(n13736), .A(n13690), .ZN(n13722) );
  INV_X1 U15818 ( .A(n13722), .ZN(n13691) );
  NAND2_X1 U15819 ( .A1(n13692), .A2(n13691), .ZN(n13704) );
  INV_X1 U15820 ( .A(n13693), .ZN(n13696) );
  INV_X1 U15821 ( .A(n13694), .ZN(n13695) );
  AND2_X1 U15822 ( .A1(n13696), .A2(n13695), .ZN(n13701) );
  INV_X1 U15823 ( .A(n13697), .ZN(n13700) );
  INV_X1 U15824 ( .A(n13698), .ZN(n13699) );
  AOI22_X1 U15825 ( .A1(n13702), .A2(n13701), .B1(n13700), .B2(n13699), .ZN(
        n13703) );
  OAI211_X1 U15826 ( .C1(n13706), .C2(n13705), .A(n13704), .B(n13703), .ZN(
        n13707) );
  INV_X1 U15827 ( .A(n13707), .ZN(n13708) );
  INV_X1 U15828 ( .A(n13808), .ZN(n13710) );
  OAI22_X1 U15829 ( .A1(n14314), .A2(n13738), .B1(n13710), .B2(n13736), .ZN(
        n13733) );
  NAND2_X1 U15830 ( .A1(n13807), .A2(n13736), .ZN(n13737) );
  NOR2_X1 U15831 ( .A1(n13748), .A2(n13761), .ZN(n13712) );
  NOR2_X1 U15832 ( .A1(n13712), .A2(n13711), .ZN(n13713) );
  NAND2_X1 U15833 ( .A1(n13737), .A2(n13713), .ZN(n13714) );
  AND2_X1 U15834 ( .A1(n13809), .A2(n13736), .ZN(n13715) );
  AOI21_X1 U15835 ( .B1(n13955), .B2(n13738), .A(n13715), .ZN(n13725) );
  NAND2_X1 U15836 ( .A1(n13955), .A2(n13736), .ZN(n13717) );
  NAND2_X1 U15837 ( .A1(n13809), .A2(n13738), .ZN(n13716) );
  NAND2_X1 U15838 ( .A1(n13717), .A2(n13716), .ZN(n13724) );
  XNOR2_X1 U15839 ( .A(n13718), .B(n13807), .ZN(n13790) );
  OAI22_X1 U15840 ( .A1(n13966), .A2(n13736), .B1(n13719), .B2(n13738), .ZN(
        n13727) );
  AOI22_X1 U15841 ( .A1(n13720), .A2(n13736), .B1(n13530), .B2(n13810), .ZN(
        n13726) );
  AOI22_X1 U15842 ( .A1(n13727), .A2(n13726), .B1(n13722), .B2(n13721), .ZN(
        n13723) );
  INV_X1 U15843 ( .A(n13724), .ZN(n13729) );
  INV_X1 U15844 ( .A(n13725), .ZN(n13728) );
  NAND2_X1 U15845 ( .A1(n13737), .A2(n13736), .ZN(n13740) );
  NAND2_X1 U15846 ( .A1(n13807), .A2(n13738), .ZN(n13739) );
  MUX2_X1 U15847 ( .A(n13740), .B(n13739), .S(n13943), .Z(n13741) );
  INV_X1 U15848 ( .A(n13742), .ZN(n13746) );
  OAI21_X1 U15849 ( .B1(n13936), .B2(n13744), .A(n13743), .ZN(n13745) );
  AOI21_X1 U15850 ( .B1(n13746), .B2(n8559), .A(n13745), .ZN(n13747) );
  INV_X1 U15851 ( .A(n13747), .ZN(n13752) );
  INV_X1 U15852 ( .A(n13748), .ZN(n13749) );
  OAI211_X1 U15853 ( .C1(n13749), .C2(n13761), .A(n8610), .B(n13936), .ZN(
        n13750) );
  XNOR2_X1 U15854 ( .A(n13946), .B(n13808), .ZN(n13788) );
  INV_X1 U15855 ( .A(n14000), .ZN(n13783) );
  XNOR2_X1 U15856 ( .A(n14047), .B(n13754), .ZN(n14036) );
  INV_X1 U15857 ( .A(n13755), .ZN(n13756) );
  OR2_X1 U15858 ( .A1(n13757), .A2(n13756), .ZN(n14066) );
  NAND2_X1 U15859 ( .A1(n13759), .A2(n13758), .ZN(n14132) );
  XNOR2_X1 U15860 ( .A(n14184), .B(n14160), .ZN(n14176) );
  NAND4_X1 U15861 ( .A1(n8563), .A2(n13761), .A3(n13760), .A4(n15519), .ZN(
        n13764) );
  XNOR2_X1 U15862 ( .A(n15544), .B(n13762), .ZN(n15486) );
  NOR3_X1 U15863 ( .A1(n13764), .A2(n13763), .A3(n15486), .ZN(n13767) );
  XNOR2_X1 U15864 ( .A(n13826), .B(n15826), .ZN(n15553) );
  NAND4_X1 U15865 ( .A1(n13767), .A2(n13766), .A3(n13765), .A4(n15553), .ZN(
        n13770) );
  NAND2_X1 U15866 ( .A1(n8571), .A2(n13768), .ZN(n13769) );
  NOR2_X1 U15867 ( .A1(n13770), .A2(n13769), .ZN(n13774) );
  NAND4_X1 U15868 ( .A1(n13774), .A2(n13773), .A3(n13772), .A4(n13771), .ZN(
        n13776) );
  XNOR2_X1 U15869 ( .A(n14296), .B(n13775), .ZN(n14198) );
  OR3_X1 U15870 ( .A1(n14176), .A2(n13776), .A3(n14198), .ZN(n13777) );
  NOR2_X1 U15871 ( .A1(n14152), .A2(n13777), .ZN(n13778) );
  XNOR2_X1 U15872 ( .A(n14166), .B(n13818), .ZN(n14150) );
  NAND3_X1 U15873 ( .A1(n14132), .A2(n13778), .A3(n14150), .ZN(n13779) );
  NOR2_X1 U15874 ( .A1(n14111), .A2(n13779), .ZN(n13780) );
  XNOR2_X1 U15875 ( .A(n14105), .B(n13814), .ZN(n14097) );
  NAND4_X1 U15876 ( .A1(n14066), .A2(n13780), .A3(n14077), .A4(n14097), .ZN(
        n13781) );
  NOR4_X1 U15877 ( .A1(n14020), .A2(n14036), .A3(n14052), .A4(n13781), .ZN(
        n13782) );
  NAND3_X1 U15878 ( .A1(n7500), .A2(n13783), .A3(n13782), .ZN(n13784) );
  NOR3_X1 U15879 ( .A1(n13786), .A2(n13785), .A3(n13784), .ZN(n13787) );
  NAND4_X1 U15880 ( .A1(n13790), .A2(n13789), .A3(n13788), .A4(n13787), .ZN(
        n13801) );
  NOR2_X1 U15881 ( .A1(n8610), .A2(n13805), .ZN(n13792) );
  NAND2_X1 U15882 ( .A1(n13792), .A2(n13791), .ZN(n13800) );
  NAND2_X1 U15883 ( .A1(n14188), .A2(n13793), .ZN(n13797) );
  INV_X1 U15884 ( .A(n13805), .ZN(n13795) );
  AOI21_X1 U15885 ( .B1(n8559), .B2(n13795), .A(n13794), .ZN(n13796) );
  OAI21_X1 U15886 ( .B1(n13798), .B2(n13797), .A(n13796), .ZN(n13799) );
  OAI21_X1 U15887 ( .B1(n13801), .B2(n13800), .A(n13799), .ZN(n13802) );
  OAI21_X1 U15888 ( .B1(n13806), .B2(n13805), .A(n13804), .ZN(P2_U3328) );
  MUX2_X1 U15889 ( .A(n13807), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13830), .Z(
        P2_U3562) );
  MUX2_X1 U15890 ( .A(n13808), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13830), .Z(
        P2_U3561) );
  MUX2_X1 U15891 ( .A(n13809), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13830), .Z(
        P2_U3560) );
  MUX2_X1 U15892 ( .A(n13810), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13830), .Z(
        P2_U3559) );
  MUX2_X1 U15893 ( .A(n13811), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13830), .Z(
        P2_U3558) );
  MUX2_X1 U15894 ( .A(n14004), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13830), .Z(
        P2_U3557) );
  MUX2_X1 U15895 ( .A(n14026), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13830), .Z(
        P2_U3556) );
  MUX2_X1 U15896 ( .A(n14041), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13830), .Z(
        P2_U3555) );
  MUX2_X1 U15897 ( .A(n14024), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13830), .Z(
        P2_U3554) );
  MUX2_X1 U15898 ( .A(n14039), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13830), .Z(
        P2_U3553) );
  MUX2_X1 U15899 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13812), .S(P2_U3947), .Z(
        P2_U3552) );
  MUX2_X1 U15900 ( .A(n13813), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13830), .Z(
        P2_U3551) );
  MUX2_X1 U15901 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13814), .S(P2_U3947), .Z(
        P2_U3550) );
  MUX2_X1 U15902 ( .A(n13815), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13830), .Z(
        P2_U3549) );
  MUX2_X1 U15903 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13816), .S(P2_U3947), .Z(
        P2_U3548) );
  MUX2_X1 U15904 ( .A(n13817), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13830), .Z(
        P2_U3547) );
  MUX2_X1 U15905 ( .A(n13818), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13830), .Z(
        P2_U3546) );
  MUX2_X1 U15906 ( .A(n14191), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13830), .Z(
        P2_U3545) );
  MUX2_X1 U15907 ( .A(n13819), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13830), .Z(
        P2_U3544) );
  MUX2_X1 U15908 ( .A(n14189), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13830), .Z(
        P2_U3543) );
  MUX2_X1 U15909 ( .A(n13820), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13830), .Z(
        P2_U3542) );
  MUX2_X1 U15910 ( .A(n13821), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13830), .Z(
        P2_U3541) );
  MUX2_X1 U15911 ( .A(n13822), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13830), .Z(
        P2_U3540) );
  MUX2_X1 U15912 ( .A(n13823), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13830), .Z(
        P2_U3539) );
  MUX2_X1 U15913 ( .A(n13824), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13830), .Z(
        P2_U3538) );
  MUX2_X1 U15914 ( .A(n13825), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13830), .Z(
        P2_U3537) );
  MUX2_X1 U15915 ( .A(n13826), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13830), .Z(
        P2_U3536) );
  MUX2_X1 U15916 ( .A(n13827), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13830), .Z(
        P2_U3535) );
  MUX2_X1 U15917 ( .A(n13828), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13830), .Z(
        P2_U3534) );
  MUX2_X1 U15918 ( .A(n13829), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13830), .Z(
        P2_U3533) );
  MUX2_X1 U15919 ( .A(n13508), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13830), .Z(
        P2_U3532) );
  MUX2_X1 U15920 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6966), .S(n13838), .Z(
        n13831) );
  OAI21_X1 U15921 ( .B1(n8127), .B2(n13832), .A(n13831), .ZN(n13833) );
  NAND3_X1 U15922 ( .A1(n15470), .A2(n13834), .A3(n13833), .ZN(n13843) );
  AOI22_X1 U15923 ( .A1(n15468), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n13842) );
  AND2_X1 U15924 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n13837) );
  OAI211_X1 U15925 ( .C1(n13837), .C2(n13836), .A(n15475), .B(n13835), .ZN(
        n13841) );
  INV_X1 U15926 ( .A(n13838), .ZN(n13839) );
  NAND2_X1 U15927 ( .A1(n15447), .A2(n13839), .ZN(n13840) );
  NAND4_X1 U15928 ( .A1(n13843), .A2(n13842), .A3(n13841), .A4(n13840), .ZN(
        P2_U3215) );
  MUX2_X1 U15929 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10584), .S(n13851), .Z(
        n13844) );
  INV_X1 U15930 ( .A(n13844), .ZN(n13847) );
  OAI211_X1 U15931 ( .C1(n13847), .C2(n13846), .A(n15470), .B(n13845), .ZN(
        n13856) );
  AOI22_X1 U15932 ( .A1(n15468), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n13855) );
  OAI211_X1 U15933 ( .C1(n13850), .C2(n13849), .A(n15475), .B(n13848), .ZN(
        n13854) );
  INV_X1 U15934 ( .A(n13851), .ZN(n13852) );
  NAND2_X1 U15935 ( .A1(n15447), .A2(n13852), .ZN(n13853) );
  NAND4_X1 U15936 ( .A1(n13856), .A2(n13855), .A3(n13854), .A4(n13853), .ZN(
        P2_U3216) );
  INV_X1 U15937 ( .A(n13861), .ZN(n13860) );
  OAI21_X1 U15938 ( .B1(n13938), .B2(n13858), .A(n13857), .ZN(n13859) );
  AOI21_X1 U15939 ( .B1(n13860), .B2(n15447), .A(n13859), .ZN(n13873) );
  MUX2_X1 U15940 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10589), .S(n13861), .Z(
        n13862) );
  NAND3_X1 U15941 ( .A1(n15454), .A2(n13863), .A3(n13862), .ZN(n13864) );
  NAND3_X1 U15942 ( .A1(n15470), .A2(n13865), .A3(n13864), .ZN(n13872) );
  INV_X1 U15943 ( .A(n13866), .ZN(n13870) );
  NAND3_X1 U15944 ( .A1(n15457), .A2(n13868), .A3(n13867), .ZN(n13869) );
  NAND3_X1 U15945 ( .A1(n15475), .A2(n13870), .A3(n13869), .ZN(n13871) );
  NAND3_X1 U15946 ( .A1(n13873), .A2(n13872), .A3(n13871), .ZN(P2_U3218) );
  INV_X1 U15947 ( .A(n13874), .ZN(n13890) );
  OR2_X1 U15948 ( .A1(n13885), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n13875) );
  NAND2_X1 U15949 ( .A1(n13885), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n13899) );
  AND2_X1 U15950 ( .A1(n13875), .A2(n13899), .ZN(n13882) );
  NAND2_X1 U15951 ( .A1(n13876), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n13880) );
  INV_X1 U15952 ( .A(n13877), .ZN(n13878) );
  NAND2_X1 U15953 ( .A1(n13878), .A2(n13884), .ZN(n13879) );
  NAND2_X1 U15954 ( .A1(n13880), .A2(n13879), .ZN(n13881) );
  NAND2_X1 U15955 ( .A1(n13881), .A2(n13882), .ZN(n13900) );
  OAI211_X1 U15956 ( .C1(n13882), .C2(n13881), .A(n15470), .B(n13900), .ZN(
        n13888) );
  XNOR2_X1 U15957 ( .A(n13885), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n13894) );
  XOR2_X1 U15958 ( .A(n13895), .B(n13894), .Z(n13886) );
  NAND2_X1 U15959 ( .A1(n15475), .A2(n13886), .ZN(n13887) );
  NAND2_X1 U15960 ( .A1(n13888), .A2(n13887), .ZN(n13889) );
  AOI211_X1 U15961 ( .C1(n15468), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n13890), 
        .B(n13889), .ZN(n13891) );
  OAI21_X1 U15962 ( .B1(n15465), .B2(n13893), .A(n13891), .ZN(P2_U3230) );
  XOR2_X1 U15963 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13915), .Z(n13916) );
  INV_X1 U15964 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n13892) );
  XOR2_X1 U15965 ( .A(n13916), .B(n13917), .Z(n13896) );
  NAND2_X1 U15966 ( .A1(n13896), .A2(n15475), .ZN(n13907) );
  INV_X1 U15967 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13897) );
  NAND2_X1 U15968 ( .A1(n13908), .A2(n13897), .ZN(n13898) );
  NAND2_X1 U15969 ( .A1(n13915), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13909) );
  AND2_X1 U15970 ( .A1(n13898), .A2(n13909), .ZN(n13902) );
  NAND2_X1 U15971 ( .A1(n13900), .A2(n13899), .ZN(n13901) );
  OAI211_X1 U15972 ( .C1(n13902), .C2(n13901), .A(n15470), .B(n13910), .ZN(
        n13903) );
  NAND2_X1 U15973 ( .A1(n13904), .A2(n13903), .ZN(n13905) );
  AOI21_X1 U15974 ( .B1(n15468), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n13905), 
        .ZN(n13906) );
  OAI211_X1 U15975 ( .C1(n15465), .C2(n13908), .A(n13907), .B(n13906), .ZN(
        P2_U3231) );
  NAND2_X1 U15976 ( .A1(n13911), .A2(n13927), .ZN(n13912) );
  INV_X1 U15977 ( .A(n13932), .ZN(n13913) );
  AOI21_X1 U15978 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n13914), .A(n13913), 
        .ZN(n13924) );
  AOI22_X1 U15979 ( .A1(n13917), .A2(n13916), .B1(n13915), .B2(
        P2_REG1_REG_17__SCAN_IN), .ZN(n13925) );
  XOR2_X1 U15980 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13928), .Z(n13922) );
  NAND2_X1 U15981 ( .A1(n15468), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n13918) );
  OAI211_X1 U15982 ( .C1(n15465), .C2(n13920), .A(n13919), .B(n13918), .ZN(
        n13921) );
  AOI21_X1 U15983 ( .B1(n13922), .B2(n15475), .A(n13921), .ZN(n13923) );
  OAI21_X1 U15984 ( .B1(n13924), .B2(n15444), .A(n13923), .ZN(P2_U3232) );
  INV_X1 U15985 ( .A(n13925), .ZN(n13926) );
  XNOR2_X1 U15986 ( .A(n13930), .B(n13929), .ZN(n13935) );
  NAND2_X1 U15987 ( .A1(n13932), .A2(n13931), .ZN(n13933) );
  NAND2_X1 U15988 ( .A1(n13939), .A2(n15484), .ZN(n13942) );
  INV_X1 U15989 ( .A(n14204), .ZN(n13940) );
  NOR2_X1 U15990 ( .A1(n14180), .A2(n13940), .ZN(n13947) );
  AOI21_X1 U15991 ( .B1(n14180), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13947), 
        .ZN(n13941) );
  OAI211_X1 U15992 ( .C1(n13943), .C2(n15504), .A(n13942), .B(n13941), .ZN(
        P2_U3234) );
  NAND2_X1 U15993 ( .A1(n14205), .A2(n15484), .ZN(n13949) );
  AOI21_X1 U15994 ( .B1(n14180), .B2(P2_REG2_REG_30__SCAN_IN), .A(n13947), 
        .ZN(n13948) );
  OAI211_X1 U15995 ( .C1(n14314), .C2(n15504), .A(n13949), .B(n13948), .ZN(
        P2_U3235) );
  NAND2_X1 U15996 ( .A1(n13951), .A2(n13950), .ZN(n13953) );
  XNOR2_X1 U15997 ( .A(n13953), .B(n13952), .ZN(n13963) );
  NAND2_X1 U15998 ( .A1(n13954), .A2(n15831), .ZN(n13962) );
  NAND2_X1 U15999 ( .A1(n13955), .A2(n15827), .ZN(n13957) );
  NAND2_X1 U16000 ( .A1(n14180), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n13956) );
  OAI211_X1 U16001 ( .C1(n15503), .C2(n13958), .A(n13957), .B(n13956), .ZN(
        n13959) );
  AOI21_X1 U16002 ( .B1(n13960), .B2(n15484), .A(n13959), .ZN(n13961) );
  OAI211_X1 U16003 ( .C1(n13963), .C2(n14200), .A(n13962), .B(n13961), .ZN(
        P2_U3236) );
  AOI22_X1 U16004 ( .A1(n13964), .A2(n15825), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n14180), .ZN(n13965) );
  OAI21_X1 U16005 ( .B1(n13966), .B2(n15504), .A(n13965), .ZN(n13967) );
  AOI21_X1 U16006 ( .B1(n13968), .B2(n15484), .A(n13967), .ZN(n13971) );
  NAND2_X1 U16007 ( .A1(n13969), .A2(n14134), .ZN(n13970) );
  OAI211_X1 U16008 ( .C1(n6491), .C2(n14180), .A(n13971), .B(n13970), .ZN(
        P2_U3237) );
  INV_X1 U16009 ( .A(n13972), .ZN(n13979) );
  AOI22_X1 U16010 ( .A1(n13973), .A2(n15825), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n14180), .ZN(n13976) );
  NAND2_X1 U16011 ( .A1(n13974), .A2(n15827), .ZN(n13975) );
  OAI211_X1 U16012 ( .C1(n13977), .C2(n15829), .A(n13976), .B(n13975), .ZN(
        n13978) );
  AOI21_X1 U16013 ( .B1(n13979), .B2(n15831), .A(n13978), .ZN(n13980) );
  OAI21_X1 U16014 ( .B1(n13981), .B2(n14200), .A(n13980), .ZN(P2_U3238) );
  XNOR2_X1 U16015 ( .A(n13982), .B(n7500), .ZN(n14211) );
  INV_X1 U16016 ( .A(n14011), .ZN(n13987) );
  NAND2_X1 U16017 ( .A1(n13987), .A2(n14210), .ZN(n13989) );
  NAND2_X1 U16018 ( .A1(n14209), .A2(n15484), .ZN(n13992) );
  AOI22_X1 U16019 ( .A1(n13990), .A2(n15825), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14180), .ZN(n13991) );
  OAI211_X1 U16020 ( .C1(n13993), .C2(n15504), .A(n13992), .B(n13991), .ZN(
        n13994) );
  AOI21_X1 U16021 ( .B1(n14208), .B2(n15831), .A(n13994), .ZN(n13995) );
  OAI21_X1 U16022 ( .B1(n14211), .B2(n14200), .A(n13995), .ZN(P2_U3239) );
  XNOR2_X1 U16023 ( .A(n13996), .B(n14000), .ZN(n14212) );
  INV_X1 U16024 ( .A(n14212), .ZN(n14017) );
  NAND2_X1 U16025 ( .A1(n13998), .A2(n13997), .ZN(n14019) );
  NAND3_X1 U16026 ( .A1(n14021), .A2(n14000), .A3(n13999), .ZN(n14002) );
  NAND2_X1 U16027 ( .A1(n14002), .A2(n14001), .ZN(n14003) );
  NAND2_X1 U16028 ( .A1(n14003), .A2(n15556), .ZN(n14006) );
  AOI22_X1 U16029 ( .A1(n14004), .A2(n14190), .B1(n14188), .B2(n14041), .ZN(
        n14005) );
  NAND2_X1 U16030 ( .A1(n14006), .A2(n14005), .ZN(n14214) );
  NAND2_X1 U16031 ( .A1(n14007), .A2(n14008), .ZN(n14009) );
  NAND2_X1 U16032 ( .A1(n14009), .A2(n14181), .ZN(n14010) );
  NOR2_X1 U16033 ( .A1(n14011), .A2(n14010), .ZN(n14213) );
  NAND2_X1 U16034 ( .A1(n14213), .A2(n15484), .ZN(n14014) );
  AOI22_X1 U16035 ( .A1(n14012), .A2(n15825), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n14180), .ZN(n14013) );
  OAI211_X1 U16036 ( .C1(n14321), .C2(n15504), .A(n14014), .B(n14013), .ZN(
        n14015) );
  AOI21_X1 U16037 ( .B1(n14214), .B2(n15831), .A(n14015), .ZN(n14016) );
  OAI21_X1 U16038 ( .B1(n14200), .B2(n14017), .A(n14016), .ZN(P2_U3240) );
  XNOR2_X1 U16039 ( .A(n14018), .B(n14020), .ZN(n14224) );
  INV_X1 U16040 ( .A(n14019), .ZN(n14022) );
  OAI21_X1 U16041 ( .B1(n14022), .B2(n6743), .A(n14021), .ZN(n14222) );
  AOI21_X1 U16042 ( .B1(n14038), .B2(n14217), .A(n15561), .ZN(n14023) );
  NAND2_X1 U16043 ( .A1(n14023), .A2(n14007), .ZN(n14219) );
  AND2_X1 U16044 ( .A1(n14024), .A2(n14188), .ZN(n14025) );
  AOI21_X1 U16045 ( .B1(n14026), .B2(n14190), .A(n14025), .ZN(n14218) );
  INV_X1 U16046 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n14027) );
  OAI22_X1 U16047 ( .A1(n14028), .A2(n15503), .B1(n14027), .B2(n15831), .ZN(
        n14029) );
  INV_X1 U16048 ( .A(n14029), .ZN(n14030) );
  OAI21_X1 U16049 ( .B1(n14218), .B2(n14180), .A(n14030), .ZN(n14031) );
  AOI21_X1 U16050 ( .B1(n14217), .B2(n15827), .A(n14031), .ZN(n14032) );
  OAI21_X1 U16051 ( .B1(n14219), .B2(n15829), .A(n14032), .ZN(n14033) );
  AOI21_X1 U16052 ( .B1(n14222), .B2(n14177), .A(n14033), .ZN(n14034) );
  OAI21_X1 U16053 ( .B1(n14200), .B2(n14224), .A(n14034), .ZN(P2_U3241) );
  XNOR2_X1 U16054 ( .A(n14035), .B(n14036), .ZN(n14231) );
  XNOR2_X1 U16055 ( .A(n14037), .B(n14036), .ZN(n14229) );
  OAI211_X1 U16056 ( .C1(n14058), .C2(n14227), .A(n14038), .B(n14181), .ZN(
        n14226) );
  AND2_X1 U16057 ( .A1(n14039), .A2(n14188), .ZN(n14040) );
  AOI21_X1 U16058 ( .B1(n14041), .B2(n14190), .A(n14040), .ZN(n14225) );
  INV_X1 U16059 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n14042) );
  OAI22_X1 U16060 ( .A1(n14043), .A2(n15503), .B1(n14042), .B2(n15831), .ZN(
        n14044) );
  INV_X1 U16061 ( .A(n14044), .ZN(n14045) );
  OAI21_X1 U16062 ( .B1(n14225), .B2(n14180), .A(n14045), .ZN(n14046) );
  AOI21_X1 U16063 ( .B1(n14047), .B2(n15827), .A(n14046), .ZN(n14048) );
  OAI21_X1 U16064 ( .B1(n14226), .B2(n15829), .A(n14048), .ZN(n14049) );
  AOI21_X1 U16065 ( .B1(n14229), .B2(n14177), .A(n14049), .ZN(n14050) );
  OAI21_X1 U16066 ( .B1(n14231), .B2(n14200), .A(n14050), .ZN(P2_U3242) );
  OAI21_X1 U16067 ( .B1(n14053), .B2(n14052), .A(n14051), .ZN(n14232) );
  OAI211_X1 U16068 ( .C1(n6466), .C2(n14055), .A(n14054), .B(n15556), .ZN(
        n14057) );
  NAND2_X1 U16069 ( .A1(n14057), .A2(n14056), .ZN(n14233) );
  NAND2_X1 U16070 ( .A1(n14233), .A2(n15831), .ZN(n14064) );
  AOI211_X1 U16071 ( .C1(n14059), .C2(n14068), .A(n15561), .B(n14058), .ZN(
        n14234) );
  AOI22_X1 U16072 ( .A1(n14060), .A2(n15825), .B1(P2_REG2_REG_22__SCAN_IN), 
        .B2(n14180), .ZN(n14061) );
  OAI21_X1 U16073 ( .B1(n14327), .B2(n15504), .A(n14061), .ZN(n14062) );
  AOI21_X1 U16074 ( .B1(n14234), .B2(n15484), .A(n14062), .ZN(n14063) );
  OAI211_X1 U16075 ( .C1(n14232), .C2(n14200), .A(n14064), .B(n14063), .ZN(
        P2_U3243) );
  XNOR2_X1 U16076 ( .A(n14065), .B(n14066), .ZN(n14243) );
  XNOR2_X1 U16077 ( .A(n14067), .B(n14066), .ZN(n14238) );
  AOI21_X1 U16078 ( .B1(n14085), .B2(n14073), .A(n15561), .ZN(n14069) );
  NAND2_X1 U16079 ( .A1(n14069), .A2(n14068), .ZN(n14240) );
  AOI22_X1 U16080 ( .A1(n14070), .A2(n15825), .B1(P2_REG2_REG_21__SCAN_IN), 
        .B2(n14180), .ZN(n14071) );
  OAI21_X1 U16081 ( .B1(n14239), .B2(n14180), .A(n14071), .ZN(n14072) );
  AOI21_X1 U16082 ( .B1(n14073), .B2(n15827), .A(n14072), .ZN(n14074) );
  OAI21_X1 U16083 ( .B1(n14240), .B2(n15829), .A(n14074), .ZN(n14075) );
  AOI21_X1 U16084 ( .B1(n14238), .B2(n14177), .A(n14075), .ZN(n14076) );
  OAI21_X1 U16085 ( .B1(n14200), .B2(n14243), .A(n14076), .ZN(P2_U3244) );
  NAND2_X1 U16086 ( .A1(n14078), .A2(n14077), .ZN(n14079) );
  NAND2_X1 U16087 ( .A1(n14082), .A2(n14081), .ZN(n14083) );
  NAND2_X1 U16088 ( .A1(n14084), .A2(n14083), .ZN(n14246) );
  AOI21_X1 U16089 ( .B1(n14100), .B2(n14092), .A(n15561), .ZN(n14086) );
  NAND2_X1 U16090 ( .A1(n14086), .A2(n14085), .ZN(n14248) );
  INV_X1 U16091 ( .A(n14087), .ZN(n14247) );
  INV_X1 U16092 ( .A(n14088), .ZN(n14089) );
  AOI22_X1 U16093 ( .A1(n14089), .A2(n15825), .B1(P2_REG2_REG_20__SCAN_IN), 
        .B2(n14180), .ZN(n14090) );
  OAI21_X1 U16094 ( .B1(n14247), .B2(n14180), .A(n14090), .ZN(n14091) );
  AOI21_X1 U16095 ( .B1(n14092), .B2(n15827), .A(n14091), .ZN(n14093) );
  OAI21_X1 U16096 ( .B1(n14248), .B2(n15829), .A(n14093), .ZN(n14094) );
  AOI21_X1 U16097 ( .B1(n14246), .B2(n14177), .A(n14094), .ZN(n14095) );
  OAI21_X1 U16098 ( .B1(n14251), .B2(n14200), .A(n14095), .ZN(P2_U3245) );
  XNOR2_X1 U16099 ( .A(n14096), .B(n14097), .ZN(n14260) );
  XNOR2_X1 U16100 ( .A(n14098), .B(n14097), .ZN(n14258) );
  OAI211_X1 U16101 ( .C1(n14099), .C2(n14256), .A(n14181), .B(n14100), .ZN(
        n14255) );
  INV_X1 U16102 ( .A(n14254), .ZN(n14104) );
  INV_X1 U16103 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n14101) );
  OAI22_X1 U16104 ( .A1(n14102), .A2(n15503), .B1(n14101), .B2(n15831), .ZN(
        n14103) );
  AOI21_X1 U16105 ( .B1(n14104), .B2(n15831), .A(n14103), .ZN(n14107) );
  NAND2_X1 U16106 ( .A1(n14105), .A2(n15827), .ZN(n14106) );
  OAI211_X1 U16107 ( .C1(n14255), .C2(n15829), .A(n14107), .B(n14106), .ZN(
        n14108) );
  AOI21_X1 U16108 ( .B1(n14258), .B2(n14177), .A(n14108), .ZN(n14109) );
  OAI21_X1 U16109 ( .B1(n14200), .B2(n14260), .A(n14109), .ZN(P2_U3246) );
  XOR2_X1 U16110 ( .A(n14110), .B(n14111), .Z(n14267) );
  XNOR2_X1 U16111 ( .A(n14112), .B(n14111), .ZN(n14265) );
  OAI21_X1 U16112 ( .B1(n14126), .B2(n14262), .A(n14181), .ZN(n14113) );
  NOR2_X1 U16113 ( .A1(n14113), .A2(n14099), .ZN(n14264) );
  NAND2_X1 U16114 ( .A1(n14264), .A2(n15484), .ZN(n14119) );
  INV_X1 U16115 ( .A(n14261), .ZN(n14117) );
  INV_X1 U16116 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n14114) );
  OAI22_X1 U16117 ( .A1(n14115), .A2(n15503), .B1(n15831), .B2(n14114), .ZN(
        n14116) );
  AOI21_X1 U16118 ( .B1(n14117), .B2(n15831), .A(n14116), .ZN(n14118) );
  OAI211_X1 U16119 ( .C1(n14262), .C2(n15504), .A(n14119), .B(n14118), .ZN(
        n14120) );
  AOI21_X1 U16120 ( .B1(n14265), .B2(n14177), .A(n14120), .ZN(n14121) );
  OAI21_X1 U16121 ( .B1(n14267), .B2(n14200), .A(n14121), .ZN(P2_U3247) );
  NAND2_X1 U16122 ( .A1(n14123), .A2(n14122), .ZN(n14138) );
  NAND2_X1 U16123 ( .A1(n14140), .A2(n14124), .ZN(n14125) );
  XNOR2_X1 U16124 ( .A(n14125), .B(n14132), .ZN(n14275) );
  INV_X1 U16125 ( .A(n14177), .ZN(n14137) );
  AOI211_X1 U16126 ( .C1(n14127), .C2(n14146), .A(n15561), .B(n14126), .ZN(
        n14269) );
  NAND2_X1 U16127 ( .A1(n14127), .A2(n15827), .ZN(n14130) );
  AOI22_X1 U16128 ( .A1(n14180), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n14128), 
        .B2(n15825), .ZN(n14129) );
  OAI211_X1 U16129 ( .C1(n14180), .C2(n14268), .A(n14130), .B(n14129), .ZN(
        n14131) );
  AOI21_X1 U16130 ( .B1(n14269), .B2(n15484), .A(n14131), .ZN(n14136) );
  XOR2_X1 U16131 ( .A(n14133), .B(n14132), .Z(n14272) );
  NAND2_X1 U16132 ( .A1(n14272), .A2(n14134), .ZN(n14135) );
  OAI211_X1 U16133 ( .C1(n14275), .C2(n14137), .A(n14136), .B(n14135), .ZN(
        P2_U3248) );
  NAND2_X1 U16134 ( .A1(n14138), .A2(n14152), .ZN(n14139) );
  NAND3_X1 U16135 ( .A1(n14140), .A2(n15556), .A3(n14139), .ZN(n14142) );
  AND2_X1 U16136 ( .A1(n14142), .A2(n14141), .ZN(n14277) );
  INV_X1 U16137 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n14144) );
  OAI22_X1 U16138 ( .A1(n15831), .A2(n14144), .B1(n14143), .B2(n15503), .ZN(
        n14149) );
  AOI21_X1 U16139 ( .B1(n14145), .B2(n14341), .A(n15561), .ZN(n14147) );
  NAND2_X1 U16140 ( .A1(n14147), .A2(n14146), .ZN(n14276) );
  NOR2_X1 U16141 ( .A1(n14276), .A2(n15829), .ZN(n14148) );
  AOI211_X1 U16142 ( .C1(n15827), .C2(n14341), .A(n14149), .B(n14148), .ZN(
        n14156) );
  INV_X1 U16143 ( .A(n14150), .ZN(n14158) );
  NAND2_X1 U16144 ( .A1(n6487), .A2(n14158), .ZN(n14157) );
  NAND2_X1 U16145 ( .A1(n14157), .A2(n14151), .ZN(n14154) );
  INV_X1 U16146 ( .A(n14152), .ZN(n14153) );
  XNOR2_X1 U16147 ( .A(n14154), .B(n14153), .ZN(n14278) );
  OR2_X1 U16148 ( .A1(n14278), .A2(n14200), .ZN(n14155) );
  OAI211_X1 U16149 ( .C1(n14277), .C2(n14180), .A(n14156), .B(n14155), .ZN(
        P2_U3249) );
  OAI21_X1 U16150 ( .B1(n6487), .B2(n14158), .A(n14157), .ZN(n14284) );
  INV_X1 U16151 ( .A(n14284), .ZN(n14173) );
  XNOR2_X1 U16152 ( .A(n14159), .B(n14158), .ZN(n14164) );
  OAI22_X1 U16153 ( .A1(n14161), .A2(n15493), .B1(n14160), .B2(n15495), .ZN(
        n14162) );
  AOI21_X1 U16154 ( .B1(n14284), .B2(n15550), .A(n14162), .ZN(n14163) );
  OAI21_X1 U16155 ( .B1(n14164), .B2(n14274), .A(n14163), .ZN(n14282) );
  NAND2_X1 U16156 ( .A1(n14282), .A2(n15831), .ZN(n14171) );
  INV_X1 U16157 ( .A(n14145), .ZN(n14165) );
  AOI211_X1 U16158 ( .C1(n14166), .C2(n6637), .A(n15561), .B(n14165), .ZN(
        n14283) );
  AOI22_X1 U16159 ( .A1(n14180), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n14167), 
        .B2(n15825), .ZN(n14168) );
  OAI21_X1 U16160 ( .B1(n14346), .B2(n15504), .A(n14168), .ZN(n14169) );
  AOI21_X1 U16161 ( .B1(n14283), .B2(n15484), .A(n14169), .ZN(n14170) );
  OAI211_X1 U16162 ( .C1(n14173), .C2(n14172), .A(n14171), .B(n14170), .ZN(
        P2_U3250) );
  XOR2_X1 U16163 ( .A(n14174), .B(n14176), .Z(n14289) );
  XOR2_X1 U16164 ( .A(n14176), .B(n14175), .Z(n14291) );
  NAND2_X1 U16165 ( .A1(n14291), .A2(n14177), .ZN(n14186) );
  AOI22_X1 U16166 ( .A1(n14180), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n14178), 
        .B2(n15825), .ZN(n14179) );
  OAI21_X1 U16167 ( .B1(n14180), .B2(n14288), .A(n14179), .ZN(n14183) );
  OAI211_X1 U16168 ( .C1(n14351), .C2(n14193), .A(n6637), .B(n14181), .ZN(
        n14287) );
  NOR2_X1 U16169 ( .A1(n14287), .A2(n15829), .ZN(n14182) );
  AOI211_X1 U16170 ( .C1(n15827), .C2(n14184), .A(n14183), .B(n14182), .ZN(
        n14185) );
  OAI211_X1 U16171 ( .C1(n14289), .C2(n14200), .A(n14186), .B(n14185), .ZN(
        P2_U3251) );
  XNOR2_X1 U16172 ( .A(n14187), .B(n14198), .ZN(n14192) );
  AOI222_X1 U16173 ( .A1(n15556), .A2(n14192), .B1(n14191), .B2(n14190), .C1(
        n14189), .C2(n14188), .ZN(n14298) );
  AOI211_X1 U16174 ( .C1(n14296), .C2(n14194), .A(n15561), .B(n14193), .ZN(
        n14295) );
  AOI22_X1 U16175 ( .A1(n14180), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n14195), 
        .B2(n15825), .ZN(n14196) );
  OAI21_X1 U16176 ( .B1(n14197), .B2(n15504), .A(n14196), .ZN(n14202) );
  XNOR2_X1 U16177 ( .A(n14199), .B(n14198), .ZN(n14299) );
  NOR2_X1 U16178 ( .A1(n14299), .A2(n14200), .ZN(n14201) );
  AOI211_X1 U16179 ( .C1(n14295), .C2(n15484), .A(n14202), .B(n14201), .ZN(
        n14203) );
  OAI21_X1 U16180 ( .B1(n14298), .B2(n14180), .A(n14203), .ZN(P2_U3252) );
  NOR2_X1 U16181 ( .A1(n14205), .A2(n14204), .ZN(n14311) );
  MUX2_X1 U16182 ( .A(n14206), .B(n14311), .S(n15580), .Z(n14207) );
  OAI21_X1 U16183 ( .B1(n14314), .B2(n14294), .A(n14207), .ZN(P2_U3529) );
  MUX2_X1 U16184 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14319), .S(n15580), .Z(
        P2_U3525) );
  MUX2_X1 U16185 ( .A(n14320), .B(P2_REG1_REG_25__SCAN_IN), .S(n15578), .Z(
        n14215) );
  INV_X1 U16186 ( .A(n14215), .ZN(n14216) );
  OAI21_X1 U16187 ( .B1(n14321), .B2(n14294), .A(n14216), .ZN(P2_U3524) );
  INV_X1 U16188 ( .A(n14217), .ZN(n14220) );
  OAI211_X1 U16189 ( .C1(n14220), .C2(n15565), .A(n14219), .B(n14218), .ZN(
        n14221) );
  AOI21_X1 U16190 ( .B1(n14222), .B2(n15556), .A(n14221), .ZN(n14223) );
  OAI21_X1 U16191 ( .B1(n14310), .B2(n14224), .A(n14223), .ZN(n14322) );
  MUX2_X1 U16192 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14322), .S(n15580), .Z(
        P2_U3523) );
  OAI211_X1 U16193 ( .C1(n14227), .C2(n15565), .A(n14226), .B(n14225), .ZN(
        n14228) );
  AOI21_X1 U16194 ( .B1(n14229), .B2(n15556), .A(n14228), .ZN(n14230) );
  OAI21_X1 U16195 ( .B1(n14310), .B2(n14231), .A(n14230), .ZN(n14323) );
  MUX2_X1 U16196 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14323), .S(n15580), .Z(
        P2_U3522) );
  INV_X1 U16197 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n14236) );
  INV_X1 U16198 ( .A(n14232), .ZN(n14235) );
  AOI211_X1 U16199 ( .C1(n14235), .C2(n14271), .A(n14234), .B(n14233), .ZN(
        n14324) );
  MUX2_X1 U16200 ( .A(n14236), .B(n14324), .S(n15580), .Z(n14237) );
  OAI21_X1 U16201 ( .B1(n14327), .B2(n14294), .A(n14237), .ZN(P2_U3521) );
  NAND2_X1 U16202 ( .A1(n14238), .A2(n15556), .ZN(n14242) );
  AND2_X1 U16203 ( .A1(n14240), .A2(n14239), .ZN(n14241) );
  OAI211_X1 U16204 ( .C1(n14310), .C2(n14243), .A(n14242), .B(n14241), .ZN(
        n14328) );
  MUX2_X1 U16205 ( .A(n14328), .B(P2_REG1_REG_21__SCAN_IN), .S(n15578), .Z(
        n14244) );
  INV_X1 U16206 ( .A(n14244), .ZN(n14245) );
  OAI21_X1 U16207 ( .B1(n7918), .B2(n14294), .A(n14245), .ZN(P2_U3520) );
  NAND2_X1 U16208 ( .A1(n14246), .A2(n15556), .ZN(n14250) );
  AND2_X1 U16209 ( .A1(n14248), .A2(n14247), .ZN(n14249) );
  OAI211_X1 U16210 ( .C1(n14310), .C2(n14251), .A(n14250), .B(n14249), .ZN(
        n14331) );
  MUX2_X1 U16211 ( .A(n14331), .B(P2_REG1_REG_20__SCAN_IN), .S(n15578), .Z(
        n14252) );
  INV_X1 U16212 ( .A(n14252), .ZN(n14253) );
  OAI21_X1 U16213 ( .B1(n14335), .B2(n14294), .A(n14253), .ZN(P2_U3519) );
  OAI211_X1 U16214 ( .C1(n14256), .C2(n15565), .A(n14255), .B(n14254), .ZN(
        n14257) );
  AOI21_X1 U16215 ( .B1(n14258), .B2(n15556), .A(n14257), .ZN(n14259) );
  OAI21_X1 U16216 ( .B1(n14310), .B2(n14260), .A(n14259), .ZN(n14336) );
  MUX2_X1 U16217 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n14336), .S(n15580), .Z(
        P2_U3518) );
  OAI21_X1 U16218 ( .B1(n14262), .B2(n15565), .A(n14261), .ZN(n14263) );
  AOI211_X1 U16219 ( .C1(n14265), .C2(n15556), .A(n14264), .B(n14263), .ZN(
        n14266) );
  OAI21_X1 U16220 ( .B1(n14310), .B2(n14267), .A(n14266), .ZN(n14337) );
  MUX2_X1 U16221 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14337), .S(n15580), .Z(
        P2_U3517) );
  OAI21_X1 U16222 ( .B1(n7923), .B2(n15565), .A(n14268), .ZN(n14270) );
  AOI211_X1 U16223 ( .C1(n14272), .C2(n14271), .A(n14270), .B(n14269), .ZN(
        n14273) );
  OAI21_X1 U16224 ( .B1(n14275), .B2(n14274), .A(n14273), .ZN(n14338) );
  MUX2_X1 U16225 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n14338), .S(n15580), .Z(
        P2_U3516) );
  OAI211_X1 U16226 ( .C1(n14310), .C2(n14278), .A(n14277), .B(n14276), .ZN(
        n14339) );
  MUX2_X1 U16227 ( .A(n14339), .B(P2_REG1_REG_16__SCAN_IN), .S(n15578), .Z(
        n14279) );
  AOI21_X1 U16228 ( .B1(n14280), .B2(n14341), .A(n14279), .ZN(n14281) );
  INV_X1 U16229 ( .A(n14281), .ZN(P2_U3515) );
  AOI211_X1 U16230 ( .C1(n15560), .C2(n14284), .A(n14283), .B(n14282), .ZN(
        n14343) );
  MUX2_X1 U16231 ( .A(n14285), .B(n14343), .S(n15580), .Z(n14286) );
  OAI21_X1 U16232 ( .B1(n14346), .B2(n14294), .A(n14286), .ZN(P2_U3514) );
  OAI211_X1 U16233 ( .C1(n14289), .C2(n14310), .A(n14288), .B(n14287), .ZN(
        n14290) );
  AOI21_X1 U16234 ( .B1(n15556), .B2(n14291), .A(n14290), .ZN(n14347) );
  MUX2_X1 U16235 ( .A(n14292), .B(n14347), .S(n15580), .Z(n14293) );
  OAI21_X1 U16236 ( .B1(n14351), .B2(n14294), .A(n14293), .ZN(P2_U3513) );
  AOI21_X1 U16237 ( .B1(n15525), .B2(n14296), .A(n14295), .ZN(n14297) );
  OAI211_X1 U16238 ( .C1(n14310), .C2(n14299), .A(n14298), .B(n14297), .ZN(
        n14352) );
  MUX2_X1 U16239 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n14352), .S(n15580), .Z(
        P2_U3512) );
  AOI21_X1 U16240 ( .B1(n15525), .B2(n14301), .A(n14300), .ZN(n14302) );
  OAI211_X1 U16241 ( .C1(n14310), .C2(n14304), .A(n14303), .B(n14302), .ZN(
        n14353) );
  MUX2_X1 U16242 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n14353), .S(n15580), .Z(
        P2_U3508) );
  AOI211_X1 U16243 ( .C1(n15525), .C2(n14307), .A(n14306), .B(n14305), .ZN(
        n14308) );
  OAI21_X1 U16244 ( .B1(n14310), .B2(n14309), .A(n14308), .ZN(n14354) );
  MUX2_X1 U16245 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n14354), .S(n15580), .Z(
        P2_U3505) );
  INV_X1 U16246 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n14312) );
  MUX2_X1 U16247 ( .A(n14312), .B(n14311), .S(n15571), .Z(n14313) );
  OAI21_X1 U16248 ( .B1(n14314), .B2(n14350), .A(n14313), .ZN(P2_U3497) );
  OAI21_X1 U16249 ( .B1(n14318), .B2(n14350), .A(n14317), .ZN(P2_U3494) );
  MUX2_X1 U16250 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14319), .S(n15571), .Z(
        P2_U3493) );
  MUX2_X1 U16251 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14322), .S(n15571), .Z(
        P2_U3491) );
  MUX2_X1 U16252 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14323), .S(n15571), .Z(
        P2_U3490) );
  MUX2_X1 U16253 ( .A(n14325), .B(n14324), .S(n15571), .Z(n14326) );
  OAI21_X1 U16254 ( .B1(n14327), .B2(n14350), .A(n14326), .ZN(P2_U3489) );
  MUX2_X1 U16255 ( .A(n14328), .B(P2_REG0_REG_21__SCAN_IN), .S(n15569), .Z(
        n14329) );
  INV_X1 U16256 ( .A(n14329), .ZN(n14330) );
  OAI21_X1 U16257 ( .B1(n7918), .B2(n14350), .A(n14330), .ZN(P2_U3488) );
  INV_X1 U16258 ( .A(n14331), .ZN(n14333) );
  MUX2_X1 U16259 ( .A(n14333), .B(n14332), .S(n15569), .Z(n14334) );
  OAI21_X1 U16260 ( .B1(n14335), .B2(n14350), .A(n14334), .ZN(P2_U3487) );
  MUX2_X1 U16261 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n14336), .S(n15571), .Z(
        P2_U3486) );
  MUX2_X1 U16262 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14337), .S(n15571), .Z(
        P2_U3484) );
  MUX2_X1 U16263 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n14338), .S(n15571), .Z(
        P2_U3481) );
  MUX2_X1 U16264 ( .A(n14339), .B(P2_REG0_REG_16__SCAN_IN), .S(n15569), .Z(
        n14340) );
  AOI21_X1 U16265 ( .B1(n10258), .B2(n14341), .A(n14340), .ZN(n14342) );
  INV_X1 U16266 ( .A(n14342), .ZN(P2_U3478) );
  MUX2_X1 U16267 ( .A(n14344), .B(n14343), .S(n15571), .Z(n14345) );
  OAI21_X1 U16268 ( .B1(n14346), .B2(n14350), .A(n14345), .ZN(P2_U3475) );
  MUX2_X1 U16269 ( .A(n14348), .B(n14347), .S(n15571), .Z(n14349) );
  OAI21_X1 U16270 ( .B1(n14351), .B2(n14350), .A(n14349), .ZN(P2_U3472) );
  MUX2_X1 U16271 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n14352), .S(n15571), .Z(
        P2_U3469) );
  MUX2_X1 U16272 ( .A(P2_REG0_REG_9__SCAN_IN), .B(n14353), .S(n15571), .Z(
        P2_U3457) );
  MUX2_X1 U16273 ( .A(P2_REG0_REG_6__SCAN_IN), .B(n14354), .S(n15571), .Z(
        P2_U3448) );
  INV_X1 U16274 ( .A(n14355), .ZN(n15157) );
  NOR4_X1 U16275 ( .A1(n14357), .A2(P2_IR_REG_30__SCAN_IN), .A3(n14356), .A4(
        P2_U3088), .ZN(n14358) );
  AOI21_X1 U16276 ( .B1(n14359), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n14358), 
        .ZN(n14360) );
  OAI21_X1 U16277 ( .B1(n15157), .B2(n14374), .A(n14360), .ZN(P2_U3296) );
  INV_X1 U16278 ( .A(n14361), .ZN(n15161) );
  OAI222_X1 U16279 ( .A1(n14363), .A2(P2_U3088), .B1(n14372), .B2(n14362), 
        .C1(n14367), .C2(n15161), .ZN(P2_U3298) );
  OAI222_X1 U16280 ( .A1(P2_U3088), .A2(n14366), .B1(n14374), .B2(n14365), 
        .C1(n14364), .C2(n14372), .ZN(P2_U3300) );
  OAI222_X1 U16281 ( .A1(P2_U3088), .A2(n14369), .B1(n14372), .B2(n14368), 
        .C1(n14367), .C2(n15168), .ZN(P2_U3301) );
  INV_X1 U16282 ( .A(n14370), .ZN(n14375) );
  INV_X1 U16283 ( .A(n14371), .ZN(n15172) );
  OAI222_X1 U16284 ( .A1(n14375), .A2(P2_U3088), .B1(n14374), .B2(n15172), 
        .C1(n14373), .C2(n14372), .ZN(P2_U3302) );
  MUX2_X1 U16285 ( .A(n14376), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  INV_X1 U16286 ( .A(n14377), .ZN(n14378) );
  AOI21_X1 U16287 ( .B1(n14380), .B2(n14379), .A(n14378), .ZN(n14388) );
  INV_X1 U16288 ( .A(n14381), .ZN(n14385) );
  AOI21_X1 U16289 ( .B1(n14491), .B2(n14383), .A(n14382), .ZN(n14384) );
  OAI21_X1 U16290 ( .B1(n14494), .B2(n14385), .A(n14384), .ZN(n14386) );
  AOI21_X1 U16291 ( .B1(n14496), .B2(n15107), .A(n14386), .ZN(n14387) );
  OAI21_X1 U16292 ( .B1(n14388), .B2(n14498), .A(n14387), .ZN(P1_U3215) );
  XOR2_X1 U16293 ( .A(n14390), .B(n14389), .Z(n14395) );
  NAND2_X1 U16294 ( .A1(n14830), .A2(n14473), .ZN(n14392) );
  AOI22_X1 U16295 ( .A1(n14831), .A2(n14478), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14391) );
  OAI211_X1 U16296 ( .C1(n14494), .C2(n14836), .A(n14392), .B(n14391), .ZN(
        n14393) );
  AOI21_X1 U16297 ( .B1(n15051), .B2(n14496), .A(n14393), .ZN(n14394) );
  OAI21_X1 U16298 ( .B1(n14395), .B2(n14498), .A(n14394), .ZN(P1_U3216) );
  AOI21_X1 U16299 ( .B1(n14397), .B2(n14396), .A(n14498), .ZN(n14399) );
  NAND2_X1 U16300 ( .A1(n14399), .A2(n14398), .ZN(n14403) );
  NAND2_X1 U16301 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14647)
         );
  OAI21_X1 U16302 ( .B1(n14482), .B2(n14869), .A(n14647), .ZN(n14401) );
  NOR2_X1 U16303 ( .A1(n14494), .A2(n14896), .ZN(n14400) );
  AOI211_X1 U16304 ( .C1(n14478), .C2(n14902), .A(n14401), .B(n14400), .ZN(
        n14402) );
  OAI211_X1 U16305 ( .C1(n14899), .C2(n14468), .A(n14403), .B(n14402), .ZN(
        P1_U3219) );
  INV_X1 U16306 ( .A(n14404), .ZN(n14405) );
  AOI21_X1 U16307 ( .B1(n14407), .B2(n14406), .A(n14405), .ZN(n14412) );
  INV_X1 U16308 ( .A(n14478), .ZN(n14471) );
  AOI22_X1 U16309 ( .A1(n14831), .A2(n14473), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14409) );
  NAND2_X1 U16310 ( .A1(n14479), .A2(n14873), .ZN(n14408) );
  OAI211_X1 U16311 ( .C1(n14869), .C2(n14471), .A(n14409), .B(n14408), .ZN(
        n14410) );
  AOI21_X1 U16312 ( .B1(n15066), .B2(n14496), .A(n14410), .ZN(n14411) );
  OAI21_X1 U16313 ( .B1(n14412), .B2(n14498), .A(n14411), .ZN(P1_U3223) );
  AOI21_X1 U16314 ( .B1(n14414), .B2(n14413), .A(n14498), .ZN(n14416) );
  NAND2_X1 U16315 ( .A1(n14416), .A2(n14415), .ZN(n14423) );
  NOR2_X1 U16316 ( .A1(n14417), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14580) );
  INV_X1 U16317 ( .A(n14418), .ZN(n14419) );
  NOR2_X1 U16318 ( .A1(n14494), .A2(n14419), .ZN(n14420) );
  AOI211_X1 U16319 ( .C1(n14491), .C2(n14421), .A(n14580), .B(n14420), .ZN(
        n14422) );
  OAI211_X1 U16320 ( .C1(n7770), .C2(n14468), .A(n14423), .B(n14422), .ZN(
        P1_U3224) );
  XNOR2_X1 U16321 ( .A(n14424), .B(n14425), .ZN(n14488) );
  NOR2_X1 U16322 ( .A1(n14488), .A2(n14487), .ZN(n14486) );
  AOI21_X1 U16323 ( .B1(n14425), .B2(n14424), .A(n14486), .ZN(n14429) );
  XNOR2_X1 U16324 ( .A(n14427), .B(n14426), .ZN(n14428) );
  XNOR2_X1 U16325 ( .A(n14429), .B(n14428), .ZN(n14436) );
  OR2_X1 U16326 ( .A1(n14921), .A2(n14980), .ZN(n14431) );
  NAND2_X1 U16327 ( .A1(n14690), .A2(n14982), .ZN(n14430) );
  AND2_X1 U16328 ( .A1(n14431), .A2(n14430), .ZN(n15093) );
  NAND2_X1 U16329 ( .A1(n14479), .A2(n14947), .ZN(n14432) );
  NAND2_X1 U16330 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14604)
         );
  OAI211_X1 U16331 ( .C1(n15093), .C2(n14433), .A(n14432), .B(n14604), .ZN(
        n14434) );
  AOI21_X1 U16332 ( .B1(n14692), .B2(n14496), .A(n14434), .ZN(n14435) );
  OAI21_X1 U16333 ( .B1(n14436), .B2(n14498), .A(n14435), .ZN(P1_U3226) );
  XOR2_X1 U16334 ( .A(n14438), .B(n14437), .Z(n14443) );
  NAND2_X1 U16335 ( .A1(n14478), .A2(n14691), .ZN(n14439) );
  NAND2_X1 U16336 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14616)
         );
  OAI211_X1 U16337 ( .C1(n14933), .C2(n14482), .A(n14439), .B(n14616), .ZN(
        n14440) );
  AOI21_X1 U16338 ( .B1(n14479), .B2(n14934), .A(n14440), .ZN(n14442) );
  NAND2_X1 U16339 ( .A1(n15088), .A2(n14496), .ZN(n14441) );
  OAI211_X1 U16340 ( .C1(n14443), .C2(n14498), .A(n14442), .B(n14441), .ZN(
        P1_U3228) );
  XOR2_X1 U16341 ( .A(n14444), .B(n14445), .Z(n14450) );
  AOI22_X1 U16342 ( .A1(n14856), .A2(n14478), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14447) );
  NAND2_X1 U16343 ( .A1(n14479), .A2(n14820), .ZN(n14446) );
  OAI211_X1 U16344 ( .C1(n14812), .C2(n14482), .A(n14447), .B(n14446), .ZN(
        n14448) );
  AOI21_X1 U16345 ( .B1(n15046), .B2(n14496), .A(n14448), .ZN(n14449) );
  OAI21_X1 U16346 ( .B1(n14450), .B2(n14498), .A(n14449), .ZN(P1_U3229) );
  OAI211_X1 U16347 ( .C1(n14453), .C2(n14452), .A(n14451), .B(n14462), .ZN(
        n14458) );
  NAND2_X1 U16348 ( .A1(n14478), .A2(n14983), .ZN(n14455) );
  OAI211_X1 U16349 ( .C1(n14981), .C2(n14482), .A(n14455), .B(n14454), .ZN(
        n14456) );
  AOI21_X1 U16350 ( .B1(n14479), .B2(n14975), .A(n14456), .ZN(n14457) );
  OAI211_X1 U16351 ( .C1(n14977), .C2(n14468), .A(n14458), .B(n14457), .ZN(
        P1_U3234) );
  OAI21_X1 U16352 ( .B1(n14461), .B2(n14460), .A(n14459), .ZN(n14463) );
  NAND2_X1 U16353 ( .A1(n14463), .A2(n14462), .ZN(n14467) );
  INV_X1 U16354 ( .A(n14855), .ZN(n14703) );
  AOI22_X1 U16355 ( .A1(n14856), .A2(n14473), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14464) );
  OAI21_X1 U16356 ( .B1(n14703), .B2(n14471), .A(n14464), .ZN(n14465) );
  AOI21_X1 U16357 ( .B1(n14857), .B2(n14479), .A(n14465), .ZN(n14466) );
  OAI211_X1 U16358 ( .C1(n14468), .C2(n15058), .A(n14467), .B(n14466), .ZN(
        P1_U3235) );
  XOR2_X1 U16359 ( .A(n14469), .B(n14470), .Z(n14477) );
  NAND2_X1 U16360 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14629)
         );
  OAI21_X1 U16361 ( .B1(n14471), .B2(n14921), .A(n14629), .ZN(n14472) );
  AOI21_X1 U16362 ( .B1(n14473), .B2(n14698), .A(n14472), .ZN(n14474) );
  OAI21_X1 U16363 ( .B1(n14914), .B2(n14494), .A(n14474), .ZN(n14475) );
  AOI21_X1 U16364 ( .B1(n15083), .B2(n14496), .A(n14475), .ZN(n14476) );
  OAI21_X1 U16365 ( .B1(n14477), .B2(n14498), .A(n14476), .ZN(P1_U3238) );
  AOI22_X1 U16366 ( .A1(n14711), .A2(n14478), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14481) );
  NAND2_X1 U16367 ( .A1(n14782), .A2(n14479), .ZN(n14480) );
  OAI211_X1 U16368 ( .C1(n14783), .C2(n14482), .A(n14481), .B(n14480), .ZN(
        n14483) );
  AOI21_X1 U16369 ( .B1(n15033), .B2(n14496), .A(n14483), .ZN(n14484) );
  OAI21_X1 U16370 ( .B1(n14485), .B2(n14498), .A(n14484), .ZN(P1_U3240) );
  AOI21_X1 U16371 ( .B1(n14488), .B2(n14487), .A(n14486), .ZN(n14499) );
  OR2_X1 U16372 ( .A1(n14932), .A2(n14980), .ZN(n14490) );
  OR2_X1 U16373 ( .A1(n14981), .A2(n14931), .ZN(n14489) );
  NAND2_X1 U16374 ( .A1(n14490), .A2(n14489), .ZN(n15102) );
  NAND2_X1 U16375 ( .A1(n14491), .A2(n15102), .ZN(n14492) );
  OAI211_X1 U16376 ( .C1(n14494), .C2(n14962), .A(n14493), .B(n14492), .ZN(
        n14495) );
  AOI21_X1 U16377 ( .B1(n15103), .B2(n14496), .A(n14495), .ZN(n14497) );
  OAI21_X1 U16378 ( .B1(n14499), .B2(n14498), .A(n14497), .ZN(P1_U3241) );
  MUX2_X1 U16379 ( .A(n14653), .B(P1_DATAO_REG_31__SCAN_IN), .S(n14525), .Z(
        P1_U3591) );
  MUX2_X1 U16380 ( .A(n14727), .B(P1_DATAO_REG_30__SCAN_IN), .S(n14525), .Z(
        P1_U3590) );
  MUX2_X1 U16381 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14740), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16382 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14758), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16383 ( .A(n14741), .B(P1_DATAO_REG_27__SCAN_IN), .S(n14525), .Z(
        P1_U3587) );
  MUX2_X1 U16384 ( .A(n14800), .B(P1_DATAO_REG_26__SCAN_IN), .S(n14525), .Z(
        P1_U3586) );
  MUX2_X1 U16385 ( .A(n14711), .B(P1_DATAO_REG_25__SCAN_IN), .S(n14525), .Z(
        P1_U3585) );
  MUX2_X1 U16386 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14830), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16387 ( .A(n14856), .B(P1_DATAO_REG_23__SCAN_IN), .S(n14525), .Z(
        P1_U3583) );
  MUX2_X1 U16388 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14831), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16389 ( .A(n14855), .B(P1_DATAO_REG_21__SCAN_IN), .S(n14525), .Z(
        P1_U3581) );
  MUX2_X1 U16390 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14904), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16391 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14698), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16392 ( .A(n14902), .B(P1_DATAO_REG_18__SCAN_IN), .S(n14525), .Z(
        P1_U3578) );
  MUX2_X1 U16393 ( .A(n14500), .B(P1_DATAO_REG_17__SCAN_IN), .S(n14525), .Z(
        P1_U3577) );
  MUX2_X1 U16394 ( .A(n14691), .B(P1_DATAO_REG_16__SCAN_IN), .S(n14525), .Z(
        P1_U3576) );
  MUX2_X1 U16395 ( .A(n14690), .B(P1_DATAO_REG_15__SCAN_IN), .S(n14525), .Z(
        P1_U3575) );
  MUX2_X1 U16396 ( .A(n14689), .B(P1_DATAO_REG_14__SCAN_IN), .S(n14525), .Z(
        P1_U3574) );
  MUX2_X1 U16397 ( .A(n14501), .B(P1_DATAO_REG_13__SCAN_IN), .S(n14525), .Z(
        P1_U3573) );
  MUX2_X1 U16398 ( .A(n14983), .B(P1_DATAO_REG_12__SCAN_IN), .S(n14525), .Z(
        P1_U3572) );
  MUX2_X1 U16399 ( .A(n14502), .B(P1_DATAO_REG_11__SCAN_IN), .S(n14525), .Z(
        P1_U3571) );
  MUX2_X1 U16400 ( .A(n14503), .B(P1_DATAO_REG_10__SCAN_IN), .S(n14525), .Z(
        P1_U3570) );
  MUX2_X1 U16401 ( .A(n14504), .B(P1_DATAO_REG_9__SCAN_IN), .S(n14525), .Z(
        P1_U3569) );
  MUX2_X1 U16402 ( .A(n14505), .B(P1_DATAO_REG_8__SCAN_IN), .S(n14525), .Z(
        P1_U3568) );
  MUX2_X1 U16403 ( .A(n14506), .B(P1_DATAO_REG_7__SCAN_IN), .S(n14525), .Z(
        P1_U3567) );
  MUX2_X1 U16404 ( .A(n14507), .B(P1_DATAO_REG_6__SCAN_IN), .S(n14525), .Z(
        P1_U3566) );
  MUX2_X1 U16405 ( .A(n14508), .B(P1_DATAO_REG_5__SCAN_IN), .S(n14525), .Z(
        P1_U3565) );
  MUX2_X1 U16406 ( .A(n14509), .B(P1_DATAO_REG_4__SCAN_IN), .S(n14525), .Z(
        P1_U3564) );
  MUX2_X1 U16407 ( .A(n14510), .B(P1_DATAO_REG_3__SCAN_IN), .S(n14525), .Z(
        P1_U3563) );
  MUX2_X1 U16408 ( .A(n14511), .B(P1_DATAO_REG_2__SCAN_IN), .S(n14525), .Z(
        P1_U3562) );
  MUX2_X1 U16409 ( .A(n14512), .B(P1_DATAO_REG_1__SCAN_IN), .S(n14525), .Z(
        P1_U3561) );
  MUX2_X1 U16410 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9435), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI22_X1 U16411 ( .A1(n15287), .A2(n14513), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7003), .ZN(n14514) );
  AOI21_X1 U16412 ( .B1(n15279), .B2(n14517), .A(n14514), .ZN(n14522) );
  OAI211_X1 U16413 ( .C1(n14516), .C2(n14515), .A(n15270), .B(n14534), .ZN(
        n14521) );
  NAND2_X1 U16414 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14524) );
  MUX2_X1 U16415 ( .A(n10460), .B(P1_REG2_REG_1__SCAN_IN), .S(n14517), .Z(
        n14518) );
  INV_X1 U16416 ( .A(n14518), .ZN(n14519) );
  OAI211_X1 U16417 ( .C1(n10461), .C2(n14519), .A(n15277), .B(n14540), .ZN(
        n14520) );
  NAND3_X1 U16418 ( .A1(n14522), .A2(n14521), .A3(n14520), .ZN(P1_U3244) );
  MUX2_X1 U16419 ( .A(n14524), .B(n14523), .S(n14651), .Z(n14529) );
  AOI21_X1 U16420 ( .B1(n14527), .B2(n14526), .A(n14525), .ZN(n14528) );
  OAI21_X1 U16421 ( .B1(n14529), .B2(n15167), .A(n14528), .ZN(n15283) );
  OAI22_X1 U16422 ( .A1(n15287), .A2(n14531), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14530), .ZN(n14532) );
  AOI21_X1 U16423 ( .B1(n15279), .B2(n14537), .A(n14532), .ZN(n14545) );
  MUX2_X1 U16424 ( .A(n10445), .B(P1_REG1_REG_2__SCAN_IN), .S(n14537), .Z(
        n14535) );
  NAND3_X1 U16425 ( .A1(n14535), .A2(n14534), .A3(n14533), .ZN(n14536) );
  NAND3_X1 U16426 ( .A1(n15270), .A2(n14551), .A3(n14536), .ZN(n14544) );
  MUX2_X1 U16427 ( .A(n14538), .B(P1_REG2_REG_2__SCAN_IN), .S(n14537), .Z(
        n14541) );
  NAND3_X1 U16428 ( .A1(n14541), .A2(n14540), .A3(n14539), .ZN(n14542) );
  NAND3_X1 U16429 ( .A1(n15277), .A2(n14556), .A3(n14542), .ZN(n14543) );
  NAND4_X1 U16430 ( .A1(n15283), .A2(n14545), .A3(n14544), .A4(n14543), .ZN(
        P1_U3245) );
  INV_X1 U16431 ( .A(n14553), .ZN(n14548) );
  OAI22_X1 U16432 ( .A1(n15287), .A2(n14546), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9457), .ZN(n14547) );
  AOI21_X1 U16433 ( .B1(n15279), .B2(n14548), .A(n14547), .ZN(n14560) );
  MUX2_X1 U16434 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10449), .S(n14553), .Z(
        n14550) );
  NAND3_X1 U16435 ( .A1(n14551), .A2(n14550), .A3(n14549), .ZN(n14552) );
  NAND3_X1 U16436 ( .A1(n15270), .A2(n15267), .A3(n14552), .ZN(n14559) );
  MUX2_X1 U16437 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n11311), .S(n14553), .Z(
        n14555) );
  NAND3_X1 U16438 ( .A1(n14556), .A2(n14555), .A3(n14554), .ZN(n14557) );
  NAND3_X1 U16439 ( .A1(n15277), .A2(n15274), .A3(n14557), .ZN(n14558) );
  NAND3_X1 U16440 ( .A1(n14560), .A2(n14559), .A3(n14558), .ZN(P1_U3246) );
  NAND2_X1 U16441 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n14561) );
  OAI21_X1 U16442 ( .B1(n15287), .B2(n10387), .A(n14561), .ZN(n14562) );
  AOI21_X1 U16443 ( .B1(n15279), .B2(n14563), .A(n14562), .ZN(n14575) );
  OAI21_X1 U16444 ( .B1(n14566), .B2(n14565), .A(n14564), .ZN(n14567) );
  NAND2_X1 U16445 ( .A1(n15270), .A2(n14567), .ZN(n14574) );
  INV_X1 U16446 ( .A(n14568), .ZN(n14572) );
  NAND3_X1 U16447 ( .A1(n14570), .A2(n15276), .A3(n14569), .ZN(n14571) );
  NAND3_X1 U16448 ( .A1(n15277), .A2(n14572), .A3(n14571), .ZN(n14573) );
  NAND3_X1 U16449 ( .A1(n14575), .A2(n14574), .A3(n14573), .ZN(P1_U3248) );
  OAI21_X1 U16450 ( .B1(n14578), .B2(n14577), .A(n14576), .ZN(n14579) );
  NAND2_X1 U16451 ( .A1(n14579), .A2(n15270), .ZN(n14589) );
  AOI21_X1 U16452 ( .B1(n14631), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n14580), 
        .ZN(n14588) );
  OAI21_X1 U16453 ( .B1(n14583), .B2(n14582), .A(n14581), .ZN(n14584) );
  NAND2_X1 U16454 ( .A1(n14584), .A2(n15277), .ZN(n14587) );
  NAND2_X1 U16455 ( .A1(n15279), .A2(n14585), .ZN(n14586) );
  NAND4_X1 U16456 ( .A1(n14589), .A2(n14588), .A3(n14587), .A4(n14586), .ZN(
        P1_U3255) );
  INV_X1 U16457 ( .A(n14590), .ZN(n14591) );
  NAND2_X1 U16458 ( .A1(n14612), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n14593) );
  OAI21_X1 U16459 ( .B1(n14612), .B2(P1_REG2_REG_16__SCAN_IN), .A(n14593), 
        .ZN(n14595) );
  INV_X1 U16460 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n14594) );
  OAI211_X1 U16461 ( .C1(n14596), .C2(n14595), .A(n14608), .B(n15277), .ZN(
        n14607) );
  XNOR2_X1 U16462 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14612), .ZN(n14602) );
  INV_X1 U16463 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14599) );
  OAI211_X1 U16464 ( .C1(n14602), .C2(n14601), .A(n15270), .B(n14610), .ZN(
        n14603) );
  NAND2_X1 U16465 ( .A1(n14604), .A2(n14603), .ZN(n14605) );
  AOI21_X1 U16466 ( .B1(n14631), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n14605), 
        .ZN(n14606) );
  OAI211_X1 U16467 ( .C1(n14644), .C2(n14612), .A(n14607), .B(n14606), .ZN(
        P1_U3259) );
  INV_X1 U16468 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n15778) );
  MUX2_X1 U16469 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n15778), .S(n14625), .Z(
        n14620) );
  XNOR2_X1 U16470 ( .A(n14622), .B(n14620), .ZN(n14609) );
  NAND2_X1 U16471 ( .A1(n14609), .A2(n15277), .ZN(n14619) );
  XNOR2_X1 U16472 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14625), .ZN(n14614) );
  INV_X1 U16473 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14611) );
  OAI21_X1 U16474 ( .B1(n14612), .B2(n14611), .A(n14610), .ZN(n14613) );
  NAND2_X1 U16475 ( .A1(n14614), .A2(n14613), .ZN(n14624) );
  OAI211_X1 U16476 ( .C1(n14614), .C2(n14613), .A(n15270), .B(n14624), .ZN(
        n14615) );
  NAND2_X1 U16477 ( .A1(n14616), .A2(n14615), .ZN(n14617) );
  AOI21_X1 U16478 ( .B1(n14631), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n14617), 
        .ZN(n14618) );
  OAI211_X1 U16479 ( .C1(n14644), .C2(n14625), .A(n14619), .B(n14618), .ZN(
        P1_U3260) );
  INV_X1 U16480 ( .A(n14620), .ZN(n14621) );
  NAND2_X1 U16481 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14623), .ZN(n14641) );
  OAI211_X1 U16482 ( .C1(n14623), .C2(P1_REG2_REG_18__SCAN_IN), .A(n15277), 
        .B(n14641), .ZN(n14633) );
  XNOR2_X1 U16483 ( .A(n14635), .B(n14634), .ZN(n14627) );
  NAND2_X1 U16484 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n14627), .ZN(n14637) );
  OAI211_X1 U16485 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n14627), .A(n15270), 
        .B(n14637), .ZN(n14628) );
  NAND2_X1 U16486 ( .A1(n14629), .A2(n14628), .ZN(n14630) );
  AOI21_X1 U16487 ( .B1(n14631), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n14630), 
        .ZN(n14632) );
  OAI211_X1 U16488 ( .C1(n14644), .C2(n14634), .A(n14633), .B(n14632), .ZN(
        P1_U3261) );
  NAND2_X1 U16489 ( .A1(n14640), .A2(n14635), .ZN(n14636) );
  NAND2_X1 U16490 ( .A1(n14640), .A2(n14639), .ZN(n14642) );
  NAND2_X1 U16491 ( .A1(n14642), .A2(n14641), .ZN(n14643) );
  XOR2_X1 U16492 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n14643), .Z(n14646) );
  NOR2_X2 U16493 ( .A1(n14929), .A2(n15083), .ZN(n14912) );
  NAND2_X1 U16494 ( .A1(n14894), .A2(n15071), .ZN(n14885) );
  INV_X1 U16495 ( .A(n15027), .ZN(n14769) );
  NAND2_X1 U16496 ( .A1(n15009), .A2(n14725), .ZN(n14649) );
  XNOR2_X1 U16497 ( .A(n14649), .B(n15004), .ZN(n14650) );
  INV_X1 U16498 ( .A(P1_B_REG_SCAN_IN), .ZN(n15720) );
  OR2_X1 U16499 ( .A1(n14651), .A2(n15720), .ZN(n14652) );
  AND2_X1 U16500 ( .A1(n14903), .A2(n14652), .ZN(n14728) );
  NAND2_X1 U16501 ( .A1(n14728), .A2(n14653), .ZN(n15007) );
  NOR2_X1 U16502 ( .A1(n15336), .A2(n15007), .ZN(n14659) );
  NOR2_X1 U16503 ( .A1(n15004), .A2(n15311), .ZN(n14654) );
  AOI211_X1 U16504 ( .C1(n15336), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14659), 
        .B(n14654), .ZN(n14655) );
  OAI21_X1 U16505 ( .B1(n15003), .B2(n14952), .A(n14655), .ZN(P1_U3263) );
  XNOR2_X1 U16506 ( .A(n14656), .B(n14725), .ZN(n14657) );
  NAND2_X1 U16507 ( .A1(n14657), .A2(n15328), .ZN(n15008) );
  NOR2_X1 U16508 ( .A1(n15009), .A2(n15311), .ZN(n14658) );
  AOI211_X1 U16509 ( .C1(n15336), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14659), 
        .B(n14658), .ZN(n14660) );
  OAI21_X1 U16510 ( .B1(n15008), .B2(n14952), .A(n14660), .ZN(P1_U3264) );
  NAND2_X1 U16511 ( .A1(n15116), .A2(n14661), .ZN(n14662) );
  AND2_X1 U16512 ( .A1(n14665), .A2(n14662), .ZN(n14663) );
  NAND2_X1 U16513 ( .A1(n14665), .A2(n14664), .ZN(n14667) );
  AND2_X1 U16514 ( .A1(n14667), .A2(n14666), .ZN(n14668) );
  AOI21_X1 U16515 ( .B1(n14692), .B2(n14932), .A(n14669), .ZN(n14670) );
  NAND2_X1 U16516 ( .A1(n14943), .A2(n14932), .ZN(n14672) );
  AOI22_X1 U16517 ( .A1(n15095), .A2(n14672), .B1(n14671), .B2(n14691), .ZN(
        n14673) );
  NAND2_X1 U16518 ( .A1(n15088), .A2(n14921), .ZN(n14674) );
  NAND2_X1 U16519 ( .A1(n14926), .A2(n14674), .ZN(n14676) );
  OR2_X1 U16520 ( .A1(n15088), .A2(n14921), .ZN(n14675) );
  OR2_X1 U16521 ( .A1(n15083), .A2(n14933), .ZN(n14677) );
  NAND2_X1 U16522 ( .A1(n15071), .A2(n14904), .ZN(n14679) );
  OR2_X1 U16523 ( .A1(n15066), .A2(n14703), .ZN(n14680) );
  NAND2_X1 U16524 ( .A1(n14827), .A2(n14829), .ZN(n14828) );
  NAND2_X1 U16525 ( .A1(n15051), .A2(n14811), .ZN(n14682) );
  NAND2_X1 U16526 ( .A1(n14822), .A2(n14830), .ZN(n14683) );
  INV_X1 U16527 ( .A(n14800), .ZN(n14684) );
  NAND2_X1 U16528 ( .A1(n15033), .A2(n14684), .ZN(n14685) );
  INV_X1 U16529 ( .A(n14748), .ZN(n15020) );
  NAND2_X1 U16530 ( .A1(n15020), .A2(n14758), .ZN(n14687) );
  NAND2_X1 U16531 ( .A1(n15107), .A2(n14689), .ZN(n14957) );
  OR2_X1 U16532 ( .A1(n14692), .A2(n14691), .ZN(n14693) );
  OR2_X1 U16533 ( .A1(n15083), .A2(n14902), .ZN(n14696) );
  NOR2_X1 U16534 ( .A1(n15066), .A2(n14855), .ZN(n14848) );
  INV_X1 U16535 ( .A(n14848), .ZN(n14699) );
  NAND2_X1 U16536 ( .A1(n14702), .A2(n14904), .ZN(n14847) );
  NAND2_X1 U16537 ( .A1(n14847), .A2(n14703), .ZN(n14705) );
  INV_X1 U16538 ( .A(n14847), .ZN(n14704) );
  AOI22_X1 U16539 ( .A1(n15066), .A2(n14705), .B1(n14704), .B2(n14855), .ZN(
        n14706) );
  NAND2_X1 U16540 ( .A1(n14849), .A2(n14706), .ZN(n14707) );
  NAND2_X1 U16541 ( .A1(n14707), .A2(n6532), .ZN(n14708) );
  NAND2_X1 U16542 ( .A1(n15051), .A2(n14856), .ZN(n14710) );
  NAND2_X1 U16543 ( .A1(n14795), .A2(n14711), .ZN(n14712) );
  NAND2_X1 U16544 ( .A1(n14792), .A2(n14712), .ZN(n14775) );
  INV_X1 U16545 ( .A(n14779), .ZN(n14774) );
  NAND2_X1 U16546 ( .A1(n15033), .A2(n14800), .ZN(n14713) );
  INV_X1 U16547 ( .A(n14716), .ZN(n14770) );
  OR2_X1 U16548 ( .A1(n15027), .A2(n14741), .ZN(n14749) );
  NAND2_X1 U16549 ( .A1(n14714), .A2(n14749), .ZN(n14718) );
  INV_X1 U16550 ( .A(n14718), .ZN(n14715) );
  NAND3_X1 U16551 ( .A1(n14716), .A2(n14715), .A3(n14717), .ZN(n14724) );
  AOI21_X1 U16552 ( .B1(n14719), .B2(n14718), .A(n14717), .ZN(n14723) );
  INV_X1 U16553 ( .A(n14719), .ZN(n14720) );
  NOR2_X1 U16554 ( .A1(n14721), .A2(n14720), .ZN(n14722) );
  INV_X1 U16555 ( .A(n14726), .ZN(n15012) );
  NAND2_X1 U16556 ( .A1(n15014), .A2(n15332), .ZN(n14735) );
  NAND2_X1 U16557 ( .A1(n15324), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n14730) );
  NAND2_X1 U16558 ( .A1(n14728), .A2(n14727), .ZN(n15010) );
  OAI22_X1 U16559 ( .A1(n14731), .A2(n14730), .B1(n15010), .B2(n14729), .ZN(
        n14733) );
  NAND2_X1 U16560 ( .A1(n14758), .A2(n14982), .ZN(n15011) );
  NOR2_X1 U16561 ( .A1(n15011), .A2(n15336), .ZN(n14732) );
  AOI211_X1 U16562 ( .C1(n15336), .C2(P1_REG2_REG_29__SCAN_IN), .A(n14733), 
        .B(n14732), .ZN(n14734) );
  OAI211_X1 U16563 ( .C1(n15012), .C2(n15311), .A(n14735), .B(n14734), .ZN(
        n14736) );
  AOI21_X1 U16564 ( .B1(n14992), .B2(n15016), .A(n14736), .ZN(n14737) );
  OAI21_X1 U16565 ( .B1(n15017), .B2(n14970), .A(n14737), .ZN(P1_U3356) );
  XNOR2_X1 U16566 ( .A(n14738), .B(n14752), .ZN(n14739) );
  AOI22_X1 U16567 ( .A1(n14741), .A2(n14982), .B1(n14903), .B2(n14740), .ZN(
        n14742) );
  OAI22_X1 U16568 ( .A1(n14744), .A2(n14997), .B1(n14743), .B2(n14935), .ZN(
        n14747) );
  NAND2_X1 U16569 ( .A1(n14748), .A2(n14763), .ZN(n14745) );
  NOR2_X1 U16570 ( .A1(n15021), .A2(n14840), .ZN(n14746) );
  AOI211_X1 U16571 ( .C1(n14995), .C2(n14748), .A(n14747), .B(n14746), .ZN(
        n14755) );
  INV_X1 U16572 ( .A(n14752), .ZN(n14750) );
  NAND2_X1 U16573 ( .A1(n14751), .A2(n14750), .ZN(n15019) );
  NAND2_X1 U16574 ( .A1(n14753), .A2(n14752), .ZN(n15018) );
  NAND3_X1 U16575 ( .A1(n15019), .A2(n14992), .A3(n15018), .ZN(n14754) );
  OAI211_X1 U16576 ( .C1(n7927), .C2(n15336), .A(n14755), .B(n14754), .ZN(
        P1_U3265) );
  OAI21_X1 U16577 ( .B1(n14757), .B2(n14772), .A(n14756), .ZN(n14762) );
  INV_X1 U16578 ( .A(n14781), .ZN(n14765) );
  INV_X1 U16579 ( .A(n14763), .ZN(n14764) );
  AOI211_X1 U16580 ( .C1(n15027), .C2(n14765), .A(n15344), .B(n14764), .ZN(
        n15026) );
  INV_X1 U16581 ( .A(n14766), .ZN(n14767) );
  AOI22_X1 U16582 ( .A1(n14767), .A2(n15324), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n15336), .ZN(n14768) );
  OAI21_X1 U16583 ( .B1(n14769), .B2(n15311), .A(n14768), .ZN(n14773) );
  OR2_X1 U16584 ( .A1(n14775), .A2(n14774), .ZN(n14776) );
  NAND2_X1 U16585 ( .A1(n14777), .A2(n14776), .ZN(n15036) );
  OAI21_X1 U16586 ( .B1(n14780), .B2(n14779), .A(n14778), .ZN(n15030) );
  NAND2_X1 U16587 ( .A1(n15030), .A2(n14993), .ZN(n14789) );
  AOI211_X1 U16588 ( .C1(n15033), .C2(n14796), .A(n15344), .B(n14781), .ZN(
        n15031) );
  INV_X1 U16589 ( .A(n15033), .ZN(n14786) );
  AOI22_X1 U16590 ( .A1(n14782), .A2(n15324), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n15336), .ZN(n14785) );
  OAI22_X1 U16591 ( .A1(n14783), .A2(n14980), .B1(n14812), .B2(n14931), .ZN(
        n15032) );
  NAND2_X1 U16592 ( .A1(n15032), .A2(n14935), .ZN(n14784) );
  OAI211_X1 U16593 ( .C1(n14786), .C2(n15311), .A(n14785), .B(n14784), .ZN(
        n14787) );
  AOI21_X1 U16594 ( .B1(n15031), .B2(n15332), .A(n14787), .ZN(n14788) );
  OAI211_X1 U16595 ( .C1(n15036), .C2(n14990), .A(n14789), .B(n14788), .ZN(
        P1_U3267) );
  XNOR2_X1 U16596 ( .A(n14791), .B(n14790), .ZN(n15044) );
  OAI21_X1 U16597 ( .B1(n14794), .B2(n14793), .A(n14792), .ZN(n15037) );
  AOI22_X1 U16598 ( .A1(n14795), .A2(n14995), .B1(n15336), .B2(
        P1_REG2_REG_25__SCAN_IN), .ZN(n14805) );
  AOI21_X1 U16599 ( .B1(n14795), .B2(n14808), .A(n15344), .ZN(n14797) );
  NAND2_X1 U16600 ( .A1(n14797), .A2(n14796), .ZN(n15039) );
  NOR2_X1 U16601 ( .A1(n14798), .A2(n14931), .ZN(n14799) );
  AOI21_X1 U16602 ( .B1(n14800), .B2(n14903), .A(n14799), .ZN(n15038) );
  OR2_X1 U16603 ( .A1(n14801), .A2(n14997), .ZN(n14802) );
  OAI211_X1 U16604 ( .C1(n15039), .C2(n9940), .A(n15038), .B(n14802), .ZN(
        n14803) );
  NAND2_X1 U16605 ( .A1(n14803), .A2(n14935), .ZN(n14804) );
  OAI211_X1 U16606 ( .C1(n15037), .C2(n14990), .A(n14805), .B(n14804), .ZN(
        n14806) );
  INV_X1 U16607 ( .A(n14806), .ZN(n14807) );
  OAI21_X1 U16608 ( .B1(n15044), .B2(n14970), .A(n14807), .ZN(P1_U3268) );
  INV_X1 U16609 ( .A(n14835), .ZN(n14809) );
  AOI211_X1 U16610 ( .C1(n15046), .C2(n14809), .A(n15344), .B(n7754), .ZN(
        n15045) );
  AOI21_X1 U16611 ( .B1(n14810), .B2(n14818), .A(n15400), .ZN(n14814) );
  OAI22_X1 U16612 ( .A1(n14812), .A2(n14980), .B1(n14811), .B2(n14931), .ZN(
        n14813) );
  AOI21_X1 U16613 ( .B1(n14815), .B2(n14814), .A(n14813), .ZN(n15048) );
  INV_X1 U16614 ( .A(n15048), .ZN(n14816) );
  AOI21_X1 U16615 ( .B1(n15045), .B2(n14817), .A(n14816), .ZN(n14826) );
  XNOR2_X1 U16616 ( .A(n14819), .B(n14818), .ZN(n15049) );
  INV_X1 U16617 ( .A(n15049), .ZN(n14824) );
  AOI22_X1 U16618 ( .A1(n14820), .A2(n15324), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n15336), .ZN(n14821) );
  OAI21_X1 U16619 ( .B1(n14822), .B2(n15311), .A(n14821), .ZN(n14823) );
  AOI21_X1 U16620 ( .B1(n14824), .B2(n14992), .A(n14823), .ZN(n14825) );
  OAI21_X1 U16621 ( .B1(n14826), .B2(n15336), .A(n14825), .ZN(P1_U3269) );
  OAI21_X1 U16622 ( .B1(n14827), .B2(n14829), .A(n14828), .ZN(n14832) );
  AOI222_X1 U16623 ( .A1(n15359), .A2(n14832), .B1(n14831), .B2(n14982), .C1(
        n14830), .C2(n14903), .ZN(n15056) );
  NOR2_X1 U16624 ( .A1(n14853), .A2(n14833), .ZN(n14834) );
  OR2_X1 U16625 ( .A1(n14835), .A2(n14834), .ZN(n15050) );
  INV_X1 U16626 ( .A(n14836), .ZN(n14837) );
  AOI22_X1 U16627 ( .A1(n14837), .A2(n15324), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n15336), .ZN(n14839) );
  NAND2_X1 U16628 ( .A1(n15051), .A2(n14995), .ZN(n14838) );
  OAI211_X1 U16629 ( .C1(n15050), .C2(n14840), .A(n14839), .B(n14838), .ZN(
        n14841) );
  INV_X1 U16630 ( .A(n14841), .ZN(n14846) );
  OR2_X1 U16631 ( .A1(n14843), .A2(n14842), .ZN(n15053) );
  NAND3_X1 U16632 ( .A1(n15053), .A2(n14844), .A3(n14992), .ZN(n14845) );
  OAI211_X1 U16633 ( .C1(n15056), .C2(n15336), .A(n14846), .B(n14845), .ZN(
        P1_U3270) );
  NAND2_X1 U16634 ( .A1(n14880), .A2(n14884), .ZN(n14879) );
  NAND2_X1 U16635 ( .A1(n14879), .A2(n14847), .ZN(n14865) );
  NOR2_X1 U16636 ( .A1(n14865), .A2(n14867), .ZN(n14864) );
  NOR2_X1 U16637 ( .A1(n14864), .A2(n14848), .ZN(n14850) );
  XNOR2_X1 U16638 ( .A(n14850), .B(n14849), .ZN(n15063) );
  OAI21_X1 U16639 ( .B1(n6534), .B2(n14852), .A(n14851), .ZN(n15061) );
  AOI211_X1 U16640 ( .C1(n14854), .C2(n14871), .A(n15344), .B(n14853), .ZN(
        n15060) );
  NAND2_X1 U16641 ( .A1(n15060), .A2(n15332), .ZN(n14861) );
  AOI22_X1 U16642 ( .A1(n14856), .A2(n14903), .B1(n14982), .B2(n14855), .ZN(
        n15057) );
  INV_X1 U16643 ( .A(n14857), .ZN(n14858) );
  OAI22_X1 U16644 ( .A1(n15057), .A2(n15336), .B1(n14858), .B2(n14997), .ZN(
        n14859) );
  AOI21_X1 U16645 ( .B1(P1_REG2_REG_22__SCAN_IN), .B2(n15336), .A(n14859), 
        .ZN(n14860) );
  OAI211_X1 U16646 ( .C1(n15311), .C2(n15058), .A(n14861), .B(n14860), .ZN(
        n14862) );
  AOI21_X1 U16647 ( .B1(n15061), .B2(n14993), .A(n14862), .ZN(n14863) );
  OAI21_X1 U16648 ( .B1(n15063), .B2(n14990), .A(n14863), .ZN(P1_U3271) );
  AOI21_X1 U16649 ( .B1(n14867), .B2(n14865), .A(n14864), .ZN(n15068) );
  XNOR2_X1 U16650 ( .A(n14866), .B(n14867), .ZN(n14868) );
  OAI222_X1 U16651 ( .A1(n14980), .A2(n14870), .B1(n14931), .B2(n14869), .C1(
        n14868), .C2(n15400), .ZN(n15064) );
  INV_X1 U16652 ( .A(n15066), .ZN(n14876) );
  AOI21_X1 U16653 ( .B1(n14885), .B2(n15066), .A(n15344), .ZN(n14872) );
  AND2_X1 U16654 ( .A1(n14872), .A2(n14871), .ZN(n15065) );
  NAND2_X1 U16655 ( .A1(n15065), .A2(n15332), .ZN(n14875) );
  AOI22_X1 U16656 ( .A1(n15336), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n14873), 
        .B2(n15324), .ZN(n14874) );
  OAI211_X1 U16657 ( .C1(n14876), .C2(n15311), .A(n14875), .B(n14874), .ZN(
        n14877) );
  AOI21_X1 U16658 ( .B1(n15064), .B2(n14935), .A(n14877), .ZN(n14878) );
  OAI21_X1 U16659 ( .B1(n15068), .B2(n14990), .A(n14878), .ZN(P1_U3272) );
  OAI21_X1 U16660 ( .B1(n14880), .B2(n14884), .A(n14879), .ZN(n15075) );
  INV_X1 U16661 ( .A(n14881), .ZN(n14882) );
  AOI21_X1 U16662 ( .B1(n14884), .B2(n14883), .A(n14882), .ZN(n15073) );
  OAI211_X1 U16663 ( .C1(n14894), .C2(n15071), .A(n15328), .B(n14885), .ZN(
        n15070) );
  INV_X1 U16664 ( .A(n14886), .ZN(n14887) );
  OAI22_X1 U16665 ( .A1(n15069), .A2(n15336), .B1(n14887), .B2(n14997), .ZN(
        n14889) );
  NOR2_X1 U16666 ( .A1(n15071), .A2(n15311), .ZN(n14888) );
  AOI211_X1 U16667 ( .C1(n15336), .C2(P1_REG2_REG_20__SCAN_IN), .A(n14889), 
        .B(n14888), .ZN(n14890) );
  OAI21_X1 U16668 ( .B1(n14952), .B2(n15070), .A(n14890), .ZN(n14891) );
  AOI21_X1 U16669 ( .B1(n15073), .B2(n14993), .A(n14891), .ZN(n14892) );
  OAI21_X1 U16670 ( .B1(n14990), .B2(n15075), .A(n14892), .ZN(P1_U3273) );
  XNOR2_X1 U16671 ( .A(n14893), .B(n14901), .ZN(n15080) );
  INV_X1 U16672 ( .A(n14912), .ZN(n14895) );
  AOI21_X1 U16673 ( .B1(n15076), .B2(n14895), .A(n14894), .ZN(n15077) );
  INV_X1 U16674 ( .A(n14896), .ZN(n14897) );
  AOI22_X1 U16675 ( .A1(n15336), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14897), 
        .B2(n15324), .ZN(n14898) );
  OAI21_X1 U16676 ( .B1(n14899), .B2(n15311), .A(n14898), .ZN(n14907) );
  OAI21_X1 U16677 ( .B1(n6535), .B2(n14901), .A(n14900), .ZN(n14905) );
  AOI222_X1 U16678 ( .A1(n15359), .A2(n14905), .B1(n14904), .B2(n14903), .C1(
        n14902), .C2(n14982), .ZN(n15079) );
  NOR2_X1 U16679 ( .A1(n15079), .A2(n15336), .ZN(n14906) );
  AOI211_X1 U16680 ( .C1(n15077), .C2(n14996), .A(n14907), .B(n14906), .ZN(
        n14908) );
  OAI21_X1 U16681 ( .B1(n15080), .B2(n14990), .A(n14908), .ZN(P1_U3274) );
  XOR2_X1 U16682 ( .A(n14909), .B(n14919), .Z(n15085) );
  INV_X1 U16683 ( .A(n14910), .ZN(n14911) );
  AOI21_X1 U16684 ( .B1(n15332), .B2(n14911), .A(n15333), .ZN(n14925) );
  AOI211_X1 U16685 ( .C1(n15083), .C2(n14929), .A(n15344), .B(n14912), .ZN(
        n15082) );
  INV_X1 U16686 ( .A(n15083), .ZN(n14913) );
  NOR2_X1 U16687 ( .A1(n14913), .A2(n15311), .ZN(n14917) );
  INV_X1 U16688 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14915) );
  OAI22_X1 U16689 ( .A1(n14935), .A2(n14915), .B1(n14914), .B2(n14997), .ZN(
        n14916) );
  AOI211_X1 U16690 ( .C1(n15082), .C2(n15332), .A(n14917), .B(n14916), .ZN(
        n14924) );
  XNOR2_X1 U16691 ( .A(n14918), .B(n14919), .ZN(n14920) );
  OAI222_X1 U16692 ( .A1(n14980), .A2(n14922), .B1(n14931), .B2(n14921), .C1(
        n14920), .C2(n15400), .ZN(n15081) );
  NAND2_X1 U16693 ( .A1(n15081), .A2(n14935), .ZN(n14923) );
  OAI211_X1 U16694 ( .C1(n15085), .C2(n14925), .A(n14924), .B(n14923), .ZN(
        P1_U3275) );
  XNOR2_X1 U16695 ( .A(n14926), .B(n14928), .ZN(n15092) );
  XOR2_X1 U16696 ( .A(n14927), .B(n14928), .Z(n15089) );
  NAND2_X1 U16697 ( .A1(n15089), .A2(n14992), .ZN(n14940) );
  INV_X1 U16698 ( .A(n14929), .ZN(n14930) );
  AOI211_X1 U16699 ( .C1(n15088), .C2(n14946), .A(n15344), .B(n14930), .ZN(
        n15086) );
  OAI22_X1 U16700 ( .A1(n14933), .A2(n14980), .B1(n14932), .B2(n14931), .ZN(
        n15087) );
  AOI22_X1 U16701 ( .A1(n14935), .A2(n15087), .B1(n14934), .B2(n15324), .ZN(
        n14937) );
  NAND2_X1 U16702 ( .A1(n15336), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14936) );
  OAI211_X1 U16703 ( .C1(n7755), .C2(n15311), .A(n14937), .B(n14936), .ZN(
        n14938) );
  AOI21_X1 U16704 ( .B1(n15086), .B2(n15332), .A(n14938), .ZN(n14939) );
  OAI211_X1 U16705 ( .C1(n15092), .C2(n14970), .A(n14940), .B(n14939), .ZN(
        P1_U3276) );
  XNOR2_X1 U16706 ( .A(n14941), .B(n6927), .ZN(n15099) );
  INV_X1 U16707 ( .A(n14959), .ZN(n14956) );
  NAND2_X1 U16708 ( .A1(n14942), .A2(n14956), .ZN(n14955) );
  NAND2_X1 U16709 ( .A1(n14955), .A2(n14943), .ZN(n14945) );
  XNOR2_X1 U16710 ( .A(n14945), .B(n14944), .ZN(n15097) );
  OAI211_X1 U16711 ( .C1(n14960), .C2(n15095), .A(n14946), .B(n15328), .ZN(
        n15094) );
  INV_X1 U16712 ( .A(n14947), .ZN(n14948) );
  OAI22_X1 U16713 ( .A1(n15336), .A2(n15093), .B1(n14948), .B2(n14997), .ZN(
        n14950) );
  NOR2_X1 U16714 ( .A1(n15095), .A2(n15311), .ZN(n14949) );
  AOI211_X1 U16715 ( .C1(n15336), .C2(P1_REG2_REG_16__SCAN_IN), .A(n14950), 
        .B(n14949), .ZN(n14951) );
  OAI21_X1 U16716 ( .B1(n15094), .B2(n14952), .A(n14951), .ZN(n14953) );
  AOI21_X1 U16717 ( .B1(n15097), .B2(n14993), .A(n14953), .ZN(n14954) );
  OAI21_X1 U16718 ( .B1(n14990), .B2(n15099), .A(n14954), .ZN(P1_U3277) );
  OAI21_X1 U16719 ( .B1(n14942), .B2(n14956), .A(n14955), .ZN(n15106) );
  NAND2_X1 U16720 ( .A1(n15110), .A2(n14957), .ZN(n14958) );
  XOR2_X1 U16721 ( .A(n14959), .B(n14958), .Z(n15100) );
  NAND2_X1 U16722 ( .A1(n15100), .A2(n14992), .ZN(n14969) );
  AOI211_X1 U16723 ( .C1(n15103), .C2(n14961), .A(n15344), .B(n14960), .ZN(
        n15101) );
  INV_X1 U16724 ( .A(n15102), .ZN(n14963) );
  OAI22_X1 U16725 ( .A1(n15336), .A2(n14963), .B1(n14962), .B2(n14997), .ZN(
        n14964) );
  AOI21_X1 U16726 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n15336), .A(n14964), 
        .ZN(n14965) );
  OAI21_X1 U16727 ( .B1(n14966), .B2(n15311), .A(n14965), .ZN(n14967) );
  AOI21_X1 U16728 ( .B1(n15101), .B2(n15332), .A(n14967), .ZN(n14968) );
  OAI211_X1 U16729 ( .C1(n15106), .C2(n14970), .A(n14969), .B(n14968), .ZN(
        P1_U3278) );
  XNOR2_X1 U16730 ( .A(n14971), .B(n7695), .ZN(n15119) );
  INV_X1 U16731 ( .A(n14973), .ZN(n14974) );
  AOI211_X1 U16732 ( .C1(n15116), .C2(n7768), .A(n15344), .B(n14974), .ZN(
        n15114) );
  AOI22_X1 U16733 ( .A1(n15336), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n14975), 
        .B2(n15324), .ZN(n14976) );
  OAI21_X1 U16734 ( .B1(n14977), .B2(n15311), .A(n14976), .ZN(n14988) );
  OAI211_X1 U16735 ( .C1(n7695), .C2(n14979), .A(n14978), .B(n15359), .ZN(
        n15118) );
  OR2_X1 U16736 ( .A1(n14981), .A2(n14980), .ZN(n14985) );
  NAND2_X1 U16737 ( .A1(n14983), .A2(n14982), .ZN(n14984) );
  NAND2_X1 U16738 ( .A1(n14985), .A2(n14984), .ZN(n15115) );
  INV_X1 U16739 ( .A(n15115), .ZN(n14986) );
  AOI21_X1 U16740 ( .B1(n15118), .B2(n14986), .A(n15336), .ZN(n14987) );
  AOI211_X1 U16741 ( .C1(n15114), .C2(n15332), .A(n14988), .B(n14987), .ZN(
        n14989) );
  OAI21_X1 U16742 ( .B1(n14990), .B2(n15119), .A(n14989), .ZN(P1_U3280) );
  OAI21_X1 U16743 ( .B1(n14993), .B2(n14992), .A(n14991), .ZN(n15002) );
  OAI21_X1 U16744 ( .B1(n14996), .B2(n14995), .A(n14994), .ZN(n15001) );
  INV_X1 U16745 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n15681) );
  OAI22_X1 U16746 ( .A1(n15336), .A2(n14998), .B1(n15681), .B2(n14997), .ZN(
        n14999) );
  AOI21_X1 U16747 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n15336), .A(n14999), .ZN(
        n15000) );
  NAND3_X1 U16748 ( .A1(n15002), .A2(n15001), .A3(n15000), .ZN(P1_U3293) );
  OAI211_X1 U16749 ( .C1(n15004), .C2(n15406), .A(n15003), .B(n15007), .ZN(
        n15131) );
  MUX2_X1 U16750 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15131), .S(n15443), .Z(
        P1_U3559) );
  OAI211_X1 U16751 ( .C1(n15009), .C2(n15406), .A(n15008), .B(n15007), .ZN(
        n15132) );
  MUX2_X1 U16752 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15132), .S(n15443), .Z(
        P1_U3558) );
  OAI211_X1 U16753 ( .C1(n15012), .C2(n15406), .A(n15011), .B(n15010), .ZN(
        n15013) );
  NAND3_X1 U16754 ( .A1(n15019), .A2(n15018), .A3(n15402), .ZN(n15024) );
  OAI22_X1 U16755 ( .A1(n15021), .A2(n15344), .B1(n15020), .B2(n15406), .ZN(
        n15022) );
  INV_X1 U16756 ( .A(n15022), .ZN(n15023) );
  NAND3_X1 U16757 ( .A1(n7927), .A2(n15024), .A3(n15023), .ZN(n15134) );
  MUX2_X1 U16758 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15134), .S(n15443), .Z(
        P1_U3556) );
  AOI21_X1 U16759 ( .B1(n15418), .B2(n15027), .A(n15026), .ZN(n15028) );
  NAND3_X1 U16760 ( .A1(n7936), .A2(n15029), .A3(n15028), .ZN(n15135) );
  MUX2_X1 U16761 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15135), .S(n15443), .Z(
        P1_U3555) );
  NAND2_X1 U16762 ( .A1(n15030), .A2(n15359), .ZN(n15035) );
  AOI211_X1 U16763 ( .C1(n15418), .C2(n15033), .A(n15032), .B(n15031), .ZN(
        n15034) );
  OAI211_X1 U16764 ( .C1(n15422), .C2(n15036), .A(n15035), .B(n15034), .ZN(
        n15136) );
  MUX2_X1 U16765 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15136), .S(n15443), .Z(
        P1_U3554) );
  INV_X1 U16766 ( .A(n15037), .ZN(n15042) );
  OAI211_X1 U16767 ( .C1(n15040), .C2(n15406), .A(n15039), .B(n15038), .ZN(
        n15041) );
  AOI21_X1 U16768 ( .B1(n15042), .B2(n15402), .A(n15041), .ZN(n15043) );
  OAI21_X1 U16769 ( .B1(n15044), .B2(n15400), .A(n15043), .ZN(n15137) );
  MUX2_X1 U16770 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15137), .S(n15443), .Z(
        P1_U3553) );
  AOI21_X1 U16771 ( .B1(n15418), .B2(n15046), .A(n15045), .ZN(n15047) );
  OAI211_X1 U16772 ( .C1(n15422), .C2(n15049), .A(n15048), .B(n15047), .ZN(
        n15138) );
  MUX2_X1 U16773 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15138), .S(n15443), .Z(
        P1_U3552) );
  INV_X1 U16774 ( .A(n15050), .ZN(n15052) );
  AOI22_X1 U16775 ( .A1(n15052), .A2(n15328), .B1(n15418), .B2(n15051), .ZN(
        n15055) );
  NAND3_X1 U16776 ( .A1(n15053), .A2(n15402), .A3(n14844), .ZN(n15054) );
  NAND3_X1 U16777 ( .A1(n15056), .A2(n15055), .A3(n15054), .ZN(n15139) );
  MUX2_X1 U16778 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15139), .S(n15443), .Z(
        P1_U3551) );
  OAI21_X1 U16779 ( .B1(n15058), .B2(n15406), .A(n15057), .ZN(n15059) );
  AOI211_X1 U16780 ( .C1(n15061), .C2(n15359), .A(n15060), .B(n15059), .ZN(
        n15062) );
  OAI21_X1 U16781 ( .B1(n15063), .B2(n15422), .A(n15062), .ZN(n15140) );
  MUX2_X1 U16782 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15140), .S(n15443), .Z(
        P1_U3550) );
  AOI211_X1 U16783 ( .C1(n15418), .C2(n15066), .A(n15065), .B(n15064), .ZN(
        n15067) );
  OAI21_X1 U16784 ( .B1(n15422), .B2(n15068), .A(n15067), .ZN(n15141) );
  MUX2_X1 U16785 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15141), .S(n15443), .Z(
        P1_U3549) );
  OAI211_X1 U16786 ( .C1(n15071), .C2(n15406), .A(n15070), .B(n15069), .ZN(
        n15072) );
  AOI21_X1 U16787 ( .B1(n15073), .B2(n15359), .A(n15072), .ZN(n15074) );
  OAI21_X1 U16788 ( .B1(n15422), .B2(n15075), .A(n15074), .ZN(n15142) );
  MUX2_X1 U16789 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15142), .S(n15443), .Z(
        P1_U3548) );
  AOI22_X1 U16790 ( .A1(n15077), .A2(n15328), .B1(n15418), .B2(n15076), .ZN(
        n15078) );
  OAI211_X1 U16791 ( .C1(n15422), .C2(n15080), .A(n15079), .B(n15078), .ZN(
        n15143) );
  INV_X2 U16792 ( .A(n15440), .ZN(n15443) );
  MUX2_X1 U16793 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15143), .S(n15443), .Z(
        P1_U3547) );
  AOI211_X1 U16794 ( .C1(n15418), .C2(n15083), .A(n15082), .B(n15081), .ZN(
        n15084) );
  OAI21_X1 U16795 ( .B1(n15422), .B2(n15085), .A(n15084), .ZN(n15144) );
  MUX2_X1 U16796 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15144), .S(n15443), .Z(
        P1_U3546) );
  AOI211_X1 U16797 ( .C1(n15418), .C2(n15088), .A(n15087), .B(n15086), .ZN(
        n15091) );
  NAND2_X1 U16798 ( .A1(n15089), .A2(n15402), .ZN(n15090) );
  OAI211_X1 U16799 ( .C1(n15400), .C2(n15092), .A(n15091), .B(n15090), .ZN(
        n15145) );
  MUX2_X1 U16800 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15145), .S(n15443), .Z(
        P1_U3545) );
  OAI211_X1 U16801 ( .C1(n15095), .C2(n15406), .A(n15094), .B(n15093), .ZN(
        n15096) );
  AOI21_X1 U16802 ( .B1(n15097), .B2(n15359), .A(n15096), .ZN(n15098) );
  OAI21_X1 U16803 ( .B1(n15422), .B2(n15099), .A(n15098), .ZN(n15146) );
  MUX2_X1 U16804 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15146), .S(n15443), .Z(
        P1_U3544) );
  NAND2_X1 U16805 ( .A1(n15100), .A2(n15402), .ZN(n15105) );
  AOI211_X1 U16806 ( .C1(n15418), .C2(n15103), .A(n15102), .B(n15101), .ZN(
        n15104) );
  OAI211_X1 U16807 ( .C1(n15400), .C2(n15106), .A(n15105), .B(n15104), .ZN(
        n15147) );
  MUX2_X1 U16808 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15147), .S(n15443), .Z(
        P1_U3543) );
  AOI22_X1 U16809 ( .A1(n15108), .A2(n15328), .B1(n15418), .B2(n15107), .ZN(
        n15112) );
  NAND3_X1 U16810 ( .A1(n15110), .A2(n15109), .A3(n15402), .ZN(n15111) );
  NAND3_X1 U16811 ( .A1(n15113), .A2(n15112), .A3(n15111), .ZN(n15148) );
  MUX2_X1 U16812 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15148), .S(n15443), .Z(
        P1_U3542) );
  AOI211_X1 U16813 ( .C1(n15418), .C2(n15116), .A(n15115), .B(n15114), .ZN(
        n15117) );
  OAI211_X1 U16814 ( .C1(n15422), .C2(n15119), .A(n15118), .B(n15117), .ZN(
        n15150) );
  MUX2_X1 U16815 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n15150), .S(n15443), .Z(
        P1_U3541) );
  AOI21_X1 U16816 ( .B1(n15418), .B2(n15121), .A(n15120), .ZN(n15122) );
  OAI211_X1 U16817 ( .C1(n15422), .C2(n15124), .A(n15123), .B(n15122), .ZN(
        n15151) );
  MUX2_X1 U16818 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n15151), .S(n15443), .Z(
        P1_U3540) );
  AOI21_X1 U16819 ( .B1(n15418), .B2(n15126), .A(n15125), .ZN(n15127) );
  OAI211_X1 U16820 ( .C1(n15422), .C2(n15129), .A(n15128), .B(n15127), .ZN(
        n15152) );
  MUX2_X1 U16821 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n15152), .S(n15443), .Z(
        P1_U3539) );
  MUX2_X1 U16822 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n15130), .S(n15443), .Z(
        P1_U3528) );
  MUX2_X1 U16823 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15131), .S(n15149), .Z(
        P1_U3527) );
  MUX2_X1 U16824 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15132), .S(n15425), .Z(
        P1_U3526) );
  MUX2_X1 U16825 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n15133), .S(n15425), .Z(
        P1_U3525) );
  MUX2_X1 U16826 ( .A(n15134), .B(P1_REG0_REG_28__SCAN_IN), .S(n15424), .Z(
        P1_U3524) );
  MUX2_X1 U16827 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15135), .S(n15425), .Z(
        P1_U3523) );
  MUX2_X1 U16828 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15136), .S(n15425), .Z(
        P1_U3522) );
  MUX2_X1 U16829 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15137), .S(n15425), .Z(
        P1_U3521) );
  MUX2_X1 U16830 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15138), .S(n15425), .Z(
        P1_U3520) );
  MUX2_X1 U16831 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15139), .S(n15425), .Z(
        P1_U3519) );
  MUX2_X1 U16832 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15140), .S(n15425), .Z(
        P1_U3518) );
  MUX2_X1 U16833 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15141), .S(n15425), .Z(
        P1_U3517) );
  MUX2_X1 U16834 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15142), .S(n15425), .Z(
        P1_U3516) );
  MUX2_X1 U16835 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15143), .S(n15149), .Z(
        P1_U3515) );
  MUX2_X1 U16836 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15144), .S(n15149), .Z(
        P1_U3513) );
  MUX2_X1 U16837 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15145), .S(n15149), .Z(
        P1_U3510) );
  MUX2_X1 U16838 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15146), .S(n15149), .Z(
        P1_U3507) );
  MUX2_X1 U16839 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15147), .S(n15149), .Z(
        P1_U3504) );
  MUX2_X1 U16840 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15148), .S(n15149), .Z(
        P1_U3501) );
  MUX2_X1 U16841 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n15150), .S(n15149), .Z(
        P1_U3498) );
  MUX2_X1 U16842 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n15151), .S(n15425), .Z(
        P1_U3495) );
  MUX2_X1 U16843 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n15152), .S(n15425), .Z(
        P1_U3492) );
  NOR4_X1 U16844 ( .A1(n9347), .A2(P1_IR_REG_30__SCAN_IN), .A3(n15153), .A4(
        P1_U3086), .ZN(n15154) );
  AOI21_X1 U16845 ( .B1(n15155), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n15154), 
        .ZN(n15156) );
  OAI21_X1 U16846 ( .B1(n15157), .B2(n15169), .A(n15156), .ZN(P1_U3324) );
  OAI222_X1 U16847 ( .A1(n15169), .A2(n15160), .B1(n15164), .B2(n15159), .C1(
        P1_U3086), .C2(n15158), .ZN(P1_U3325) );
  OAI222_X1 U16848 ( .A1(n15164), .A2(n15163), .B1(P1_U3086), .B2(n15162), 
        .C1(n15169), .C2(n15161), .ZN(P1_U3326) );
  OAI222_X1 U16849 ( .A1(n15167), .A2(P1_U3086), .B1(n15169), .B2(n15166), 
        .C1(n15165), .C2(n15164), .ZN(P1_U3327) );
  OAI222_X1 U16850 ( .A1(n15171), .A2(P1_U3086), .B1(n15164), .B2(n15170), 
        .C1(n15169), .C2(n15168), .ZN(P1_U3329) );
  OAI222_X1 U16851 ( .A1(n15164), .A2(n15175), .B1(P1_U3086), .B2(n15173), 
        .C1(n15169), .C2(n15172), .ZN(P1_U3330) );
  MUX2_X1 U16852 ( .A(n15177), .B(n15176), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  MUX2_X1 U16853 ( .A(n15178), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XOR2_X1 U16854 ( .A(n15179), .B(n15180), .Z(SUB_1596_U57) );
  XOR2_X1 U16855 ( .A(n15181), .B(n15182), .Z(SUB_1596_U56) );
  XOR2_X1 U16856 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n15183), .Z(SUB_1596_U54) );
  NAND2_X1 U16857 ( .A1(n15187), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n15188) );
  NAND2_X1 U16858 ( .A1(n15189), .A2(n15188), .ZN(n15192) );
  INV_X1 U16859 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n15190) );
  NAND2_X1 U16860 ( .A1(n15190), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n15191) );
  NAND2_X1 U16861 ( .A1(n15192), .A2(n15191), .ZN(n15201) );
  XNOR2_X1 U16862 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n15200) );
  INV_X1 U16863 ( .A(n15200), .ZN(n15193) );
  XNOR2_X1 U16864 ( .A(n15201), .B(n15193), .ZN(n15194) );
  XNOR2_X1 U16865 ( .A(n15196), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  NAND2_X1 U16866 ( .A1(n15201), .A2(n15200), .ZN(n15203) );
  NAND2_X1 U16867 ( .A1(n11345), .A2(P3_ADDR_REG_14__SCAN_IN), .ZN(n15202) );
  NAND2_X1 U16868 ( .A1(n15203), .A2(n15202), .ZN(n15216) );
  XNOR2_X1 U16869 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n15204) );
  XNOR2_X1 U16870 ( .A(n15216), .B(n15204), .ZN(n15208) );
  INV_X1 U16871 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15209) );
  XNOR2_X1 U16872 ( .A(n15208), .B(n15209), .ZN(n15205) );
  XNOR2_X1 U16873 ( .A(n15207), .B(n15205), .ZN(SUB_1596_U65) );
  NAND2_X1 U16874 ( .A1(n15208), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n15206) );
  INV_X1 U16875 ( .A(n15208), .ZN(n15210) );
  NAND2_X1 U16876 ( .A1(n15210), .A2(n15209), .ZN(n15211) );
  NAND2_X1 U16877 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n15213), .ZN(n15215) );
  NOR2_X1 U16878 ( .A1(n15213), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n15214) );
  AOI21_X1 U16879 ( .B1(n15216), .B2(n15215), .A(n15214), .ZN(n15229) );
  INV_X1 U16880 ( .A(n15229), .ZN(n15219) );
  AND2_X1 U16881 ( .A1(n15226), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n15227) );
  INV_X1 U16882 ( .A(n15227), .ZN(n15217) );
  OAI21_X1 U16883 ( .B1(n15226), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n15217), 
        .ZN(n15218) );
  XNOR2_X1 U16884 ( .A(n15219), .B(n15218), .ZN(n15220) );
  NAND2_X1 U16885 ( .A1(n15224), .A2(n15225), .ZN(n15222) );
  XNOR2_X1 U16886 ( .A(n15222), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  INV_X1 U16887 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15223) );
  OR2_X1 U16888 ( .A1(n15226), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n15228) );
  AOI21_X1 U16889 ( .B1(n15229), .B2(n15228), .A(n15227), .ZN(n15242) );
  XNOR2_X1 U16890 ( .A(n15242), .B(P1_ADDR_REG_17__SCAN_IN), .ZN(n15240) );
  INV_X1 U16891 ( .A(n15240), .ZN(n15230) );
  XNOR2_X1 U16892 ( .A(n15230), .B(P3_ADDR_REG_17__SCAN_IN), .ZN(n15231) );
  NAND2_X1 U16893 ( .A1(n15232), .A2(n15231), .ZN(n15238) );
  INV_X1 U16894 ( .A(n15238), .ZN(n15237) );
  INV_X1 U16895 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15233) );
  INV_X1 U16896 ( .A(n15234), .ZN(n15235) );
  OAI21_X1 U16897 ( .B1(n15235), .B2(n15237), .A(P2_ADDR_REG_17__SCAN_IN), 
        .ZN(n15236) );
  OAI21_X1 U16898 ( .B1(n15237), .B2(n15239), .A(n15236), .ZN(SUB_1596_U63) );
  NAND2_X1 U16899 ( .A1(n15240), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n15244) );
  INV_X1 U16900 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n15241) );
  NAND2_X1 U16901 ( .A1(n15242), .A2(n15241), .ZN(n15243) );
  NAND2_X1 U16902 ( .A1(n15244), .A2(n15243), .ZN(n15250) );
  XNOR2_X1 U16903 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n15251) );
  INV_X1 U16904 ( .A(n15251), .ZN(n15245) );
  AOI21_X1 U16905 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n15247), .A(n15249), 
        .ZN(n15248) );
  INV_X1 U16906 ( .A(n15248), .ZN(SUB_1596_U62) );
  NOR2_X1 U16907 ( .A1(n15249), .A2(n6527), .ZN(n15258) );
  INV_X1 U16908 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15253) );
  NAND2_X1 U16909 ( .A1(n15251), .A2(n15250), .ZN(n15252) );
  OAI21_X1 U16910 ( .B1(n15253), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n15252), 
        .ZN(n15256) );
  XNOR2_X1 U16911 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n15254) );
  XNOR2_X1 U16912 ( .A(n15254), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n15255) );
  XNOR2_X1 U16913 ( .A(n15256), .B(n15255), .ZN(n15257) );
  XNOR2_X1 U16914 ( .A(n15258), .B(n15257), .ZN(SUB_1596_U4) );
  AOI21_X1 U16915 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15259) );
  OAI21_X1 U16916 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n15259), 
        .ZN(U28) );
  AOI21_X1 U16917 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n15260) );
  OAI21_X1 U16918 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n15260), 
        .ZN(U29) );
  AND2_X1 U16919 ( .A1(n15262), .A2(n15261), .ZN(n15263) );
  XOR2_X1 U16920 ( .A(n15263), .B(P2_ADDR_REG_2__SCAN_IN), .Z(SUB_1596_U61) );
  INV_X1 U16921 ( .A(n15264), .ZN(n15269) );
  NAND3_X1 U16922 ( .A1(n15267), .A2(n15266), .A3(n15265), .ZN(n15268) );
  NAND3_X1 U16923 ( .A1(n15270), .A2(n15269), .A3(n15268), .ZN(n15282) );
  MUX2_X1 U16924 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10467), .S(n15271), .Z(
        n15272) );
  NAND3_X1 U16925 ( .A1(n15274), .A2(n15273), .A3(n15272), .ZN(n15275) );
  NAND3_X1 U16926 ( .A1(n15277), .A2(n15276), .A3(n15275), .ZN(n15281) );
  NAND2_X1 U16927 ( .A1(n15279), .A2(n15278), .ZN(n15280) );
  AND4_X1 U16928 ( .A1(n15283), .A2(n15282), .A3(n15281), .A4(n15280), .ZN(
        n15285) );
  OAI211_X1 U16929 ( .C1(n15287), .C2(n15286), .A(n15285), .B(n15284), .ZN(
        P1_U3247) );
  INV_X1 U16930 ( .A(n15305), .ZN(n15386) );
  INV_X1 U16931 ( .A(n15288), .ZN(n15292) );
  NAND2_X1 U16932 ( .A1(n15290), .A2(n15289), .ZN(n15291) );
  AOI21_X1 U16933 ( .B1(n15292), .B2(n15291), .A(n15400), .ZN(n15293) );
  AOI211_X1 U16934 ( .C1(n15386), .C2(n15411), .A(n15294), .B(n15293), .ZN(
        n15408) );
  AOI22_X1 U16935 ( .A1(n15336), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n15295), 
        .B2(n15324), .ZN(n15296) );
  OAI21_X1 U16936 ( .B1(n15311), .B2(n15407), .A(n15296), .ZN(n15297) );
  INV_X1 U16937 ( .A(n15297), .ZN(n15301) );
  OAI211_X1 U16938 ( .C1(n6478), .C2(n15407), .A(n15328), .B(n15298), .ZN(
        n15405) );
  INV_X1 U16939 ( .A(n15405), .ZN(n15299) );
  AOI22_X1 U16940 ( .A1(n15411), .A2(n15333), .B1(n15332), .B2(n15299), .ZN(
        n15300) );
  OAI211_X1 U16941 ( .C1(n15336), .C2(n15408), .A(n15301), .B(n15300), .ZN(
        P1_U3284) );
  XNOR2_X1 U16942 ( .A(n15304), .B(n15302), .ZN(n15308) );
  XNOR2_X1 U16943 ( .A(n15304), .B(n15303), .ZN(n15392) );
  NOR2_X1 U16944 ( .A1(n15392), .A2(n15305), .ZN(n15306) );
  AOI211_X1 U16945 ( .C1(n15359), .C2(n15308), .A(n15307), .B(n15306), .ZN(
        n15391) );
  AOI22_X1 U16946 ( .A1(n15336), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n15309), 
        .B2(n15324), .ZN(n15310) );
  OAI21_X1 U16947 ( .B1(n15311), .B2(n7762), .A(n15310), .ZN(n15312) );
  INV_X1 U16948 ( .A(n15312), .ZN(n15317) );
  INV_X1 U16949 ( .A(n15392), .ZN(n15315) );
  AOI211_X1 U16950 ( .C1(n15389), .C2(n15314), .A(n15344), .B(n15313), .ZN(
        n15388) );
  AOI22_X1 U16951 ( .A1(n15315), .A2(n15333), .B1(n15332), .B2(n15388), .ZN(
        n15316) );
  OAI211_X1 U16952 ( .C1(n15336), .C2(n15391), .A(n15317), .B(n15316), .ZN(
        P1_U3286) );
  XNOR2_X1 U16953 ( .A(n15318), .B(n15320), .ZN(n15377) );
  XNOR2_X1 U16954 ( .A(n15319), .B(n15320), .ZN(n15321) );
  NOR2_X1 U16955 ( .A1(n15321), .A2(n15400), .ZN(n15322) );
  AOI211_X1 U16956 ( .C1(n15386), .C2(n15377), .A(n15323), .B(n15322), .ZN(
        n15374) );
  AOI22_X1 U16957 ( .A1(n15336), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n15325), 
        .B2(n15324), .ZN(n15326) );
  OAI21_X1 U16958 ( .B1(n15311), .B2(n15373), .A(n15326), .ZN(n15327) );
  INV_X1 U16959 ( .A(n15327), .ZN(n15335) );
  OAI211_X1 U16960 ( .C1(n15330), .C2(n15373), .A(n15329), .B(n15328), .ZN(
        n15372) );
  INV_X1 U16961 ( .A(n15372), .ZN(n15331) );
  AOI22_X1 U16962 ( .A1(n15377), .A2(n15333), .B1(n15332), .B2(n15331), .ZN(
        n15334) );
  OAI211_X1 U16963 ( .C1(n15336), .C2(n15374), .A(n15335), .B(n15334), .ZN(
        P1_U3288) );
  AND2_X1 U16964 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15338), .ZN(P1_U3294) );
  AND2_X1 U16965 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15338), .ZN(P1_U3295) );
  AND2_X1 U16966 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15338), .ZN(P1_U3296) );
  AND2_X1 U16967 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15338), .ZN(P1_U3297) );
  AND2_X1 U16968 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15338), .ZN(P1_U3298) );
  AND2_X1 U16969 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15338), .ZN(P1_U3299) );
  INV_X1 U16970 ( .A(n15338), .ZN(n15337) );
  INV_X1 U16971 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n15711) );
  NOR2_X1 U16972 ( .A1(n15337), .A2(n15711), .ZN(P1_U3300) );
  AND2_X1 U16973 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15338), .ZN(P1_U3301) );
  AND2_X1 U16974 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15338), .ZN(P1_U3302) );
  AND2_X1 U16975 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15338), .ZN(P1_U3303) );
  AND2_X1 U16976 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15338), .ZN(P1_U3304) );
  AND2_X1 U16977 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15338), .ZN(P1_U3305) );
  AND2_X1 U16978 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15338), .ZN(P1_U3306) );
  AND2_X1 U16979 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15338), .ZN(P1_U3307) );
  AND2_X1 U16980 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15338), .ZN(P1_U3308) );
  AND2_X1 U16981 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15338), .ZN(P1_U3309) );
  AND2_X1 U16982 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15338), .ZN(P1_U3310) );
  AND2_X1 U16983 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15338), .ZN(P1_U3311) );
  AND2_X1 U16984 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15338), .ZN(P1_U3312) );
  AND2_X1 U16985 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15338), .ZN(P1_U3313) );
  AND2_X1 U16986 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15338), .ZN(P1_U3314) );
  AND2_X1 U16987 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15338), .ZN(P1_U3315) );
  AND2_X1 U16988 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15338), .ZN(P1_U3316) );
  AND2_X1 U16989 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15338), .ZN(P1_U3317) );
  INV_X1 U16990 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n15735) );
  NOR2_X1 U16991 ( .A1(n15337), .A2(n15735), .ZN(P1_U3318) );
  AND2_X1 U16992 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15338), .ZN(P1_U3319) );
  AND2_X1 U16993 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15338), .ZN(P1_U3320) );
  AND2_X1 U16994 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15338), .ZN(P1_U3321) );
  AND2_X1 U16995 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15338), .ZN(P1_U3322) );
  AND2_X1 U16996 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15338), .ZN(P1_U3323) );
  INV_X1 U16997 ( .A(n15393), .ZN(n15412) );
  INV_X1 U16998 ( .A(n15339), .ZN(n15347) );
  AOI21_X1 U16999 ( .B1(n15418), .B2(n15341), .A(n15340), .ZN(n15342) );
  OAI21_X1 U17000 ( .B1(n15344), .B2(n15343), .A(n15342), .ZN(n15346) );
  AOI211_X1 U17001 ( .C1(n15412), .C2(n15347), .A(n15346), .B(n15345), .ZN(
        n15426) );
  AOI22_X1 U17002 ( .A1(n15425), .A2(n15426), .B1(n7005), .B2(n15424), .ZN(
        P1_U3462) );
  INV_X1 U17003 ( .A(n15353), .ZN(n15348) );
  NOR2_X1 U17004 ( .A1(n15348), .A2(n15393), .ZN(n15352) );
  OAI211_X1 U17005 ( .C1(n9891), .C2(n15406), .A(n15350), .B(n15349), .ZN(
        n15351) );
  AOI211_X1 U17006 ( .C1(n15386), .C2(n15353), .A(n15352), .B(n15351), .ZN(
        n15427) );
  INV_X1 U17007 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n15354) );
  AOI22_X1 U17008 ( .A1(n15425), .A2(n15427), .B1(n15354), .B2(n15424), .ZN(
        P1_U3465) );
  INV_X1 U17009 ( .A(n15362), .ZN(n15364) );
  OAI21_X1 U17010 ( .B1(n15356), .B2(n15406), .A(n15355), .ZN(n15358) );
  AOI211_X1 U17011 ( .C1(n15360), .C2(n15359), .A(n15358), .B(n15357), .ZN(
        n15361) );
  OAI21_X1 U17012 ( .B1(n15362), .B2(n15393), .A(n15361), .ZN(n15363) );
  AOI21_X1 U17013 ( .B1(n15386), .B2(n15364), .A(n15363), .ZN(n15428) );
  INV_X1 U17014 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n15365) );
  AOI22_X1 U17015 ( .A1(n15425), .A2(n15428), .B1(n15365), .B2(n15424), .ZN(
        P1_U3468) );
  OAI211_X1 U17016 ( .C1(n15368), .C2(n15406), .A(n15367), .B(n15366), .ZN(
        n15369) );
  AOI21_X1 U17017 ( .B1(n15370), .B2(n15402), .A(n15369), .ZN(n15430) );
  INV_X1 U17018 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n15371) );
  AOI22_X1 U17019 ( .A1(n15425), .A2(n15430), .B1(n15371), .B2(n15424), .ZN(
        P1_U3471) );
  OAI21_X1 U17020 ( .B1(n15373), .B2(n15406), .A(n15372), .ZN(n15376) );
  INV_X1 U17021 ( .A(n15374), .ZN(n15375) );
  AOI211_X1 U17022 ( .C1(n15412), .C2(n15377), .A(n15376), .B(n15375), .ZN(
        n15432) );
  INV_X1 U17023 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15378) );
  AOI22_X1 U17024 ( .A1(n15425), .A2(n15432), .B1(n15378), .B2(n15424), .ZN(
        P1_U3474) );
  INV_X1 U17025 ( .A(n15383), .ZN(n15385) );
  AOI21_X1 U17026 ( .B1(n15418), .B2(n15380), .A(n15379), .ZN(n15382) );
  OAI211_X1 U17027 ( .C1(n15383), .C2(n15393), .A(n15382), .B(n15381), .ZN(
        n15384) );
  AOI21_X1 U17028 ( .B1(n15386), .B2(n15385), .A(n15384), .ZN(n15434) );
  INV_X1 U17029 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n15387) );
  AOI22_X1 U17030 ( .A1(n15425), .A2(n15434), .B1(n15387), .B2(n15424), .ZN(
        P1_U3477) );
  AOI21_X1 U17031 ( .B1(n15418), .B2(n15389), .A(n15388), .ZN(n15390) );
  OAI211_X1 U17032 ( .C1(n15393), .C2(n15392), .A(n15391), .B(n15390), .ZN(
        n15394) );
  INV_X1 U17033 ( .A(n15394), .ZN(n15436) );
  AOI22_X1 U17034 ( .A1(n15425), .A2(n15436), .B1(n7183), .B2(n15424), .ZN(
        P1_U3480) );
  AOI211_X1 U17035 ( .C1(n15418), .C2(n15397), .A(n15396), .B(n15395), .ZN(
        n15398) );
  OAI21_X1 U17036 ( .B1(n15400), .B2(n15399), .A(n15398), .ZN(n15401) );
  AOI21_X1 U17037 ( .B1(n15403), .B2(n15402), .A(n15401), .ZN(n15437) );
  INV_X1 U17038 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15404) );
  AOI22_X1 U17039 ( .A1(n15425), .A2(n15437), .B1(n15404), .B2(n15424), .ZN(
        P1_U3483) );
  OAI21_X1 U17040 ( .B1(n15407), .B2(n15406), .A(n15405), .ZN(n15410) );
  INV_X1 U17041 ( .A(n15408), .ZN(n15409) );
  AOI211_X1 U17042 ( .C1(n15412), .C2(n15411), .A(n15410), .B(n15409), .ZN(
        n15439) );
  INV_X1 U17043 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15413) );
  AOI22_X1 U17044 ( .A1(n15425), .A2(n15439), .B1(n15413), .B2(n15424), .ZN(
        P1_U3486) );
  INV_X1 U17045 ( .A(n15414), .ZN(n15416) );
  AOI211_X1 U17046 ( .C1(n15418), .C2(n15417), .A(n15416), .B(n15415), .ZN(
        n15419) );
  OAI211_X1 U17047 ( .C1(n15422), .C2(n15421), .A(n15420), .B(n15419), .ZN(
        n15423) );
  INV_X1 U17048 ( .A(n15423), .ZN(n15442) );
  INV_X1 U17049 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n15790) );
  AOI22_X1 U17050 ( .A1(n15425), .A2(n15442), .B1(n15790), .B2(n15424), .ZN(
        P1_U3489) );
  AOI22_X1 U17051 ( .A1(n15443), .A2(n15426), .B1(n10446), .B2(n15440), .ZN(
        P1_U3529) );
  AOI22_X1 U17052 ( .A1(n15443), .A2(n15427), .B1(n10445), .B2(n15440), .ZN(
        P1_U3530) );
  AOI22_X1 U17053 ( .A1(n15443), .A2(n15428), .B1(n10449), .B2(n15440), .ZN(
        P1_U3531) );
  AOI22_X1 U17054 ( .A1(n15443), .A2(n15430), .B1(n15429), .B2(n15440), .ZN(
        P1_U3532) );
  AOI22_X1 U17055 ( .A1(n15443), .A2(n15432), .B1(n15431), .B2(n15440), .ZN(
        P1_U3533) );
  AOI22_X1 U17056 ( .A1(n15443), .A2(n15434), .B1(n15433), .B2(n15440), .ZN(
        P1_U3534) );
  AOI22_X1 U17057 ( .A1(n15443), .A2(n15436), .B1(n15435), .B2(n15440), .ZN(
        P1_U3535) );
  AOI22_X1 U17058 ( .A1(n15443), .A2(n15437), .B1(n10444), .B2(n15440), .ZN(
        P1_U3536) );
  AOI22_X1 U17059 ( .A1(n15443), .A2(n15439), .B1(n15438), .B2(n15440), .ZN(
        P1_U3537) );
  AOI22_X1 U17060 ( .A1(n15443), .A2(n15442), .B1(n15441), .B2(n15440), .ZN(
        P1_U3538) );
  NOR2_X1 U17061 ( .A1(n15468), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U17062 ( .A1(n15470), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n15475), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n15450) );
  AOI22_X1 U17063 ( .A1(n15468), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n15449) );
  OAI22_X1 U17064 ( .A1(n15445), .A2(P2_REG1_REG_0__SCAN_IN), .B1(
        P2_REG2_REG_0__SCAN_IN), .B2(n15444), .ZN(n15446) );
  OAI21_X1 U17065 ( .B1(n15447), .B2(n15446), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n15448) );
  OAI211_X1 U17066 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n15450), .A(n15449), .B(
        n15448), .ZN(P2_U3214) );
  OAI22_X1 U17067 ( .A1(n15465), .A2(n15452), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15451), .ZN(n15453) );
  AOI21_X1 U17068 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n15468), .A(n15453), .ZN(
        n15462) );
  OAI211_X1 U17069 ( .C1(n15456), .C2(n15455), .A(n15470), .B(n15454), .ZN(
        n15461) );
  OAI211_X1 U17070 ( .C1(n15459), .C2(n15458), .A(n15475), .B(n15457), .ZN(
        n15460) );
  NAND3_X1 U17071 ( .A1(n15462), .A2(n15461), .A3(n15460), .ZN(P2_U3217) );
  INV_X1 U17072 ( .A(n15463), .ZN(n15467) );
  NOR2_X1 U17073 ( .A1(n15465), .A2(n15464), .ZN(n15466) );
  AOI211_X1 U17074 ( .C1(n15468), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n15467), .B(
        n15466), .ZN(n15479) );
  OAI211_X1 U17075 ( .C1(n15472), .C2(n15471), .A(n15470), .B(n15469), .ZN(
        n15478) );
  XOR2_X1 U17076 ( .A(n15474), .B(n15473), .Z(n15476) );
  NAND2_X1 U17077 ( .A1(n15476), .A2(n15475), .ZN(n15477) );
  NAND3_X1 U17078 ( .A1(n15479), .A2(n15478), .A3(n15477), .ZN(P2_U3220) );
  INV_X1 U17079 ( .A(n15486), .ZN(n15489) );
  XNOR2_X1 U17080 ( .A(n15480), .B(n15489), .ZN(n15500) );
  INV_X1 U17081 ( .A(n15500), .ZN(n15542) );
  OAI211_X1 U17082 ( .C1(n7178), .C2(n15545), .A(n14181), .B(n15562), .ZN(
        n15539) );
  INV_X1 U17083 ( .A(n15539), .ZN(n15483) );
  AOI22_X1 U17084 ( .A1(n15542), .A2(n15835), .B1(n15484), .B2(n15483), .ZN(
        n15508) );
  NAND2_X1 U17085 ( .A1(n15486), .A2(n15485), .ZN(n15491) );
  NAND2_X1 U17086 ( .A1(n15488), .A2(n15487), .ZN(n15490) );
  NAND2_X1 U17087 ( .A1(n15490), .A2(n15489), .ZN(n15552) );
  OAI21_X1 U17088 ( .B1(n15492), .B2(n15491), .A(n15552), .ZN(n15498) );
  OAI22_X1 U17089 ( .A1(n15496), .A2(n15495), .B1(n15494), .B2(n15493), .ZN(
        n15497) );
  AOI21_X1 U17090 ( .B1(n15498), .B2(n15556), .A(n15497), .ZN(n15499) );
  OAI21_X1 U17091 ( .B1(n15501), .B2(n15500), .A(n15499), .ZN(n15540) );
  MUX2_X1 U17092 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n15540), .S(n15831), .Z(
        n15506) );
  OAI22_X1 U17093 ( .A1(n15504), .A2(n15545), .B1(n15503), .B2(n15502), .ZN(
        n15505) );
  NOR2_X1 U17094 ( .A1(n15506), .A2(n15505), .ZN(n15507) );
  NAND2_X1 U17095 ( .A1(n15508), .A2(n15507), .ZN(P2_U3261) );
  INV_X1 U17096 ( .A(n15517), .ZN(n15514) );
  NOR2_X1 U17097 ( .A1(n15514), .A2(n15509), .ZN(n15510) );
  AND2_X1 U17098 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15511), .ZN(P2_U3266) );
  AND2_X1 U17099 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15511), .ZN(P2_U3267) );
  INV_X1 U17100 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n15746) );
  NOR2_X1 U17101 ( .A1(n15510), .A2(n15746), .ZN(P2_U3268) );
  AND2_X1 U17102 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15511), .ZN(P2_U3269) );
  AND2_X1 U17103 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15511), .ZN(P2_U3270) );
  AND2_X1 U17104 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15511), .ZN(P2_U3271) );
  AND2_X1 U17105 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15511), .ZN(P2_U3272) );
  AND2_X1 U17106 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15511), .ZN(P2_U3273) );
  AND2_X1 U17107 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15511), .ZN(P2_U3274) );
  AND2_X1 U17108 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15511), .ZN(P2_U3275) );
  AND2_X1 U17109 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15511), .ZN(P2_U3276) );
  AND2_X1 U17110 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15511), .ZN(P2_U3277) );
  AND2_X1 U17111 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15511), .ZN(P2_U3278) );
  AND2_X1 U17112 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15511), .ZN(P2_U3279) );
  AND2_X1 U17113 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15511), .ZN(P2_U3280) );
  AND2_X1 U17114 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15511), .ZN(P2_U3281) );
  INV_X1 U17115 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n15810) );
  NOR2_X1 U17116 ( .A1(n15510), .A2(n15810), .ZN(P2_U3282) );
  AND2_X1 U17117 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15511), .ZN(P2_U3283) );
  AND2_X1 U17118 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15511), .ZN(P2_U3284) );
  AND2_X1 U17119 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15511), .ZN(P2_U3285) );
  AND2_X1 U17120 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15511), .ZN(P2_U3286) );
  AND2_X1 U17121 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15511), .ZN(P2_U3287) );
  AND2_X1 U17122 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15511), .ZN(P2_U3288) );
  AND2_X1 U17123 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15511), .ZN(P2_U3289) );
  AND2_X1 U17124 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15511), .ZN(P2_U3290) );
  AND2_X1 U17125 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15511), .ZN(P2_U3291) );
  AND2_X1 U17126 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15511), .ZN(P2_U3292) );
  AND2_X1 U17127 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15511), .ZN(P2_U3293) );
  AND2_X1 U17128 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15511), .ZN(P2_U3294) );
  AND2_X1 U17129 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15511), .ZN(P2_U3295) );
  AOI22_X1 U17130 ( .A1(n15517), .A2(n15513), .B1(n15512), .B2(n15514), .ZN(
        P2_U3416) );
  AOI22_X1 U17131 ( .A1(n15517), .A2(n15516), .B1(n15515), .B2(n15514), .ZN(
        P2_U3417) );
  OAI22_X1 U17132 ( .A1(n15519), .A2(n15528), .B1(n15518), .B2(n7237), .ZN(
        n15520) );
  OR2_X1 U17133 ( .A1(n15521), .A2(n15520), .ZN(n15572) );
  OAI22_X1 U17134 ( .A1(n15569), .A2(n15572), .B1(P2_REG0_REG_0__SCAN_IN), 
        .B2(n15571), .ZN(n15522) );
  INV_X1 U17135 ( .A(n15522), .ZN(P2_U3430) );
  AOI21_X1 U17136 ( .B1(n15525), .B2(n15524), .A(n15523), .ZN(n15526) );
  OAI211_X1 U17137 ( .C1(n15529), .C2(n15528), .A(n15527), .B(n15526), .ZN(
        n15530) );
  INV_X1 U17138 ( .A(n15530), .ZN(n15574) );
  INV_X1 U17139 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n15531) );
  AOI22_X1 U17140 ( .A1(n15571), .A2(n15574), .B1(n15531), .B2(n15569), .ZN(
        P2_U3433) );
  OAI21_X1 U17141 ( .B1(n15533), .B2(n15565), .A(n15532), .ZN(n15536) );
  INV_X1 U17142 ( .A(n15534), .ZN(n15535) );
  AOI211_X1 U17143 ( .C1(n15560), .C2(n15537), .A(n15536), .B(n15535), .ZN(
        n15575) );
  INV_X1 U17144 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15538) );
  AOI22_X1 U17145 ( .A1(n15571), .A2(n15575), .B1(n15538), .B2(n15569), .ZN(
        P2_U3436) );
  OAI21_X1 U17146 ( .B1(n15545), .B2(n15565), .A(n15539), .ZN(n15541) );
  AOI211_X1 U17147 ( .C1(n15560), .C2(n15542), .A(n15541), .B(n15540), .ZN(
        n15577) );
  INV_X1 U17148 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15543) );
  AOI22_X1 U17149 ( .A1(n15571), .A2(n15577), .B1(n15543), .B2(n15569), .ZN(
        P2_U3442) );
  OAI21_X1 U17150 ( .B1(n15480), .B2(n15545), .A(n15544), .ZN(n15547) );
  NAND2_X1 U17151 ( .A1(n15480), .A2(n15545), .ZN(n15546) );
  NAND2_X1 U17152 ( .A1(n15547), .A2(n15546), .ZN(n15549) );
  INV_X1 U17153 ( .A(n15553), .ZN(n15548) );
  XNOR2_X1 U17154 ( .A(n15549), .B(n15548), .ZN(n15836) );
  NAND2_X1 U17155 ( .A1(n15836), .A2(n15550), .ZN(n15559) );
  NAND2_X1 U17156 ( .A1(n15552), .A2(n15551), .ZN(n15554) );
  XNOR2_X1 U17157 ( .A(n15554), .B(n15553), .ZN(n15557) );
  AOI21_X1 U17158 ( .B1(n15557), .B2(n15556), .A(n15555), .ZN(n15558) );
  NAND2_X1 U17159 ( .A1(n15559), .A2(n15558), .ZN(n15832) );
  AND2_X1 U17160 ( .A1(n15836), .A2(n15560), .ZN(n15568) );
  AOI21_X1 U17161 ( .B1(n15562), .B2(n15826), .A(n15561), .ZN(n15564) );
  NAND2_X1 U17162 ( .A1(n15564), .A2(n15563), .ZN(n15830) );
  OAI21_X1 U17163 ( .B1(n15566), .B2(n15565), .A(n15830), .ZN(n15567) );
  NOR3_X1 U17164 ( .A1(n15832), .A2(n15568), .A3(n15567), .ZN(n15579) );
  INV_X1 U17165 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n15570) );
  AOI22_X1 U17166 ( .A1(n15571), .A2(n15579), .B1(n15570), .B2(n15569), .ZN(
        P2_U3445) );
  OAI22_X1 U17167 ( .A1(n15578), .A2(n15572), .B1(P2_REG1_REG_0__SCAN_IN), 
        .B2(n15580), .ZN(n15573) );
  INV_X1 U17168 ( .A(n15573), .ZN(P2_U3499) );
  AOI22_X1 U17169 ( .A1(n15580), .A2(n15574), .B1(n10567), .B2(n15578), .ZN(
        P2_U3500) );
  AOI22_X1 U17170 ( .A1(n15580), .A2(n15575), .B1(n10568), .B2(n15578), .ZN(
        P2_U3501) );
  AOI22_X1 U17171 ( .A1(n15580), .A2(n15577), .B1(n15576), .B2(n15578), .ZN(
        P2_U3503) );
  AOI22_X1 U17172 ( .A1(n15580), .A2(n15579), .B1(n10672), .B2(n15578), .ZN(
        P2_U3504) );
  NOR2_X1 U17173 ( .A1(P3_U3897), .A2(n15581), .ZN(P3_U3150) );
  INV_X1 U17174 ( .A(n15582), .ZN(n15598) );
  XNOR2_X1 U17175 ( .A(n15584), .B(n15583), .ZN(n15596) );
  INV_X1 U17176 ( .A(n15596), .ZN(n15614) );
  AND2_X1 U17177 ( .A1(n15585), .A2(n15637), .ZN(n15613) );
  NAND2_X1 U17178 ( .A1(n15613), .A2(n15586), .ZN(n15587) );
  OAI21_X1 U17179 ( .B1(n15588), .B2(n10900), .A(n15587), .ZN(n15597) );
  XNOR2_X1 U17180 ( .A(n15590), .B(n15589), .ZN(n15594) );
  OAI22_X1 U17181 ( .A1(n15592), .A2(n15652), .B1(n15591), .B2(n15642), .ZN(
        n15593) );
  AOI21_X1 U17182 ( .B1(n15594), .B2(n15611), .A(n15593), .ZN(n15595) );
  OAI21_X1 U17183 ( .B1(n15644), .B2(n15596), .A(n15595), .ZN(n15612) );
  AOI211_X1 U17184 ( .C1(n15598), .C2(n15614), .A(n15597), .B(n15612), .ZN(
        n15600) );
  AOI22_X1 U17185 ( .A1(n15601), .A2(n10203), .B1(n15600), .B2(n15599), .ZN(
        P3_U3231) );
  NAND2_X1 U17186 ( .A1(n15603), .A2(n15602), .ZN(n15607) );
  AOI21_X1 U17187 ( .B1(n15638), .B2(n15605), .A(n15604), .ZN(n15606) );
  OAI211_X1 U17188 ( .C1(n15608), .C2(n15642), .A(n15607), .B(n15606), .ZN(
        n15609) );
  AOI21_X1 U17189 ( .B1(n15611), .B2(n15610), .A(n15609), .ZN(n15667) );
  AOI22_X1 U17190 ( .A1(n15666), .A2(n15667), .B1(n8832), .B2(n15664), .ZN(
        P3_U3393) );
  AOI211_X1 U17191 ( .C1(n15648), .C2(n15614), .A(n15613), .B(n15612), .ZN(
        n15668) );
  AOI22_X1 U17192 ( .A1(n15666), .A2(n15668), .B1(n8839), .B2(n15664), .ZN(
        P3_U3396) );
  AOI22_X1 U17193 ( .A1(n15616), .A2(n15648), .B1(n15615), .B2(n15637), .ZN(
        n15617) );
  AND2_X1 U17194 ( .A1(n15618), .A2(n15617), .ZN(n15669) );
  AOI22_X1 U17195 ( .A1(n15666), .A2(n15669), .B1(n8852), .B2(n15664), .ZN(
        P3_U3399) );
  AOI22_X1 U17196 ( .A1(n15620), .A2(n15638), .B1(n15637), .B2(n15619), .ZN(
        n15621) );
  OAI211_X1 U17197 ( .C1(n15623), .C2(n15642), .A(n15622), .B(n15621), .ZN(
        n15626) );
  AOI21_X1 U17198 ( .B1(n15644), .B2(n15659), .A(n15624), .ZN(n15625) );
  NOR2_X1 U17199 ( .A1(n15626), .A2(n15625), .ZN(n15670) );
  AOI22_X1 U17200 ( .A1(n15666), .A2(n15670), .B1(n8866), .B2(n15664), .ZN(
        P3_U3402) );
  INV_X1 U17201 ( .A(n15633), .ZN(n15635) );
  OAI22_X1 U17202 ( .A1(n15628), .A2(n15652), .B1(n15651), .B2(n15627), .ZN(
        n15629) );
  AOI21_X1 U17203 ( .B1(n15656), .B2(n15630), .A(n15629), .ZN(n15632) );
  OAI211_X1 U17204 ( .C1(n15633), .C2(n15659), .A(n15632), .B(n15631), .ZN(
        n15634) );
  AOI21_X1 U17205 ( .B1(n15635), .B2(n15662), .A(n15634), .ZN(n15671) );
  AOI22_X1 U17206 ( .A1(n15666), .A2(n15671), .B1(n8881), .B2(n15664), .ZN(
        P3_U3405) );
  INV_X1 U17207 ( .A(n15645), .ZN(n15649) );
  AOI22_X1 U17208 ( .A1(n15639), .A2(n15638), .B1(n15637), .B2(n15636), .ZN(
        n15640) );
  OAI211_X1 U17209 ( .C1(n15643), .C2(n15642), .A(n15641), .B(n15640), .ZN(
        n15647) );
  NOR2_X1 U17210 ( .A1(n15645), .A2(n15644), .ZN(n15646) );
  AOI211_X1 U17211 ( .C1(n15649), .C2(n15648), .A(n15647), .B(n15646), .ZN(
        n15673) );
  AOI22_X1 U17212 ( .A1(n15666), .A2(n15673), .B1(n8900), .B2(n15664), .ZN(
        P3_U3408) );
  INV_X1 U17213 ( .A(n15660), .ZN(n15663) );
  OAI22_X1 U17214 ( .A1(n15653), .A2(n15652), .B1(n15651), .B2(n15650), .ZN(
        n15654) );
  AOI21_X1 U17215 ( .B1(n15656), .B2(n15655), .A(n15654), .ZN(n15658) );
  OAI211_X1 U17216 ( .C1(n15660), .C2(n15659), .A(n15658), .B(n15657), .ZN(
        n15661) );
  AOI21_X1 U17217 ( .B1(n15663), .B2(n15662), .A(n15661), .ZN(n15675) );
  INV_X1 U17218 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15665) );
  AOI22_X1 U17219 ( .A1(n15666), .A2(n15675), .B1(n15665), .B2(n15664), .ZN(
        P3_U3411) );
  AOI22_X1 U17220 ( .A1(n15676), .A2(n15667), .B1(n10955), .B2(n15674), .ZN(
        P3_U3460) );
  AOI22_X1 U17221 ( .A1(n15676), .A2(n15668), .B1(n10173), .B2(n15674), .ZN(
        P3_U3461) );
  AOI22_X1 U17222 ( .A1(n15676), .A2(n15669), .B1(n10793), .B2(n15674), .ZN(
        P3_U3462) );
  AOI22_X1 U17223 ( .A1(n15676), .A2(n15670), .B1(n10180), .B2(n15674), .ZN(
        P3_U3463) );
  AOI22_X1 U17224 ( .A1(n15676), .A2(n15671), .B1(n10214), .B2(n15674), .ZN(
        P3_U3464) );
  AOI22_X1 U17225 ( .A1(n15676), .A2(n15673), .B1(n15672), .B2(n15674), .ZN(
        P3_U3465) );
  AOI22_X1 U17226 ( .A1(n15676), .A2(n15675), .B1(n10181), .B2(n15674), .ZN(
        P3_U3466) );
  NAND4_X1 U17227 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P1_REG3_REG_19__SCAN_IN), .A4(P1_REG1_REG_7__SCAN_IN), .ZN(n15685) );
  NAND4_X1 U17228 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(n15733), .A3(n15677), .A4(
        n15747), .ZN(n15678) );
  NOR2_X1 U17229 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(n15678), .ZN(n15682) );
  NAND4_X1 U17230 ( .A1(n15682), .A2(n15681), .A3(n15680), .A4(n15679), .ZN(
        n15684) );
  NAND4_X1 U17231 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .A3(
        P3_REG1_REG_0__SCAN_IN), .A4(P1_REG2_REG_28__SCAN_IN), .ZN(n15683) );
  NOR3_X1 U17232 ( .A1(n15685), .A2(n15684), .A3(n15683), .ZN(n15823) );
  INV_X1 U17233 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n15714) );
  NAND4_X1 U17234 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(n15714), .A3(n15705), .A4(
        n15704), .ZN(n15701) );
  NAND4_X1 U17235 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(P1_B_REG_SCAN_IN), .A3(
        n15703), .A4(n15719), .ZN(n15700) );
  NAND4_X1 U17236 ( .A1(n15687), .A2(n15686), .A3(P1_ADDR_REG_5__SCAN_IN), 
        .A4(n15731), .ZN(n15699) );
  NOR4_X1 U17237 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P2_RD_REG_SCAN_IN), .A4(n15774), .ZN(n15697) );
  NAND4_X1 U17238 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(n15776), .A3(n15766), .A4(
        n15778), .ZN(n15689) );
  NAND4_X1 U17239 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), 
        .A3(P1_REG3_REG_9__SCAN_IN), .A4(P1_REG2_REG_16__SCAN_IN), .ZN(n15688)
         );
  OR4_X1 U17240 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(n15689), .A3(n15688), .A4(
        P2_REG2_REG_6__SCAN_IN), .ZN(n15690) );
  NOR3_X1 U17241 ( .A1(n15690), .A2(P3_REG3_REG_0__SCAN_IN), .A3(
        P2_REG3_REG_12__SCAN_IN), .ZN(n15696) );
  INV_X1 U17242 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n15788) );
  NOR4_X1 U17243 ( .A1(P1_REG0_REG_10__SCAN_IN), .A2(P3_IR_REG_29__SCAN_IN), 
        .A3(P1_REG3_REG_1__SCAN_IN), .A4(n15788), .ZN(n15695) );
  NAND4_X1 U17244 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), 
        .A3(P3_DATAO_REG_23__SCAN_IN), .A4(n15763), .ZN(n15693) );
  INV_X1 U17245 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n15811) );
  NAND4_X1 U17246 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .A3(P2_IR_REG_29__SCAN_IN), .A4(n15811), .ZN(n15692) );
  NAND3_X1 U17247 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P1_REG1_REG_26__SCAN_IN), 
        .A3(n8912), .ZN(n15691) );
  NOR4_X1 U17248 ( .A1(P3_REG3_REG_20__SCAN_IN), .A2(n15693), .A3(n15692), 
        .A4(n15691), .ZN(n15694) );
  NAND4_X1 U17249 ( .A1(n15697), .A2(n15696), .A3(n15695), .A4(n15694), .ZN(
        n15698) );
  NOR4_X1 U17250 ( .A1(n15701), .A2(n15700), .A3(n15699), .A4(n15698), .ZN(
        n15822) );
  AOI22_X1 U17251 ( .A1(n15704), .A2(keyinput35), .B1(n15703), .B2(keyinput36), 
        .ZN(n15702) );
  OAI221_X1 U17252 ( .B1(n15704), .B2(keyinput35), .C1(n15703), .C2(keyinput36), .A(n15702), .ZN(n15709) );
  XNOR2_X1 U17253 ( .A(n15705), .B(keyinput46), .ZN(n15708) );
  XNOR2_X1 U17254 ( .A(n15706), .B(keyinput49), .ZN(n15707) );
  OR3_X1 U17255 ( .A1(n15709), .A2(n15708), .A3(n15707), .ZN(n15717) );
  AOI22_X1 U17256 ( .A1(n15711), .A2(keyinput33), .B1(keyinput3), .B2(n10387), 
        .ZN(n15710) );
  OAI221_X1 U17257 ( .B1(n15711), .B2(keyinput33), .C1(n10387), .C2(keyinput3), 
        .A(n15710), .ZN(n15716) );
  INV_X1 U17258 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n15713) );
  AOI22_X1 U17259 ( .A1(n15714), .A2(keyinput4), .B1(n15713), .B2(keyinput7), 
        .ZN(n15712) );
  OAI221_X1 U17260 ( .B1(n15714), .B2(keyinput4), .C1(n15713), .C2(keyinput7), 
        .A(n15712), .ZN(n15715) );
  NOR3_X1 U17261 ( .A1(n15717), .A2(n15716), .A3(n15715), .ZN(n15759) );
  AOI22_X1 U17262 ( .A1(n15720), .A2(keyinput40), .B1(n15719), .B2(keyinput16), 
        .ZN(n15718) );
  OAI221_X1 U17263 ( .B1(n15720), .B2(keyinput40), .C1(n15719), .C2(keyinput16), .A(n15718), .ZN(n15729) );
  XOR2_X1 U17264 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput60), .Z(n15728) );
  XNOR2_X1 U17265 ( .A(P3_REG0_REG_25__SCAN_IN), .B(keyinput37), .ZN(n15724)
         );
  XNOR2_X1 U17266 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput9), .ZN(n15723) );
  XNOR2_X1 U17267 ( .A(P1_REG3_REG_0__SCAN_IN), .B(keyinput34), .ZN(n15722) );
  XNOR2_X1 U17268 ( .A(P3_REG3_REG_3__SCAN_IN), .B(keyinput41), .ZN(n15721) );
  NAND4_X1 U17269 ( .A1(n15724), .A2(n15723), .A3(n15722), .A4(n15721), .ZN(
        n15727) );
  XNOR2_X1 U17270 ( .A(keyinput28), .B(n15725), .ZN(n15726) );
  NOR4_X1 U17271 ( .A1(n15729), .A2(n15728), .A3(n15727), .A4(n15726), .ZN(
        n15758) );
  AOI22_X1 U17272 ( .A1(n15731), .A2(keyinput18), .B1(n14743), .B2(keyinput63), 
        .ZN(n15730) );
  OAI221_X1 U17273 ( .B1(n15731), .B2(keyinput18), .C1(n14743), .C2(keyinput63), .A(n15730), .ZN(n15742) );
  INV_X1 U17274 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n15734) );
  AOI22_X1 U17275 ( .A1(n15734), .A2(keyinput57), .B1(keyinput59), .B2(n15733), 
        .ZN(n15732) );
  OAI221_X1 U17276 ( .B1(n15734), .B2(keyinput57), .C1(n15733), .C2(keyinput59), .A(n15732), .ZN(n15741) );
  XNOR2_X1 U17277 ( .A(n15735), .B(keyinput8), .ZN(n15740) );
  XNOR2_X1 U17278 ( .A(P3_REG1_REG_24__SCAN_IN), .B(keyinput29), .ZN(n15738)
         );
  XNOR2_X1 U17279 ( .A(P3_IR_REG_2__SCAN_IN), .B(keyinput31), .ZN(n15737) );
  XNOR2_X1 U17280 ( .A(P2_IR_REG_15__SCAN_IN), .B(keyinput45), .ZN(n15736) );
  NAND3_X1 U17281 ( .A1(n15738), .A2(n15737), .A3(n15736), .ZN(n15739) );
  NOR4_X1 U17282 ( .A1(n15742), .A2(n15741), .A3(n15740), .A4(n15739), .ZN(
        n15757) );
  AOI22_X1 U17283 ( .A1(n15744), .A2(keyinput2), .B1(n10889), .B2(keyinput55), 
        .ZN(n15743) );
  OAI221_X1 U17284 ( .B1(n15744), .B2(keyinput2), .C1(n10889), .C2(keyinput55), 
        .A(n15743), .ZN(n15755) );
  AOI22_X1 U17285 ( .A1(n15747), .A2(keyinput51), .B1(n15746), .B2(keyinput47), 
        .ZN(n15745) );
  OAI221_X1 U17286 ( .B1(n15747), .B2(keyinput51), .C1(n15746), .C2(keyinput47), .A(n15745), .ZN(n15754) );
  AOI22_X1 U17287 ( .A1(n11357), .A2(keyinput19), .B1(n15749), .B2(keyinput62), 
        .ZN(n15748) );
  OAI221_X1 U17288 ( .B1(n11357), .B2(keyinput19), .C1(n15749), .C2(keyinput62), .A(n15748), .ZN(n15753) );
  XNOR2_X1 U17289 ( .A(P3_IR_REG_1__SCAN_IN), .B(keyinput39), .ZN(n15751) );
  XNOR2_X1 U17290 ( .A(keyinput32), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n15750) );
  NAND2_X1 U17291 ( .A1(n15751), .A2(n15750), .ZN(n15752) );
  NOR4_X1 U17292 ( .A1(n15755), .A2(n15754), .A3(n15753), .A4(n15752), .ZN(
        n15756) );
  NAND4_X1 U17293 ( .A1(n15759), .A2(n15758), .A3(n15757), .A4(n15756), .ZN(
        n15821) );
  AOI22_X1 U17294 ( .A1(n8370), .A2(keyinput0), .B1(keyinput21), .B2(n14594), 
        .ZN(n15760) );
  OAI221_X1 U17295 ( .B1(n8370), .B2(keyinput0), .C1(n14594), .C2(keyinput21), 
        .A(n15760), .ZN(n15772) );
  AOI22_X1 U17296 ( .A1(n15763), .A2(keyinput27), .B1(keyinput44), .B2(n15762), 
        .ZN(n15761) );
  OAI221_X1 U17297 ( .B1(n15763), .B2(keyinput27), .C1(n15762), .C2(keyinput44), .A(n15761), .ZN(n15771) );
  AOI22_X1 U17298 ( .A1(n15766), .A2(keyinput42), .B1(n15765), .B2(keyinput50), 
        .ZN(n15764) );
  OAI221_X1 U17299 ( .B1(n15766), .B2(keyinput42), .C1(n15765), .C2(keyinput50), .A(n15764), .ZN(n15770) );
  XNOR2_X1 U17300 ( .A(P1_REG3_REG_9__SCAN_IN), .B(keyinput5), .ZN(n15768) );
  XNOR2_X1 U17301 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput30), .ZN(n15767) );
  NAND2_X1 U17302 ( .A1(n15768), .A2(n15767), .ZN(n15769) );
  NOR4_X1 U17303 ( .A1(n15772), .A2(n15771), .A3(n15770), .A4(n15769), .ZN(
        n15819) );
  AOI22_X1 U17304 ( .A1(n15774), .A2(keyinput52), .B1(keyinput12), .B2(n7563), 
        .ZN(n15773) );
  OAI221_X1 U17305 ( .B1(n15774), .B2(keyinput52), .C1(n7563), .C2(keyinput12), 
        .A(n15773), .ZN(n15785) );
  INV_X1 U17306 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n15777) );
  AOI22_X1 U17307 ( .A1(n15777), .A2(keyinput26), .B1(keyinput13), .B2(n15776), 
        .ZN(n15775) );
  OAI221_X1 U17308 ( .B1(n15777), .B2(keyinput26), .C1(n15776), .C2(keyinput13), .A(n15775), .ZN(n15784) );
  XOR2_X1 U17309 ( .A(n15778), .B(keyinput11), .Z(n15782) );
  XNOR2_X1 U17310 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput53), .ZN(n15781)
         );
  XNOR2_X1 U17311 ( .A(P3_IR_REG_17__SCAN_IN), .B(keyinput24), .ZN(n15780) );
  XNOR2_X1 U17312 ( .A(P2_IR_REG_13__SCAN_IN), .B(keyinput25), .ZN(n15779) );
  NAND4_X1 U17313 ( .A1(n15782), .A2(n15781), .A3(n15780), .A4(n15779), .ZN(
        n15783) );
  NOR3_X1 U17314 ( .A1(n15785), .A2(n15784), .A3(n15783), .ZN(n15818) );
  INV_X1 U17315 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n15787) );
  AOI22_X1 U17316 ( .A1(n15788), .A2(keyinput58), .B1(n15787), .B2(keyinput6), 
        .ZN(n15786) );
  OAI221_X1 U17317 ( .B1(n15788), .B2(keyinput58), .C1(n15787), .C2(keyinput6), 
        .A(n15786), .ZN(n15800) );
  INV_X1 U17318 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n15791) );
  AOI22_X1 U17319 ( .A1(n15791), .A2(keyinput56), .B1(keyinput20), .B2(n15790), 
        .ZN(n15789) );
  OAI221_X1 U17320 ( .B1(n15791), .B2(keyinput56), .C1(n15790), .C2(keyinput20), .A(n15789), .ZN(n15799) );
  AOI22_X1 U17321 ( .A1(n15794), .A2(keyinput61), .B1(n15793), .B2(keyinput38), 
        .ZN(n15792) );
  OAI221_X1 U17322 ( .B1(n15794), .B2(keyinput61), .C1(n15793), .C2(keyinput38), .A(n15792), .ZN(n15798) );
  INV_X1 U17323 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n15796) );
  AOI22_X1 U17324 ( .A1(n15796), .A2(keyinput10), .B1(keyinput23), .B2(n8912), 
        .ZN(n15795) );
  OAI221_X1 U17325 ( .B1(n15796), .B2(keyinput10), .C1(n8912), .C2(keyinput23), 
        .A(n15795), .ZN(n15797) );
  NOR4_X1 U17326 ( .A1(n15800), .A2(n15799), .A3(n15798), .A4(n15797), .ZN(
        n15817) );
  XNOR2_X1 U17327 ( .A(n15801), .B(keyinput1), .ZN(n15808) );
  XNOR2_X1 U17328 ( .A(P3_IR_REG_29__SCAN_IN), .B(keyinput48), .ZN(n15803) );
  XNOR2_X1 U17329 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput15), .ZN(n15802) );
  NAND2_X1 U17330 ( .A1(n15803), .A2(n15802), .ZN(n15807) );
  XNOR2_X1 U17331 ( .A(n15804), .B(keyinput22), .ZN(n15806) );
  XNOR2_X1 U17332 ( .A(keyinput14), .B(n7003), .ZN(n15805) );
  OR4_X1 U17333 ( .A1(n15808), .A2(n15807), .A3(n15806), .A4(n15805), .ZN(
        n15815) );
  AOI22_X1 U17334 ( .A1(n15811), .A2(keyinput17), .B1(n15810), .B2(keyinput54), 
        .ZN(n15809) );
  OAI221_X1 U17335 ( .B1(n15811), .B2(keyinput17), .C1(n15810), .C2(keyinput54), .A(n15809), .ZN(n15814) );
  INV_X1 U17336 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n15812) );
  XNOR2_X1 U17337 ( .A(n15812), .B(keyinput43), .ZN(n15813) );
  NOR3_X1 U17338 ( .A1(n15815), .A2(n15814), .A3(n15813), .ZN(n15816) );
  NAND4_X1 U17339 ( .A1(n15819), .A2(n15818), .A3(n15817), .A4(n15816), .ZN(
        n15820) );
  AOI211_X1 U17340 ( .C1(n15823), .C2(n15822), .A(n15821), .B(n15820), .ZN(
        n15838) );
  AOI22_X1 U17341 ( .A1(n15827), .A2(n15826), .B1(n15825), .B2(n15824), .ZN(
        n15828) );
  OAI21_X1 U17342 ( .B1(n15830), .B2(n15829), .A(n15828), .ZN(n15834) );
  MUX2_X1 U17343 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n15832), .S(n15831), .Z(
        n15833) );
  AOI211_X1 U17344 ( .C1(n15836), .C2(n15835), .A(n15834), .B(n15833), .ZN(
        n15837) );
  XNOR2_X1 U17345 ( .A(n15838), .B(n15837), .ZN(P2_U3260) );
  XOR2_X1 U17346 ( .A(n15840), .B(n15839), .Z(SUB_1596_U59) );
  AOI21_X1 U17347 ( .B1(n15842), .B2(n15841), .A(n15848), .ZN(SUB_1596_U53) );
  XOR2_X1 U17348 ( .A(n15844), .B(n15843), .Z(n15846) );
  XOR2_X1 U17349 ( .A(n15846), .B(n15845), .Z(SUB_1596_U60) );
  XOR2_X1 U17350 ( .A(n15848), .B(n15847), .Z(SUB_1596_U5) );
  NAND2_X2 U7489 ( .A1(n6501), .A2(n7136), .ZN(n14651) );
  BUF_X1 U10054 ( .A(n10407), .Z(n7215) );
  INV_X2 U7420 ( .A(n9907), .ZN(n9461) );
  NAND2_X1 U11377 ( .A1(n10845), .A2(n12646), .ZN(n10853) );
  NOR2_X1 U13607 ( .A1(n7699), .A2(n14994), .ZN(n11368) );
  CLKBUF_X1 U7212 ( .A(n9425), .Z(n9690) );
  CLKBUF_X1 U7216 ( .A(n12853), .Z(n12915) );
  CLKBUF_X1 U7260 ( .A(n8938), .Z(n10166) );
  AND2_X1 U7286 ( .A1(n12261), .A2(n12259), .ZN(n12821) );
  CLKBUF_X1 U7304 ( .A(n13379), .Z(n7172) );
  INV_X1 U7318 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n15153) );
  AND2_X1 U7396 ( .A1(n8193), .A2(n15884), .ZN(n15883) );
  NAND2_X1 U7629 ( .A1(n8194), .A2(n15883), .ZN(n14307) );
  NAND2_X1 U7676 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n8403), .ZN(n15884) );
  CLKBUF_X1 U9709 ( .A(n10250), .Z(n7177) );
endmodule

