

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618;

  NAND2_X1 U4905 ( .A1(n5268), .A2(n5267), .ZN(n8636) );
  CLKBUF_X1 U4906 ( .A(n7029), .Z(n4413) );
  INV_X1 U4907 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND2_X1 U4908 ( .A1(n8022), .A2(n10017), .ZN(n8072) );
  INV_X1 U4909 ( .A(n8327), .ZN(n9039) );
  BUF_X2 U4910 ( .A(n6194), .Z(n7258) );
  AND3_X1 U4911 ( .A1(n5535), .A2(n5534), .A3(n5533), .ZN(n7848) );
  CLKBUF_X2 U4912 ( .A(n5484), .Z(n4406) );
  INV_X1 U4913 ( .A(n7287), .ZN(n5885) );
  AND2_X1 U4914 ( .A1(n5477), .A2(n5372), .ZN(n5478) );
  CLKBUF_X3 U4915 ( .A(n5553), .Z(n4408) );
  INV_X1 U4918 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n4401) );
  OAI21_X1 U4919 ( .B1(n9392), .B2(n9411), .A(n5016), .ZN(n9414) );
  INV_X1 U4920 ( .A(n6705), .ZN(n7524) );
  OR2_X1 U4921 ( .A1(n9625), .A2(n9608), .ZN(n9347) );
  INV_X1 U4922 ( .A(n5444), .ZN(n4403) );
  INV_X1 U4923 ( .A(n6185), .ZN(n5222) );
  INV_X1 U4924 ( .A(n7071), .ZN(n6441) );
  OR2_X1 U4925 ( .A1(n5713), .A2(n9087), .ZN(n5738) );
  OR2_X1 U4926 ( .A1(n9578), .A2(n6967), .ZN(n9394) );
  OAI21_X1 U4927 ( .B1(n5293), .B2(n4974), .A(n4970), .ZN(n6948) );
  INV_X1 U4928 ( .A(n6194), .ZN(n6528) );
  XNOR2_X1 U4929 ( .A(n6539), .B(n6537), .ZN(n8464) );
  OR2_X1 U4930 ( .A1(n6579), .A2(n6159), .ZN(n6160) );
  OR2_X1 U4931 ( .A1(n4912), .A2(n7882), .ZN(n4909) );
  INV_X2 U4932 ( .A(n5484), .ZN(n5777) );
  NAND2_X1 U4933 ( .A1(n9556), .A2(n9465), .ZN(n9323) );
  INV_X1 U4934 ( .A(n9490), .ZN(n6918) );
  INV_X1 U4935 ( .A(n9072), .ZN(n7581) );
  NAND2_X1 U4936 ( .A1(n5532), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4763) );
  NAND2_X1 U4937 ( .A1(n6226), .A2(n5005), .ZN(n7673) );
  OR2_X1 U4938 ( .A1(n5428), .A2(n10036), .ZN(n6106) );
  AND2_X1 U4939 ( .A1(n8332), .A2(n8331), .ZN(n9049) );
  AND4_X1 U4940 ( .A1(n5543), .A2(n5542), .A3(n5541), .A4(n5540), .ZN(n7885)
         );
  NOR2_X1 U4941 ( .A1(n9561), .A2(n9822), .ZN(n9850) );
  NAND2_X1 U4942 ( .A1(n5736), .A2(n5735), .ZN(n9941) );
  AOI21_X1 U4943 ( .B1(n7033), .B2(n9782), .A(n7032), .ZN(n8286) );
  AND2_X1 U4944 ( .A1(n5413), .A2(n5412), .ZN(n5558) );
  AND2_X1 U4945 ( .A1(n6077), .A2(n6076), .ZN(n4402) );
  NOR2_X2 U4946 ( .A1(n5997), .A2(n9008), .ZN(n4887) );
  OAI21_X2 U4947 ( .B1(n9024), .B2(n5908), .A(n5907), .ZN(n9149) );
  OAI21_X2 U4948 ( .B1(n6565), .B2(P2_D_REG_0__SCAN_IN), .A(n7352), .ZN(n6705)
         );
  INV_X4 U4949 ( .A(n6238), .ZN(n6270) );
  NAND4_X2 U4951 ( .A1(n5505), .A2(n5504), .A3(n5503), .A4(n5502), .ZN(n9489)
         );
  NAND2_X2 U4952 ( .A1(n7121), .A2(n7123), .ZN(n7602) );
  OAI211_X2 U4953 ( .C1(n5318), .C2(n4910), .A(n4909), .B(n4907), .ZN(n7874)
         );
  INV_X1 U4954 ( .A(n6176), .ZN(n8317) );
  OAI21_X2 U4955 ( .B1(n5423), .B2(P1_IR_REG_26__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n4739) );
  OAI211_X2 U4956 ( .C1(P1_IR_REG_31__SCAN_IN), .C2(P1_IR_REG_1__SCAN_IN), .A(
        n4766), .B(n4765), .ZN(n7321) );
  NAND2_X1 U4957 ( .A1(n4764), .A2(n10385), .ZN(n4766) );
  XNOR2_X2 U4958 ( .A(n6160), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7594) );
  INV_X1 U4959 ( .A(n5558), .ZN(n4404) );
  INV_X4 U4960 ( .A(n4404), .ZN(n4405) );
  NAND2_X1 U4961 ( .A1(n5410), .A2(n5409), .ZN(n5484) );
  AND2_X1 U4962 ( .A1(n4943), .A2(n7765), .ZN(n4941) );
  XNOR2_X2 U4963 ( .A(n4763), .B(P1_IR_REG_3__SCAN_IN), .ZN(n7372) );
  XNOR2_X2 U4964 ( .A(n6233), .B(n6224), .ZN(n10184) );
  NAND2_X1 U4965 ( .A1(n6598), .A2(n7247), .ZN(n4407) );
  NAND2_X1 U4966 ( .A1(n8464), .A2(n8465), .ZN(n8463) );
  NAND2_X1 U4967 ( .A1(n4640), .A2(n4986), .ZN(n9597) );
  OR2_X1 U4968 ( .A1(n9451), .A2(n9398), .ZN(n9399) );
  NAND2_X2 U4969 ( .A1(n6428), .A2(n4473), .ZN(n5310) );
  NAND2_X1 U4970 ( .A1(n9708), .A2(n9376), .ZN(n9701) );
  NAND2_X1 U4971 ( .A1(n6680), .A2(n4490), .ZN(n8735) );
  AOI21_X1 U4972 ( .B1(n4794), .B2(n4793), .A(n4491), .ZN(n4792) );
  NAND2_X1 U4973 ( .A1(n4993), .A2(n7176), .ZN(n8784) );
  NAND2_X1 U4974 ( .A1(n9359), .A2(n5036), .ZN(n8015) );
  AND2_X1 U4975 ( .A1(n6493), .A2(n6492), .ZN(n8313) );
  INV_X2 U4976 ( .A(n9036), .ZN(n8329) );
  NAND2_X2 U4977 ( .A1(n5115), .A2(n9348), .ZN(n6970) );
  NAND2_X1 U4978 ( .A1(n9486), .A2(n7812), .ZN(n9354) );
  INV_X4 U4979 ( .A(n6057), .ZN(n5822) );
  INV_X1 U4980 ( .A(n9485), .ZN(n4645) );
  INV_X1 U4981 ( .A(n7710), .ZN(n7589) );
  AND4_X2 U4982 ( .A1(n6177), .A2(n5304), .A3(n5305), .A4(n5308), .ZN(n6633)
         );
  CLKBUF_X2 U4983 ( .A(n5501), .Z(n6112) );
  INV_X2 U4984 ( .A(n6208), .ZN(n6265) );
  OR2_X1 U4985 ( .A1(n7371), .A2(n4516), .ZN(n4758) );
  OAI21_X1 U4986 ( .B1(n5425), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5427) );
  XNOR2_X1 U4987 ( .A(n7357), .B(n5066), .ZN(n7358) );
  BUF_X2 U4988 ( .A(n6598), .Z(n6910) );
  AND3_X2 U4989 ( .A1(n5337), .A2(n5338), .A3(n4949), .ZN(n5399) );
  AND4_X2 U4990 ( .A1(n4458), .A2(n6203), .A3(n4592), .A4(n4591), .ZN(n4992)
         );
  INV_X4 U4991 ( .A(n5444), .ZN(n4409) );
  INV_X1 U4992 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n10302) );
  NAND2_X1 U4993 ( .A1(n8463), .A2(n6594), .ZN(n7274) );
  AOI21_X1 U4994 ( .B1(n9572), .B2(n9959), .A(n7000), .ZN(n7015) );
  OAI21_X1 U4995 ( .B1(n6699), .B2(n10218), .A(n6698), .ZN(n8650) );
  OAI22_X1 U4996 ( .A1(n8636), .A2(n6745), .B1(n8647), .B2(n7223), .ZN(n6762)
         );
  NOR2_X1 U4997 ( .A1(n9864), .A2(n4466), .ZN(n4658) );
  NAND2_X1 U4998 ( .A1(n8382), .A2(n6525), .ZN(n6539) );
  AOI21_X1 U4999 ( .B1(n6917), .B2(n10288), .A(n4596), .ZN(n4595) );
  OAI21_X1 U5000 ( .B1(n7076), .B2(n7075), .A(n7086), .ZN(n7077) );
  AOI21_X1 U5001 ( .B1(n4746), .B2(n4743), .A(n9305), .ZN(n9307) );
  OAI21_X1 U5002 ( .B1(n9126), .B2(n5332), .A(n5329), .ZN(n8340) );
  AOI21_X1 U5003 ( .B1(n4745), .B2(n4744), .A(n4506), .ZN(n4743) );
  NAND2_X1 U5004 ( .A1(n8427), .A2(n6486), .ZN(n8298) );
  NAND2_X1 U5005 ( .A1(n8373), .A2(n4487), .ZN(n8427) );
  NAND2_X1 U5006 ( .A1(n4934), .A2(n9615), .ZN(n9606) );
  INV_X1 U5007 ( .A(n9666), .ZN(n4410) );
  NAND2_X1 U5008 ( .A1(n4838), .A2(n4836), .ZN(n8373) );
  NAND2_X1 U5009 ( .A1(n8719), .A2(n6682), .ZN(n8706) );
  NAND2_X1 U5010 ( .A1(n4564), .A2(n4419), .ZN(n4563) );
  NOR2_X1 U5011 ( .A1(n4983), .A2(n4433), .ZN(n4982) );
  NAND2_X1 U5012 ( .A1(n9709), .A2(n9710), .ZN(n9708) );
  NAND2_X1 U5013 ( .A1(n10113), .A2(n4773), .ZN(n10122) );
  NAND2_X1 U5014 ( .A1(n9076), .A2(n4489), .ZN(n9164) );
  OAI21_X1 U5015 ( .B1(n8559), .B2(n8881), .A(n5241), .ZN(n8572) );
  XNOR2_X1 U5016 ( .A(n5243), .B(n5242), .ZN(n8559) );
  NAND2_X1 U5017 ( .A1(n9764), .A2(n6978), .ZN(n6979) );
  NAND2_X1 U5018 ( .A1(n9149), .A2(n9148), .ZN(n4927) );
  AND2_X1 U5019 ( .A1(n7073), .A2(n7072), .ZN(n8901) );
  NAND2_X1 U5020 ( .A1(n9777), .A2(n9271), .ZN(n9765) );
  AOI21_X1 U5021 ( .B1(n5283), .B2(n5281), .A(n4493), .ZN(n5280) );
  AOI21_X1 U5022 ( .B1(n5245), .B2(n8887), .A(n5238), .ZN(n5237) );
  NAND2_X1 U5023 ( .A1(n6068), .A2(n6067), .ZN(n9866) );
  NAND2_X1 U5024 ( .A1(n6955), .A2(n6954), .ZN(n9859) );
  NAND2_X1 U5025 ( .A1(n7932), .A2(n6277), .ZN(n8213) );
  NOR2_X1 U5026 ( .A1(n4655), .A2(n9715), .ZN(n4654) );
  OR2_X1 U5027 ( .A1(n7930), .A2(n7929), .ZN(n7932) );
  NAND2_X1 U5028 ( .A1(n6516), .A2(n6515), .ZN(n8912) );
  NAND2_X1 U5029 ( .A1(n7790), .A2(n6260), .ZN(n7930) );
  AND2_X1 U5030 ( .A1(n8416), .A2(n8417), .ZN(n4864) );
  NAND2_X1 U5031 ( .A1(n7721), .A2(n5299), .ZN(n7790) );
  NAND2_X1 U5032 ( .A1(n9506), .A2(n4539), .ZN(n8191) );
  XNOR2_X1 U5033 ( .A(n6541), .B(n6540), .ZN(n8987) );
  NAND2_X1 U5034 ( .A1(n6742), .A2(n6731), .ZN(n6541) );
  NAND2_X1 U5035 ( .A1(n5037), .A2(n9436), .ZN(n9359) );
  NOR2_X1 U5036 ( .A1(n4502), .A2(n5342), .ZN(n5341) );
  NAND2_X1 U5037 ( .A1(n5978), .A2(n5977), .ZN(n9688) );
  NAND2_X1 U5038 ( .A1(n9502), .A2(n4559), .ZN(n8197) );
  NAND2_X1 U5039 ( .A1(n6466), .A2(n6465), .ZN(n8863) );
  XNOR2_X1 U5040 ( .A(n6038), .B(n6037), .ZN(n8990) );
  NAND2_X1 U5041 ( .A1(n6038), .A2(n6037), .ZN(n6742) );
  AND2_X1 U5042 ( .A1(n5046), .A2(n9810), .ZN(n5045) );
  XNOR2_X1 U5043 ( .A(n5936), .B(n5935), .ZN(n8080) );
  NAND2_X1 U5044 ( .A1(n5947), .A2(n5946), .ZN(n9702) );
  NAND2_X1 U5045 ( .A1(n6454), .A2(n6453), .ZN(n8927) );
  NAND2_X1 U5046 ( .A1(n6489), .A2(n6013), .ZN(n6038) );
  AOI21_X1 U5047 ( .B1(n5351), .B2(n5353), .A(n5348), .ZN(n5347) );
  INV_X1 U5048 ( .A(n9810), .ZN(n9820) );
  NAND3_X1 U5049 ( .A1(n5320), .A2(n5322), .A3(n5319), .ZN(n5318) );
  NAND2_X1 U5050 ( .A1(n5994), .A2(n5993), .ZN(n6489) );
  OAI21_X1 U5051 ( .B1(n10438), .B2(n7992), .A(n5229), .ZN(n7977) );
  OAI21_X1 U5052 ( .B1(n4942), .B2(n4945), .A(n4941), .ZN(n7760) );
  INV_X1 U5053 ( .A(n8787), .ZN(n8783) );
  NAND2_X1 U5054 ( .A1(n6829), .A2(n7996), .ZN(n5229) );
  OAI21_X1 U5055 ( .B1(n5962), .B2(n5954), .A(n5955), .ZN(n5934) );
  OR2_X1 U5056 ( .A1(n4657), .A2(n9425), .ZN(n9357) );
  NOR2_X1 U5057 ( .A1(n7814), .A2(n5325), .ZN(n5324) );
  OR2_X1 U5058 ( .A1(n9941), .A2(n9934), .ZN(n9366) );
  NAND2_X1 U5059 ( .A1(n9067), .A2(n5500), .ZN(n7699) );
  NAND2_X1 U5060 ( .A1(n5035), .A2(n5912), .ZN(n5962) );
  NAND2_X1 U5061 ( .A1(n5843), .A2(n5842), .ZN(n9755) );
  NAND2_X1 U5062 ( .A1(n4603), .A2(n6382), .ZN(n8952) );
  NAND2_X1 U5063 ( .A1(n6357), .A2(n6356), .ZN(n8964) );
  NAND2_X1 U5064 ( .A1(n6342), .A2(n6341), .ZN(n8893) );
  NAND2_X1 U5065 ( .A1(n5712), .A2(n5711), .ZN(n9093) );
  NAND2_X1 U5066 ( .A1(n5052), .A2(n5051), .ZN(n8045) );
  OR2_X1 U5067 ( .A1(n7147), .A2(n7148), .ZN(n7945) );
  NAND2_X1 U5068 ( .A1(n5810), .A2(n5809), .ZN(n9937) );
  OAI21_X1 U5069 ( .B1(n5731), .B2(n5730), .A(n5754), .ZN(n5732) );
  XNOR2_X1 U5070 ( .A(n5731), .B(n5728), .ZN(n7437) );
  AND2_X1 U5071 ( .A1(n8174), .A2(n7153), .ZN(n8132) );
  NAND2_X1 U5072 ( .A1(n6294), .A2(n6293), .ZN(n8360) );
  NAND2_X1 U5073 ( .A1(n8006), .A2(n7151), .ZN(n7950) );
  AND2_X1 U5074 ( .A1(n7140), .A2(n7916), .ZN(n7148) );
  XNOR2_X1 U5075 ( .A(n5705), .B(n5706), .ZN(n7392) );
  AND2_X1 U5076 ( .A1(n7137), .A2(n7142), .ZN(n7663) );
  NAND2_X1 U5077 ( .A1(n4998), .A2(n5752), .ZN(n5731) );
  NAND2_X1 U5078 ( .A1(n9355), .A2(n4641), .ZN(n9431) );
  OAI21_X1 U5079 ( .B1(n5680), .B2(n5024), .A(n5023), .ZN(n5805) );
  NAND2_X1 U5080 ( .A1(n6304), .A2(n6303), .ZN(n8257) );
  NOR3_X1 U5081 ( .A1(n6821), .A2(n6910), .A3(n10284), .ZN(n10191) );
  NAND2_X1 U5082 ( .A1(n5618), .A2(n4665), .ZN(n9838) );
  INV_X1 U5083 ( .A(n7573), .ZN(n4947) );
  NAND2_X1 U5084 ( .A1(n4844), .A2(n4842), .ZN(n6194) );
  INV_X1 U5085 ( .A(n9489), .ZN(n7849) );
  NAND2_X1 U5086 ( .A1(n4716), .A2(n4714), .ZN(n5272) );
  AND2_X1 U5087 ( .A1(n5071), .A2(n5070), .ZN(n7386) );
  NAND2_X2 U5088 ( .A1(n5466), .A2(n9332), .ZN(n8327) );
  XNOR2_X1 U5089 ( .A(n4666), .B(n5368), .ZN(n7338) );
  NAND2_X1 U5090 ( .A1(n6257), .A2(n4445), .ZN(n8494) );
  AND3_X1 U5091 ( .A1(n5486), .A2(n5485), .A3(n4948), .ZN(n7573) );
  INV_X1 U5092 ( .A(n7885), .ZN(n9486) );
  NAND4_X1 U5093 ( .A1(n5593), .A2(n5592), .A3(n5591), .A4(n5590), .ZN(n9483)
         );
  NAND3_X2 U5094 ( .A1(n6210), .A2(n6212), .A3(n4451), .ZN(n8497) );
  NAND4_X1 U5095 ( .A1(n6245), .A2(n6244), .A3(n6243), .A4(n6242), .ZN(n8495)
         );
  NAND4_X2 U5096 ( .A1(n5357), .A2(n5474), .A3(n5473), .A4(n5472), .ZN(n9490)
         );
  AND4_X1 U5097 ( .A1(n6183), .A2(n6181), .A3(n6180), .A4(n6182), .ZN(n7604)
         );
  AND4_X1 U5098 ( .A1(n5625), .A2(n5624), .A3(n5623), .A4(n5622), .ZN(n9063)
         );
  INV_X2 U5099 ( .A(P2_U3893), .ZN(n8606) );
  NAND2_X1 U5100 ( .A1(n4994), .A2(n5578), .ZN(n5602) );
  INV_X1 U5101 ( .A(n7450), .ZN(n10224) );
  AND2_X1 U5102 ( .A1(n4722), .A2(n4715), .ZN(n4714) );
  INV_X1 U5103 ( .A(n7607), .ZN(n7964) );
  NAND2_X1 U5104 ( .A1(n4894), .A2(n4893), .ZN(n5235) );
  INV_X1 U5105 ( .A(n4408), .ZN(n6986) );
  OR2_X1 U5106 ( .A1(n5531), .A2(n7322), .ZN(n5477) );
  NAND2_X1 U5107 ( .A1(n4758), .A2(n4757), .ZN(n5063) );
  AOI21_X1 U5108 ( .B1(n7428), .B2(P2_REG1_REG_3__SCAN_IN), .A(n4668), .ZN(
        n10186) );
  XNOR2_X1 U5109 ( .A(n5427), .B(n5426), .ZN(n10036) );
  XNOR2_X1 U5110 ( .A(n4669), .B(n5247), .ZN(n7428) );
  NAND2_X1 U5111 ( .A1(n8317), .A2(n5307), .ZN(n6208) );
  INV_X1 U5112 ( .A(n5307), .ZN(n4577) );
  XNOR2_X1 U5113 ( .A(n5431), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9464) );
  NAND2_X1 U5114 ( .A1(n4862), .A2(n4863), .ZN(n8992) );
  NAND2_X2 U5115 ( .A1(n6598), .A2(n7247), .ZN(n6185) );
  XNOR2_X1 U5116 ( .A(n5432), .B(n10302), .ZN(n9455) );
  AND2_X1 U5117 ( .A1(n6161), .A2(n6158), .ZN(n6579) );
  NAND2_X1 U5118 ( .A1(n5547), .A2(SI_4_), .ZN(n5567) );
  INV_X1 U5119 ( .A(n7372), .ZN(n7357) );
  OR2_X1 U5120 ( .A1(n5404), .A2(n10021), .ZN(n5401) );
  NOR2_X1 U5121 ( .A1(n6165), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U5122 ( .A1(n4457), .A2(n4691), .ZN(n5547) );
  AND2_X1 U5123 ( .A1(n5399), .A2(n10302), .ZN(n5429) );
  NAND2_X1 U5124 ( .A1(n4992), .A2(n5365), .ZN(n6154) );
  AND3_X1 U5125 ( .A1(n5399), .A2(n5339), .A3(n5135), .ZN(n5404) );
  INV_X2 U5126 ( .A(n8976), .ZN(n4411) );
  AND2_X1 U5127 ( .A1(n4426), .A2(n4532), .ZN(n5339) );
  AND4_X1 U5128 ( .A1(n5393), .A2(n5396), .A3(n5394), .A4(n5395), .ZN(n4949)
         );
  AND3_X1 U5129 ( .A1(n6190), .A2(n10297), .A3(n4786), .ZN(n6203) );
  AND3_X1 U5130 ( .A1(n6143), .A2(n6142), .A3(n6141), .ZN(n6151) );
  INV_X1 U5131 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6233) );
  INV_X1 U5132 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6280) );
  NOR2_X1 U5133 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n6135) );
  INV_X1 U5134 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n10317) );
  INV_X4 U5135 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5136 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5463) );
  NOR2_X1 U5137 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n6136) );
  INV_X1 U5138 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5450) );
  INV_X1 U5139 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6395) );
  INV_X1 U5140 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6190) );
  NOR2_X1 U5141 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5393) );
  NOR2_X1 U5142 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5394) );
  NOR2_X1 U5143 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5395) );
  INV_X1 U5144 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6394) );
  NOR2_X1 U5145 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5390) );
  INV_X1 U5146 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6353) );
  NOR2_X1 U5147 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5388) );
  NOR2_X1 U5148 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5389) );
  NOR2_X1 U5149 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5392) );
  INV_X2 U5150 ( .A(n9220), .ZN(n5579) );
  AOI21_X2 U5151 ( .B1(n8334), .B2(n8333), .A(n9049), .ZN(n8335) );
  OAI21_X2 U5152 ( .B1(n9597), .B2(n5291), .A(n5290), .ZN(n7017) );
  AND2_X4 U5153 ( .A1(n4606), .A2(n4605), .ZN(n5444) );
  INV_X1 U5154 ( .A(n4402), .ZN(n4412) );
  NAND2_X1 U5155 ( .A1(n5413), .A2(n5409), .ZN(n5553) );
  XNOR2_X1 U5156 ( .A(n4739), .B(n5450), .ZN(n7029) );
  AOI22_X2 U5157 ( .A1(n5579), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n5885), .B2(
        n7384), .ZN(n5569) );
  NOR2_X1 U5158 ( .A1(n6176), .A2(n5307), .ZN(n4414) );
  NOR2_X1 U5159 ( .A1(n6176), .A2(n5307), .ZN(n4415) );
  NOR2_X2 U5160 ( .A1(n6176), .A2(n5307), .ZN(n6604) );
  INV_X1 U5161 ( .A(n6238), .ZN(n4416) );
  INV_X1 U5162 ( .A(n6185), .ZN(n4417) );
  AND2_X2 U5163 ( .A1(n4810), .A2(n7275), .ZN(P1_U3973) );
  NAND2_X1 U5164 ( .A1(n4635), .A2(n4634), .ZN(n7128) );
  NAND2_X1 U5165 ( .A1(n7598), .A2(n8082), .ZN(n4634) );
  NAND2_X1 U5166 ( .A1(n4636), .A2(n7594), .ZN(n4635) );
  NAND2_X1 U5167 ( .A1(n7125), .A2(n8085), .ZN(n4636) );
  NAND2_X1 U5168 ( .A1(n7986), .A2(n5364), .ZN(n6807) );
  NOR2_X1 U5169 ( .A1(n6690), .A2(n5253), .ZN(n5252) );
  INV_X1 U5170 ( .A(n6687), .ZN(n5253) );
  NAND2_X1 U5171 ( .A1(n4407), .A2(n5444), .ZN(n6225) );
  AND2_X1 U5172 ( .A1(n7250), .A2(n7594), .ZN(n4420) );
  INV_X1 U5173 ( .A(n6139), .ZN(n4591) );
  AND2_X1 U5174 ( .A1(n4968), .A2(n4518), .ZN(n4966) );
  OAI21_X1 U5175 ( .B1(n5883), .B2(n5864), .A(n5863), .ZN(n5909) );
  NAND2_X1 U5176 ( .A1(n5869), .A2(n9455), .ZN(n9335) );
  NAND2_X1 U5177 ( .A1(n5280), .A2(n5282), .ZN(n5278) );
  AND2_X1 U5178 ( .A1(n4940), .A2(n9254), .ZN(n4939) );
  INV_X1 U5179 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4646) );
  MUX2_X1 U5180 ( .A(n7124), .B(n7123), .S(n4420), .Z(n7131) );
  NAND2_X1 U5181 ( .A1(n8132), .A2(n7150), .ZN(n7157) );
  MUX2_X1 U5182 ( .A(n7149), .B(n7152), .S(n7217), .Z(n7150) );
  AOI21_X1 U5183 ( .B1(n7184), .B2(n7182), .A(n7181), .ZN(n7186) );
  NAND3_X1 U5184 ( .A1(n4626), .A2(n4859), .A3(n4625), .ZN(n7184) );
  NAND2_X1 U5185 ( .A1(n5112), .A2(n7964), .ZN(n7121) );
  OR2_X1 U5186 ( .A1(n6730), .A2(n6729), .ZN(n6734) );
  AND2_X1 U5187 ( .A1(n5027), .A2(n5026), .ZN(n5025) );
  NAND2_X1 U5188 ( .A1(n5530), .A2(n5529), .ZN(n5038) );
  NOR2_X1 U5189 ( .A1(n7243), .A2(n4843), .ZN(n4842) );
  AND2_X1 U5190 ( .A1(n7594), .A2(n7936), .ZN(n4843) );
  OR2_X1 U5191 ( .A1(n7104), .A2(n4955), .ZN(n7112) );
  AND3_X1 U5192 ( .A1(n4701), .A2(n8661), .A3(n4431), .ZN(n4956) );
  INV_X1 U5193 ( .A(n6374), .ZN(n6209) );
  NAND2_X1 U5194 ( .A1(n4577), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5306) );
  AND2_X1 U5195 ( .A1(n5307), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5303) );
  AND2_X1 U5196 ( .A1(n4965), .A2(n4964), .ZN(n4963) );
  INV_X1 U5197 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n4964) );
  INV_X1 U5198 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6266) );
  NAND2_X1 U5199 ( .A1(n6657), .A2(n4849), .ZN(n5106) );
  AND2_X1 U5200 ( .A1(n4476), .A2(n6656), .ZN(n4849) );
  INV_X1 U5201 ( .A(n8716), .ZN(n4564) );
  AND2_X1 U5202 ( .A1(n8684), .A2(n4566), .ZN(n4565) );
  NAND2_X1 U5203 ( .A1(n4567), .A2(n4419), .ZN(n4566) );
  INV_X1 U5204 ( .A(n7187), .ZN(n4567) );
  INV_X1 U5205 ( .A(n6685), .ZN(n5257) );
  NAND2_X1 U5206 ( .A1(n8795), .A2(n6672), .ZN(n6674) );
  NAND2_X1 U5207 ( .A1(n6600), .A2(n6185), .ZN(n6695) );
  AND2_X1 U5208 ( .A1(n5333), .A2(n4919), .ZN(n4918) );
  OR2_X1 U5209 ( .A1(n9157), .A2(n4920), .ZN(n4919) );
  NOR2_X1 U5210 ( .A1(n5335), .A2(n5334), .ZN(n5333) );
  INV_X1 U5211 ( .A(n5386), .ZN(n5334) );
  NAND2_X1 U5212 ( .A1(n4726), .A2(n4724), .ZN(n5801) );
  AND2_X1 U5213 ( .A1(n5800), .A2(n4725), .ZN(n4724) );
  NAND2_X1 U5214 ( .A1(n7489), .A2(n4728), .ZN(n4726) );
  INV_X1 U5215 ( .A(n6944), .ZN(n4975) );
  AND2_X1 U5216 ( .A1(n4472), .A2(n6942), .ZN(n5292) );
  AND3_X1 U5217 ( .A1(n9431), .A2(n5378), .A3(n9427), .ZN(n6923) );
  NAND2_X1 U5218 ( .A1(n5869), .A2(n9405), .ZN(n6968) );
  NAND2_X1 U5219 ( .A1(n5381), .A2(n5987), .ZN(n5994) );
  OAI21_X1 U5220 ( .B1(n5911), .B2(n5030), .A(n5028), .ZN(n5381) );
  INV_X1 U5221 ( .A(n5032), .ZN(n5030) );
  AND2_X1 U5222 ( .A1(n4520), .A2(n5029), .ZN(n5028) );
  INV_X1 U5223 ( .A(n5856), .ZN(n5021) );
  XNOR2_X1 U5224 ( .A(n6168), .B(n6169), .ZN(n6598) );
  NAND2_X1 U5225 ( .A1(n4593), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6168) );
  AOI21_X1 U5226 ( .B1(n5009), .B2(n5008), .A(n4513), .ZN(n5007) );
  INV_X1 U5227 ( .A(n8117), .ZN(n5008) );
  NAND2_X1 U5228 ( .A1(n6178), .A2(n6633), .ZN(n6187) );
  OR2_X1 U5229 ( .A1(n8397), .A2(n8489), .ZN(n6426) );
  AOI21_X1 U5230 ( .B1(n7238), .B2(n4633), .A(n4630), .ZN(n4629) );
  NAND2_X1 U5231 ( .A1(n4632), .A2(n4631), .ZN(n4630) );
  AOI21_X1 U5232 ( .B1(n7228), .B2(n7229), .A(n4504), .ZN(n4631) );
  INV_X2 U5233 ( .A(n6209), .ZN(n7058) );
  NAND2_X1 U5234 ( .A1(n10179), .A2(n4670), .ZN(n6789) );
  NAND2_X1 U5235 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n10297), .ZN(n4670) );
  NAND2_X1 U5236 ( .A1(n6807), .A2(n4675), .ZN(n6808) );
  NAND2_X1 U5237 ( .A1(n5146), .A2(n8507), .ZN(n5145) );
  OAI211_X1 U5238 ( .C1(n8499), .C2(n4673), .A(n4671), .B(n4543), .ZN(n5246)
         );
  NAND2_X1 U5239 ( .A1(n8515), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4673) );
  NAND2_X1 U5240 ( .A1(n4672), .A2(n8515), .ZN(n4671) );
  XNOR2_X1 U5241 ( .A(n4679), .B(n6906), .ZN(n5232) );
  NAND2_X1 U5242 ( .A1(n4680), .A2(n4562), .ZN(n4679) );
  NAND2_X1 U5243 ( .A1(n8600), .A2(n8601), .ZN(n4680) );
  INV_X1 U5244 ( .A(n8484), .ZN(n7223) );
  XNOR2_X1 U5245 ( .A(n8484), .B(n8844), .ZN(n8641) );
  INV_X1 U5246 ( .A(n8670), .ZN(n8465) );
  NAND2_X1 U5247 ( .A1(n5266), .A2(n6692), .ZN(n6728) );
  OR2_X1 U5248 ( .A1(n6477), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6494) );
  AND2_X1 U5249 ( .A1(n6643), .A2(n7190), .ZN(n5219) );
  NAND2_X1 U5250 ( .A1(n4446), .A2(n4571), .ZN(n4570) );
  NAND2_X1 U5251 ( .A1(n4699), .A2(n6502), .ZN(n6650) );
  NAND2_X1 U5252 ( .A1(n8990), .A2(n6278), .ZN(n4699) );
  NAND2_X1 U5253 ( .A1(n4563), .A2(n4565), .ZN(n6649) );
  INV_X1 U5254 ( .A(n7857), .ZN(n7080) );
  INV_X1 U5255 ( .A(n8761), .ZN(n8732) );
  NOR2_X1 U5256 ( .A1(n4471), .A2(n5264), .ZN(n5263) );
  INV_X1 U5257 ( .A(n6678), .ZN(n5264) );
  OR2_X1 U5258 ( .A1(n7217), .A2(n6631), .ZN(n7517) );
  NAND2_X1 U5259 ( .A1(n8085), .A2(n8082), .ZN(n10242) );
  AND2_X1 U5260 ( .A1(n7353), .A2(n6584), .ZN(n7332) );
  AND2_X1 U5261 ( .A1(n6912), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6584) );
  NAND2_X1 U5262 ( .A1(n8970), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6174) );
  NOR2_X1 U5263 ( .A1(n7279), .A2(n5496), .ZN(n9069) );
  NOR2_X1 U5264 ( .A1(n5650), .A2(n5343), .ZN(n5342) );
  NAND2_X1 U5265 ( .A1(n4819), .A2(n4818), .ZN(n4817) );
  NAND2_X1 U5266 ( .A1(n5317), .A2(n5323), .ZN(n5316) );
  INV_X1 U5267 ( .A(n5324), .ZN(n5317) );
  INV_X1 U5268 ( .A(n4925), .ZN(n4924) );
  AOI21_X1 U5269 ( .B1(n4925), .B2(n4923), .A(n4922), .ZN(n4921) );
  INV_X1 U5270 ( .A(n9402), .ZN(n7692) );
  NAND2_X1 U5271 ( .A1(n9068), .A2(n9069), .ZN(n9067) );
  NAND2_X1 U5272 ( .A1(n9335), .A2(n5490), .ZN(n4811) );
  NOR2_X1 U5273 ( .A1(n7783), .A2(n5359), .ZN(n5319) );
  NOR2_X1 U5274 ( .A1(n6123), .A2(n7692), .ZN(n6118) );
  AND2_X1 U5275 ( .A1(n7286), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7275) );
  AND2_X1 U5276 ( .A1(n7562), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5061) );
  NOR2_X1 U5277 ( .A1(n9532), .A2(n4558), .ZN(n9543) );
  NAND2_X1 U5278 ( .A1(n4770), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n4772) );
  INV_X1 U5279 ( .A(n9533), .ZN(n4770) );
  NAND2_X1 U5280 ( .A1(n10123), .A2(n9552), .ZN(n10143) );
  NAND2_X1 U5281 ( .A1(n10120), .A2(n4551), .ZN(n10140) );
  AOI21_X1 U5282 ( .B1(n9446), .B2(n4931), .A(n4930), .ZN(n4929) );
  INV_X1 U5283 ( .A(n9342), .ZN(n4931) );
  INV_X1 U5284 ( .A(n9394), .ZN(n4930) );
  INV_X1 U5285 ( .A(n5280), .ZN(n5279) );
  NAND2_X1 U5286 ( .A1(n4410), .A2(n4429), .ZN(n4987) );
  INV_X1 U5287 ( .A(n5286), .ZN(n5284) );
  NAND2_X1 U5288 ( .A1(n6941), .A2(n4479), .ZN(n5293) );
  INV_X1 U5289 ( .A(n6940), .ZN(n5294) );
  AOI21_X1 U5290 ( .B1(n4966), .B2(n5288), .A(n4500), .ZN(n4651) );
  NAND2_X1 U5291 ( .A1(n4966), .A2(n8152), .ZN(n4650) );
  NOR2_X1 U5292 ( .A1(n5177), .A2(n9838), .ZN(n5176) );
  INV_X1 U5293 ( .A(n5178), .ZN(n5177) );
  AND2_X1 U5294 ( .A1(n9357), .A2(n9437), .ZN(n5036) );
  INV_X1 U5295 ( .A(n9804), .ZN(n9815) );
  INV_X1 U5296 ( .A(n9877), .ZN(n9943) );
  AND2_X1 U5297 ( .A1(n9335), .A2(n7619), .ZN(n10154) );
  OR2_X1 U5298 ( .A1(n9323), .A2(n9400), .ZN(n9968) );
  NAND2_X1 U5299 ( .A1(n6983), .A2(n9332), .ZN(n9782) );
  NAND2_X1 U5300 ( .A1(n7705), .A2(n9968), .ZN(n9959) );
  AND2_X1 U5301 ( .A1(n6106), .A2(n7275), .ZN(n9402) );
  MUX2_X1 U5302 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5403), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5405) );
  XNOR2_X1 U5303 ( .A(n5909), .B(n5910), .ZN(n7856) );
  NAND2_X1 U5304 ( .A1(n4599), .A2(n4598), .ZN(n7424) );
  INV_X1 U5305 ( .A(n7427), .ZN(n4598) );
  INV_X1 U5306 ( .A(n7426), .ZN(n4599) );
  INV_X1 U5307 ( .A(n10191), .ZN(n10176) );
  XNOR2_X1 U5308 ( .A(n6830), .B(n8507), .ZN(n8499) );
  OAI211_X1 U5309 ( .C1(n5366), .C2(n9462), .A(n9461), .B(n9460), .ZN(n9463)
         );
  NAND2_X1 U5310 ( .A1(n10122), .A2(n10121), .ZN(n10120) );
  NAND2_X1 U5311 ( .A1(n9222), .A2(n9221), .ZN(n9855) );
  NAND2_X1 U5312 ( .A1(n7142), .A2(n7132), .ZN(n4991) );
  NAND2_X1 U5313 ( .A1(n7134), .A2(n7217), .ZN(n4989) );
  NAND2_X1 U5314 ( .A1(n7137), .A2(n7133), .ZN(n7134) );
  AOI21_X1 U5315 ( .B1(n7146), .B2(n4477), .A(n4638), .ZN(n4637) );
  INV_X1 U5316 ( .A(n7148), .ZN(n4638) );
  NOR2_X1 U5317 ( .A1(n4465), .A2(n5083), .ZN(n5082) );
  NAND2_X1 U5318 ( .A1(n7139), .A2(n4488), .ZN(n5084) );
  NAND2_X1 U5319 ( .A1(n4732), .A2(n9228), .ZN(n9229) );
  AND2_X1 U5320 ( .A1(n9355), .A2(n9354), .ZN(n4738) );
  OR2_X1 U5321 ( .A1(n4424), .A2(n4525), .ZN(n4627) );
  OR2_X1 U5322 ( .A1(n7179), .A2(n7178), .ZN(n4859) );
  INV_X1 U5323 ( .A(n7189), .ZN(n4614) );
  INV_X1 U5324 ( .A(n7190), .ZN(n4613) );
  INV_X1 U5325 ( .A(n7193), .ZN(n4612) );
  NAND2_X1 U5326 ( .A1(n4610), .A2(n4609), .ZN(n4616) );
  AOI21_X1 U5327 ( .B1(n7187), .B2(n7188), .A(n4420), .ZN(n4609) );
  NAND2_X1 U5328 ( .A1(n7191), .A2(n7187), .ZN(n4610) );
  OAI211_X1 U5329 ( .C1(n9278), .C2(n9323), .A(n9747), .B(n4742), .ZN(n5141)
         );
  NAND2_X1 U5330 ( .A1(n4430), .A2(n9323), .ZN(n4742) );
  OAI211_X1 U5331 ( .C1(n5141), .C2(n5139), .A(n5138), .B(n5137), .ZN(n9296)
         );
  NAND2_X1 U5332 ( .A1(n5140), .A2(n9323), .ZN(n5139) );
  NOR2_X1 U5333 ( .A1(n9289), .A2(n9290), .ZN(n5137) );
  NAND2_X1 U5334 ( .A1(n4741), .A2(n4464), .ZN(n5138) );
  AND2_X1 U5335 ( .A1(n5148), .A2(n7306), .ZN(n6792) );
  INV_X1 U5336 ( .A(n4583), .ZN(n4581) );
  INV_X1 U5337 ( .A(n8574), .ZN(n4579) );
  INV_X1 U5338 ( .A(n8590), .ZN(n4582) );
  NOR2_X1 U5339 ( .A1(n6901), .A2(n4584), .ZN(n4583) );
  INV_X1 U5340 ( .A(n6897), .ZN(n4584) );
  NAND2_X1 U5341 ( .A1(n9701), .A2(n9380), .ZN(n9412) );
  NAND2_X1 U5342 ( .A1(n5047), .A2(n9364), .ZN(n5046) );
  INV_X1 U5343 ( .A(n9250), .ZN(n5047) );
  AND2_X1 U5344 ( .A1(n9252), .A2(n8045), .ZN(n9243) );
  INV_X1 U5345 ( .A(n5761), .ZN(n5020) );
  AND2_X1 U5346 ( .A1(n5707), .A2(n5656), .ZN(n5271) );
  INV_X1 U5347 ( .A(n5261), .ZN(n4723) );
  INV_X1 U5348 ( .A(n5602), .ZN(n4717) );
  NAND2_X1 U5349 ( .A1(n5260), .A2(n5368), .ZN(n4722) );
  INV_X1 U5350 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n4690) );
  AOI21_X1 U5351 ( .B1(n6514), .B2(n4829), .A(n4828), .ZN(n4827) );
  INV_X1 U5352 ( .A(n6501), .ZN(n4829) );
  INV_X1 U5353 ( .A(n6514), .ZN(n4830) );
  AND2_X1 U5354 ( .A1(n8440), .A2(n6312), .ZN(n6336) );
  AND2_X1 U5355 ( .A1(n7236), .A2(n4420), .ZN(n4633) );
  INV_X1 U5356 ( .A(n8901), .ZN(n7240) );
  NAND2_X1 U5357 ( .A1(n7429), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10190) );
  NAND2_X1 U5358 ( .A1(n10184), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5234) );
  NAND2_X1 U5359 ( .A1(n6797), .A2(n6796), .ZN(n6800) );
  NAND2_X1 U5360 ( .A1(n7545), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6796) );
  INV_X1 U5361 ( .A(n8545), .ZN(n4590) );
  AOI21_X1 U5362 ( .B1(n8550), .B2(n8549), .A(n4442), .ZN(n5153) );
  OR2_X1 U5363 ( .A1(n8536), .A2(n5152), .ZN(n5151) );
  INV_X1 U5364 ( .A(n6692), .ZN(n5270) );
  INV_X1 U5365 ( .A(n7221), .ZN(n4957) );
  AND2_X1 U5366 ( .A1(n5102), .A2(n8675), .ZN(n4848) );
  INV_X1 U5367 ( .A(n5104), .ZN(n5099) );
  INV_X1 U5368 ( .A(n6505), .ZN(n6504) );
  INV_X1 U5369 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n4962) );
  INV_X1 U5370 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6444) );
  INV_X1 U5371 ( .A(n6446), .ZN(n6445) );
  INV_X1 U5372 ( .A(n6345), .ZN(n6344) );
  OR2_X1 U5373 ( .A1(n7522), .A2(n6705), .ZN(n6702) );
  OR2_X1 U5374 ( .A1(n8313), .A2(n8681), .ZN(n7208) );
  OR2_X1 U5375 ( .A1(n8863), .A2(n6644), .ZN(n8288) );
  OR2_X1 U5376 ( .A1(n8938), .A2(n8732), .ZN(n7192) );
  AOI21_X1 U5377 ( .B1(n6652), .B2(n5207), .A(n5206), .ZN(n5205) );
  INV_X1 U5378 ( .A(n6651), .ZN(n5207) );
  INV_X1 U5379 ( .A(n7182), .ZN(n5206) );
  AND2_X1 U5380 ( .A1(n5211), .A2(n7155), .ZN(n4575) );
  NOR2_X1 U5381 ( .A1(n5213), .A2(n5212), .ZN(n5211) );
  NAND2_X1 U5382 ( .A1(n4995), .A2(n7169), .ZN(n5210) );
  NAND2_X1 U5383 ( .A1(n5216), .A2(n8833), .ZN(n4995) );
  NAND2_X1 U5384 ( .A1(n6640), .A2(n7165), .ZN(n5216) );
  NOR2_X1 U5385 ( .A1(n4501), .A2(n5108), .ZN(n5107) );
  INV_X1 U5386 ( .A(n6668), .ZN(n5108) );
  NAND2_X1 U5387 ( .A1(n5199), .A2(n7138), .ZN(n5198) );
  INV_X1 U5388 ( .A(n7137), .ZN(n5199) );
  OR2_X1 U5389 ( .A1(n7594), .A2(n7936), .ZN(n6587) );
  NOR2_X1 U5390 ( .A1(n5315), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n5314) );
  NOR2_X1 U5391 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n6150) );
  NAND2_X1 U5392 ( .A1(n5347), .A2(n5352), .ZN(n5343) );
  AND2_X1 U5393 ( .A1(n4926), .A2(n9147), .ZN(n4925) );
  OR2_X1 U5394 ( .A1(n7698), .A2(n4421), .ZN(n5322) );
  AND2_X1 U5395 ( .A1(n9128), .A2(n4903), .ZN(n4902) );
  NAND2_X1 U5396 ( .A1(n4904), .A2(n9004), .ZN(n4903) );
  INV_X1 U5397 ( .A(n9003), .ZN(n4904) );
  NAND2_X1 U5398 ( .A1(n4747), .A2(n9323), .ZN(n4746) );
  NAND2_X1 U5399 ( .A1(n6967), .A2(n9578), .ZN(n9309) );
  NOR2_X1 U5400 ( .A1(n6952), .A2(n5277), .ZN(n4985) );
  NAND2_X1 U5401 ( .A1(n9633), .A2(n9625), .ZN(n4986) );
  NAND2_X1 U5402 ( .A1(n5039), .A2(n4494), .ZN(n5382) );
  NAND2_X1 U5403 ( .A1(n5012), .A2(n9876), .ZN(n9424) );
  AND2_X1 U5404 ( .A1(n5184), .A2(n5187), .ZN(n5183) );
  NOR2_X1 U5405 ( .A1(n9789), .A2(n5185), .ZN(n5184) );
  INV_X1 U5406 ( .A(n5186), .ZN(n5185) );
  INV_X1 U5407 ( .A(n9354), .ZN(n4946) );
  NAND2_X1 U5408 ( .A1(n9226), .A2(n9354), .ZN(n9427) );
  NAND2_X1 U5409 ( .A1(n6751), .A2(n6750), .ZN(n7047) );
  OR2_X1 U5410 ( .A1(n6546), .A2(n6545), .ZN(n6729) );
  INV_X1 U5411 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5420) );
  AND2_X1 U5412 ( .A1(n6544), .A2(n6042), .ZN(n6540) );
  INV_X1 U5413 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6104) );
  NOR2_X1 U5414 ( .A1(n5961), .A2(n5033), .ZN(n5032) );
  INV_X1 U5415 ( .A(n5912), .ZN(n5033) );
  OR2_X1 U5416 ( .A1(n5909), .A2(n5910), .ZN(n5035) );
  NAND2_X1 U5417 ( .A1(n5805), .A2(n4698), .ZN(n5017) );
  NOR2_X1 U5418 ( .A1(n4418), .A2(n5804), .ZN(n4698) );
  NAND2_X1 U5419 ( .A1(n5762), .A2(n4460), .ZN(n5019) );
  INV_X1 U5420 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5457) );
  INV_X1 U5421 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4815) );
  NAND2_X1 U5422 ( .A1(n5262), .A2(n5604), .ZN(n5261) );
  INV_X1 U5423 ( .A(n5628), .ZN(n5262) );
  OAI21_X1 U5424 ( .B1(n5547), .B2(SI_4_), .A(n4688), .ZN(n4687) );
  INV_X1 U5425 ( .A(n5568), .ZN(n4688) );
  OR2_X1 U5426 ( .A1(n6389), .A2(n8771), .ZN(n6390) );
  NAND2_X1 U5427 ( .A1(n5011), .A2(n8117), .ZN(n5010) );
  AND2_X1 U5428 ( .A1(n4837), .A2(n8371), .ZN(n4836) );
  OR2_X1 U5429 ( .A1(n4864), .A2(n8372), .ZN(n4837) );
  NAND2_X1 U5430 ( .A1(n4821), .A2(n7415), .ZN(n7416) );
  INV_X1 U5431 ( .A(n7418), .ZN(n4821) );
  AND2_X1 U5432 ( .A1(n6614), .A2(n6613), .ZN(n6701) );
  OR2_X1 U5433 ( .A1(n7217), .A2(n7243), .ZN(n6613) );
  AND2_X1 U5434 ( .A1(n7936), .A2(n7857), .ZN(n7243) );
  AND4_X2 U5435 ( .A1(n6199), .A2(n6198), .A3(n6197), .A4(n6196), .ZN(n7605)
         );
  OR2_X1 U5436 ( .A1(n5306), .A2(n6176), .ZN(n5308) );
  OR2_X1 U5437 ( .A1(n6208), .A2(n6179), .ZN(n6181) );
  OR2_X1 U5438 ( .A1(n6374), .A2(n6836), .ZN(n6183) );
  AOI21_X1 U5439 ( .B1(n10190), .B2(n10188), .A(n10189), .ZN(n10193) );
  INV_X1 U5440 ( .A(n10187), .ZN(n4893) );
  NAND2_X1 U5441 ( .A1(n6800), .A2(n6798), .ZN(n6799) );
  NAND2_X1 U5442 ( .A1(n5173), .A2(n6855), .ZN(n5172) );
  INV_X1 U5443 ( .A(n6800), .ZN(n5173) );
  AND3_X1 U5444 ( .A1(n5172), .A2(n6799), .A3(P2_REG2_REG_7__SCAN_IN), .ZN(
        n7749) );
  NAND2_X1 U5445 ( .A1(n6861), .A2(n6860), .ZN(n7994) );
  OAI21_X1 U5446 ( .B1(n7743), .B2(n7744), .A(n5230), .ZN(n6829) );
  OR2_X1 U5447 ( .A1(n7333), .A2(n10426), .ZN(n5230) );
  AOI21_X1 U5448 ( .B1(n7977), .B2(n7978), .A(n5227), .ZN(n6830) );
  NOR2_X1 U5449 ( .A1(n6867), .A2(n5228), .ZN(n5227) );
  AND2_X1 U5450 ( .A1(n4443), .A2(n5145), .ZN(n8523) );
  NAND2_X1 U5451 ( .A1(n6185), .A2(P2_B_REG_SCAN_IN), .ZN(n6772) );
  OAI21_X1 U5452 ( .B1(n6765), .B2(n7221), .A(n6764), .ZN(n8642) );
  NOR2_X1 U5453 ( .A1(n7223), .A2(n10212), .ZN(n6697) );
  AND2_X1 U5454 ( .A1(n4950), .A2(n6563), .ZN(n8659) );
  NAND2_X1 U5455 ( .A1(n8651), .A2(n6270), .ZN(n4950) );
  OR2_X1 U5456 ( .A1(n6494), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6505) );
  NAND2_X1 U5457 ( .A1(n8735), .A2(n4602), .ZN(n8719) );
  AND2_X1 U5458 ( .A1(n8720), .A2(n6681), .ZN(n4602) );
  AOI21_X1 U5459 ( .B1(n8738), .B2(n6270), .A(n6450), .ZN(n8749) );
  NAND2_X1 U5460 ( .A1(n6674), .A2(n4607), .ZN(n5113) );
  NAND2_X1 U5461 ( .A1(n4719), .A2(n4718), .ZN(n7165) );
  AND2_X1 U5462 ( .A1(n8128), .A2(n7155), .ZN(n6641) );
  AND2_X1 U5463 ( .A1(n4462), .A2(n6284), .ZN(n4951) );
  NAND2_X1 U5464 ( .A1(n6267), .A2(n4462), .ZN(n6319) );
  INV_X1 U5465 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n4953) );
  NAND2_X1 U5466 ( .A1(n4954), .A2(n6239), .ZN(n6252) );
  INV_X1 U5467 ( .A(n6240), .ZN(n4954) );
  NAND2_X1 U5468 ( .A1(n10213), .A2(n7666), .ZN(n7137) );
  NAND2_X1 U5469 ( .A1(n10204), .A2(n7133), .ZN(n7661) );
  NAND2_X1 U5470 ( .A1(n7123), .A2(n7599), .ZN(n10205) );
  INV_X1 U5471 ( .A(n8497), .ZN(n10213) );
  NOR2_X1 U5472 ( .A1(n6171), .A2(n4409), .ZN(n5223) );
  OR2_X1 U5473 ( .A1(n10242), .A2(n7245), .ZN(n6706) );
  NAND4_X1 U5474 ( .A1(n6702), .A2(n6701), .A3(P2_STATE_REG_SCAN_IN), .A4(
        n6700), .ZN(n7521) );
  AND2_X1 U5475 ( .A1(n6704), .A2(n7217), .ZN(n7525) );
  NAND2_X1 U5476 ( .A1(n6527), .A2(n6526), .ZN(n8462) );
  XNOR2_X1 U5477 ( .A(n8679), .B(n8689), .ZN(n4713) );
  NAND2_X1 U5478 ( .A1(n5254), .A2(n6687), .ZN(n8679) );
  NAND2_X1 U5479 ( .A1(n6686), .A2(n5255), .ZN(n5254) );
  NAND2_X1 U5480 ( .A1(n8716), .A2(n7187), .ZN(n5218) );
  OR2_X1 U5481 ( .A1(n8933), .A2(n8749), .ZN(n8715) );
  AND2_X1 U5482 ( .A1(n6461), .A2(n6460), .ZN(n8733) );
  NAND2_X1 U5483 ( .A1(n8744), .A2(n7192), .ZN(n8729) );
  INV_X1 U5484 ( .A(n7178), .ZN(n8759) );
  AOI21_X1 U5485 ( .B1(n5205), .B2(n5208), .A(n5202), .ZN(n5201) );
  INV_X1 U5486 ( .A(n6652), .ZN(n5208) );
  INV_X1 U5487 ( .A(n7183), .ZN(n5202) );
  NAND2_X1 U5488 ( .A1(n8784), .A2(n5205), .ZN(n5203) );
  OR2_X1 U5489 ( .A1(n7217), .A2(n6695), .ZN(n10211) );
  AND2_X1 U5490 ( .A1(n7183), .A2(n7182), .ZN(n8776) );
  NAND2_X1 U5491 ( .A1(n5217), .A2(n5215), .ZN(n8832) );
  INV_X1 U5492 ( .A(n4995), .ZN(n5215) );
  NAND2_X1 U5493 ( .A1(n6641), .A2(n7165), .ZN(n5217) );
  INV_X1 U5494 ( .A(n10211), .ZN(n8825) );
  NAND2_X1 U5495 ( .A1(n6694), .A2(n6693), .ZN(n8829) );
  INV_X1 U5496 ( .A(n8989), .ZN(n6583) );
  INV_X1 U5497 ( .A(n8986), .ZN(n6566) );
  INV_X1 U5498 ( .A(n5314), .ZN(n5312) );
  NOR2_X1 U5499 ( .A1(n5313), .A2(n6159), .ZN(n4853) );
  AND2_X1 U5500 ( .A1(n6151), .A2(n6146), .ZN(n4841) );
  INV_X1 U5501 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6158) );
  INV_X1 U5502 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4896) );
  AND2_X1 U5503 ( .A1(n5824), .A2(n5823), .ZN(n8994) );
  AND2_X1 U5504 ( .A1(n9165), .A2(n9004), .ZN(n4740) );
  AND2_X1 U5505 ( .A1(n9097), .A2(n4902), .ZN(n4899) );
  NAND2_X1 U5506 ( .A1(n7874), .A2(n5345), .ZN(n5344) );
  NOR2_X1 U5507 ( .A1(n5650), .A2(n5346), .ZN(n5345) );
  INV_X1 U5508 ( .A(n5347), .ZN(n5346) );
  INV_X1 U5509 ( .A(n5844), .ZN(n5846) );
  NAND2_X1 U5510 ( .A1(n9156), .A2(n9157), .ZN(n4917) );
  NAND2_X1 U5511 ( .A1(n4887), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6046) );
  INV_X1 U5512 ( .A(n4887), .ZN(n6021) );
  NAND2_X1 U5513 ( .A1(n5537), .A2(n5328), .ZN(n5327) );
  INV_X1 U5514 ( .A(n5538), .ZN(n5328) );
  NAND2_X1 U5515 ( .A1(n5704), .A2(n4806), .ZN(n4803) );
  INV_X1 U5516 ( .A(n5344), .ZN(n4801) );
  INV_X1 U5517 ( .A(n4888), .ZN(n5812) );
  INV_X1 U5518 ( .A(n5668), .ZN(n5687) );
  AOI21_X1 U5519 ( .B1(n4918), .B2(n4920), .A(n4916), .ZN(n4915) );
  OAI21_X1 U5520 ( .B1(n5832), .B2(n5335), .A(n4510), .ZN(n4916) );
  AND2_X1 U5521 ( .A1(n5316), .A2(n4913), .ZN(n4912) );
  INV_X1 U5522 ( .A(n5316), .ZN(n4908) );
  INV_X1 U5523 ( .A(n7882), .ZN(n4911) );
  NAND2_X1 U5524 ( .A1(n4900), .A2(n4902), .ZN(n9126) );
  NAND2_X1 U5525 ( .A1(n9097), .A2(n6035), .ZN(n5331) );
  XNOR2_X1 U5526 ( .A(n4817), .B(n9107), .ZN(n9202) );
  NAND2_X1 U5527 ( .A1(n9202), .A2(n9203), .ZN(n9201) );
  AND2_X1 U5528 ( .A1(n5377), .A2(n9341), .ZN(n5134) );
  NOR2_X1 U5529 ( .A1(n5133), .A2(n9321), .ZN(n5128) );
  NAND2_X1 U5530 ( .A1(n9319), .A2(n9320), .ZN(n5131) );
  NAND2_X1 U5531 ( .A1(n9315), .A2(n9323), .ZN(n5133) );
  NOR2_X1 U5532 ( .A1(n5130), .A2(n5129), .ZN(n5126) );
  NOR2_X1 U5533 ( .A1(n9328), .A2(n9331), .ZN(n5130) );
  INV_X1 U5534 ( .A(n9327), .ZN(n5129) );
  INV_X1 U5535 ( .A(n7358), .ZN(n4776) );
  NAND2_X1 U5536 ( .A1(n5068), .A2(n5067), .ZN(n4775) );
  NAND2_X1 U5537 ( .A1(n7361), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5067) );
  INV_X1 U5538 ( .A(n10097), .ZN(n4757) );
  OR2_X1 U5539 ( .A1(n10093), .A2(n4526), .ZN(n5073) );
  NAND2_X1 U5540 ( .A1(n5073), .A2(n5072), .ZN(n5071) );
  INV_X1 U5541 ( .A(n7369), .ZN(n5072) );
  OR2_X1 U5542 ( .A1(n7396), .A2(n4879), .ZN(n4783) );
  AND2_X1 U5543 ( .A1(n7400), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n4879) );
  AND2_X1 U5544 ( .A1(n7562), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5074) );
  NAND2_X1 U5545 ( .A1(n7775), .A2(n4478), .ZN(n4845) );
  INV_X1 U5546 ( .A(n5060), .ZN(n4759) );
  OR2_X1 U5547 ( .A1(n7776), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5060) );
  NOR2_X1 U5548 ( .A1(n8190), .A2(n5069), .ZN(n9507) );
  AND2_X1 U5549 ( .A1(n8194), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5069) );
  AND2_X1 U5550 ( .A1(n8194), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5059) );
  OR2_X1 U5551 ( .A1(n9517), .A2(n4554), .ZN(n4785) );
  NAND3_X1 U5552 ( .A1(n4772), .A2(n4771), .A3(n10114), .ZN(n10113) );
  AOI21_X1 U5553 ( .B1(n10143), .B2(n4867), .A(n5057), .ZN(n5056) );
  OAI22_X1 U5554 ( .A1(n9553), .A2(n5058), .B1(n9555), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n5057) );
  NAND2_X1 U5555 ( .A1(n4987), .A2(n4985), .ZN(n4640) );
  NAND2_X1 U5556 ( .A1(n4937), .A2(n4936), .ZN(n9615) );
  NOR2_X1 U5557 ( .A1(n9445), .A2(n5373), .ZN(n4936) );
  INV_X1 U5558 ( .A(n4452), .ZN(n5281) );
  OR2_X1 U5559 ( .A1(n9673), .A2(n9688), .ZN(n5286) );
  AND2_X1 U5560 ( .A1(n5295), .A2(n4971), .ZN(n4970) );
  NAND2_X1 U5561 ( .A1(n5293), .A2(n5292), .ZN(n4976) );
  NAND2_X1 U5562 ( .A1(n6979), .A2(n5049), .ZN(n9729) );
  NOR2_X1 U5563 ( .A1(n9731), .A2(n5050), .ZN(n5049) );
  INV_X1 U5564 ( .A(n9281), .ZN(n5050) );
  AOI21_X1 U5565 ( .B1(n5287), .B2(n4423), .A(n4455), .ZN(n4968) );
  INV_X1 U5566 ( .A(n6934), .ZN(n4969) );
  OAI21_X1 U5567 ( .B1(n8149), .B2(n5048), .A(n5045), .ZN(n9811) );
  INV_X1 U5568 ( .A(n7898), .ZN(n5037) );
  INV_X1 U5569 ( .A(n4644), .ZN(n4642) );
  INV_X1 U5570 ( .A(n5569), .ZN(n4643) );
  NAND2_X1 U5571 ( .A1(n6974), .A2(n6973), .ZN(n9227) );
  NAND2_X1 U5572 ( .A1(n4947), .A2(n7695), .ZN(n7572) );
  NAND2_X1 U5573 ( .A1(n5501), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5486) );
  NOR2_X1 U5574 ( .A1(n4475), .A2(n4428), .ZN(n4948) );
  NAND2_X1 U5575 ( .A1(n5777), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5485) );
  NOR2_X1 U5576 ( .A1(n7620), .A2(n9455), .ZN(n7618) );
  NAND2_X1 U5577 ( .A1(n5887), .A2(n5886), .ZN(n9914) );
  INV_X1 U5578 ( .A(n9959), .ZN(n10157) );
  NAND2_X1 U5579 ( .A1(n6092), .A2(n10020), .ZN(n7616) );
  NAND2_X1 U5580 ( .A1(n6089), .A2(n6091), .ZN(n7611) );
  AND2_X1 U5581 ( .A1(n10340), .A2(n5136), .ZN(n5135) );
  XNOR2_X1 U5582 ( .A(n5857), .B(n5856), .ZN(n7641) );
  NAND2_X1 U5583 ( .A1(n5017), .A2(n4453), .ZN(n5857) );
  XNOR2_X1 U5584 ( .A(n4604), .B(n5788), .ZN(n7489) );
  NAND2_X1 U5585 ( .A1(n5762), .A2(n5761), .ZN(n4604) );
  OR2_X1 U5586 ( .A1(n5630), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5662) );
  OR3_X1 U5587 ( .A1(n5616), .A2(P1_IR_REG_7__SCAN_IN), .A3(
        P1_IR_REG_6__SCAN_IN), .ZN(n5630) );
  OAI211_X1 U5588 ( .C1(n5440), .C2(n5475), .A(n5441), .B(n4653), .ZN(n5529)
         );
  INV_X1 U5589 ( .A(n8492), .ZN(n8142) );
  NAND2_X1 U5590 ( .A1(n6744), .A2(n6743), .ZN(n8844) );
  AND2_X1 U5591 ( .A1(n6483), .A2(n6482), .ZN(n8708) );
  AND3_X1 U5592 ( .A1(n6425), .A2(n6424), .A3(n6423), .ZN(n8772) );
  NAND2_X1 U5593 ( .A1(n8390), .A2(n6415), .ZN(n8399) );
  OR2_X1 U5594 ( .A1(n6414), .A2(n8402), .ZN(n6415) );
  INV_X1 U5595 ( .A(n8695), .ZN(n8681) );
  NAND2_X1 U5596 ( .A1(n7509), .A2(n6215), .ZN(n7671) );
  INV_X1 U5597 ( .A(n8454), .ZN(n8473) );
  AND2_X1 U5598 ( .A1(n7791), .A2(n6247), .ZN(n5299) );
  NAND2_X1 U5599 ( .A1(n6597), .A2(n10207), .ZN(n8457) );
  INV_X1 U5600 ( .A(n8457), .ZN(n8481) );
  NAND2_X1 U5601 ( .A1(n6609), .A2(n6608), .ZN(n8484) );
  INV_X1 U5602 ( .A(n8659), .ZN(n8485) );
  NAND2_X1 U5603 ( .A1(n6536), .A2(n6535), .ZN(n8670) );
  NAND2_X1 U5604 ( .A1(n6512), .A2(n6511), .ZN(n8669) );
  INV_X1 U5605 ( .A(n8749), .ZN(n8722) );
  NAND2_X1 U5606 ( .A1(n6439), .A2(n6438), .ZN(n8761) );
  NAND2_X1 U5607 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n6172) );
  NAND2_X1 U5608 ( .A1(n7424), .A2(n6844), .ZN(n10182) );
  NAND2_X1 U5609 ( .A1(n4601), .A2(n4600), .ZN(n7535) );
  INV_X1 U5610 ( .A(n7538), .ZN(n4600) );
  INV_X1 U5611 ( .A(n7537), .ZN(n4601) );
  NAND2_X1 U5612 ( .A1(n7647), .A2(n7646), .ZN(n7645) );
  XNOR2_X1 U5613 ( .A(n6829), .B(n7996), .ZN(n7992) );
  NAND2_X1 U5614 ( .A1(n4676), .A2(n4675), .ZN(n4674) );
  INV_X1 U5615 ( .A(n6830), .ZN(n4676) );
  INV_X1 U5616 ( .A(n5246), .ZN(n6832) );
  NAND2_X1 U5617 ( .A1(n5246), .A2(n8535), .ZN(n5245) );
  OR2_X1 U5618 ( .A1(n8530), .A2(n8887), .ZN(n5240) );
  OAI21_X1 U5619 ( .B1(n8551), .B2(n8550), .A(n8549), .ZN(n8553) );
  NAND2_X1 U5620 ( .A1(n6884), .A2(n6883), .ZN(n8546) );
  OR2_X1 U5621 ( .A1(n5158), .A2(n5159), .ZN(n6820) );
  NAND2_X1 U5622 ( .A1(n5157), .A2(n5155), .ZN(n5158) );
  AOI21_X1 U5623 ( .B1(n8594), .B2(n4444), .A(n5156), .ZN(n5155) );
  NAND2_X1 U5624 ( .A1(n4883), .A2(n4597), .ZN(n4596) );
  INV_X1 U5625 ( .A(n6916), .ZN(n4597) );
  NAND2_X1 U5626 ( .A1(n5232), .A2(n5231), .ZN(n4883) );
  XNOR2_X1 U5627 ( .A(n7076), .B(n7237), .ZN(n8635) );
  NOR2_X1 U5628 ( .A1(n8672), .A2(n4538), .ZN(n4855) );
  NAND2_X1 U5629 ( .A1(n6476), .A2(n6475), .ZN(n8700) );
  AND2_X1 U5630 ( .A1(n10221), .A2(n7597), .ZN(n8804) );
  NAND2_X1 U5631 ( .A1(n7530), .A2(n10207), .ZN(n10221) );
  INV_X2 U5632 ( .A(n10221), .ZN(n10223) );
  INV_X1 U5633 ( .A(n8462), .ZN(n8909) );
  NAND2_X1 U5634 ( .A1(n5002), .A2(n7212), .ZN(n8674) );
  NAND2_X1 U5635 ( .A1(n6649), .A2(n6648), .ZN(n5002) );
  INV_X1 U5636 ( .A(n5349), .ZN(n8055) );
  OAI21_X1 U5637 ( .B1(n7874), .B2(n5350), .A(n5355), .ZN(n5349) );
  INV_X1 U5638 ( .A(n5356), .ZN(n5350) );
  NAND2_X1 U5639 ( .A1(n5871), .A2(n5870), .ZN(n9720) );
  OR2_X1 U5640 ( .A1(n6126), .A2(n6120), .ZN(n9194) );
  NAND2_X1 U5641 ( .A1(n7338), .A2(n6953), .ZN(n4665) );
  NAND2_X1 U5642 ( .A1(n5915), .A2(n5914), .ZN(n9903) );
  INV_X1 U5643 ( .A(n9213), .ZN(n9171) );
  INV_X1 U5644 ( .A(n5498), .ZN(n5499) );
  AND2_X1 U5645 ( .A1(n6118), .A2(n6107), .ZN(n9204) );
  INV_X1 U5646 ( .A(n9194), .ZN(n9210) );
  OR2_X1 U5647 ( .A1(n9601), .A2(n6985), .ZN(n6077) );
  NAND2_X1 U5648 ( .A1(n5924), .A2(n5923), .ZN(n9712) );
  NAND2_X1 U5649 ( .A1(n5878), .A2(n5877), .ZN(n9477) );
  INV_X1 U5650 ( .A(n9919), .ZN(n9780) );
  INV_X1 U5651 ( .A(n9934), .ZN(n9478) );
  NOR2_X1 U5652 ( .A1(n7363), .A2(n7362), .ZN(n7371) );
  NOR2_X1 U5653 ( .A1(n7386), .A2(n7385), .ZN(n7396) );
  AND2_X1 U5654 ( .A1(n5076), .A2(n5075), .ZN(n7554) );
  INV_X1 U5655 ( .A(n7476), .ZN(n5075) );
  NOR2_X1 U5656 ( .A1(n7773), .A2(n7774), .ZN(n7859) );
  AND2_X1 U5657 ( .A1(n4780), .A2(n4779), .ZN(n8190) );
  INV_X1 U5658 ( .A(n7860), .ZN(n4779) );
  NOR2_X1 U5659 ( .A1(n8191), .A2(n8192), .ZN(n9517) );
  NOR2_X1 U5660 ( .A1(n8197), .A2(n8198), .ZN(n9520) );
  OAI21_X1 U5661 ( .B1(n10148), .B2(n10542), .A(n10147), .ZN(n4761) );
  INV_X1 U5662 ( .A(n10144), .ZN(n4762) );
  XNOR2_X1 U5663 ( .A(n9546), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9559) );
  INV_X1 U5664 ( .A(n9567), .ZN(n5182) );
  XNOR2_X1 U5665 ( .A(n4933), .B(n9321), .ZN(n7033) );
  NAND2_X1 U5666 ( .A1(n4660), .A2(n9611), .ZN(n9864) );
  INV_X1 U5667 ( .A(n9607), .ZN(n4660) );
  OR2_X1 U5668 ( .A1(n6108), .A2(n9968), .ZN(n9785) );
  NAND2_X1 U5669 ( .A1(n9855), .A2(n9856), .ZN(n5181) );
  AND2_X1 U5670 ( .A1(n10164), .A2(n10154), .ZN(n9856) );
  NAND2_X1 U5671 ( .A1(n9854), .A2(n9853), .ZN(n9973) );
  NAND2_X1 U5672 ( .A1(n5380), .A2(n6999), .ZN(n7000) );
  INV_X1 U5673 ( .A(n6998), .ZN(n6999) );
  XNOR2_X1 U5674 ( .A(n5461), .B(n5460), .ZN(n5869) );
  INV_X1 U5675 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U5676 ( .A1(n5459), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5461) );
  NOR2_X1 U5677 ( .A1(n10067), .A2(n10066), .ZN(n10275) );
  AND2_X1 U5678 ( .A1(n4990), .A2(n4989), .ZN(n4988) );
  NAND2_X1 U5679 ( .A1(n4991), .A2(n4420), .ZN(n4990) );
  NAND2_X1 U5680 ( .A1(n7141), .A2(n4420), .ZN(n5083) );
  AND2_X1 U5681 ( .A1(n9226), .A2(n6973), .ZN(n4737) );
  MUX2_X1 U5682 ( .A(n7159), .B(n7158), .S(n7217), .Z(n7160) );
  NOR2_X1 U5683 ( .A1(n5212), .A2(n7217), .ZN(n5094) );
  NAND2_X1 U5684 ( .A1(n4425), .A2(n4495), .ZN(n4625) );
  NAND2_X1 U5685 ( .A1(n5117), .A2(n9258), .ZN(n5116) );
  NAND2_X1 U5686 ( .A1(n9259), .A2(n4498), .ZN(n5117) );
  AOI21_X1 U5687 ( .B1(n5085), .B2(n4492), .A(n4612), .ZN(n4611) );
  OR2_X1 U5688 ( .A1(n7113), .A2(n7217), .ZN(n7215) );
  NAND2_X1 U5689 ( .A1(n5141), .A2(n9375), .ZN(n4741) );
  INV_X1 U5690 ( .A(n9377), .ZN(n5140) );
  INV_X1 U5691 ( .A(n7205), .ZN(n4857) );
  INV_X1 U5692 ( .A(n8675), .ZN(n4700) );
  NAND2_X1 U5693 ( .A1(n8549), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5152) );
  NOR2_X1 U5694 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n4965) );
  NAND2_X1 U5695 ( .A1(n10224), .A2(n8498), .ZN(n7132) );
  AOI21_X1 U5696 ( .B1(n5793), .B2(n5531), .A(n5979), .ZN(n4728) );
  NAND2_X1 U5697 ( .A1(n4728), .A2(n4729), .ZN(n4725) );
  INV_X1 U5698 ( .A(n5793), .ZN(n4729) );
  NAND2_X1 U5699 ( .A1(n9294), .A2(n9667), .ZN(n4745) );
  INV_X1 U5700 ( .A(n9296), .ZN(n9295) );
  AND2_X1 U5701 ( .A1(n9631), .A2(n9330), .ZN(n4854) );
  NOR2_X1 U5702 ( .A1(n9293), .A2(n9323), .ZN(n4744) );
  NOR2_X1 U5703 ( .A1(n9859), .A2(n9866), .ZN(n5175) );
  NAND2_X1 U5704 ( .A1(n5910), .A2(n5032), .ZN(n5029) );
  INV_X1 U5705 ( .A(n5985), .ZN(n5034) );
  INV_X1 U5706 ( .A(SI_21_), .ZN(n10399) );
  INV_X1 U5707 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5860) );
  INV_X1 U5708 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5836) );
  INV_X1 U5709 ( .A(n5447), .ZN(n4703) );
  INV_X1 U5710 ( .A(n5546), .ZN(n4664) );
  NAND2_X1 U5711 ( .A1(n4687), .A2(n5447), .ZN(n4661) );
  INV_X1 U5712 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6169) );
  NOR2_X1 U5713 ( .A1(n8372), .A2(n4840), .ZN(n4839) );
  INV_X1 U5714 ( .A(n5309), .ZN(n4840) );
  AND2_X1 U5715 ( .A1(n8350), .A2(n8349), .ZN(n8352) );
  XNOR2_X1 U5716 ( .A(n8462), .B(n6528), .ZN(n6537) );
  NAND2_X1 U5717 ( .A1(n4789), .A2(n4788), .ZN(n7063) );
  AOI21_X1 U5718 ( .B1(n4792), .B2(n4795), .A(n4790), .ZN(n4789) );
  NAND2_X1 U5719 ( .A1(n6765), .A2(n4792), .ZN(n4788) );
  INV_X1 U5720 ( .A(n7086), .ZN(n4790) );
  NAND2_X1 U5721 ( .A1(n4633), .A2(n7237), .ZN(n4632) );
  NAND2_X1 U5722 ( .A1(n4622), .A2(n4619), .ZN(n7234) );
  NOR2_X1 U5723 ( .A1(n4621), .A2(n4620), .ZN(n4619) );
  INV_X1 U5724 ( .A(n7219), .ZN(n4620) );
  NAND2_X1 U5725 ( .A1(n4415), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6182) );
  INV_X1 U5726 ( .A(SI_17_), .ZN(n10409) );
  NOR2_X1 U5727 ( .A1(n6792), .A2(n5147), .ZN(n7429) );
  NOR2_X1 U5728 ( .A1(n5233), .A2(n5164), .ZN(n5163) );
  INV_X1 U5729 ( .A(n4674), .ZN(n4672) );
  INV_X1 U5730 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n4885) );
  INV_X1 U5731 ( .A(n8544), .ZN(n5238) );
  NAND2_X1 U5732 ( .A1(n4580), .A2(n4578), .ZN(n6902) );
  AOI22_X1 U5733 ( .A1(n4583), .A2(n4579), .B1(n4582), .B2(n4585), .ZN(n4578)
         );
  OR2_X1 U5734 ( .A1(n8575), .A2(n4581), .ZN(n4580) );
  NAND2_X1 U5735 ( .A1(n6504), .A2(n4965), .ZN(n6529) );
  INV_X1 U5736 ( .A(n5205), .ZN(n4571) );
  NOR2_X1 U5737 ( .A1(n6677), .A2(n5114), .ZN(n4607) );
  INV_X1 U5738 ( .A(n6673), .ZN(n5114) );
  INV_X1 U5739 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10528) );
  AND2_X1 U5740 ( .A1(n6407), .A2(n6406), .ZN(n6420) );
  NOR2_X1 U5741 ( .A1(n6383), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6407) );
  NOR2_X1 U5742 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n4959) );
  OR2_X1 U5743 ( .A1(n6645), .A2(n4861), .ZN(n6646) );
  NAND2_X1 U5744 ( .A1(n8289), .A2(n7208), .ZN(n4861) );
  INV_X1 U5745 ( .A(n7243), .ZN(n6631) );
  NAND2_X1 U5746 ( .A1(n6155), .A2(n6169), .ZN(n5315) );
  OR2_X1 U5747 ( .A1(n6366), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n6367) );
  OR2_X1 U5748 ( .A1(n6301), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n6291) );
  OR2_X1 U5749 ( .A1(n6248), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n6261) );
  INV_X1 U5750 ( .A(n8053), .ZN(n5348) );
  NOR2_X1 U5751 ( .A1(n5491), .A2(n4928), .ZN(n5495) );
  AND2_X1 U5752 ( .A1(n7695), .A2(n5490), .ZN(n5491) );
  NOR2_X1 U5753 ( .A1(n6057), .A2(n7573), .ZN(n4928) );
  NOR2_X1 U5754 ( .A1(n5738), .A2(n5737), .ZN(n4888) );
  INV_X1 U5755 ( .A(n5952), .ZN(n4922) );
  INV_X1 U5756 ( .A(n9148), .ZN(n4923) );
  NOR2_X1 U5757 ( .A1(n5685), .A2(n5684), .ZN(n5668) );
  NAND2_X1 U5758 ( .A1(n4808), .A2(n4807), .ZN(n6056) );
  NAND2_X1 U5759 ( .A1(n4812), .A2(n6968), .ZN(n4808) );
  AOI21_X1 U5760 ( .B1(n6968), .B2(n5433), .A(n4810), .ZN(n4807) );
  INV_X1 U5761 ( .A(n9335), .ZN(n4812) );
  INV_X1 U5762 ( .A(n5750), .ZN(n4920) );
  NOR2_X1 U5763 ( .A1(n5557), .A2(n5407), .ZN(n5586) );
  OR2_X1 U5764 ( .A1(n7616), .A2(n6102), .ZN(n6123) );
  AND2_X1 U5765 ( .A1(n9383), .A2(n9382), .ZN(n9395) );
  INV_X1 U5766 ( .A(n5014), .ZN(n9417) );
  NAND2_X1 U5767 ( .A1(n4753), .A2(n4754), .ZN(n4756) );
  INV_X1 U5768 ( .A(n10109), .ZN(n4754) );
  NAND2_X1 U5769 ( .A1(n9555), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5058) );
  NOR2_X1 U5770 ( .A1(n10142), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5055) );
  INV_X1 U5771 ( .A(n5058), .ZN(n4867) );
  NAND2_X1 U5772 ( .A1(n4509), .A2(n4986), .ZN(n4984) );
  NOR2_X1 U5773 ( .A1(n9641), .A2(n9625), .ZN(n9598) );
  AND2_X1 U5774 ( .A1(n9424), .A2(n9630), .ZN(n9344) );
  AND2_X1 U5775 ( .A1(n5195), .A2(n5012), .ZN(n5194) );
  INV_X1 U5776 ( .A(n5196), .ZN(n5195) );
  OR2_X1 U5777 ( .A1(n9673), .A2(n9896), .ZN(n5196) );
  NAND2_X1 U5778 ( .A1(n4973), .A2(n4972), .ZN(n4971) );
  INV_X1 U5779 ( .A(n5292), .ZN(n4972) );
  AND2_X1 U5780 ( .A1(n4470), .A2(n6946), .ZN(n5295) );
  NOR2_X1 U5781 ( .A1(n5796), .A2(n5775), .ZN(n5844) );
  NOR2_X1 U5782 ( .A1(n5889), .A2(n5888), .ZN(n4889) );
  INV_X1 U5783 ( .A(n6935), .ZN(n5289) );
  AND2_X1 U5784 ( .A1(n5043), .A2(n9262), .ZN(n5042) );
  NOR2_X1 U5785 ( .A1(n9941), .A2(n9937), .ZN(n5186) );
  NAND2_X1 U5786 ( .A1(n4656), .A2(n9247), .ZN(n9425) );
  INV_X1 U5787 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7482) );
  NOR2_X1 U5788 ( .A1(n9965), .A2(n7968), .ZN(n5178) );
  NAND2_X1 U5789 ( .A1(n6918), .A2(n9072), .ZN(n5115) );
  NAND2_X1 U5790 ( .A1(n7581), .A2(n9490), .ZN(n9348) );
  NAND2_X1 U5791 ( .A1(n9598), .A2(n5175), .ZN(n9592) );
  INV_X1 U5792 ( .A(n9421), .ZN(n6995) );
  NAND2_X1 U5793 ( .A1(n5777), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5541) );
  INV_X1 U5794 ( .A(n7611), .ZN(n7002) );
  NAND2_X1 U5795 ( .A1(n4947), .A2(n7625), .ZN(n9350) );
  OAI21_X1 U5796 ( .B1(n7047), .B2(n7046), .A(n7045), .ZN(n7066) );
  INV_X1 U5797 ( .A(SI_20_), .ZN(n5954) );
  OR2_X1 U5798 ( .A1(n4418), .A2(n4460), .ZN(n5018) );
  AOI21_X1 U5799 ( .B1(n5025), .B2(n4435), .A(n4507), .ZN(n5023) );
  INV_X1 U5800 ( .A(n5025), .ZN(n5024) );
  XNOR2_X1 U5801 ( .A(n5446), .B(SI_5_), .ZN(n5568) );
  NAND2_X1 U5802 ( .A1(n5510), .A2(n10363), .ZN(n5436) );
  OR2_X1 U5803 ( .A1(n5444), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4667) );
  OAI211_X1 U5804 ( .C1(n5444), .C2(P2_DATAO_REG_0__SCAN_IN), .A(SI_0_), .B(
        n5273), .ZN(n5476) );
  INV_X1 U5805 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4649) );
  INV_X1 U5806 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4647) );
  OR2_X1 U5807 ( .A1(n6364), .A2(n6642), .ZN(n6365) );
  AND2_X1 U5808 ( .A1(n4461), .A2(n8364), .ZN(n5309) );
  XNOR2_X1 U5809 ( .A(n7267), .B(n8659), .ZN(n6591) );
  NAND2_X1 U5810 ( .A1(n4825), .A2(n4823), .ZN(n8382) );
  AOI21_X1 U5811 ( .B1(n4827), .B2(n4830), .A(n4824), .ZN(n4823) );
  INV_X1 U5812 ( .A(n8381), .ZN(n4824) );
  NAND2_X1 U5813 ( .A1(n4820), .A2(n6231), .ZN(n7669) );
  NAND2_X1 U5814 ( .A1(n7336), .A2(n7532), .ZN(n7125) );
  INV_X1 U5815 ( .A(n4553), .ZN(n5011) );
  AND2_X1 U5816 ( .A1(n6611), .A2(n6610), .ZN(n8441) );
  OR2_X1 U5817 ( .A1(n6427), .A2(n8772), .ZN(n5361) );
  INV_X1 U5818 ( .A(n8493), .ZN(n7792) );
  INV_X1 U5819 ( .A(n8816), .ZN(n8475) );
  NAND2_X1 U5820 ( .A1(n6209), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4797) );
  NAND2_X1 U5821 ( .A1(n10289), .A2(n4560), .ZN(n10292) );
  NAND2_X1 U5822 ( .A1(n10290), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n10289) );
  NAND2_X1 U5823 ( .A1(n4866), .A2(n4865), .ZN(n6837) );
  OR2_X1 U5824 ( .A1(n6910), .A2(n10169), .ZN(n4866) );
  NAND2_X1 U5825 ( .A1(n6910), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4865) );
  NOR2_X1 U5826 ( .A1(n10167), .A2(n6791), .ZN(n7497) );
  AND2_X1 U5827 ( .A1(n4669), .A2(n7306), .ZN(n4668) );
  INV_X1 U5828 ( .A(n5235), .ZN(n10185) );
  OR2_X1 U5829 ( .A1(n10193), .A2(n6794), .ZN(n6795) );
  INV_X1 U5830 ( .A(n5234), .ZN(n4686) );
  OR2_X1 U5831 ( .A1(n7543), .A2(n7544), .ZN(n6797) );
  OAI21_X1 U5832 ( .B1(n7456), .B2(n6827), .A(n4681), .ZN(n7540) );
  INV_X1 U5833 ( .A(n4682), .ZN(n4681) );
  NAND2_X1 U5834 ( .A1(n7540), .A2(n7541), .ZN(n7539) );
  NAND2_X1 U5835 ( .A1(n7539), .A2(n4884), .ZN(n6828) );
  OR2_X1 U5836 ( .A1(n6851), .A2(n10308), .ZN(n4884) );
  NAND2_X1 U5837 ( .A1(n7750), .A2(n7748), .ZN(n5170) );
  AND2_X1 U5838 ( .A1(n7748), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5171) );
  NAND2_X1 U5839 ( .A1(n7645), .A2(n6857), .ZN(n7746) );
  NOR2_X1 U5840 ( .A1(n7998), .A2(n7999), .ZN(n7997) );
  NAND2_X1 U5841 ( .A1(n4587), .A2(n6865), .ZN(n7980) );
  NAND2_X1 U5842 ( .A1(n5143), .A2(n5145), .ZN(n5142) );
  AND2_X1 U5843 ( .A1(n6808), .A2(n4441), .ZN(n5143) );
  NAND2_X1 U5844 ( .A1(n8522), .A2(n8521), .ZN(n5144) );
  OAI21_X1 U5845 ( .B1(n6810), .B2(n8535), .A(n6811), .ZN(n8536) );
  NOR2_X1 U5846 ( .A1(n8536), .A2(n10468), .ZN(n8551) );
  NAND2_X1 U5847 ( .A1(n6815), .A2(n8579), .ZN(n8565) );
  OAI21_X1 U5848 ( .B1(n6884), .B2(n4590), .A(n4588), .ZN(n8561) );
  INV_X1 U5849 ( .A(n4589), .ZN(n4588) );
  OAI21_X1 U5850 ( .B1(n4590), .B2(n6883), .A(n6888), .ZN(n4589) );
  NAND2_X1 U5851 ( .A1(n5168), .A2(n5167), .ZN(n8581) );
  AOI21_X1 U5852 ( .B1(n8579), .B2(n8791), .A(n4552), .ZN(n5167) );
  NAND2_X1 U5853 ( .A1(n5166), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8564) );
  INV_X1 U5854 ( .A(n8565), .ZN(n5166) );
  NAND2_X1 U5855 ( .A1(n6902), .A2(n6903), .ZN(n8612) );
  INV_X1 U5856 ( .A(n6819), .ZN(n5156) );
  NAND2_X1 U5857 ( .A1(n6557), .A2(n6556), .ZN(n6602) );
  OR2_X1 U5858 ( .A1(n6602), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8624) );
  AOI21_X1 U5859 ( .B1(n5269), .B2(n4515), .A(n4436), .ZN(n5267) );
  NOR2_X1 U5860 ( .A1(n6727), .A2(n5270), .ZN(n5269) );
  AND2_X1 U5861 ( .A1(n4439), .A2(n4961), .ZN(n4960) );
  INV_X1 U5862 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n4961) );
  NAND2_X1 U5863 ( .A1(n6445), .A2(n4439), .ZN(n6467) );
  OR2_X1 U5864 ( .A1(n6432), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6446) );
  NAND2_X1 U5865 ( .A1(n6445), .A2(n6444), .ZN(n6455) );
  NAND2_X1 U5866 ( .A1(n6420), .A2(n10528), .ZN(n6432) );
  NAND2_X1 U5867 ( .A1(n6344), .A2(n6343), .ZN(n6358) );
  NAND2_X1 U5868 ( .A1(n6344), .A2(n4959), .ZN(n6372) );
  OR2_X1 U5869 ( .A1(n6296), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6345) );
  OR2_X1 U5870 ( .A1(n6306), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U5871 ( .A1(n6267), .A2(n6266), .ZN(n6317) );
  NAND2_X1 U5872 ( .A1(n6216), .A2(n6217), .ZN(n6240) );
  NAND2_X1 U5873 ( .A1(n5106), .A2(n6658), .ZN(n7631) );
  INV_X1 U5874 ( .A(n7602), .ZN(n7600) );
  NAND2_X1 U5875 ( .A1(n7600), .A2(n6634), .ZN(n7599) );
  NAND2_X1 U5876 ( .A1(n7528), .A2(n7527), .ZN(n7530) );
  INV_X1 U5877 ( .A(n6646), .ZN(n8684) );
  NAND2_X1 U5878 ( .A1(n5218), .A2(n4419), .ZN(n8287) );
  NOR2_X1 U5879 ( .A1(n8623), .A2(n8622), .ZN(n8899) );
  NAND2_X1 U5880 ( .A1(n5252), .A2(n5256), .ZN(n5250) );
  INV_X1 U5881 ( .A(n5252), .ZN(n5251) );
  NAND2_X1 U5882 ( .A1(n6674), .A2(n6673), .ZN(n8785) );
  OR2_X1 U5883 ( .A1(n8785), .A2(n8783), .ZN(n8786) );
  NAND2_X1 U5884 ( .A1(n4573), .A2(n7173), .ZN(n8803) );
  AND2_X1 U5885 ( .A1(n5210), .A2(n7172), .ZN(n5209) );
  NAND2_X1 U5886 ( .A1(n4705), .A2(n6671), .ZN(n4608) );
  NAND2_X1 U5887 ( .A1(n8231), .A2(n4474), .ZN(n4705) );
  AND2_X1 U5888 ( .A1(n7176), .A2(n7175), .ZN(n8802) );
  OR2_X1 U5889 ( .A1(n8360), .A2(n8351), .ZN(n8225) );
  NAND2_X1 U5890 ( .A1(n7166), .A2(n7165), .ZN(n8229) );
  INV_X1 U5891 ( .A(n8229), .ZN(n8234) );
  INV_X1 U5892 ( .A(n7824), .ZN(n10243) );
  OR2_X1 U5893 ( .A1(n6587), .A2(n6694), .ZN(n6714) );
  NAND2_X1 U5894 ( .A1(n6579), .A2(n6578), .ZN(n6585) );
  XNOR2_X1 U5895 ( .A(n6314), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7333) );
  OR2_X1 U5896 ( .A1(n6223), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n6232) );
  INV_X1 U5897 ( .A(n6203), .ZN(n6223) );
  NAND2_X1 U5898 ( .A1(n7872), .A2(n7871), .ZN(n5356) );
  NAND2_X1 U5899 ( .A1(n4888), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5814) );
  INV_X1 U5900 ( .A(n9688), .ZN(n9300) );
  INV_X1 U5901 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U5902 ( .A1(n4889), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5917) );
  OR2_X1 U5903 ( .A1(n5917), .A2(n5916), .ZN(n5941) );
  XNOR2_X1 U5904 ( .A(n5948), .B(n8327), .ZN(n5949) );
  NAND2_X1 U5905 ( .A1(n4927), .A2(n4925), .ZN(n9076) );
  NAND2_X1 U5906 ( .A1(n9126), .A2(n6036), .ZN(n9096) );
  INV_X1 U5907 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5775) );
  OR2_X1 U5908 ( .A1(n9104), .A2(n8994), .ZN(n5825) );
  AND2_X1 U5909 ( .A1(n5830), .A2(n5831), .ZN(n5832) );
  INV_X1 U5910 ( .A(n5327), .ZN(n5325) );
  NAND2_X1 U5911 ( .A1(n5320), .A2(n4440), .ZN(n5326) );
  OR2_X1 U5912 ( .A1(n5634), .A2(n7482), .ZN(n5636) );
  NAND2_X1 U5913 ( .A1(n9036), .A2(n4947), .ZN(n5494) );
  AND2_X1 U5914 ( .A1(n7277), .A2(n7276), .ZN(n7279) );
  XOR2_X1 U5915 ( .A(n8327), .B(n5879), .Z(n9028) );
  OAI22_X1 U5916 ( .A1(n9996), .A2(n5979), .B1(n9900), .B2(n6057), .ZN(n5879)
         );
  NAND2_X1 U5917 ( .A1(n5939), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5971) );
  INV_X1 U5918 ( .A(n5941), .ZN(n5939) );
  NAND2_X1 U5919 ( .A1(n5344), .A2(n5341), .ZN(n9176) );
  INV_X1 U5920 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5407) );
  NAND2_X1 U5921 ( .A1(n9096), .A2(n9097), .ZN(n6086) );
  AND2_X1 U5922 ( .A1(n6992), .A2(n6991), .ZN(n7020) );
  AND2_X1 U5923 ( .A1(n6966), .A2(n6965), .ZN(n6967) );
  OR2_X1 U5924 ( .A1(n9045), .A2(n6985), .ZN(n6966) );
  AND4_X1 U5925 ( .A1(n5693), .A2(n5692), .A3(n5691), .A4(n5690), .ZN(n9183)
         );
  NAND2_X1 U5926 ( .A1(n9494), .A2(n7293), .ZN(n7295) );
  XNOR2_X1 U5927 ( .A(n7316), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n7296) );
  AND2_X1 U5928 ( .A1(n7292), .A2(n7291), .ZN(n7360) );
  NAND2_X1 U5929 ( .A1(n7372), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4777) );
  OR2_X1 U5930 ( .A1(n7380), .A2(n4874), .ZN(n4873) );
  NOR2_X1 U5931 ( .A1(n4875), .A2(n5552), .ZN(n4874) );
  INV_X1 U5932 ( .A(n7384), .ZN(n4875) );
  OR2_X1 U5933 ( .A1(n7399), .A2(n4752), .ZN(n4751) );
  AND2_X1 U5934 ( .A1(n7400), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4752) );
  NAND2_X1 U5935 ( .A1(n4783), .A2(n4782), .ZN(n5078) );
  INV_X1 U5936 ( .A(n7397), .ZN(n4782) );
  OR2_X1 U5937 ( .A1(n7478), .A2(n4750), .ZN(n4749) );
  AND2_X1 U5938 ( .A1(n7479), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4750) );
  NAND2_X1 U5939 ( .A1(n5078), .A2(n5077), .ZN(n5076) );
  NAND2_X1 U5940 ( .A1(n7479), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5077) );
  AND2_X1 U5941 ( .A1(n7863), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4781) );
  NAND2_X1 U5942 ( .A1(n4845), .A2(n4541), .ZN(n4870) );
  INV_X1 U5943 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9087) );
  NAND2_X1 U5944 ( .A1(n9504), .A2(n9503), .ZN(n9502) );
  AND2_X1 U5945 ( .A1(n9535), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5065) );
  NOR2_X1 U5946 ( .A1(n9548), .A2(n5064), .ZN(n10110) );
  NOR2_X1 U5947 ( .A1(n9547), .A2(n5080), .ZN(n5064) );
  NAND2_X1 U5948 ( .A1(n4814), .A2(n4813), .ZN(n5769) );
  NOR2_X1 U5949 ( .A1(n4422), .A2(n4508), .ZN(n4813) );
  INV_X1 U5950 ( .A(n5456), .ZN(n4814) );
  NOR2_X1 U5951 ( .A1(n9543), .A2(n5080), .ZN(n5079) );
  NAND2_X1 U5952 ( .A1(n4756), .A2(n4755), .ZN(n10123) );
  AND2_X1 U5953 ( .A1(n10125), .A2(n4877), .ZN(n4755) );
  AOI21_X1 U5954 ( .B1(n4433), .B2(n9586), .A(n4499), .ZN(n5290) );
  NAND2_X1 U5955 ( .A1(n4509), .A2(n9586), .ZN(n5291) );
  AND2_X1 U5956 ( .A1(n6960), .A2(n6111), .ZN(n9588) );
  NOR2_X1 U5957 ( .A1(n4985), .A2(n4984), .ZN(n4983) );
  INV_X1 U5958 ( .A(n4984), .ZN(n4981) );
  NOR2_X1 U5959 ( .A1(n9604), .A2(n4935), .ZN(n4934) );
  INV_X1 U5960 ( .A(n9347), .ZN(n4935) );
  NAND2_X1 U5961 ( .A1(n5193), .A2(n5191), .ZN(n9641) );
  AND2_X1 U5962 ( .A1(n5192), .A2(n5194), .ZN(n5191) );
  NAND2_X1 U5963 ( .A1(n5193), .A2(n5194), .ZN(n9640) );
  NAND2_X1 U5964 ( .A1(n9380), .A2(n5041), .ZN(n5040) );
  INV_X1 U5965 ( .A(n9376), .ZN(n5041) );
  NAND2_X1 U5966 ( .A1(n9709), .A2(n4654), .ZN(n5039) );
  OR2_X1 U5967 ( .A1(n9903), .A2(n9893), .ZN(n9685) );
  NOR2_X1 U5968 ( .A1(n9695), .A2(n9896), .ZN(n9677) );
  NAND2_X1 U5969 ( .A1(n5844), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5889) );
  INV_X1 U5970 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5888) );
  INV_X1 U5971 ( .A(n4889), .ZN(n5891) );
  INV_X1 U5972 ( .A(n9279), .ZN(n9747) );
  NAND2_X1 U5973 ( .A1(n8154), .A2(n5184), .ZN(n9783) );
  NAND2_X1 U5974 ( .A1(n8154), .A2(n6996), .ZN(n9824) );
  NAND2_X1 U5975 ( .A1(n8152), .A2(n6934), .ZN(n9821) );
  NAND2_X1 U5976 ( .A1(n9821), .A2(n9820), .ZN(n9819) );
  INV_X1 U5977 ( .A(n8154), .ZN(n9823) );
  NAND2_X1 U5978 ( .A1(n4639), .A2(n6930), .ZN(n8039) );
  NAND2_X1 U5979 ( .A1(n7896), .A2(n5178), .ZN(n8110) );
  NAND2_X1 U5980 ( .A1(n7896), .A2(n8058), .ZN(n8112) );
  NAND2_X1 U5981 ( .A1(n7888), .A2(n4645), .ZN(n9223) );
  NAND2_X1 U5982 ( .A1(n9227), .A2(n9354), .ZN(n9225) );
  NAND2_X1 U5983 ( .A1(n4944), .A2(n4946), .ZN(n4943) );
  OR2_X1 U5984 ( .A1(n7888), .A2(n7710), .ZN(n5189) );
  NAND2_X1 U5985 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5555) );
  NAND2_X1 U5986 ( .A1(n7576), .A2(n5115), .ZN(n7590) );
  AND4_X1 U5987 ( .A1(n5528), .A2(n5527), .A3(n5526), .A4(n5525), .ZN(n6922)
         );
  NAND2_X1 U5988 ( .A1(n4731), .A2(n4730), .ZN(n7576) );
  INV_X1 U5989 ( .A(n7574), .ZN(n4730) );
  INV_X1 U5990 ( .A(n6970), .ZN(n4731) );
  NAND2_X1 U5991 ( .A1(n9217), .A2(n9216), .ZN(n9331) );
  NOR2_X1 U5992 ( .A1(n6120), .A2(n6995), .ZN(n9877) );
  NAND2_X1 U5993 ( .A1(n8165), .A2(n6953), .ZN(n5013) );
  NAND2_X1 U5994 ( .A1(n7489), .A2(n6953), .ZN(n4727) );
  AND4_X1 U5995 ( .A1(n5720), .A2(n5719), .A3(n5718), .A4(n5717), .ZN(n9944)
         );
  AND4_X1 U5996 ( .A1(n5418), .A2(n5417), .A3(n5416), .A4(n5415), .ZN(n7897)
         );
  INV_X1 U5997 ( .A(n4978), .ZN(n4977) );
  NAND2_X1 U5998 ( .A1(n6953), .A2(n7308), .ZN(n4979) );
  XNOR2_X1 U5999 ( .A(n7066), .B(n7065), .ZN(n9218) );
  XNOR2_X1 U6000 ( .A(n7047), .B(n6752), .ZN(n8974) );
  AOI21_X1 U6001 ( .B1(n6742), .B2(n6741), .A(n5358), .ZN(n6747) );
  INV_X1 U6002 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5340) );
  XNOR2_X1 U6003 ( .A(n6552), .B(n6735), .ZN(n8980) );
  XNOR2_X1 U6004 ( .A(n5424), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U6005 ( .A1(n5423), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5424) );
  XNOR2_X1 U6006 ( .A(n6066), .B(n6065), .ZN(n8984) );
  XNOR2_X1 U6007 ( .A(n5422), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6087) );
  INV_X1 U6008 ( .A(n5994), .ZN(n5991) );
  XNOR2_X1 U6009 ( .A(n6105), .B(n6104), .ZN(n7286) );
  AND2_X1 U6010 ( .A1(n6103), .A2(n5465), .ZN(n9405) );
  NAND2_X1 U6011 ( .A1(n5031), .A2(n5960), .ZN(n5986) );
  NAND2_X1 U6012 ( .A1(n5035), .A2(n5032), .ZN(n5031) );
  OAI21_X1 U6013 ( .B1(n5840), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5884) );
  OR2_X1 U6014 ( .A1(n5769), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U6015 ( .A1(n5019), .A2(n5022), .ZN(n5833) );
  NOR2_X1 U6016 ( .A1(n5456), .A2(n4422), .ZN(n5789) );
  NOR2_X1 U6017 ( .A1(n5456), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5733) );
  NAND2_X1 U6018 ( .A1(n5272), .A2(n5656), .ZN(n5705) );
  OAI21_X1 U6019 ( .B1(n5602), .B2(n5261), .A(n5259), .ZN(n4666) );
  NAND2_X1 U6020 ( .A1(n5258), .A2(n5604), .ZN(n5629) );
  NAND2_X1 U6021 ( .A1(n5602), .A2(n5601), .ZN(n5258) );
  INV_X1 U6022 ( .A(n4687), .ZN(n5445) );
  OR2_X1 U6023 ( .A1(n5451), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5563) );
  OR2_X1 U6024 ( .A1(n5444), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5434) );
  NAND2_X1 U6025 ( .A1(n5444), .A2(n4721), .ZN(n4720) );
  NAND2_X1 U6026 ( .A1(n4897), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5053) );
  NAND2_X1 U6027 ( .A1(n5053), .A2(n5507), .ZN(n5532) );
  NAND2_X1 U6028 ( .A1(n7446), .A2(n4895), .ZN(n7509) );
  AND2_X1 U6029 ( .A1(n7510), .A2(n6202), .ZN(n4895) );
  XNOR2_X1 U6030 ( .A(n6213), .B(n8497), .ZN(n7510) );
  NAND2_X1 U6031 ( .A1(n5310), .A2(n5309), .ZN(n8418) );
  AND2_X1 U6032 ( .A1(n7263), .A2(n7262), .ZN(n7264) );
  AND2_X1 U6033 ( .A1(n7268), .A2(n8470), .ZN(n7262) );
  AND4_X1 U6034 ( .A1(n6311), .A2(n6310), .A3(n6309), .A4(n6308), .ZN(n8180)
         );
  NAND2_X1 U6035 ( .A1(n7598), .A2(n6186), .ZN(n7415) );
  INV_X1 U6036 ( .A(n8669), .ZN(n8386) );
  INV_X1 U6037 ( .A(n4832), .ZN(n4831) );
  OAI21_X1 U6038 ( .B1(n5007), .B2(n4834), .A(n6390), .ZN(n4832) );
  NAND2_X1 U6039 ( .A1(n8298), .A2(n6501), .ZN(n4826) );
  OR2_X1 U6040 ( .A1(n6601), .A2(n6610), .ZN(n8454) );
  NAND2_X1 U6041 ( .A1(n5006), .A2(n5009), .ZN(n8167) );
  NAND2_X1 U6042 ( .A1(n8119), .A2(n8117), .ZN(n5006) );
  OAI21_X1 U6043 ( .B1(n8119), .B2(n5011), .A(n8117), .ZN(n8169) );
  NAND2_X1 U6044 ( .A1(n8373), .A2(n6474), .ZN(n8426) );
  INV_X1 U6045 ( .A(n8441), .ZN(n8476) );
  NAND2_X1 U6046 ( .A1(n7447), .A2(n7448), .ZN(n7446) );
  NAND2_X1 U6047 ( .A1(n5301), .A2(n5300), .ZN(n8471) );
  XNOR2_X1 U6048 ( .A(n6586), .B(P2_IR_REG_22__SCAN_IN), .ZN(n7250) );
  NAND2_X1 U6049 ( .A1(n6585), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6586) );
  NAND2_X1 U6050 ( .A1(n4628), .A2(n4629), .ZN(n7242) );
  AND2_X1 U6051 ( .A1(n5087), .A2(n4695), .ZN(n4693) );
  INV_X1 U6052 ( .A(n7244), .ZN(n5087) );
  INV_X1 U6053 ( .A(n7241), .ZN(n4696) );
  NAND2_X1 U6054 ( .A1(n6500), .A2(n6499), .ZN(n8695) );
  INV_X1 U6055 ( .A(n8733), .ZN(n8488) );
  OAI211_X1 U6056 ( .C1(n7058), .C2(n6816), .A(n6413), .B(n6412), .ZN(n8789)
         );
  INV_X1 U6057 ( .A(n8180), .ZN(n8491) );
  NAND4_X1 U6058 ( .A1(n6323), .A2(n6322), .A3(n6321), .A4(n6320), .ZN(n8492)
         );
  NAND2_X1 U6059 ( .A1(n7508), .A2(n10250), .ZN(n5248) );
  OR2_X1 U6060 ( .A1(n7508), .A2(n10250), .ZN(n5249) );
  NAND2_X1 U6061 ( .A1(n7503), .A2(n6841), .ZN(n7426) );
  OAI21_X1 U6062 ( .B1(n10182), .B2(n10183), .A(n6846), .ZN(n7465) );
  OAI211_X1 U6063 ( .C1(n5235), .C2(n6847), .A(n4685), .B(n4683), .ZN(n7456)
         );
  NAND2_X1 U6064 ( .A1(n5233), .A2(n4686), .ZN(n4685) );
  NAND2_X1 U6065 ( .A1(n5235), .A2(n4684), .ZN(n4683) );
  NOR2_X1 U6066 ( .A1(n5233), .A2(n4686), .ZN(n4684) );
  NAND2_X1 U6067 ( .A1(n7535), .A2(n6853), .ZN(n7647) );
  NAND2_X1 U6068 ( .A1(n5172), .A2(n6799), .ZN(n7648) );
  AND2_X1 U6069 ( .A1(n5170), .A2(n5169), .ZN(n7752) );
  OAI21_X1 U6070 ( .B1(n7997), .B2(n7984), .A(n7983), .ZN(n7986) );
  NAND2_X1 U6071 ( .A1(n6808), .A2(n5145), .ZN(n8502) );
  XNOR2_X1 U6072 ( .A(n6833), .B(n6899), .ZN(n8587) );
  NAND2_X1 U6073 ( .A1(n4586), .A2(n6897), .ZN(n8591) );
  NAND2_X1 U6074 ( .A1(n8575), .A2(n8574), .ZN(n4586) );
  OR2_X1 U6075 ( .A1(n4528), .A2(n5159), .ZN(n8605) );
  OR2_X1 U6076 ( .A1(n6899), .A2(n10436), .ZN(n4678) );
  AND2_X1 U6077 ( .A1(n6899), .A2(n10436), .ZN(n4677) );
  OAI211_X1 U6078 ( .C1(n8177), .C2(n8635), .A(n6775), .B(n6774), .ZN(n8628)
         );
  INV_X1 U6079 ( .A(n4791), .ZN(n8644) );
  AOI21_X1 U6080 ( .B1(n6765), .B2(n6764), .A(n4795), .ZN(n4791) );
  NOR2_X1 U6081 ( .A1(n6697), .A2(n6696), .ZN(n6698) );
  XNOR2_X1 U6082 ( .A(n6728), .B(n4621), .ZN(n6699) );
  NOR2_X1 U6083 ( .A1(n8465), .A2(n10211), .ZN(n6696) );
  NAND2_X1 U6084 ( .A1(n5000), .A2(n4434), .ZN(n8660) );
  NAND2_X1 U6085 ( .A1(n5001), .A2(n4427), .ZN(n5000) );
  INV_X1 U6086 ( .A(n6649), .ZN(n5001) );
  AND2_X1 U6087 ( .A1(n8735), .A2(n6681), .ZN(n8721) );
  NAND2_X1 U6088 ( .A1(n5220), .A2(n7190), .ZN(n8742) );
  NAND2_X1 U6089 ( .A1(n5203), .A2(n4446), .ZN(n5220) );
  NAND2_X1 U6090 ( .A1(n5265), .A2(n6678), .ZN(n8748) );
  NAND2_X1 U6091 ( .A1(n5214), .A2(n7165), .ZN(n8834) );
  OR2_X1 U6092 ( .A1(n6641), .A2(n6640), .ZN(n5214) );
  NAND2_X1 U6093 ( .A1(n5200), .A2(n7137), .ZN(n7636) );
  NAND2_X1 U6094 ( .A1(n7661), .A2(n7663), .ZN(n5200) );
  NAND2_X1 U6095 ( .A1(n6206), .A2(n5004), .ZN(n7666) );
  OR2_X1 U6096 ( .A1(n10242), .A2(n7595), .ZN(n10206) );
  NAND2_X1 U6097 ( .A1(n6185), .A2(n4467), .ZN(n5224) );
  INV_X1 U6098 ( .A(n8711), .ZN(n8838) );
  INV_X1 U6099 ( .A(n6653), .ZN(n7532) );
  NAND2_X1 U6100 ( .A1(n6596), .A2(n7332), .ZN(n10207) );
  OR2_X1 U6101 ( .A1(n7530), .A2(n10206), .ZN(n8711) );
  AND2_X1 U6102 ( .A1(n6264), .A2(n6263), .ZN(n7957) );
  NOR2_X1 U6103 ( .A1(n7521), .A2(n6711), .ZN(n10254) );
  AOI21_X1 U6104 ( .B1(n10245), .B2(n8654), .A(n8650), .ZN(n6721) );
  INV_X1 U6105 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n4708) );
  NAND2_X1 U6106 ( .A1(n4712), .A2(n4710), .ZN(n8916) );
  AOI21_X1 U6107 ( .B1(n8486), .B2(n8826), .A(n4711), .ZN(n4710) );
  NAND2_X1 U6108 ( .A1(n4713), .A2(n8829), .ZN(n4712) );
  NOR2_X1 U6109 ( .A1(n8681), .A2(n10211), .ZN(n4711) );
  NAND2_X1 U6110 ( .A1(n6686), .A2(n6685), .ZN(n8291) );
  NAND2_X1 U6111 ( .A1(n5218), .A2(n7195), .ZN(n8704) );
  NAND2_X1 U6112 ( .A1(n6443), .A2(n6442), .ZN(n8933) );
  NAND2_X1 U6113 ( .A1(n6680), .A2(n6679), .ZN(n8730) );
  NAND2_X1 U6114 ( .A1(n6431), .A2(n6430), .ZN(n8938) );
  NAND2_X1 U6115 ( .A1(n6419), .A2(n6418), .ZN(n8941) );
  NAND2_X1 U6116 ( .A1(n7641), .A2(n6278), .ZN(n6419) );
  NAND2_X1 U6117 ( .A1(n5203), .A2(n5201), .ZN(n8755) );
  NAND2_X1 U6118 ( .A1(n5204), .A2(n6652), .ZN(n8777) );
  NAND2_X1 U6119 ( .A1(n8784), .A2(n6651), .ZN(n5204) );
  NAND2_X1 U6120 ( .A1(n7489), .A2(n6278), .ZN(n4603) );
  NAND2_X1 U6121 ( .A1(n8832), .A2(n7169), .ZN(n8808) );
  NAND2_X1 U6122 ( .A1(n10247), .A2(n10245), .ZN(n8967) );
  INV_X1 U6123 ( .A(n7957), .ZN(n8033) );
  OAI22_X1 U6124 ( .A1(n6565), .A2(P2_D_REG_1__SCAN_IN), .B1(n6583), .B2(n6566), .ZN(n7522) );
  XNOR2_X1 U6125 ( .A(n6581), .B(n6580), .ZN(n7353) );
  INV_X1 U6126 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6580) );
  OAI21_X1 U6127 ( .B1(n6585), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6581) );
  NOR2_X1 U6128 ( .A1(n5090), .A2(n5089), .ZN(n5088) );
  NOR2_X1 U6129 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5089) );
  NOR2_X1 U6130 ( .A1(n5444), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8982) );
  XNOR2_X1 U6131 ( .A(n6156), .B(n6155), .ZN(n8986) );
  NAND2_X1 U6132 ( .A1(n6154), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6156) );
  NAND2_X1 U6133 ( .A1(n6152), .A2(n6154), .ZN(n8989) );
  MUX2_X1 U6134 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6148), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6152) );
  AND2_X1 U6135 ( .A1(n6147), .A2(n4535), .ZN(n4862) );
  OR2_X1 U6136 ( .A1(n6145), .A2(n6146), .ZN(n4863) );
  INV_X1 U6137 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n10520) );
  AND2_X1 U6138 ( .A1(P2_U3151), .A2(n5444), .ZN(n8976) );
  INV_X1 U6139 ( .A(n7250), .ZN(n8085) );
  INV_X1 U6140 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8087) );
  INV_X1 U6141 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8081) );
  NAND2_X1 U6142 ( .A1(n6164), .A2(n6163), .ZN(n7936) );
  MUX2_X1 U6143 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6162), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n6164) );
  OR2_X1 U6144 ( .A1(n6161), .A2(n6159), .ZN(n6162) );
  XNOR2_X1 U6145 ( .A(n6167), .B(n6166), .ZN(n7857) );
  INV_X1 U6146 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6166) );
  INV_X1 U6147 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10487) );
  INV_X1 U6148 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7691) );
  INV_X1 U6149 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7516) );
  INV_X1 U6150 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7438) );
  INV_X1 U6151 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10330) );
  INV_X1 U6152 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7341) );
  INV_X1 U6153 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7335) );
  NAND2_X1 U6154 ( .A1(n5444), .A2(SI_0_), .ZN(n6184) );
  NAND2_X1 U6155 ( .A1(n8339), .A2(n5330), .ZN(n4905) );
  AND2_X1 U6156 ( .A1(n5643), .A2(n5642), .ZN(n9058) );
  XNOR2_X1 U6157 ( .A(n5949), .B(n4850), .ZN(n9079) );
  INV_X1 U6158 ( .A(n5950), .ZN(n4850) );
  NAND2_X1 U6159 ( .A1(n4927), .A2(n9147), .ZN(n9078) );
  AND4_X1 U6160 ( .A1(n5675), .A2(n5674), .A3(n5673), .A4(n5672), .ZN(n9091)
         );
  OAI21_X1 U6161 ( .B1(n5341), .B2(n4806), .A(n5704), .ZN(n4804) );
  NAND2_X1 U6162 ( .A1(n9201), .A2(n4816), .ZN(n9111) );
  AND2_X1 U6163 ( .A1(n5318), .A2(n4912), .ZN(n7881) );
  NAND2_X1 U6164 ( .A1(n5318), .A2(n5316), .ZN(n4906) );
  NAND2_X1 U6165 ( .A1(n5336), .A2(n5832), .ZN(n9118) );
  NAND2_X1 U6166 ( .A1(n8995), .A2(n5386), .ZN(n5336) );
  NAND2_X1 U6167 ( .A1(n4901), .A2(n9004), .ZN(n9127) );
  NAND2_X1 U6168 ( .A1(n9005), .A2(n9003), .ZN(n4901) );
  AND2_X1 U6169 ( .A1(n6046), .A2(n6022), .ZN(n9637) );
  NAND2_X1 U6170 ( .A1(n5326), .A2(n5327), .ZN(n7813) );
  AOI21_X1 U6171 ( .B1(n4801), .B2(n4505), .A(n4798), .ZN(n5727) );
  NOR2_X1 U6172 ( .A1(n5571), .A2(n4911), .ZN(n4910) );
  NAND2_X1 U6173 ( .A1(n4908), .A2(n5571), .ZN(n4907) );
  AND2_X1 U6174 ( .A1(n5121), .A2(n5126), .ZN(n4886) );
  INV_X1 U6175 ( .A(n6967), .ZN(n9584) );
  INV_X1 U6176 ( .A(n9609), .ZN(n9476) );
  OR2_X1 U6177 ( .A1(n9622), .A2(n6985), .ZN(n6052) );
  OR2_X1 U6178 ( .A1(n5799), .A2(n5798), .ZN(n9803) );
  INV_X1 U6179 ( .A(n9944), .ZN(n9479) );
  INV_X1 U6180 ( .A(n9183), .ZN(n9481) );
  INV_X1 U6181 ( .A(n7897), .ZN(n9484) );
  NAND2_X1 U6182 ( .A1(n5501), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U6183 ( .A1(n5777), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5560) );
  INV_X1 U6184 ( .A(n6922), .ZN(n9487) );
  AOI21_X1 U6185 ( .B1(n7361), .B2(P1_REG2_REG_2__SCAN_IN), .A(n7360), .ZN(
        n7363) );
  XNOR2_X1 U6186 ( .A(n7372), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n7362) );
  INV_X1 U6187 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5066) );
  INV_X1 U6188 ( .A(n4775), .ZN(n7359) );
  INV_X1 U6189 ( .A(n4758), .ZN(n10098) );
  INV_X1 U6190 ( .A(n5063), .ZN(n10096) );
  AND2_X1 U6191 ( .A1(n5063), .A2(n5062), .ZN(n7375) );
  NAND2_X1 U6192 ( .A1(n7373), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5062) );
  INV_X1 U6193 ( .A(n5071), .ZN(n7383) );
  INV_X1 U6194 ( .A(n5073), .ZN(n7370) );
  NAND2_X1 U6195 ( .A1(n7384), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5070) );
  AND2_X1 U6196 ( .A1(n4873), .A2(n4872), .ZN(n7399) );
  INV_X1 U6197 ( .A(n7381), .ZN(n4872) );
  INV_X1 U6198 ( .A(n4873), .ZN(n7382) );
  AND2_X1 U6199 ( .A1(n4751), .A2(n7402), .ZN(n7478) );
  INV_X1 U6200 ( .A(n4751), .ZN(n7404) );
  INV_X1 U6201 ( .A(n5078), .ZN(n7475) );
  INV_X1 U6202 ( .A(n4783), .ZN(n7398) );
  AND2_X1 U6203 ( .A1(n4749), .A2(n4748), .ZN(n7561) );
  INV_X1 U6204 ( .A(n7480), .ZN(n4748) );
  INV_X1 U6205 ( .A(n4749), .ZN(n7481) );
  INV_X1 U6206 ( .A(n5076), .ZN(n7477) );
  INV_X1 U6207 ( .A(n4845), .ZN(n7862) );
  NAND2_X1 U6208 ( .A1(n7775), .A2(n5060), .ZN(n7777) );
  INV_X1 U6209 ( .A(n4780), .ZN(n7861) );
  AND2_X1 U6210 ( .A1(n4870), .A2(n4869), .ZN(n8193) );
  INV_X1 U6211 ( .A(n7864), .ZN(n4869) );
  INV_X1 U6212 ( .A(n4870), .ZN(n7865) );
  INV_X1 U6213 ( .A(n9518), .ZN(n4784) );
  INV_X1 U6214 ( .A(n4785), .ZN(n9519) );
  NOR2_X1 U6215 ( .A1(n9520), .A2(n4550), .ZN(n9525) );
  XNOR2_X1 U6216 ( .A(n9543), .B(n5080), .ZN(n9533) );
  INV_X1 U6217 ( .A(n4772), .ZN(n9544) );
  NOR2_X1 U6218 ( .A1(n9536), .A2(n9787), .ZN(n9548) );
  INV_X1 U6219 ( .A(n10100), .ZN(n10146) );
  NAND2_X1 U6220 ( .A1(n9550), .A2(n4774), .ZN(n4773) );
  INV_X1 U6221 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n4774) );
  NAND2_X1 U6222 ( .A1(n4987), .A2(n5276), .ZN(n9614) );
  AND2_X1 U6223 ( .A1(n4937), .A2(n4938), .ZN(n9617) );
  NAND2_X1 U6224 ( .A1(n9666), .A2(n5283), .ZN(n5275) );
  NAND2_X1 U6225 ( .A1(n5285), .A2(n5286), .ZN(n9654) );
  NAND2_X1 U6226 ( .A1(n4410), .A2(n4452), .ZN(n5285) );
  NAND2_X1 U6227 ( .A1(n4976), .A2(n4973), .ZN(n5296) );
  NAND2_X1 U6228 ( .A1(n4976), .A2(n6944), .ZN(n9693) );
  NAND2_X1 U6229 ( .A1(n5293), .A2(n6942), .ZN(n9716) );
  NAND2_X1 U6230 ( .A1(n6979), .A2(n9281), .ZN(n9732) );
  AND3_X1 U6231 ( .A1(n5781), .A2(n5780), .A3(n5779), .ZN(n9919) );
  NAND2_X1 U6232 ( .A1(n4652), .A2(n5287), .ZN(n4967) );
  AND4_X1 U6233 ( .A1(n5744), .A2(n5743), .A3(n5742), .A4(n5741), .ZN(n9934)
         );
  NAND2_X1 U6234 ( .A1(n8149), .A2(n9250), .ZN(n9813) );
  INV_X1 U6235 ( .A(n9837), .ZN(n9763) );
  INV_X1 U6236 ( .A(n9847), .ZN(n9809) );
  NAND2_X1 U6237 ( .A1(n9842), .A2(n5869), .ZN(n9840) );
  INV_X1 U6238 ( .A(n9785), .ZN(n9836) );
  INV_X1 U6239 ( .A(n9840), .ZN(n9807) );
  NAND2_X1 U6240 ( .A1(n7617), .A2(n9785), .ZN(n9842) );
  NAND2_X1 U6241 ( .A1(n4644), .A2(n5569), .ZN(n7888) );
  INV_X1 U6242 ( .A(n9331), .ZN(n9972) );
  OAI21_X1 U6243 ( .B1(n9867), .B2(n10157), .A(n4658), .ZN(n9978) );
  AND2_X1 U6244 ( .A1(n9866), .A2(n10154), .ZN(n4659) );
  INV_X1 U6245 ( .A(n9720), .ZN(n9996) );
  INV_X1 U6246 ( .A(n8074), .ZN(n10017) );
  INV_X1 U6247 ( .A(n7888), .ZN(n7840) );
  XNOR2_X1 U6248 ( .A(n6747), .B(n6746), .ZN(n8977) );
  INV_X1 U6249 ( .A(n6091), .ZN(n10033) );
  INV_X1 U6250 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5426) );
  INV_X1 U6251 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10038) );
  INV_X1 U6252 ( .A(n6087), .ZN(n10041) );
  OR2_X1 U6253 ( .A1(n7286), .A2(P1_U3086), .ZN(n9456) );
  INV_X1 U6254 ( .A(n9405), .ZN(n9465) );
  INV_X1 U6255 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8090) );
  INV_X1 U6256 ( .A(n9464), .ZN(n8088) );
  INV_X1 U6257 ( .A(n5399), .ZN(n5419) );
  INV_X1 U6258 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7962) );
  INV_X1 U6259 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8319) );
  XNOR2_X1 U6260 ( .A(n5665), .B(P1_IR_REG_11__SCAN_IN), .ZN(n8194) );
  XNOR2_X1 U6261 ( .A(n5617), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7776) );
  XNOR2_X1 U6262 ( .A(n5631), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7562) );
  NAND2_X1 U6263 ( .A1(n4871), .A2(n5532), .ZN(n7316) );
  OR2_X1 U6264 ( .A1(n5053), .A2(n5507), .ZN(n4871) );
  NAND2_X1 U6265 ( .A1(n5444), .A2(n4401), .ZN(n10037) );
  NOR2_X1 U6266 ( .A1(n5444), .A2(n5487), .ZN(n5489) );
  NOR2_X1 U6267 ( .A1(n10061), .A2(n10060), .ZN(n10281) );
  NOR2_X1 U6268 ( .A1(n10065), .A2(n10064), .ZN(n10277) );
  NOR2_X1 U6269 ( .A1(n10069), .A2(n10068), .ZN(n10273) );
  INV_X1 U6270 ( .A(n4891), .ZN(n4890) );
  OAI21_X1 U6271 ( .B1(n8909), .B2(n8481), .A(n8469), .ZN(n4891) );
  OAI21_X1 U6272 ( .B1(n8499), .B2(n6831), .A(n4674), .ZN(n8514) );
  NAND2_X1 U6273 ( .A1(n5245), .A2(n5240), .ZN(n8543) );
  NAND2_X1 U6274 ( .A1(n4595), .A2(n4497), .ZN(P2_U3201) );
  AND2_X1 U6275 ( .A1(n8910), .A2(n4855), .ZN(n8678) );
  NAND2_X1 U6276 ( .A1(n4709), .A2(n4706), .ZN(P2_U3451) );
  NOR2_X1 U6277 ( .A1(n8919), .A2(n4707), .ZN(n4706) );
  NAND2_X1 U6278 ( .A1(n8916), .A2(n10247), .ZN(n4709) );
  NOR2_X1 U6279 ( .A1(n10247), .A2(n4708), .ZN(n4707) );
  AOI21_X1 U6280 ( .B1(n7699), .B2(n7698), .A(n4421), .ZN(n7784) );
  AOI22_X1 U6281 ( .A1(n9210), .A2(n4947), .B1(n9489), .B2(n9192), .ZN(n9073)
         );
  NAND2_X1 U6282 ( .A1(P1_U3973), .A2(n4947), .ZN(n7471) );
  OAI211_X1 U6283 ( .C1(n4456), .C2(n4846), .A(n4762), .B(n4760), .ZN(P1_U3261) );
  NOR2_X1 U6284 ( .A1(n4556), .A2(n4761), .ZN(n4760) );
  NAND2_X1 U6285 ( .A1(n4847), .A2(n10127), .ZN(n4846) );
  NAND2_X1 U6286 ( .A1(n9559), .A2(n4557), .ZN(n4767) );
  NAND2_X1 U6287 ( .A1(n5181), .A2(n5180), .ZN(n5179) );
  NAND2_X1 U6288 ( .A1(n10162), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5180) );
  OAI22_X1 U6289 ( .A1(n5174), .A2(n9962), .B1(n10164), .B2(n10496), .ZN(n7007) );
  OAI21_X1 U6290 ( .B1(n7038), .B2(n10016), .A(n7037), .ZN(n7039) );
  NOR2_X1 U6291 ( .A1(n5174), .A2(n10016), .ZN(n7011) );
  NAND2_X1 U6292 ( .A1(n5022), .A2(n4519), .ZN(n4418) );
  INV_X1 U6293 ( .A(n9321), .ZN(n5132) );
  INV_X1 U6294 ( .A(n7165), .ZN(n5212) );
  AND2_X1 U6295 ( .A1(n6369), .A2(n6380), .ZN(n6886) );
  AND2_X1 U6296 ( .A1(n7200), .A2(n7195), .ZN(n4419) );
  AND2_X1 U6297 ( .A1(n5522), .A2(n5521), .ZN(n4421) );
  INV_X1 U6298 ( .A(n9119), .ZN(n5335) );
  NAND2_X1 U6299 ( .A1(n5457), .A2(n4815), .ZN(n4422) );
  OR2_X1 U6300 ( .A1(n5289), .A2(n4969), .ZN(n4423) );
  NAND2_X1 U6301 ( .A1(n7174), .A2(n8802), .ZN(n4424) );
  INV_X1 U6302 ( .A(n9625), .ZN(n9982) );
  NAND2_X1 U6303 ( .A1(n6044), .A2(n6043), .ZN(n9625) );
  OAI21_X1 U6304 ( .B1(n5601), .B2(n5261), .A(n5610), .ZN(n5260) );
  INV_X1 U6305 ( .A(n9313), .ZN(n5120) );
  INV_X1 U6306 ( .A(n6764), .ZN(n4793) );
  AND3_X1 U6307 ( .A1(n8759), .A2(n7177), .A3(n8783), .ZN(n4425) );
  AND4_X1 U6308 ( .A1(n5398), .A2(n5397), .A3(n10302), .A4(n5463), .ZN(n4426)
         );
  AND2_X1 U6309 ( .A1(n7213), .A2(n7212), .ZN(n4427) );
  NAND2_X1 U6310 ( .A1(n5013), .A2(n5996), .ZN(n9656) );
  INV_X1 U6311 ( .A(n9656), .ZN(n5012) );
  AND2_X1 U6312 ( .A1(n5558), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n4428) );
  NOR2_X1 U6313 ( .A1(n5279), .A2(n6950), .ZN(n4429) );
  AND3_X1 U6314 ( .A1(n9267), .A2(n9742), .A3(n9266), .ZN(n4430) );
  AND4_X1 U6315 ( .A1(n7103), .A2(n8689), .A3(n5103), .A4(n4700), .ZN(n4431)
         );
  AND4_X1 U6316 ( .A1(n6290), .A2(n6289), .A3(n6288), .A4(n6287), .ZN(n8357)
         );
  INV_X1 U6317 ( .A(n8357), .ZN(n4718) );
  AND4_X1 U6318 ( .A1(n5641), .A2(n5640), .A3(n5639), .A4(n5638), .ZN(n9142)
         );
  INV_X1 U6319 ( .A(n9142), .ZN(n5051) );
  AND2_X1 U6320 ( .A1(n5175), .A2(n5174), .ZN(n4432) );
  NOR2_X1 U6321 ( .A1(n9866), .A2(n4412), .ZN(n4433) );
  AND2_X1 U6322 ( .A1(n8168), .A2(n5010), .ZN(n5009) );
  AND2_X1 U6323 ( .A1(n4787), .A2(n7113), .ZN(n4434) );
  AND2_X1 U6324 ( .A1(n4957), .A2(n6764), .ZN(n7220) );
  INV_X1 U6325 ( .A(n7220), .ZN(n4621) );
  NAND2_X1 U6326 ( .A1(n5271), .A2(n5754), .ZN(n4435) );
  AND2_X1 U6327 ( .A1(n6726), .A2(n8659), .ZN(n4436) );
  INV_X1 U6328 ( .A(n8070), .ZN(n4940) );
  NAND2_X1 U6329 ( .A1(n6379), .A2(n8475), .ZN(n4437) );
  AND2_X1 U6330 ( .A1(n7241), .A2(n7595), .ZN(n4438) );
  INV_X1 U6331 ( .A(n4945), .ZN(n4944) );
  OAI21_X1 U6332 ( .B1(n6973), .B2(n4946), .A(n9226), .ZN(n4945) );
  INV_X1 U6333 ( .A(n7306), .ZN(n5247) );
  INV_X1 U6334 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10583) );
  AND2_X1 U6335 ( .A1(n6444), .A2(n4962), .ZN(n4439) );
  AND2_X1 U6336 ( .A1(n5321), .A2(n5322), .ZN(n4440) );
  AND2_X1 U6337 ( .A1(n6523), .A2(n6522), .ZN(n8680) );
  INV_X1 U6338 ( .A(n8680), .ZN(n8486) );
  AND2_X1 U6339 ( .A1(n8521), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4441) );
  AND2_X1 U6340 ( .A1(n5154), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4442) );
  AND2_X1 U6341 ( .A1(n6808), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4443) );
  NAND2_X1 U6342 ( .A1(n7682), .A2(n7848), .ZN(n7681) );
  AND2_X1 U6343 ( .A1(n5161), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4444) );
  OR2_X1 U6344 ( .A1(n7620), .A2(n9400), .ZN(n9822) );
  INV_X1 U6345 ( .A(n9822), .ZN(n9784) );
  INV_X1 U6346 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6503) );
  INV_X1 U6347 ( .A(n5869), .ZN(n9556) );
  AND3_X1 U6348 ( .A1(n6256), .A2(n6255), .A3(n6254), .ZN(n4445) );
  NAND2_X1 U6349 ( .A1(n5984), .A2(n9165), .ZN(n9005) );
  INV_X1 U6350 ( .A(n4795), .ZN(n4794) );
  NAND2_X1 U6351 ( .A1(n4796), .A2(n8641), .ZN(n4795) );
  NAND2_X1 U6352 ( .A1(n4915), .A2(n4914), .ZN(n9024) );
  INV_X1 U6353 ( .A(n8694), .ZN(n5103) );
  AND2_X1 U6354 ( .A1(n5201), .A2(n7180), .ZN(n4446) );
  AND2_X1 U6355 ( .A1(n9735), .A2(n9739), .ZN(n9717) );
  AND2_X1 U6356 ( .A1(n8418), .A2(n4864), .ZN(n4447) );
  INV_X1 U6357 ( .A(n9297), .ZN(n9667) );
  AND2_X1 U6358 ( .A1(n4826), .A2(n6514), .ZN(n4448) );
  OR2_X1 U6359 ( .A1(n9695), .A2(n5196), .ZN(n4449) );
  NAND2_X1 U6360 ( .A1(n4432), .A2(n9598), .ZN(n4450) );
  AND2_X1 U6361 ( .A1(n6211), .A2(n4797), .ZN(n4451) );
  NAND2_X1 U6362 ( .A1(n9673), .A2(n9688), .ZN(n4452) );
  INV_X1 U6363 ( .A(n5288), .ZN(n5287) );
  INV_X1 U6364 ( .A(n9364), .ZN(n5048) );
  INV_X1 U6365 ( .A(n5352), .ZN(n5351) );
  OAI21_X1 U6366 ( .B1(n5353), .B2(n5356), .A(n4555), .ZN(n5352) );
  NAND2_X1 U6367 ( .A1(n5572), .A2(n5573), .ZN(n5355) );
  AND2_X1 U6368 ( .A1(n5018), .A2(n5835), .ZN(n4453) );
  OR2_X1 U6369 ( .A1(n6817), .A2(n8594), .ZN(n5160) );
  INV_X1 U6370 ( .A(n6847), .ZN(n5233) );
  NAND2_X1 U6371 ( .A1(n5399), .A2(n4426), .ZN(n5423) );
  OR2_X1 U6372 ( .A1(n7157), .A2(n7950), .ZN(n4454) );
  NOR2_X1 U6373 ( .A1(n9937), .A2(n9779), .ZN(n4455) );
  AND2_X1 U6374 ( .A1(n8715), .A2(n7193), .ZN(n8731) );
  AND2_X1 U6375 ( .A1(n9554), .A2(n9553), .ZN(n4456) );
  OR2_X1 U6376 ( .A1(n4403), .A2(n4860), .ZN(n4457) );
  INV_X1 U6377 ( .A(n9633), .ZN(n9608) );
  NAND2_X1 U6378 ( .A1(n6052), .A2(n6051), .ZN(n9633) );
  AND4_X1 U6379 ( .A1(n6135), .A2(n6134), .A3(n6233), .A4(n6204), .ZN(n4458)
         );
  AND3_X1 U6380 ( .A1(n9136), .A2(n9058), .A3(n9056), .ZN(n4459) );
  NOR2_X1 U6381 ( .A1(n5766), .A2(n5020), .ZN(n4460) );
  NAND2_X1 U6382 ( .A1(n6440), .A2(n8732), .ZN(n4461) );
  AND2_X1 U6383 ( .A1(n6266), .A2(n4952), .ZN(n4462) );
  AND2_X1 U6384 ( .A1(n5405), .A2(n10022), .ZN(n5412) );
  AND2_X1 U6385 ( .A1(n7812), .A2(n7848), .ZN(n4463) );
  NAND2_X1 U6386 ( .A1(n9819), .A2(n6935), .ZN(n9794) );
  NAND2_X1 U6387 ( .A1(n5275), .A2(n5280), .ZN(n9635) );
  AND3_X1 U6388 ( .A1(n9376), .A2(n9330), .A3(n9284), .ZN(n4464) );
  NAND2_X1 U6389 ( .A1(n5296), .A2(n6946), .ZN(n9676) );
  NAND2_X1 U6390 ( .A1(n4967), .A2(n4968), .ZN(n9772) );
  INV_X1 U6391 ( .A(n9097), .ZN(n5332) );
  NAND2_X1 U6392 ( .A1(n6957), .A2(n6956), .ZN(n9578) );
  INV_X1 U6393 ( .A(n9578), .ZN(n5174) );
  AND2_X1 U6394 ( .A1(n7915), .A2(n7140), .ZN(n4465) );
  OR2_X1 U6395 ( .A1(n9865), .A2(n4659), .ZN(n4466) );
  AND2_X1 U6396 ( .A1(n4409), .A2(n4997), .ZN(n4467) );
  OR2_X1 U6397 ( .A1(n6185), .A2(n7306), .ZN(n4468) );
  INV_X1 U6398 ( .A(n5979), .ZN(n9041) );
  NAND2_X1 U6399 ( .A1(n6106), .A2(n7704), .ZN(n5979) );
  NAND2_X1 U6400 ( .A1(n8232), .A2(n6670), .ZN(n8231) );
  INV_X1 U6401 ( .A(n7594), .ZN(n8082) );
  AND2_X1 U6402 ( .A1(n4805), .A2(n9086), .ZN(n4469) );
  OR2_X1 U6403 ( .A1(n9694), .A2(n9903), .ZN(n9695) );
  INV_X1 U6404 ( .A(n9695), .ZN(n5193) );
  AND2_X1 U6405 ( .A1(n5585), .A2(n5584), .ZN(n8058) );
  INV_X1 U6406 ( .A(n8058), .ZN(n7968) );
  OR2_X1 U6407 ( .A1(n9896), .A2(n9702), .ZN(n4470) );
  AND2_X1 U6408 ( .A1(n8938), .A2(n8761), .ZN(n4471) );
  NAND2_X1 U6409 ( .A1(n6003), .A2(n6002), .ZN(n9876) );
  OR2_X1 U6410 ( .A1(n9720), .A2(n9477), .ZN(n4472) );
  NOR2_X1 U6411 ( .A1(n8453), .A2(n5311), .ZN(n4473) );
  NAND2_X1 U6412 ( .A1(n4727), .A2(n5793), .ZN(n9789) );
  AND2_X1 U6413 ( .A1(n8810), .A2(n8809), .ZN(n4474) );
  NOR2_X1 U6414 ( .A1(n4408), .A2(n5483), .ZN(n4475) );
  INV_X1 U6415 ( .A(n9393), .ZN(n5016) );
  OR2_X1 U6416 ( .A1(n8497), .A2(n7666), .ZN(n4476) );
  INV_X1 U6417 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n10340) );
  AND2_X1 U6418 ( .A1(n7144), .A2(n7145), .ZN(n4477) );
  NOR2_X1 U6419 ( .A1(n7778), .A2(n4759), .ZN(n4478) );
  NOR2_X1 U6420 ( .A1(n6943), .A2(n5294), .ZN(n4479) );
  AND2_X1 U6421 ( .A1(n9385), .A2(n9667), .ZN(n4480) );
  NAND2_X1 U6422 ( .A1(n5016), .A2(n9311), .ZN(n4481) );
  INV_X1 U6423 ( .A(n5283), .ZN(n5282) );
  NOR2_X1 U6424 ( .A1(n6949), .A2(n5284), .ZN(n5283) );
  AND2_X1 U6425 ( .A1(n5160), .A2(n8603), .ZN(n4482) );
  AND2_X1 U6426 ( .A1(n9447), .A2(n9394), .ZN(n4483) );
  INV_X1 U6427 ( .A(n7169), .ZN(n5213) );
  OR2_X1 U6428 ( .A1(n6839), .A2(n10250), .ZN(n4484) );
  AND2_X1 U6429 ( .A1(n5463), .A2(n6104), .ZN(n4485) );
  INV_X1 U6430 ( .A(n5355), .ZN(n5353) );
  NAND2_X1 U6431 ( .A1(n8494), .A2(n8064), .ZN(n4486) );
  NAND2_X1 U6432 ( .A1(n4917), .A2(n5750), .ZN(n8995) );
  AND2_X1 U6433 ( .A1(n6484), .A2(n6474), .ZN(n4487) );
  AND2_X1 U6434 ( .A1(n7148), .A2(n7138), .ZN(n4488) );
  AND2_X1 U6435 ( .A1(n5981), .A2(n5952), .ZN(n4489) );
  INV_X1 U6436 ( .A(n5979), .ZN(n5490) );
  AND2_X1 U6437 ( .A1(n4852), .A2(n6679), .ZN(n4490) );
  AND2_X1 U6438 ( .A1(n8844), .A2(n7223), .ZN(n4491) );
  OR2_X1 U6439 ( .A1(n4614), .A2(n4613), .ZN(n4492) );
  AND2_X1 U6440 ( .A1(n9656), .A2(n9876), .ZN(n4493) );
  AND2_X1 U6441 ( .A1(n5040), .A2(n4480), .ZN(n4494) );
  AND2_X1 U6442 ( .A1(n4627), .A2(n4424), .ZN(n4495) );
  AND4_X1 U6443 ( .A1(n7215), .A2(n7214), .A3(n7213), .A4(n7212), .ZN(n4496)
         );
  NAND2_X1 U6444 ( .A1(n6822), .A2(n10191), .ZN(n4497) );
  NAND2_X1 U6445 ( .A1(n9256), .A2(n9255), .ZN(n4498) );
  AND2_X1 U6446 ( .A1(n9280), .A2(n9376), .ZN(n9710) );
  INV_X1 U6447 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5313) );
  INV_X1 U6448 ( .A(n9445), .ZN(n9616) );
  NAND2_X1 U6449 ( .A1(n9347), .A2(n9388), .ZN(n9445) );
  INV_X1 U6450 ( .A(n5330), .ZN(n5329) );
  NAND2_X1 U6451 ( .A1(n6085), .A2(n5331), .ZN(n5330) );
  INV_X1 U6452 ( .A(n5277), .ZN(n5276) );
  OAI21_X1 U6453 ( .B1(n6950), .B2(n5278), .A(n6951), .ZN(n5277) );
  NOR2_X1 U6454 ( .A1(n9859), .A2(n9476), .ZN(n4499) );
  INV_X1 U6455 ( .A(n5256), .ZN(n5255) );
  OR2_X1 U6456 ( .A1(n6688), .A2(n5257), .ZN(n5256) );
  AND2_X1 U6457 ( .A1(n9789), .A2(n9803), .ZN(n4500) );
  AND2_X1 U6458 ( .A1(n8360), .A2(n8490), .ZN(n4501) );
  OR2_X1 U6459 ( .A1(n5354), .A2(n4459), .ZN(n4502) );
  INV_X1 U6460 ( .A(n5359), .ZN(n5323) );
  OR2_X1 U6461 ( .A1(n4407), .A2(n10184), .ZN(n4503) );
  AND2_X1 U6462 ( .A1(n8901), .A2(n7239), .ZN(n4504) );
  AND2_X1 U6463 ( .A1(n4803), .A2(n9086), .ZN(n4505) );
  OR2_X1 U6464 ( .A1(n9636), .A2(n4854), .ZN(n4506) );
  AND2_X1 U6465 ( .A1(n5758), .A2(SI_13_), .ZN(n4507) );
  OR2_X1 U6466 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4508) );
  INV_X1 U6467 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U6468 ( .A1(n9866), .A2(n4412), .ZN(n4509) );
  INV_X1 U6469 ( .A(n4974), .ZN(n4973) );
  OR2_X1 U6470 ( .A1(n6945), .A2(n4975), .ZN(n4974) );
  NAND2_X1 U6471 ( .A1(n5855), .A2(n5854), .ZN(n4510) );
  INV_X1 U6472 ( .A(n5086), .ZN(n5085) );
  NAND2_X1 U6473 ( .A1(n8715), .A2(n7192), .ZN(n5086) );
  INV_X1 U6474 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10021) );
  AND2_X1 U6475 ( .A1(n5314), .A2(n5313), .ZN(n4511) );
  NAND2_X1 U6476 ( .A1(n9972), .A2(n9419), .ZN(n4512) );
  NAND2_X1 U6477 ( .A1(n5302), .A2(n6365), .ZN(n4513) );
  NAND2_X1 U6478 ( .A1(n9598), .A2(n9600), .ZN(n9590) );
  XOR2_X1 U6479 ( .A(n7240), .B(n8623), .Z(n4514) );
  NOR2_X1 U6480 ( .A1(n8462), .A2(n8670), .ZN(n4515) );
  AND2_X1 U6481 ( .A1(n7372), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4516) );
  INV_X1 U6482 ( .A(n7229), .ZN(n4701) );
  XNOR2_X1 U6483 ( .A(n8893), .B(n8815), .ZN(n8833) );
  OR2_X1 U6484 ( .A1(n9310), .A2(n9393), .ZN(n4517) );
  OR2_X1 U6485 ( .A1(n9789), .A2(n9803), .ZN(n4518) );
  OR2_X1 U6486 ( .A1(n5834), .A2(SI_16_), .ZN(n4519) );
  AND2_X1 U6487 ( .A1(n5034), .A2(n5960), .ZN(n4520) );
  NOR2_X1 U6488 ( .A1(n4408), .A2(n5552), .ZN(n4521) );
  INV_X1 U6489 ( .A(n9673), .ZN(n9990) );
  NAND2_X1 U6490 ( .A1(n5968), .A2(n5967), .ZN(n9673) );
  NOR2_X1 U6491 ( .A1(n9544), .A2(n5079), .ZN(n4522) );
  NAND2_X1 U6492 ( .A1(n8659), .A2(n6725), .ZN(n6764) );
  AND2_X1 U6493 ( .A1(n9259), .A2(n9254), .ZN(n4523) );
  NOR2_X1 U6494 ( .A1(n5163), .A2(n5233), .ZN(n4524) );
  AND2_X1 U6495 ( .A1(n7170), .A2(n8814), .ZN(n4525) );
  AND2_X1 U6496 ( .A1(n9394), .A2(n9309), .ZN(n9446) );
  INV_X1 U6497 ( .A(n9446), .ZN(n4932) );
  AND2_X1 U6498 ( .A1(n7373), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n4526) );
  NAND2_X1 U6499 ( .A1(n8462), .A2(n8465), .ZN(n4527) );
  AND2_X1 U6500 ( .A1(n5160), .A2(n4444), .ZN(n4528) );
  NAND3_X1 U6501 ( .A1(n5562), .A2(n5561), .A3(n5560), .ZN(n9485) );
  NAND2_X1 U6502 ( .A1(n8496), .A2(n7673), .ZN(n4529) );
  INV_X1 U6503 ( .A(n5699), .ZN(n4806) );
  NOR2_X1 U6504 ( .A1(n5376), .A2(n5698), .ZN(n5699) );
  NOR2_X1 U6505 ( .A1(n5251), .A2(n5103), .ZN(n5102) );
  AND2_X1 U6506 ( .A1(n5310), .A2(n4461), .ZN(n4530) );
  NAND2_X1 U6507 ( .A1(n9855), .A2(n9566), .ZN(n4531) );
  AND2_X1 U6508 ( .A1(n5450), .A2(n5340), .ZN(n4532) );
  OR2_X1 U6509 ( .A1(n6185), .A2(n7508), .ZN(n4533) );
  NAND2_X1 U6510 ( .A1(n4979), .A2(n4977), .ZN(n10153) );
  INV_X1 U6511 ( .A(n10153), .ZN(n7812) );
  AND2_X1 U6512 ( .A1(n4453), .A2(n5021), .ZN(n4534) );
  INV_X1 U6513 ( .A(n5300), .ZN(n4834) );
  AND2_X1 U6514 ( .A1(n8472), .A2(n4437), .ZN(n5300) );
  INV_X1 U6515 ( .A(n5373), .ZN(n4938) );
  OR2_X1 U6516 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4535) );
  NOR2_X1 U6517 ( .A1(n6847), .A2(n5164), .ZN(n4536) );
  INV_X1 U6518 ( .A(n6106), .ZN(n4810) );
  AND2_X1 U6519 ( .A1(n5250), .A2(n6689), .ZN(n5104) );
  INV_X1 U6520 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10297) );
  INV_X1 U6521 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6155) );
  INV_X1 U6522 ( .A(n8283), .ZN(n7038) );
  NAND2_X1 U6523 ( .A1(n7019), .A2(n7018), .ZN(n8283) );
  INV_X2 U6524 ( .A(n9842), .ZN(n9827) );
  INV_X1 U6525 ( .A(n6891), .ZN(n5242) );
  OR2_X1 U6526 ( .A1(n7010), .A2(n7616), .ZN(n10162) );
  NAND2_X1 U6527 ( .A1(n4835), .A2(n5007), .ZN(n5301) );
  NAND2_X1 U6528 ( .A1(n6338), .A2(n6337), .ZN(n8119) );
  OAI21_X1 U6529 ( .B1(n7874), .B2(n5352), .A(n5347), .ZN(n9055) );
  INV_X1 U6530 ( .A(n10179), .ZN(n5221) );
  AND2_X1 U6531 ( .A1(n8154), .A2(n5186), .ZN(n4537) );
  NAND2_X1 U6532 ( .A1(n6555), .A2(n6554), .ZN(n6725) );
  INV_X1 U6533 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4721) );
  INV_X1 U6534 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n4860) );
  AND2_X1 U6535 ( .A1(n8673), .A2(n8821), .ZN(n4538) );
  NAND2_X1 U6536 ( .A1(n4608), .A2(n7089), .ZN(n8795) );
  NAND2_X1 U6537 ( .A1(n5109), .A2(n6668), .ZN(n8178) );
  OR2_X1 U6538 ( .A1(n4802), .A2(n4804), .ZN(n9085) );
  INV_X1 U6539 ( .A(n6644), .ZN(n8723) );
  INV_X1 U6540 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5164) );
  XNOR2_X1 U6541 ( .A(n6340), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6876) );
  NAND2_X1 U6542 ( .A1(n6513), .A2(n8386), .ZN(n8380) );
  INV_X1 U6543 ( .A(n8380), .ZN(n4828) );
  INV_X1 U6544 ( .A(n6980), .ZN(n5192) );
  AND2_X1 U6545 ( .A1(n7062), .A2(n7061), .ZN(n8623) );
  OR2_X1 U6546 ( .A1(n9513), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n4539) );
  AND2_X1 U6547 ( .A1(n8015), .A2(n9254), .ZN(n4540) );
  NAND2_X1 U6548 ( .A1(n7863), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4541) );
  INV_X1 U6549 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4997) );
  AND2_X1 U6550 ( .A1(n4906), .A2(n5571), .ZN(n4542) );
  INV_X1 U6551 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6343) );
  INV_X1 U6552 ( .A(n5704), .ZN(n4805) );
  OR2_X1 U6553 ( .A1(n6876), .A2(n4885), .ZN(n4543) );
  OR2_X1 U6554 ( .A1(n7699), .A2(n4421), .ZN(n5320) );
  INV_X2 U6555 ( .A(n4420), .ZN(n7217) );
  AND2_X1 U6556 ( .A1(n4959), .A2(n4958), .ZN(n4544) );
  AND2_X1 U6557 ( .A1(n5326), .A2(n5324), .ZN(n4545) );
  AND2_X1 U6558 ( .A1(n5144), .A2(n5142), .ZN(n4546) );
  INV_X1 U6559 ( .A(n4992), .ZN(n6149) );
  AND2_X1 U6560 ( .A1(n7721), .A2(n6247), .ZN(n4547) );
  AND2_X1 U6561 ( .A1(n5301), .A2(n4437), .ZN(n4548) );
  INV_X1 U6562 ( .A(n9549), .ZN(n5080) );
  INV_X1 U6563 ( .A(n10197), .ZN(n5231) );
  NAND2_X1 U6564 ( .A1(n6590), .A2(n6589), .ZN(n8470) );
  NAND2_X1 U6565 ( .A1(n6283), .A2(n6282), .ZN(n8447) );
  INV_X1 U6566 ( .A(n8447), .ZN(n4719) );
  AND2_X1 U6567 ( .A1(n7682), .A2(n4463), .ZN(n4549) );
  AND2_X1 U6568 ( .A1(n9521), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4550) );
  OR2_X1 U6569 ( .A1(n10092), .A2(n7294), .ZN(n10137) );
  OR2_X1 U6570 ( .A1(n10092), .A2(n7289), .ZN(n10141) );
  INV_X1 U6571 ( .A(n8829), .ZN(n10218) );
  OR2_X1 U6572 ( .A1(n10128), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n4551) );
  INV_X1 U6573 ( .A(n8826), .ZN(n10212) );
  AND2_X1 U6574 ( .A1(n4420), .A2(n6695), .ZN(n8826) );
  XOR2_X1 U6575 ( .A(n8578), .B(n6816), .Z(n4552) );
  OR2_X1 U6576 ( .A1(n6351), .A2(n8815), .ZN(n4553) );
  NAND2_X1 U6577 ( .A1(n5773), .A2(n5772), .ZN(n9925) );
  INV_X1 U6578 ( .A(n9925), .ZN(n5187) );
  AND2_X1 U6579 ( .A1(n9521), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n4554) );
  OR2_X1 U6580 ( .A1(n5599), .A2(n5598), .ZN(n4555) );
  NAND2_X1 U6581 ( .A1(n5633), .A2(n5632), .ZN(n9965) );
  INV_X1 U6582 ( .A(n9965), .ZN(n5052) );
  AND2_X1 U6583 ( .A1(n10146), .A2(n10145), .ZN(n4556) );
  AND2_X1 U6584 ( .A1(n10131), .A2(n9556), .ZN(n4557) );
  AND2_X1 U6585 ( .A1(n9535), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n4558) );
  OR2_X1 U6586 ( .A1(n9513), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4559) );
  OR2_X1 U6587 ( .A1(n10290), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n4560) );
  INV_X1 U6588 ( .A(n6901), .ZN(n4585) );
  OAI21_X1 U6589 ( .B1(n10148), .B2(n4648), .A(n9560), .ZN(n4868) );
  INV_X1 U6590 ( .A(n5190), .ZN(n7682) );
  OR2_X1 U6591 ( .A1(n7587), .A2(n7710), .ZN(n5190) );
  AND2_X1 U6592 ( .A1(n5771), .A2(n5840), .ZN(n10112) );
  INV_X2 U6593 ( .A(n10162), .ZN(n10164) );
  AND2_X1 U6594 ( .A1(n7446), .A2(n6202), .ZN(n4561) );
  INV_X1 U6595 ( .A(n8602), .ZN(n5161) );
  INV_X1 U6596 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6217) );
  INV_X1 U6597 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5136) );
  INV_X1 U6598 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n4958) );
  INV_X1 U6599 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n4952) );
  NAND2_X1 U6600 ( .A1(n7295), .A2(n7296), .ZN(n5068) );
  OR2_X1 U6601 ( .A1(n8610), .A2(n6436), .ZN(n4562) );
  INV_X1 U6602 ( .A(n4877), .ZN(n4876) );
  NAND2_X1 U6603 ( .A1(n10112), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4877) );
  INV_X1 U6604 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4764) );
  NAND3_X1 U6605 ( .A1(n4511), .A2(n4992), .A3(n5365), .ZN(n8970) );
  INV_X1 U6606 ( .A(n8970), .ZN(n5090) );
  INV_X1 U6607 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n4851) );
  INV_X1 U6608 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5274) );
  INV_X1 U6609 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4648) );
  INV_X1 U6610 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5228) );
  NAND3_X1 U6611 ( .A1(n4563), .A2(n4565), .A3(n4427), .ZN(n4568) );
  NAND3_X1 U6612 ( .A1(n4568), .A2(n4434), .A3(n4527), .ZN(n4999) );
  INV_X1 U6613 ( .A(n8784), .ZN(n4569) );
  NAND2_X1 U6614 ( .A1(n4569), .A2(n4446), .ZN(n4572) );
  NAND3_X1 U6615 ( .A1(n4572), .A2(n5219), .A3(n4570), .ZN(n8744) );
  NAND2_X1 U6616 ( .A1(n8803), .A2(n7175), .ZN(n4993) );
  NAND2_X1 U6617 ( .A1(n4574), .A2(n5209), .ZN(n4573) );
  NAND2_X1 U6618 ( .A1(n8128), .A2(n4575), .ZN(n4574) );
  NAND2_X1 U6619 ( .A1(n7661), .A2(n4576), .ZN(n5197) );
  AND2_X1 U6620 ( .A1(n7663), .A2(n7138), .ZN(n4576) );
  NAND2_X1 U6621 ( .A1(n8496), .A2(n10235), .ZN(n7138) );
  NAND2_X2 U6622 ( .A1(n5091), .A2(n5088), .ZN(n5307) );
  OAI21_X2 U6623 ( .B1(n6765), .B2(n4795), .A(n4792), .ZN(n7076) );
  NAND2_X1 U6624 ( .A1(n7980), .A2(n7979), .ZN(n6870) );
  NAND2_X1 U6625 ( .A1(n7994), .A2(n7993), .ZN(n4587) );
  NAND2_X1 U6626 ( .A1(n8561), .A2(n8560), .ZN(n6893) );
  AND2_X1 U6627 ( .A1(n4458), .A2(n6203), .ZN(n6279) );
  NOR2_X1 U6628 ( .A1(n6140), .A2(n6139), .ZN(n4594) );
  INV_X1 U6629 ( .A(n6140), .ZN(n4592) );
  NAND4_X1 U6630 ( .A1(n5365), .A2(n6279), .A3(n4594), .A4(n6155), .ZN(n4593)
         );
  NOR2_X1 U6631 ( .A1(n8628), .A2(n6776), .ZN(n6782) );
  MUX2_X1 U6632 ( .A(n5611), .B(n7341), .S(n5444), .Z(n5613) );
  NAND3_X1 U6633 ( .A1(n4646), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4605) );
  NAND3_X1 U6634 ( .A1(n4648), .A2(n4649), .A3(n4647), .ZN(n4606) );
  NAND3_X1 U6635 ( .A1(n4722), .A2(n4716), .A3(n5651), .ZN(n5680) );
  NAND3_X1 U6636 ( .A1(n5368), .A2(n4717), .A3(n4723), .ZN(n4716) );
  OAI21_X1 U6637 ( .B1(n7191), .B2(n5086), .A(n4611), .ZN(n4618) );
  NAND2_X1 U6638 ( .A1(n4615), .A2(n7199), .ZN(n7207) );
  NAND3_X1 U6639 ( .A1(n4617), .A2(n7195), .A3(n4616), .ZN(n4615) );
  NAND2_X1 U6640 ( .A1(n4618), .A2(n4420), .ZN(n4617) );
  NAND2_X1 U6641 ( .A1(n4623), .A2(n8661), .ZN(n4622) );
  NAND2_X1 U6642 ( .A1(n4624), .A2(n7216), .ZN(n4623) );
  NAND2_X1 U6643 ( .A1(n4856), .A2(n4496), .ZN(n4624) );
  NAND3_X1 U6644 ( .A1(n5092), .A2(n4425), .A3(n4627), .ZN(n4626) );
  NAND3_X1 U6645 ( .A1(n4628), .A2(n4629), .A3(n7243), .ZN(n4694) );
  NAND2_X1 U6646 ( .A1(n7230), .A2(n7228), .ZN(n4628) );
  INV_X1 U6647 ( .A(n7604), .ZN(n7336) );
  OAI21_X1 U6648 ( .B1(n4637), .B2(n7147), .A(n7217), .ZN(n4882) );
  OAI21_X1 U6649 ( .B1(n8100), .B2(n8102), .A(n4639), .ZN(n9963) );
  NAND2_X1 U6650 ( .A1(n8100), .A2(n8102), .ZN(n4639) );
  NAND2_X2 U6651 ( .A1(n6948), .A2(n6947), .ZN(n9666) );
  OAI21_X1 U6652 ( .B1(n4642), .B2(n4643), .A(n4645), .ZN(n4641) );
  NAND3_X1 U6653 ( .A1(n4644), .A2(n9485), .A3(n5569), .ZN(n9355) );
  NAND2_X1 U6654 ( .A1(n7311), .A2(n6953), .ZN(n4644) );
  INV_X1 U6655 ( .A(n8152), .ZN(n4652) );
  NAND2_X1 U6656 ( .A1(n4651), .A2(n4650), .ZN(n9758) );
  NAND3_X1 U6657 ( .A1(n5438), .A2(n5439), .A3(n5508), .ZN(n4653) );
  NAND2_X2 U6658 ( .A1(n9765), .A2(n9766), .ZN(n9764) );
  INV_X1 U6659 ( .A(n9380), .ZN(n4655) );
  NAND2_X1 U6660 ( .A1(n9243), .A2(n9237), .ZN(n4656) );
  NOR2_X1 U6661 ( .A1(n9433), .A2(n6976), .ZN(n4657) );
  NAND2_X1 U6662 ( .A1(n9239), .A2(n9252), .ZN(n9433) );
  AND2_X1 U6663 ( .A1(n8045), .A2(n6975), .ZN(n9239) );
  NAND3_X1 U6664 ( .A1(n5575), .A2(n4662), .A3(n4661), .ZN(n4994) );
  NAND3_X1 U6665 ( .A1(n5038), .A2(n4663), .A3(n5567), .ZN(n4662) );
  NAND3_X1 U6666 ( .A1(n5038), .A2(n5567), .A3(n5546), .ZN(n4704) );
  NOR2_X1 U6667 ( .A1(n4703), .A2(n4664), .ZN(n4663) );
  NAND3_X1 U6668 ( .A1(n4667), .A2(SI_1_), .A3(n4996), .ZN(n5510) );
  NAND2_X1 U6669 ( .A1(n4667), .A2(n4996), .ZN(n5475) );
  NAND2_X1 U6670 ( .A1(n7493), .A2(n4484), .ZN(n4669) );
  NAND2_X1 U6671 ( .A1(n7494), .A2(n7495), .ZN(n7493) );
  MUX2_X1 U6672 ( .A(n8993), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  MUX2_X1 U6673 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8993), .S(n6185), .Z(n6653) );
  INV_X1 U6674 ( .A(n8507), .ZN(n4675) );
  AOI21_X2 U6675 ( .B1(n6833), .B2(n4678), .A(n4677), .ZN(n8600) );
  AOI21_X1 U6676 ( .B1(n5235), .B2(n5234), .A(n6847), .ZN(n4682) );
  OAI21_X1 U6677 ( .B1(n5444), .B2(n4690), .A(n4689), .ZN(n5446) );
  NAND2_X1 U6678 ( .A1(n5444), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n4689) );
  NAND2_X1 U6679 ( .A1(n4409), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4691) );
  NAND2_X1 U6680 ( .A1(n4692), .A2(n7253), .ZN(P2_U3296) );
  NAND4_X1 U6681 ( .A1(n7246), .A2(n4694), .A3(n4693), .A4(n4697), .ZN(n4692)
         );
  NAND2_X1 U6682 ( .A1(n4696), .A2(n7243), .ZN(n4695) );
  NAND2_X1 U6683 ( .A1(n7242), .A2(n4438), .ZN(n4697) );
  NAND2_X1 U6684 ( .A1(n5805), .A2(n5759), .ZN(n5762) );
  NAND2_X1 U6685 ( .A1(n5017), .A2(n4534), .ZN(n5859) );
  NAND2_X1 U6686 ( .A1(n4702), .A2(n5447), .ZN(n5576) );
  NAND2_X1 U6687 ( .A1(n4704), .A2(n5445), .ZN(n4702) );
  AND2_X1 U6688 ( .A1(n5679), .A2(n5651), .ZN(n4715) );
  NAND2_X1 U6689 ( .A1(n5434), .A2(n4720), .ZN(n5512) );
  NAND2_X1 U6690 ( .A1(n8693), .A2(n8694), .ZN(n6686) );
  NAND2_X2 U6691 ( .A1(n6684), .A2(n6683), .ZN(n8693) );
  OR2_X1 U6692 ( .A1(n7683), .A2(n4736), .ZN(n4735) );
  NAND3_X1 U6693 ( .A1(n4735), .A2(n4738), .A3(n4733), .ZN(n4732) );
  NAND2_X1 U6694 ( .A1(n7683), .A2(n9428), .ZN(n6974) );
  NAND2_X1 U6695 ( .A1(n4734), .A2(n4737), .ZN(n4733) );
  INV_X1 U6696 ( .A(n9428), .ZN(n4734) );
  INV_X1 U6697 ( .A(n4737), .ZN(n4736) );
  NAND2_X4 U6698 ( .A1(n6120), .A2(n7029), .ZN(n7287) );
  NAND2_X1 U6699 ( .A1(n5984), .A2(n4740), .ZN(n4900) );
  NAND3_X1 U6700 ( .A1(n4900), .A2(n8339), .A3(n4899), .ZN(n4898) );
  OAI21_X1 U6701 ( .B1(n9302), .B2(n9384), .A(n9424), .ZN(n4747) );
  MUX2_X1 U6702 ( .A(n5605), .B(n7335), .S(n5444), .Z(n5607) );
  INV_X1 U6703 ( .A(n10110), .ZN(n4753) );
  INV_X1 U6704 ( .A(n4756), .ZN(n10108) );
  NOR2_X1 U6705 ( .A1(n10108), .A2(n4876), .ZN(n10124) );
  NAND3_X1 U6706 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_IR_REG_1__SCAN_IN), .ZN(n4765) );
  NAND2_X1 U6707 ( .A1(n4880), .A2(n5869), .ZN(n4768) );
  AOI21_X1 U6708 ( .B1(n9558), .B2(n9556), .A(n4868), .ZN(n4769) );
  NAND3_X1 U6709 ( .A1(n4769), .A2(n4768), .A3(n4767), .ZN(P1_U3262) );
  INV_X1 U6710 ( .A(n5079), .ZN(n4771) );
  NAND2_X1 U6711 ( .A1(n4776), .A2(n4775), .ZN(n4778) );
  AND2_X1 U6712 ( .A1(n4778), .A2(n4777), .ZN(n10095) );
  INV_X1 U6713 ( .A(n4778), .ZN(n7367) );
  OR2_X2 U6714 ( .A1(n7859), .A2(n4781), .ZN(n4780) );
  AND2_X2 U6715 ( .A1(n4785), .A2(n4784), .ZN(n9532) );
  INV_X1 U6716 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4786) );
  NOR2_X2 U6717 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6188) );
  INV_X1 U6718 ( .A(n6647), .ZN(n6648) );
  NAND2_X1 U6719 ( .A1(n6647), .A2(n4427), .ZN(n4787) );
  NAND2_X1 U6720 ( .A1(n7221), .A2(n6764), .ZN(n4796) );
  OAI21_X1 U6721 ( .B1(n5341), .B2(n4800), .A(n4799), .ZN(n4798) );
  NAND2_X1 U6722 ( .A1(n4803), .A2(n4469), .ZN(n4799) );
  NAND2_X1 U6723 ( .A1(n5699), .A2(n9086), .ZN(n4800) );
  NOR2_X1 U6724 ( .A1(n5344), .A2(n4806), .ZN(n4802) );
  NAND3_X1 U6725 ( .A1(n6106), .A2(n5869), .A3(n9405), .ZN(n4809) );
  NAND2_X2 U6726 ( .A1(n4811), .A2(n4809), .ZN(n9036) );
  NAND2_X1 U6727 ( .A1(n4817), .A2(n9105), .ZN(n4816) );
  NAND2_X1 U6728 ( .A1(n8995), .A2(n9104), .ZN(n4818) );
  INV_X1 U6729 ( .A(n9103), .ZN(n4819) );
  NAND2_X1 U6730 ( .A1(n7669), .A2(n7717), .ZN(n5003) );
  INV_X1 U6731 ( .A(n7671), .ZN(n4820) );
  NAND2_X1 U6732 ( .A1(n6187), .A2(n4822), .ZN(n7418) );
  OR2_X1 U6733 ( .A1(n6178), .A2(n6633), .ZN(n4822) );
  NAND2_X1 U6734 ( .A1(n8298), .A2(n4827), .ZN(n4825) );
  NAND2_X1 U6735 ( .A1(n4833), .A2(n4831), .ZN(n8392) );
  NAND4_X1 U6736 ( .A1(n6338), .A2(n6337), .A3(n5009), .A4(n5300), .ZN(n4833)
         );
  NAND3_X1 U6737 ( .A1(n6338), .A2(n5009), .A3(n6337), .ZN(n4835) );
  NAND2_X1 U6738 ( .A1(n5310), .A2(n4839), .ZN(n4838) );
  NAND2_X1 U6739 ( .A1(n4992), .A2(n6151), .ZN(n6144) );
  NAND2_X1 U6740 ( .A1(n4992), .A2(n4841), .ZN(n6147) );
  XNOR2_X1 U6741 ( .A(n6194), .B(n7607), .ZN(n6178) );
  NAND2_X1 U6742 ( .A1(n7524), .A2(n4878), .ZN(n4844) );
  NAND2_X1 U6743 ( .A1(n7416), .A2(n6187), .ZN(n7447) );
  NAND2_X1 U6744 ( .A1(n8399), .A2(n6426), .ZN(n6428) );
  NAND2_X1 U6745 ( .A1(n5003), .A2(n7718), .ZN(n7721) );
  NAND2_X1 U6746 ( .A1(n8392), .A2(n8391), .ZN(n8390) );
  XNOR2_X1 U6747 ( .A(n6194), .B(n10224), .ZN(n6200) );
  NAND3_X1 U6748 ( .A1(n6192), .A2(n4533), .A3(n6193), .ZN(n7450) );
  XNOR2_X1 U6749 ( .A(n7316), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n7292) );
  NOR2_X1 U6750 ( .A1(n7375), .A2(n7374), .ZN(n7380) );
  NOR2_X2 U6751 ( .A1(n7561), .A2(n5061), .ZN(n7565) );
  NAND2_X1 U6752 ( .A1(n5056), .A2(n5054), .ZN(n9557) );
  OAI21_X1 U6753 ( .B1(n9559), .B2(n10137), .A(n4881), .ZN(n4880) );
  XNOR2_X1 U6754 ( .A(n9547), .B(n5080), .ZN(n9536) );
  NOR2_X1 U6755 ( .A1(n9534), .A2(n5065), .ZN(n9547) );
  NAND2_X1 U6756 ( .A1(n7565), .A2(n7564), .ZN(n7775) );
  NOR2_X1 U6757 ( .A1(n9525), .A2(n9524), .ZN(n9534) );
  NAND2_X1 U6758 ( .A1(n10143), .A2(n10142), .ZN(n4847) );
  NAND2_X1 U6759 ( .A1(n5113), .A2(n5375), .ZN(n5265) );
  NAND2_X1 U6760 ( .A1(n8693), .A2(n4848), .ZN(n5100) );
  NAND2_X1 U6761 ( .A1(n5044), .A2(n5042), .ZN(n9774) );
  NAND2_X1 U6762 ( .A1(n6984), .A2(n9446), .ZN(n7024) );
  NAND3_X1 U6763 ( .A1(n5106), .A2(n4529), .A3(n6658), .ZN(n5105) );
  OAI22_X2 U6764 ( .A1(n7821), .A2(n6660), .B1(n10243), .B2(n7793), .ZN(n7920)
         );
  AND2_X2 U6765 ( .A1(n9366), .A2(n9799), .ZN(n9810) );
  NAND2_X1 U6766 ( .A1(n6157), .A2(n6566), .ZN(n6565) );
  NAND2_X1 U6767 ( .A1(n6633), .A2(n7607), .ZN(n7123) );
  AND3_X2 U6768 ( .A1(n5226), .A2(n5225), .A3(n5224), .ZN(n7607) );
  NAND2_X1 U6769 ( .A1(n7949), .A2(n7950), .ZN(n6665) );
  NAND2_X1 U6770 ( .A1(n10209), .A2(n7127), .ZN(n6657) );
  INV_X1 U6771 ( .A(n8731), .ZN(n4852) );
  OAI21_X1 U6772 ( .B1(n6154), .B2(n5312), .A(n4853), .ZN(n5091) );
  INV_X1 U6773 ( .A(n6633), .ZN(n5112) );
  NAND2_X1 U6774 ( .A1(n5105), .A2(n6659), .ZN(n7821) );
  NOR2_X1 U6775 ( .A1(n8603), .A2(n8602), .ZN(n5159) );
  NAND2_X1 U6776 ( .A1(n5150), .A2(n5149), .ZN(n5148) );
  INV_X1 U6777 ( .A(n5260), .ZN(n5259) );
  MUX2_X1 U6778 ( .A(n9261), .B(n9260), .S(n9330), .Z(n9269) );
  NAND2_X1 U6779 ( .A1(n5272), .A2(n5271), .ZN(n4998) );
  NAND2_X1 U6780 ( .A1(n4858), .A2(n4857), .ZN(n4856) );
  NAND2_X1 U6781 ( .A1(n7207), .A2(n7206), .ZN(n4858) );
  NAND2_X1 U6782 ( .A1(n5095), .A2(n5094), .ZN(n5093) );
  INV_X1 U6783 ( .A(n7085), .ZN(n7246) );
  AOI21_X1 U6784 ( .B1(n6635), .B2(n5370), .A(n5369), .ZN(n7943) );
  OAI21_X1 U6785 ( .B1(n7678), .B2(n7731), .A(n6923), .ZN(n6926) );
  OR2_X2 U6786 ( .A1(n7017), .A2(n7016), .ZN(n8275) );
  INV_X1 U6787 ( .A(n6587), .ZN(n4878) );
  NAND2_X1 U6788 ( .A1(n4992), .A2(n4896), .ZN(n6165) );
  NAND2_X1 U6789 ( .A1(n9615), .A2(n9347), .ZN(n9605) );
  NAND2_X1 U6790 ( .A1(n8149), .A2(n5045), .ZN(n5044) );
  AOI21_X1 U6791 ( .B1(n9606), .B2(n5379), .A(n9817), .ZN(n9607) );
  NAND2_X1 U6792 ( .A1(n9557), .A2(n10127), .ZN(n4881) );
  NAND2_X2 U6793 ( .A1(n5479), .A2(n5478), .ZN(n9072) );
  AOI21_X1 U6794 ( .B1(n5118), .B2(n4523), .A(n5116), .ZN(n9260) );
  MUX2_X1 U6795 ( .A(n7186), .B(n7185), .S(n4420), .Z(n7191) );
  NAND2_X1 U6796 ( .A1(n7163), .A2(n7165), .ZN(n5097) );
  AOI21_X1 U6797 ( .B1(n7136), .B2(n4988), .A(n7135), .ZN(n7143) );
  OR2_X2 U6798 ( .A1(n10139), .A2(n10140), .ZN(n10136) );
  INV_X1 U6799 ( .A(n5506), .ZN(n4897) );
  NOR2_X1 U6800 ( .A1(n7554), .A2(n5074), .ZN(n7555) );
  NAND2_X1 U6801 ( .A1(n9507), .A2(n9508), .ZN(n9506) );
  NOR2_X2 U6802 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5506) );
  INV_X1 U6803 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6204) );
  NAND2_X1 U6804 ( .A1(n4882), .A2(n5081), .ZN(n7162) );
  NAND2_X1 U6805 ( .A1(n7167), .A2(n7166), .ZN(n5095) );
  NAND2_X1 U6806 ( .A1(n5249), .A2(n5248), .ZN(n7495) );
  AOI22_X2 U6807 ( .A1(n8572), .A2(n8573), .B1(P2_REG1_REG_16__SCAN_IN), .B2(
        n8578), .ZN(n6833) );
  NOR2_X1 U6808 ( .A1(n5128), .A2(n5131), .ZN(n5127) );
  NAND3_X1 U6809 ( .A1(n4886), .A2(n5122), .A3(n5123), .ZN(n9466) );
  NAND2_X1 U6810 ( .A1(n4892), .A2(n4890), .ZN(P2_U3180) );
  NAND2_X1 U6811 ( .A1(n8466), .A2(n8470), .ZN(n4892) );
  INV_X1 U6812 ( .A(n10186), .ZN(n4894) );
  NAND2_X1 U6813 ( .A1(n7132), .A2(n7133), .ZN(n7127) );
  NAND2_X1 U6814 ( .A1(n6665), .A2(n5110), .ZN(n5109) );
  NAND2_X1 U6815 ( .A1(n5265), .A2(n5263), .ZN(n6680) );
  NAND2_X1 U6816 ( .A1(n5097), .A2(n7217), .ZN(n5096) );
  AOI21_X1 U6817 ( .B1(n7225), .B2(n7224), .A(n7237), .ZN(n7230) );
  NAND2_X1 U6818 ( .A1(n4905), .A2(n4898), .ZN(n9044) );
  INV_X1 U6819 ( .A(n5571), .ZN(n4913) );
  NAND2_X1 U6820 ( .A1(n9156), .A2(n4918), .ZN(n4914) );
  OAI21_X1 U6821 ( .B1(n9149), .B2(n4924), .A(n4921), .ZN(n5983) );
  INV_X1 U6822 ( .A(n9079), .ZN(n4926) );
  OAI21_X1 U6823 ( .B1(n6982), .B2(n4932), .A(n4929), .ZN(n4933) );
  NAND2_X1 U6824 ( .A1(n6982), .A2(n9342), .ZN(n6984) );
  NAND2_X1 U6825 ( .A1(n5382), .A2(n5374), .ZN(n4937) );
  NAND2_X2 U6826 ( .A1(n8015), .A2(n4939), .ZN(n8149) );
  INV_X1 U6827 ( .A(n6974), .ZN(n4942) );
  INV_X1 U6828 ( .A(n5451), .ZN(n5337) );
  AND4_X2 U6829 ( .A1(n5391), .A2(n5389), .A3(n5388), .A4(n5390), .ZN(n5338)
         );
  NAND2_X1 U6830 ( .A1(n6267), .A2(n4951), .ZN(n6306) );
  NAND4_X1 U6831 ( .A1(n4953), .A2(n6217), .A3(n6216), .A4(n6239), .ZN(n6268)
         );
  NAND4_X1 U6832 ( .A1(n7220), .A2(n4956), .A3(n4514), .A4(n8641), .ZN(n4955)
         );
  NAND2_X1 U6833 ( .A1(n6344), .A2(n4544), .ZN(n6383) );
  NAND2_X1 U6834 ( .A1(n6445), .A2(n4960), .ZN(n6477) );
  NAND2_X1 U6835 ( .A1(n6504), .A2(n4963), .ZN(n6558) );
  NAND2_X1 U6836 ( .A1(n6504), .A2(n6503), .ZN(n6517) );
  OAI22_X1 U6837 ( .A1(n9220), .A2(n7320), .B1(n7287), .B2(n10099), .ZN(n4978)
         );
  NAND2_X4 U6838 ( .A1(n7287), .A2(n5444), .ZN(n9220) );
  XNOR2_X1 U6839 ( .A(n5566), .B(n5565), .ZN(n7308) );
  INV_X2 U6840 ( .A(n5531), .ZN(n6953) );
  OAI21_X1 U6841 ( .B1(n9666), .B2(n4980), .A(n4982), .ZN(n9587) );
  NAND2_X1 U6842 ( .A1(n4981), .A2(n4429), .ZN(n4980) );
  NAND2_X1 U6843 ( .A1(n5444), .A2(n4997), .ZN(n4996) );
  MUX2_X1 U6844 ( .A(n10329), .B(n7307), .S(n5444), .Z(n5442) );
  NAND2_X1 U6845 ( .A1(n4999), .A2(n7218), .ZN(n6765) );
  OAI21_X2 U6846 ( .B1(n6154), .B2(n5315), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6170) );
  AND2_X1 U6847 ( .A1(n6207), .A2(n4468), .ZN(n5004) );
  AND2_X1 U6848 ( .A1(n6227), .A2(n4503), .ZN(n5005) );
  NAND2_X1 U6849 ( .A1(n10286), .A2(n4407), .ZN(n6788) );
  OAI21_X1 U6850 ( .B1(n9414), .B2(n5015), .A(n4483), .ZN(n5014) );
  AND2_X1 U6851 ( .A1(n9383), .A2(n9415), .ZN(n5015) );
  OR2_X1 U6852 ( .A1(n5787), .A2(SI_15_), .ZN(n5022) );
  NAND3_X1 U6853 ( .A1(n5271), .A2(n5653), .A3(n5754), .ZN(n5026) );
  AND2_X1 U6854 ( .A1(n5756), .A2(n5757), .ZN(n5027) );
  NAND2_X1 U6855 ( .A1(n5038), .A2(n5546), .ZN(n5566) );
  NAND3_X1 U6856 ( .A1(n5040), .A2(n9385), .A3(n5039), .ZN(n9664) );
  NAND3_X1 U6857 ( .A1(n9810), .A2(n5046), .A3(n5048), .ZN(n5043) );
  NAND2_X1 U6858 ( .A1(n9729), .A2(n9284), .ZN(n9709) );
  NAND2_X1 U6859 ( .A1(n9554), .A2(n5055), .ZN(n5054) );
  NOR2_X2 U6860 ( .A1(n8193), .A2(n5059), .ZN(n9504) );
  AOI21_X1 U6861 ( .B1(n5084), .B2(n5082), .A(n4454), .ZN(n5081) );
  NAND2_X1 U6862 ( .A1(n5307), .A2(n6176), .ZN(n6374) );
  NAND3_X1 U6863 ( .A1(n5096), .A2(n5093), .A3(n8833), .ZN(n5092) );
  NAND3_X1 U6864 ( .A1(n5100), .A2(n5098), .A3(n6691), .ZN(n8657) );
  NAND2_X1 U6865 ( .A1(n5099), .A2(n8675), .ZN(n5098) );
  NAND2_X1 U6866 ( .A1(n5101), .A2(n5104), .ZN(n8668) );
  NAND2_X1 U6867 ( .A1(n8693), .A2(n5102), .ZN(n5101) );
  NAND2_X1 U6868 ( .A1(n6657), .A2(n6656), .ZN(n7662) );
  NAND2_X1 U6869 ( .A1(n5109), .A2(n5107), .ZN(n8232) );
  NAND2_X1 U6870 ( .A1(n6665), .A2(n6664), .ZN(n8009) );
  NOR2_X1 U6871 ( .A1(n6669), .A2(n5111), .ZN(n5110) );
  INV_X1 U6872 ( .A(n6664), .ZN(n5111) );
  NAND2_X1 U6873 ( .A1(n9253), .A2(n9252), .ZN(n5118) );
  NAND3_X1 U6874 ( .A1(n4481), .A2(n5120), .A3(n5132), .ZN(n5125) );
  NAND3_X1 U6875 ( .A1(n5120), .A2(n5119), .A3(n4481), .ZN(n5124) );
  AND2_X1 U6876 ( .A1(n5132), .A2(n4517), .ZN(n5119) );
  NAND3_X1 U6877 ( .A1(n5127), .A2(n5124), .A3(n5125), .ZN(n5121) );
  NAND3_X1 U6878 ( .A1(n9306), .A2(n5127), .A3(n5134), .ZN(n5122) );
  NAND3_X1 U6879 ( .A1(n9314), .A2(n5124), .A3(n5127), .ZN(n5123) );
  NAND2_X1 U6880 ( .A1(n5399), .A2(n5339), .ZN(n5448) );
  NAND3_X1 U6881 ( .A1(n5399), .A2(n5339), .A3(n10340), .ZN(n5402) );
  AOI21_X1 U6882 ( .B1(n9299), .B2(n9298), .A(n9297), .ZN(n9302) );
  OR2_X1 U6883 ( .A1(n5553), .A2(n5470), .ZN(n5474) );
  NAND2_X1 U6884 ( .A1(n4417), .A2(n5221), .ZN(n5226) );
  NAND2_X1 U6885 ( .A1(n5501), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5473) );
  NAND2_X1 U6886 ( .A1(n7234), .A2(n7222), .ZN(n7225) );
  NAND3_X1 U6887 ( .A1(n5144), .A2(n6809), .A3(n5142), .ZN(n6810) );
  INV_X1 U6888 ( .A(n6807), .ZN(n5146) );
  NOR2_X1 U6889 ( .A1(n5148), .A2(n7306), .ZN(n5147) );
  NAND2_X1 U6890 ( .A1(n7508), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5149) );
  INV_X1 U6891 ( .A(n7496), .ZN(n5150) );
  NAND2_X1 U6892 ( .A1(n5153), .A2(n5151), .ZN(n6813) );
  INV_X1 U6893 ( .A(n6813), .ZN(n6814) );
  INV_X1 U6894 ( .A(n6886), .ZN(n5154) );
  NAND3_X1 U6895 ( .A1(n5160), .A2(P2_REG2_REG_17__SCAN_IN), .A3(n8603), .ZN(
        n8588) );
  NAND2_X1 U6896 ( .A1(n6817), .A2(n4444), .ZN(n5157) );
  NAND2_X1 U6897 ( .A1(n6795), .A2(n4524), .ZN(n5162) );
  OAI21_X1 U6898 ( .B1(n6795), .B2(n4536), .A(n5162), .ZN(n7543) );
  XNOR2_X1 U6899 ( .A(n6795), .B(n6847), .ZN(n7457) );
  INV_X1 U6900 ( .A(n6797), .ZN(n7542) );
  INV_X1 U6901 ( .A(n6815), .ZN(n5165) );
  NAND2_X1 U6902 ( .A1(n5165), .A2(n8579), .ZN(n5168) );
  NAND3_X1 U6903 ( .A1(n5170), .A2(n6803), .A3(n5169), .ZN(n6804) );
  NAND3_X1 U6904 ( .A1(n5172), .A2(n6799), .A3(n5171), .ZN(n5169) );
  NAND3_X1 U6905 ( .A1(n4432), .A2(n7038), .A3(n9598), .ZN(n9566) );
  AND2_X2 U6906 ( .A1(n7896), .A2(n5176), .ZN(n8023) );
  AOI21_X1 U6907 ( .B1(n9973), .B2(n10164), .A(n5179), .ZN(n9857) );
  NAND3_X1 U6908 ( .A1(n5182), .A2(n4531), .A3(n9784), .ZN(n9854) );
  NAND2_X1 U6909 ( .A1(n5183), .A2(n8154), .ZN(n9751) );
  NAND2_X1 U6910 ( .A1(n4463), .A2(n5188), .ZN(n7805) );
  NOR2_X1 U6911 ( .A1(n5189), .A2(n7587), .ZN(n5188) );
  NAND3_X1 U6912 ( .A1(n5197), .A2(n5198), .A3(n7145), .ZN(n7819) );
  NAND2_X2 U6913 ( .A1(n4407), .A2(n4409), .ZN(n7071) );
  NAND2_X1 U6914 ( .A1(n6185), .A2(n5223), .ZN(n5225) );
  NAND2_X1 U6915 ( .A1(n5236), .A2(n5244), .ZN(n5243) );
  NAND2_X1 U6916 ( .A1(n5239), .A2(n5237), .ZN(n5236) );
  NAND2_X1 U6917 ( .A1(n8530), .A2(n5245), .ZN(n5239) );
  NAND2_X1 U6918 ( .A1(n5243), .A2(n5242), .ZN(n5241) );
  NAND2_X1 U6919 ( .A1(n5154), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5244) );
  OR2_X1 U6920 ( .A1(n8657), .A2(n4515), .ZN(n5266) );
  NAND2_X1 U6921 ( .A1(n8657), .A2(n5269), .ZN(n5268) );
  NAND2_X1 U6922 ( .A1(n5444), .A2(n5274), .ZN(n5273) );
  OAI21_X1 U6923 ( .B1(n9820), .B2(n5289), .A(n6936), .ZN(n5288) );
  NAND2_X1 U6924 ( .A1(n6941), .A2(n6940), .ZN(n9728) );
  MUX2_X1 U6925 ( .A(n9219), .B(n10346), .S(n5444), .Z(n7049) );
  MUX2_X1 U6926 ( .A(n9215), .B(n7070), .S(n5444), .Z(n7067) );
  XNOR2_X1 U6927 ( .A(n5297), .B(n5568), .ZN(n7311) );
  OAI21_X1 U6928 ( .B1(n5565), .B2(n5298), .A(n5567), .ZN(n5297) );
  INV_X1 U6929 ( .A(n5566), .ZN(n5298) );
  NAND2_X1 U6930 ( .A1(n8167), .A2(n6365), .ZN(n8244) );
  INV_X1 U6931 ( .A(n5301), .ZN(n8243) );
  INV_X1 U6932 ( .A(n8245), .ZN(n5302) );
  NAND2_X1 U6933 ( .A1(n5303), .A2(n8317), .ZN(n5304) );
  NAND3_X1 U6934 ( .A1(n5307), .A2(n6176), .A3(P2_REG2_REG_1__SCAN_IN), .ZN(
        n5305) );
  NAND2_X1 U6935 ( .A1(n6428), .A2(n5361), .ZN(n8452) );
  INV_X1 U6936 ( .A(n5310), .ZN(n8451) );
  INV_X1 U6937 ( .A(n5361), .ZN(n5311) );
  INV_X1 U6938 ( .A(n7783), .ZN(n5321) );
  NAND2_X1 U6939 ( .A1(n5338), .A2(n5337), .ZN(n5456) );
  INV_X1 U6940 ( .A(n5649), .ZN(n5354) );
  NAND2_X1 U6941 ( .A1(n4405), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5357) );
  INV_X1 U6942 ( .A(n9866), .ZN(n9600) );
  NAND2_X1 U6943 ( .A1(n10205), .A2(n10210), .ZN(n10204) );
  NOR2_X1 U6944 ( .A1(n4521), .A2(n5387), .ZN(n5562) );
  NAND2_X1 U6945 ( .A1(n9072), .A2(n5490), .ZN(n5480) );
  NOR2_X1 U6946 ( .A1(n9490), .A2(n9072), .ZN(n7584) );
  NAND2_X1 U6947 ( .A1(n9307), .A2(n9347), .ZN(n9314) );
  NAND2_X1 U6948 ( .A1(n6972), .A2(n6971), .ZN(n7683) );
  AOI21_X1 U6949 ( .B1(n6132), .B2(n6131), .A(n6130), .ZN(n6133) );
  NAND2_X1 U6950 ( .A1(n8021), .A2(n8020), .ZN(n8019) );
  NAND2_X1 U6951 ( .A1(n9490), .A2(n5822), .ZN(n5481) );
  NAND2_X1 U6952 ( .A1(n5448), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5449) );
  AND2_X1 U6953 ( .A1(n8340), .A2(n9204), .ZN(n6131) );
  INV_X1 U6954 ( .A(n4405), .ZN(n6985) );
  XNOR2_X1 U6955 ( .A(n5497), .B(n5498), .ZN(n9068) );
  NAND2_X1 U6956 ( .A1(n5497), .A2(n5499), .ZN(n5500) );
  NOR2_X1 U6957 ( .A1(n6740), .A2(n6739), .ZN(n5358) );
  INV_X1 U6958 ( .A(n10228), .ZN(n8137) );
  INV_X1 U6959 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5995) );
  AND2_X1 U6960 ( .A1(n5551), .A2(n5550), .ZN(n5359) );
  AND2_X1 U6961 ( .A1(n6784), .A2(n6783), .ZN(n5360) );
  OR2_X1 U6962 ( .A1(n8082), .A2(n7105), .ZN(n5362) );
  AND2_X1 U6963 ( .A1(n6780), .A2(n6779), .ZN(n5363) );
  INV_X1 U6964 ( .A(n6725), .ZN(n6726) );
  OR2_X1 U6965 ( .A1(n6867), .A2(n6806), .ZN(n5364) );
  AND2_X1 U6966 ( .A1(n6151), .A2(n6150), .ZN(n5365) );
  NAND2_X1 U6967 ( .A1(n10259), .A2(n8892), .ZN(n8884) );
  OR2_X1 U6968 ( .A1(n9335), .A2(n9456), .ZN(n5366) );
  INV_X2 U6969 ( .A(n10160), .ZN(n10161) );
  XNOR2_X1 U6970 ( .A(n5482), .B(n8327), .ZN(n5497) );
  INV_X1 U6971 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6452) );
  OR2_X1 U6972 ( .A1(n7227), .A2(n8623), .ZN(n5367) );
  AND2_X1 U6973 ( .A1(n5651), .A2(n5615), .ZN(n5368) );
  INV_X1 U6974 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6578) );
  INV_X1 U6975 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8163) );
  NOR2_X1 U6976 ( .A1(n7950), .A2(n7945), .ZN(n5369) );
  NOR2_X1 U6977 ( .A1(n7944), .A2(n7950), .ZN(n5370) );
  AND2_X1 U6978 ( .A1(n7804), .A2(n8043), .ZN(n5371) );
  OR2_X1 U6979 ( .A1(n7287), .A2(n7321), .ZN(n5372) );
  INV_X1 U6980 ( .A(n7333), .ZN(n6802) );
  AND2_X1 U6981 ( .A1(n6981), .A2(n9343), .ZN(n5373) );
  AND2_X1 U6982 ( .A1(n9344), .A2(n9343), .ZN(n5374) );
  INV_X1 U6983 ( .A(n8623), .ZN(n7239) );
  INV_X1 U6984 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5400) );
  AND2_X1 U6985 ( .A1(n7178), .A2(n6676), .ZN(n5375) );
  INV_X1 U6986 ( .A(n6855), .ZN(n6798) );
  AND2_X1 U6987 ( .A1(n9177), .A2(n5700), .ZN(n5376) );
  INV_X1 U6988 ( .A(n6777), .ZN(n8629) );
  AND2_X1 U6989 ( .A1(n9347), .A2(n9323), .ZN(n5377) );
  OR2_X1 U6990 ( .A1(n6922), .A2(n7848), .ZN(n5378) );
  NAND2_X1 U6991 ( .A1(n9605), .A2(n9604), .ZN(n5379) );
  AND2_X1 U6992 ( .A1(n6994), .A2(n6993), .ZN(n5380) );
  OR2_X1 U6993 ( .A1(n8949), .A2(n8948), .ZN(P2_U3438) );
  OR2_X1 U6994 ( .A1(n8880), .A2(n8879), .ZN(P2_U3475) );
  OR2_X1 U6995 ( .A1(n8782), .A2(n8781), .ZN(P2_U3217) );
  AND2_X1 U6996 ( .A1(n5826), .A2(n5825), .ZN(n5386) );
  AND2_X1 U6997 ( .A1(n4405), .A2(n7889), .ZN(n5387) );
  INV_X1 U6998 ( .A(n10257), .ZN(n10259) );
  INV_X1 U6999 ( .A(n10254), .ZN(n10257) );
  AND2_X1 U7000 ( .A1(n7332), .A2(n6565), .ZN(n7351) );
  INV_X2 U7001 ( .A(n10249), .ZN(n10247) );
  AND2_X1 U7002 ( .A1(n6720), .A2(n6719), .ZN(n10249) );
  INV_X1 U7003 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6134) );
  NAND2_X1 U7004 ( .A1(n7233), .A2(n7223), .ZN(n7224) );
  INV_X1 U7005 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6138) );
  OR2_X1 U7006 ( .A1(n8297), .A2(n8695), .ZN(n6501) );
  AND2_X1 U7007 ( .A1(n7087), .A2(n7086), .ZN(n7236) );
  INV_X1 U7008 ( .A(n10184), .ZN(n6793) );
  INV_X1 U7009 ( .A(n7237), .ZN(n6761) );
  OR2_X1 U7010 ( .A1(n5701), .A2(n9177), .ZN(n5703) );
  INV_X1 U7011 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5916) );
  OR2_X1 U7012 ( .A1(n6738), .A2(n6737), .ZN(n6739) );
  OR2_X1 U7013 ( .A1(n6485), .A2(n8708), .ZN(n6486) );
  OR2_X1 U7014 ( .A1(n8212), .A2(n8142), .ZN(n6324) );
  NAND2_X1 U7015 ( .A1(n7240), .A2(n8623), .ZN(n7241) );
  NAND2_X1 U7016 ( .A1(n6804), .A2(n7996), .ZN(n6805) );
  INV_X1 U7017 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6406) );
  OR2_X1 U7018 ( .A1(n7915), .A2(n7147), .ZN(n7944) );
  OR2_X1 U7019 ( .A1(n6650), .A2(n8669), .ZN(n6689) );
  NAND2_X1 U7020 ( .A1(n5481), .A2(n5480), .ZN(n5482) );
  INV_X1 U7021 ( .A(n5982), .ZN(n5981) );
  NAND2_X1 U7022 ( .A1(n8101), .A2(n7968), .ZN(n8042) );
  INV_X1 U7023 ( .A(SI_25_), .ZN(n6039) );
  INV_X1 U7024 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5458) );
  AND2_X1 U7025 ( .A1(n6336), .A2(n6324), .ZN(n6325) );
  INV_X1 U7026 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6284) );
  INV_X1 U7027 ( .A(n6604), .ZN(n6769) );
  INV_X1 U7028 ( .A(n10294), .ZN(n10170) );
  INV_X1 U7029 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10488) );
  INV_X1 U7030 ( .A(n8957), .ZN(n6778) );
  NAND2_X1 U7031 ( .A1(n7336), .A2(n6653), .ZN(n7601) );
  INV_X1 U7032 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6393) );
  OAI22_X1 U7033 ( .A1(n6918), .A2(n6056), .B1(n7581), .B2(n6057), .ZN(n5498)
         );
  INV_X1 U7034 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5737) );
  OR2_X1 U7035 ( .A1(n6119), .A2(n9404), .ZN(n6126) );
  NAND2_X1 U7036 ( .A1(n6045), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6071) );
  NAND2_X1 U7037 ( .A1(n5969), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5997) );
  NAND2_X1 U7038 ( .A1(n5774), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5796) );
  OR2_X1 U7039 ( .A1(n9914), .A2(n9744), .ZN(n6942) );
  AND2_X1 U7040 ( .A1(n9405), .A2(n9464), .ZN(n9421) );
  OR2_X1 U7041 ( .A1(n9335), .A2(n6995), .ZN(n9404) );
  INV_X1 U7042 ( .A(n8797), .ZN(n8771) );
  AOI21_X1 U7043 ( .B1(n6336), .B2(n6335), .A(n6334), .ZN(n6337) );
  INV_X1 U7044 ( .A(n8425), .ZN(n6484) );
  INV_X1 U7045 ( .A(n8578), .ZN(n6895) );
  AND2_X1 U7046 ( .A1(n4527), .A2(n7218), .ZN(n8661) );
  INV_X1 U7047 ( .A(n8741), .ZN(n6643) );
  INV_X1 U7048 ( .A(n6706), .ZN(n6596) );
  OAI21_X1 U7049 ( .B1(n6576), .B2(n6575), .A(n6574), .ZN(n6700) );
  NAND2_X1 U7050 ( .A1(n10249), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6779) );
  AND2_X1 U7051 ( .A1(n7212), .A2(n7088), .ZN(n8689) );
  NOR2_X1 U7052 ( .A1(n6620), .A2(n7315), .ZN(n6718) );
  INV_X1 U7053 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6146) );
  AND2_X1 U7054 ( .A1(n6398), .A2(n6397), .ZN(n6402) );
  INV_X1 U7055 ( .A(n9197), .ZN(n9206) );
  INV_X1 U7056 ( .A(n9610), .ZN(n9611) );
  NAND2_X1 U7057 ( .A1(n6019), .A2(n6018), .ZN(n6980) );
  INV_X1 U7058 ( .A(n9477), .ZN(n9900) );
  NAND2_X1 U7059 ( .A1(n10160), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7037) );
  NAND2_X1 U7060 ( .A1(n8153), .A2(n9439), .ZN(n8152) );
  INV_X1 U7061 ( .A(n9455), .ZN(n9400) );
  INV_X1 U7062 ( .A(n7912), .ZN(n7909) );
  INV_X1 U7063 ( .A(n9782), .ZN(n9817) );
  NAND2_X1 U7064 ( .A1(n9465), .A2(n8088), .ZN(n7620) );
  AND2_X1 U7065 ( .A1(n6731), .A2(n6017), .ZN(n6037) );
  NAND2_X1 U7066 ( .A1(n6583), .A2(n6582), .ZN(n6912) );
  NAND2_X1 U7067 ( .A1(n6624), .A2(n6623), .ZN(n8478) );
  AND2_X1 U7068 ( .A1(P2_U3893), .A2(n7247), .ZN(n10288) );
  INV_X1 U7069 ( .A(n10207), .ZN(n8821) );
  INV_X1 U7070 ( .A(n8884), .ZN(n8888) );
  NAND2_X1 U7071 ( .A1(n6710), .A2(n6709), .ZN(n6711) );
  INV_X1 U7072 ( .A(n10242), .ZN(n8892) );
  INV_X1 U7073 ( .A(n7091), .ZN(n8008) );
  AND2_X1 U7074 ( .A1(n8085), .A2(n7595), .ZN(n10228) );
  NAND2_X1 U7075 ( .A1(n8177), .A2(n8137), .ZN(n10245) );
  INV_X1 U7076 ( .A(n9207), .ZN(n9192) );
  NAND2_X1 U7077 ( .A1(n6125), .A2(n9456), .ZN(n9197) );
  INV_X1 U7078 ( .A(n10141), .ZN(n10127) );
  INV_X1 U7079 ( .A(n10137), .ZN(n10131) );
  NOR2_X2 U7080 ( .A1(n7300), .A2(n6995), .ZN(n9804) );
  AND2_X1 U7081 ( .A1(n9842), .A2(n7706), .ZN(n9847) );
  AND2_X1 U7082 ( .A1(n9842), .A2(n7618), .ZN(n9837) );
  INV_X1 U7083 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10572) );
  INV_X1 U7084 ( .A(n7848), .ZN(n9349) );
  NOR2_X1 U7085 ( .A1(n10161), .A2(n7012), .ZN(n7013) );
  AND2_X1 U7086 ( .A1(n5808), .A2(n5807), .ZN(n9535) );
  XNOR2_X1 U7087 ( .A(n5442), .B(SI_3_), .ZN(n5530) );
  INV_X1 U7088 ( .A(n6628), .ZN(n6629) );
  INV_X1 U7089 ( .A(n6650), .ZN(n8917) );
  INV_X1 U7090 ( .A(n8470), .ZN(n8460) );
  AND2_X1 U7091 ( .A1(n7062), .A2(n6760), .ZN(n8638) );
  INV_X1 U7092 ( .A(n8708), .ZN(n8487) );
  OR2_X1 U7093 ( .A1(P2_U3150), .A2(n6914), .ZN(n10294) );
  NAND2_X1 U7094 ( .A1(n10286), .A2(n6834), .ZN(n10197) );
  INV_X1 U7095 ( .A(n8804), .ZN(n8835) );
  NAND2_X1 U7096 ( .A1(n10259), .A2(n10245), .ZN(n8891) );
  NAND2_X1 U7097 ( .A1(n10247), .A2(n8892), .ZN(n8957) );
  INV_X1 U7098 ( .A(n7351), .ZN(n7340) );
  INV_X1 U7099 ( .A(n7332), .ZN(n7315) );
  INV_X1 U7100 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8985) );
  INV_X1 U7101 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7858) );
  INV_X1 U7102 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7395) );
  AND2_X1 U7103 ( .A1(n7299), .A2(n7298), .ZN(n10089) );
  INV_X1 U7104 ( .A(n9204), .ZN(n9199) );
  INV_X1 U7105 ( .A(n7020), .ZN(n9475) );
  INV_X1 U7106 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10567) );
  INV_X1 U7107 ( .A(n9856), .ZN(n9962) );
  INV_X1 U7108 ( .A(n9789), .ZN(n10006) );
  NAND2_X1 U7109 ( .A1(n10161), .A2(n10154), .ZN(n10016) );
  OR2_X1 U7110 ( .A1(n7010), .A2(n7009), .ZN(n10160) );
  INV_X1 U7111 ( .A(n10150), .ZN(n10149) );
  NAND2_X1 U7112 ( .A1(n7611), .A2(n9402), .ZN(n10150) );
  INV_X1 U7113 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9219) );
  INV_X1 U7114 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10030) );
  INV_X1 U7115 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8084) );
  INV_X1 U7116 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7444) );
  NAND2_X1 U7117 ( .A1(n4409), .A2(P1_U3086), .ZN(n10040) );
  NOR2_X1 U7118 ( .A1(n10059), .A2(n10058), .ZN(n10283) );
  NOR2_X1 U7119 ( .A1(n10063), .A2(n10062), .ZN(n10279) );
  AND2_X1 U7120 ( .A1(n7353), .A2(n6786), .ZN(P2_U3893) );
  NOR2_X1 U7121 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5391) );
  NAND2_X1 U7122 ( .A1(n5506), .A2(n5392), .ZN(n5451) );
  NOR2_X1 U7123 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5396) );
  NOR2_X1 U7124 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5398) );
  NOR2_X1 U7125 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5397) );
  XNOR2_X2 U7126 ( .A(n5401), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5413) );
  NAND2_X1 U7127 ( .A1(n5402), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5403) );
  INV_X1 U7128 ( .A(n5404), .ZN(n10022) );
  INV_X1 U7129 ( .A(n5555), .ZN(n5406) );
  NAND2_X1 U7130 ( .A1(n5406), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5557) );
  INV_X1 U7131 ( .A(n5586), .ZN(n5588) );
  NAND2_X1 U7132 ( .A1(n5557), .A2(n5407), .ZN(n5408) );
  AND2_X1 U7133 ( .A1(n5588), .A2(n5408), .ZN(n7878) );
  NAND2_X1 U7134 ( .A1(n4405), .A2(n7878), .ZN(n5418) );
  NOR2_X2 U7135 ( .A1(n5413), .A2(n5409), .ZN(n5501) );
  NAND2_X1 U7136 ( .A1(n5501), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5417) );
  INV_X1 U7137 ( .A(n5413), .ZN(n5410) );
  INV_X1 U7138 ( .A(n5412), .ZN(n5409) );
  INV_X1 U7139 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5411) );
  OR2_X1 U7140 ( .A1(n4406), .A2(n5411), .ZN(n5416) );
  INV_X1 U7141 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5414) );
  OR2_X1 U7142 ( .A1(n4408), .A2(n5414), .ZN(n5415) );
  NAND2_X1 U7143 ( .A1(n5429), .A2(n5420), .ZN(n5462) );
  INV_X1 U7144 ( .A(n5462), .ZN(n5421) );
  NAND2_X1 U7145 ( .A1(n5421), .A2(n4485), .ZN(n5425) );
  NAND2_X1 U7146 ( .A1(n5425), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5422) );
  NAND2_X1 U7147 ( .A1(n6087), .A2(n6091), .ZN(n5428) );
  INV_X1 U7148 ( .A(n5429), .ZN(n5430) );
  NAND2_X1 U7149 ( .A1(n5430), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U7150 ( .A1(n5419), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5432) );
  NAND2_X1 U7151 ( .A1(n9464), .A2(n9455), .ZN(n7704) );
  INV_X1 U7152 ( .A(n7704), .ZN(n5433) );
  AND2_X2 U7153 ( .A1(n6106), .A2(n5433), .ZN(n5468) );
  INV_X1 U7154 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7323) );
  INV_X1 U7155 ( .A(SI_2_), .ZN(n10363) );
  INV_X1 U7156 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10306) );
  INV_X1 U7157 ( .A(n5512), .ZN(n5435) );
  NAND2_X1 U7158 ( .A1(n5436), .A2(n5435), .ZN(n5441) );
  NAND2_X1 U7159 ( .A1(n5512), .A2(n10363), .ZN(n5439) );
  INV_X1 U7160 ( .A(n5476), .ZN(n5508) );
  INV_X1 U7161 ( .A(SI_1_), .ZN(n5437) );
  NAND2_X1 U7162 ( .A1(n5475), .A2(n5437), .ZN(n5438) );
  NAND2_X1 U7163 ( .A1(SI_1_), .A2(SI_2_), .ZN(n5440) );
  INV_X1 U7164 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7307) );
  INV_X1 U7165 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10329) );
  INV_X1 U7166 ( .A(n5442), .ZN(n5443) );
  NAND2_X1 U7167 ( .A1(n5443), .A2(SI_3_), .ZN(n5546) );
  NAND2_X1 U7168 ( .A1(n5446), .A2(SI_5_), .ZN(n5447) );
  MUX2_X1 U7169 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n4403), .Z(n5577) );
  XNOR2_X1 U7170 ( .A(n5577), .B(SI_6_), .ZN(n5574) );
  XNOR2_X1 U7171 ( .A(n5576), .B(n5574), .ZN(n7309) );
  XNOR2_X2 U7172 ( .A(n5449), .B(n10340), .ZN(n6120) );
  NAND2_X2 U7173 ( .A1(n7287), .A2(n4409), .ZN(n5531) );
  NAND2_X1 U7174 ( .A1(n7309), .A2(n6953), .ZN(n5455) );
  INV_X1 U7175 ( .A(n5563), .ZN(n5453) );
  INV_X1 U7176 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U7177 ( .A1(n5453), .A2(n5452), .ZN(n5616) );
  NAND2_X1 U7178 ( .A1(n5616), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5581) );
  XNOR2_X1 U7179 ( .A(n5581), .B(P1_IR_REG_6__SCAN_IN), .ZN(n7400) );
  AOI22_X1 U7180 ( .A1(n5579), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5885), .B2(
        n7400), .ZN(n5454) );
  NAND2_X1 U7181 ( .A1(n5455), .A2(n5454), .ZN(n7912) );
  OAI22_X1 U7182 ( .A1(n7897), .A2(n6057), .B1(n7909), .B2(n5979), .ZN(n5467)
         );
  NAND2_X1 U7183 ( .A1(n5884), .A2(n5458), .ZN(n5459) );
  NAND2_X1 U7184 ( .A1(n5462), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U7185 ( .A1(n5464), .A2(n5463), .ZN(n6103) );
  OR2_X1 U7186 ( .A1(n5464), .A2(n5463), .ZN(n5465) );
  NAND2_X1 U7187 ( .A1(n6968), .A2(n8088), .ZN(n5466) );
  NAND2_X1 U7188 ( .A1(n9464), .A2(n9400), .ZN(n9332) );
  XNOR2_X1 U7189 ( .A(n5467), .B(n8327), .ZN(n7872) );
  INV_X1 U7190 ( .A(n7872), .ZN(n5573) );
  INV_X2 U7191 ( .A(n5468), .ZN(n6057) );
  AND2_X1 U7192 ( .A1(n7912), .A2(n5468), .ZN(n5469) );
  AOI21_X1 U7193 ( .B1(n9484), .B2(n9036), .A(n5469), .ZN(n7871) );
  INV_X1 U7194 ( .A(n7871), .ZN(n5572) );
  INV_X1 U7195 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5470) );
  INV_X1 U7196 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5471) );
  OR2_X1 U7197 ( .A1(n5484), .A2(n5471), .ZN(n5472) );
  OR2_X1 U7198 ( .A1(n9220), .A2(n7323), .ZN(n5479) );
  XNOR2_X1 U7199 ( .A(n5475), .B(SI_1_), .ZN(n5509) );
  XNOR2_X1 U7200 ( .A(n5476), .B(n5509), .ZN(n6171) );
  INV_X1 U7201 ( .A(n6171), .ZN(n7322) );
  INV_X1 U7202 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5483) );
  INV_X1 U7203 ( .A(SI_0_), .ZN(n5487) );
  INV_X1 U7204 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5488) );
  XNOR2_X1 U7205 ( .A(n5489), .B(n5488), .ZN(n10042) );
  MUX2_X1 U7206 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10042), .S(n7287), .Z(n7695)
         );
  NAND2_X1 U7207 ( .A1(n4810), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5492) );
  NAND2_X1 U7208 ( .A1(n5495), .A2(n5492), .ZN(n7277) );
  AOI22_X1 U7209 ( .A1(n7695), .A2(n5822), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n4810), .ZN(n5493) );
  NAND2_X1 U7210 ( .A1(n5494), .A2(n5493), .ZN(n7276) );
  AND2_X1 U7211 ( .A1(n5495), .A2(n8327), .ZN(n5496) );
  NAND2_X1 U7212 ( .A1(n5777), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U7213 ( .A1(n4405), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5504) );
  NAND2_X1 U7214 ( .A1(n6986), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U7215 ( .A1(n5501), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5502) );
  NAND2_X1 U7216 ( .A1(n9489), .A2(n5822), .ZN(n5518) );
  INV_X1 U7217 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U7218 ( .A1(n5509), .A2(n5508), .ZN(n5511) );
  NAND2_X1 U7219 ( .A1(n5511), .A2(n5510), .ZN(n5514) );
  XNOR2_X1 U7220 ( .A(n5512), .B(SI_2_), .ZN(n5513) );
  XNOR2_X1 U7221 ( .A(n5514), .B(n5513), .ZN(n7317) );
  OR2_X1 U7222 ( .A1(n7317), .A2(n5531), .ZN(n5516) );
  OR2_X1 U7223 ( .A1(n9220), .A2(n10306), .ZN(n5515) );
  OAI211_X1 U7224 ( .C1(n7287), .C2(n7316), .A(n5516), .B(n5515), .ZN(n7710)
         );
  NAND2_X1 U7225 ( .A1(n7710), .A2(n9041), .ZN(n5517) );
  NAND2_X1 U7226 ( .A1(n5518), .A2(n5517), .ZN(n5519) );
  XNOR2_X1 U7227 ( .A(n5519), .B(n8327), .ZN(n5521) );
  OAI22_X1 U7228 ( .A1(n7849), .A2(n6056), .B1(n7589), .B2(n6057), .ZN(n5520)
         );
  XNOR2_X1 U7229 ( .A(n5521), .B(n5520), .ZN(n7698) );
  INV_X1 U7230 ( .A(n5520), .ZN(n5522) );
  NAND2_X1 U7231 ( .A1(n5501), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5528) );
  INV_X1 U7232 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7846) );
  NAND2_X1 U7233 ( .A1(n4405), .A2(n7846), .ZN(n5527) );
  INV_X1 U7234 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5523) );
  OR2_X1 U7235 ( .A1(n4406), .A2(n5523), .ZN(n5526) );
  INV_X1 U7236 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5524) );
  OR2_X1 U7237 ( .A1(n4408), .A2(n5524), .ZN(n5525) );
  XNOR2_X1 U7238 ( .A(n5529), .B(n5530), .ZN(n7318) );
  OR2_X1 U7239 ( .A1(n7318), .A2(n5531), .ZN(n5535) );
  OR2_X1 U7240 ( .A1(n9220), .A2(n10329), .ZN(n5534) );
  OR2_X1 U7241 ( .A1(n7287), .A2(n7357), .ZN(n5533) );
  OAI22_X1 U7242 ( .A1(n6922), .A2(n8329), .B1(n7848), .B2(n6057), .ZN(n5538)
         );
  OAI22_X1 U7243 ( .A1(n6922), .A2(n6057), .B1(n7848), .B2(n5979), .ZN(n5536)
         );
  XNOR2_X1 U7244 ( .A(n5536), .B(n8327), .ZN(n5537) );
  XOR2_X1 U7245 ( .A(n5538), .B(n5537), .Z(n7783) );
  NAND2_X1 U7246 ( .A1(n5501), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5543) );
  OAI21_X1 U7247 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(P1_REG3_REG_4__SCAN_IN), 
        .A(n5555), .ZN(n7737) );
  INV_X1 U7248 ( .A(n7737), .ZN(n7817) );
  NAND2_X1 U7249 ( .A1(n4405), .A2(n7817), .ZN(n5542) );
  INV_X1 U7250 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5539) );
  INV_X1 U7251 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7736) );
  OR2_X1 U7252 ( .A1(n4408), .A2(n7736), .ZN(n5540) );
  NAND2_X1 U7253 ( .A1(n5451), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5544) );
  MUX2_X1 U7254 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5544), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5545) );
  NAND2_X1 U7255 ( .A1(n5545), .A2(n5563), .ZN(n10099) );
  XNOR2_X1 U7256 ( .A(n5547), .B(SI_4_), .ZN(n5565) );
  INV_X1 U7257 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7320) );
  OAI22_X1 U7258 ( .A1(n7885), .A2(n8329), .B1(n7812), .B2(n6057), .ZN(n5550)
         );
  OAI22_X1 U7259 ( .A1(n7885), .A2(n6057), .B1(n7812), .B2(n5979), .ZN(n5548)
         );
  XNOR2_X1 U7260 ( .A(n5548), .B(n8327), .ZN(n5549) );
  XOR2_X1 U7261 ( .A(n5550), .B(n5549), .Z(n7814) );
  INV_X1 U7262 ( .A(n5549), .ZN(n5551) );
  INV_X1 U7263 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5552) );
  INV_X1 U7264 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5554) );
  NAND2_X1 U7265 ( .A1(n5555), .A2(n5554), .ZN(n5556) );
  AND2_X1 U7266 ( .A1(n5557), .A2(n5556), .ZN(n7889) );
  INV_X1 U7267 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U7268 ( .A1(n5563), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5564) );
  XNOR2_X1 U7269 ( .A(n5564), .B(P1_IR_REG_5__SCAN_IN), .ZN(n7384) );
  OAI22_X1 U7270 ( .A1(n4645), .A2(n6057), .B1(n7840), .B2(n5979), .ZN(n5570)
         );
  XNOR2_X1 U7271 ( .A(n5570), .B(n8327), .ZN(n5571) );
  OAI22_X1 U7272 ( .A1(n4645), .A2(n8329), .B1(n7840), .B2(n6057), .ZN(n7882)
         );
  INV_X1 U7273 ( .A(n5574), .ZN(n5575) );
  NAND2_X1 U7274 ( .A1(n5577), .A2(SI_6_), .ZN(n5578) );
  MUX2_X1 U7275 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4409), .Z(n5603) );
  XNOR2_X1 U7276 ( .A(n5603), .B(SI_7_), .ZN(n5600) );
  XNOR2_X1 U7277 ( .A(n5602), .B(n5600), .ZN(n7326) );
  NAND2_X1 U7278 ( .A1(n7326), .A2(n6953), .ZN(n5585) );
  INV_X1 U7279 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U7280 ( .A1(n5581), .A2(n5580), .ZN(n5582) );
  NAND2_X1 U7281 ( .A1(n5582), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5583) );
  XNOR2_X1 U7282 ( .A(n5583), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7479) );
  AOI22_X1 U7283 ( .A1(n5579), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5885), .B2(
        n7479), .ZN(n5584) );
  NAND2_X1 U7284 ( .A1(n5501), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U7285 ( .A1(n5777), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U7286 ( .A1(n5586), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5634) );
  INV_X1 U7287 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U7288 ( .A1(n5588), .A2(n5587), .ZN(n5589) );
  AND2_X1 U7289 ( .A1(n5634), .A2(n5589), .ZN(n8060) );
  NAND2_X1 U7290 ( .A1(n4405), .A2(n8060), .ZN(n5591) );
  NAND2_X1 U7291 ( .A1(n6986), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5590) );
  NAND2_X1 U7292 ( .A1(n9483), .A2(n5822), .ZN(n5594) );
  OAI21_X1 U7293 ( .B1(n8058), .B2(n5979), .A(n5594), .ZN(n5595) );
  XNOR2_X1 U7294 ( .A(n5595), .B(n9039), .ZN(n5599) );
  OR2_X1 U7295 ( .A1(n8058), .A2(n6057), .ZN(n5597) );
  NAND2_X1 U7296 ( .A1(n9036), .A2(n9483), .ZN(n5596) );
  NAND2_X1 U7297 ( .A1(n5597), .A2(n5596), .ZN(n5598) );
  NAND2_X1 U7298 ( .A1(n5599), .A2(n5598), .ZN(n8053) );
  INV_X1 U7299 ( .A(n5600), .ZN(n5601) );
  NAND2_X1 U7300 ( .A1(n5603), .A2(SI_7_), .ZN(n5604) );
  INV_X1 U7301 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5605) );
  INV_X1 U7302 ( .A(SI_8_), .ZN(n5606) );
  NAND2_X1 U7303 ( .A1(n5607), .A2(n5606), .ZN(n5610) );
  INV_X1 U7304 ( .A(n5607), .ZN(n5608) );
  NAND2_X1 U7305 ( .A1(n5608), .A2(SI_8_), .ZN(n5609) );
  NAND2_X1 U7306 ( .A1(n5610), .A2(n5609), .ZN(n5628) );
  INV_X1 U7307 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5611) );
  INV_X1 U7308 ( .A(SI_9_), .ZN(n5612) );
  NAND2_X1 U7309 ( .A1(n5613), .A2(n5612), .ZN(n5651) );
  INV_X1 U7310 ( .A(n5613), .ZN(n5614) );
  NAND2_X1 U7311 ( .A1(n5614), .A2(SI_9_), .ZN(n5615) );
  NAND2_X1 U7312 ( .A1(n5662), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5617) );
  AOI22_X1 U7313 ( .A1(n5579), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5885), .B2(
        n7776), .ZN(n5618) );
  NAND2_X1 U7314 ( .A1(n6112), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5625) );
  INV_X1 U7315 ( .A(n5636), .ZN(n5619) );
  NAND2_X1 U7316 ( .A1(n5619), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5685) );
  INV_X1 U7317 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10362) );
  NAND2_X1 U7318 ( .A1(n5636), .A2(n10362), .ZN(n5620) );
  AND2_X1 U7319 ( .A1(n5685), .A2(n5620), .ZN(n9835) );
  NAND2_X1 U7320 ( .A1(n4405), .A2(n9835), .ZN(n5624) );
  INV_X1 U7321 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10397) );
  OR2_X1 U7322 ( .A1(n4406), .A2(n10397), .ZN(n5623) );
  INV_X1 U7323 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n5621) );
  OR2_X1 U7324 ( .A1(n4408), .A2(n5621), .ZN(n5622) );
  INV_X1 U7325 ( .A(n9063), .ZN(n9482) );
  AOI22_X1 U7326 ( .A1(n9838), .A2(n9041), .B1(n5822), .B2(n9482), .ZN(n5626)
         );
  XOR2_X1 U7327 ( .A(n8327), .B(n5626), .Z(n9137) );
  NOR2_X1 U7328 ( .A1(n9063), .A2(n8329), .ZN(n5627) );
  AOI21_X1 U7329 ( .B1(n9838), .B2(n5822), .A(n5627), .ZN(n9136) );
  XNOR2_X1 U7330 ( .A(n5628), .B(n5629), .ZN(n7330) );
  NAND2_X1 U7331 ( .A1(n7330), .A2(n6953), .ZN(n5633) );
  NAND2_X1 U7332 ( .A1(n5630), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5631) );
  AOI22_X1 U7333 ( .A1(n5579), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5885), .B2(
        n7562), .ZN(n5632) );
  NAND2_X1 U7334 ( .A1(n9965), .A2(n5822), .ZN(n5643) );
  NAND2_X1 U7335 ( .A1(n6112), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U7336 ( .A1(n5634), .A2(n7482), .ZN(n5635) );
  AND2_X1 U7337 ( .A1(n5636), .A2(n5635), .ZN(n9059) );
  NAND2_X1 U7338 ( .A1(n4405), .A2(n9059), .ZN(n5640) );
  INV_X1 U7339 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10525) );
  OR2_X1 U7340 ( .A1(n4406), .A2(n10525), .ZN(n5639) );
  INV_X1 U7341 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5637) );
  OR2_X1 U7342 ( .A1(n4408), .A2(n5637), .ZN(n5638) );
  NAND2_X1 U7343 ( .A1(n5051), .A2(n9036), .ZN(n5642) );
  NAND2_X1 U7344 ( .A1(n9965), .A2(n9041), .ZN(n5645) );
  NAND2_X1 U7345 ( .A1(n5051), .A2(n5822), .ZN(n5644) );
  NAND2_X1 U7346 ( .A1(n5645), .A2(n5644), .ZN(n5646) );
  XNOR2_X1 U7347 ( .A(n5646), .B(n8327), .ZN(n9056) );
  OAI22_X1 U7348 ( .A1(n9137), .A2(n9136), .B1(n9058), .B2(n9056), .ZN(n5650)
         );
  INV_X1 U7349 ( .A(n9056), .ZN(n9135) );
  INV_X1 U7350 ( .A(n9058), .ZN(n5647) );
  NOR2_X1 U7351 ( .A1(n9135), .A2(n5647), .ZN(n5648) );
  OAI21_X1 U7352 ( .B1(n9136), .B2(n5648), .A(n9137), .ZN(n5649) );
  INV_X1 U7353 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5652) );
  MUX2_X1 U7354 ( .A(n10330), .B(n5652), .S(n4409), .Z(n5654) );
  XNOR2_X1 U7355 ( .A(n5654), .B(SI_10_), .ZN(n5679) );
  INV_X1 U7356 ( .A(n5679), .ZN(n5653) );
  INV_X1 U7357 ( .A(n5654), .ZN(n5655) );
  NAND2_X1 U7358 ( .A1(n5655), .A2(SI_10_), .ZN(n5656) );
  INV_X1 U7359 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5657) );
  MUX2_X1 U7360 ( .A(n7395), .B(n5657), .S(n4409), .Z(n5659) );
  INV_X1 U7361 ( .A(SI_11_), .ZN(n5658) );
  NAND2_X1 U7362 ( .A1(n5659), .A2(n5658), .ZN(n5752) );
  INV_X1 U7363 ( .A(n5659), .ZN(n5660) );
  NAND2_X1 U7364 ( .A1(n5660), .A2(SI_11_), .ZN(n5661) );
  NAND2_X1 U7365 ( .A1(n5752), .A2(n5661), .ZN(n5706) );
  NAND2_X1 U7366 ( .A1(n7392), .A2(n6953), .ZN(n5667) );
  OAI21_X1 U7367 ( .B1(n5662), .B2(P1_IR_REG_9__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5681) );
  INV_X1 U7368 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U7369 ( .A1(n5681), .A2(n5663), .ZN(n5664) );
  NAND2_X1 U7370 ( .A1(n5664), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5665) );
  AOI22_X1 U7371 ( .A1(n5579), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5885), .B2(
        n8194), .ZN(n5666) );
  NAND2_X1 U7372 ( .A1(n5667), .A2(n5666), .ZN(n8074) );
  NAND2_X1 U7373 ( .A1(n8074), .A2(n9041), .ZN(n5677) );
  NAND2_X1 U7374 ( .A1(n5668), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5713) );
  INV_X1 U7375 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5669) );
  NAND2_X1 U7376 ( .A1(n5687), .A2(n5669), .ZN(n5670) );
  AND2_X1 U7377 ( .A1(n5713), .A2(n5670), .ZN(n9186) );
  NAND2_X1 U7378 ( .A1(n4405), .A2(n9186), .ZN(n5675) );
  NAND2_X1 U7379 ( .A1(n6112), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5674) );
  INV_X1 U7380 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10014) );
  OR2_X1 U7381 ( .A1(n4406), .A2(n10014), .ZN(n5673) );
  INV_X1 U7382 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n5671) );
  OR2_X1 U7383 ( .A1(n4408), .A2(n5671), .ZN(n5672) );
  INV_X1 U7384 ( .A(n9091), .ZN(n9480) );
  NAND2_X1 U7385 ( .A1(n9480), .A2(n5822), .ZN(n5676) );
  NAND2_X1 U7386 ( .A1(n5677), .A2(n5676), .ZN(n5678) );
  XNOR2_X1 U7387 ( .A(n5678), .B(n9039), .ZN(n9177) );
  OAI22_X1 U7388 ( .A1(n10017), .A2(n6057), .B1(n9091), .B2(n6056), .ZN(n5700)
         );
  XNOR2_X1 U7389 ( .A(n5680), .B(n5679), .ZN(n7343) );
  NAND2_X1 U7390 ( .A1(n7343), .A2(n6953), .ZN(n5683) );
  XNOR2_X1 U7391 ( .A(n5681), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7863) );
  AOI22_X1 U7392 ( .A1(n5579), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5885), .B2(
        n7863), .ZN(n5682) );
  NAND2_X1 U7393 ( .A1(n5683), .A2(n5682), .ZN(n8097) );
  NAND2_X1 U7394 ( .A1(n8097), .A2(n9041), .ZN(n5695) );
  NAND2_X1 U7395 ( .A1(n5685), .A2(n5684), .ZN(n5686) );
  AND2_X1 U7396 ( .A1(n5687), .A2(n5686), .ZN(n9021) );
  NAND2_X1 U7397 ( .A1(n4405), .A2(n9021), .ZN(n5693) );
  NAND2_X1 U7398 ( .A1(n6112), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5692) );
  INV_X1 U7399 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5688) );
  OR2_X1 U7400 ( .A1(n4406), .A2(n5688), .ZN(n5691) );
  INV_X1 U7401 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n5689) );
  OR2_X1 U7402 ( .A1(n4408), .A2(n5689), .ZN(n5690) );
  NAND2_X1 U7403 ( .A1(n9481), .A2(n5822), .ZN(n5694) );
  NAND2_X1 U7404 ( .A1(n5695), .A2(n5694), .ZN(n5696) );
  XNOR2_X1 U7405 ( .A(n5696), .B(n8327), .ZN(n9175) );
  NOR2_X1 U7406 ( .A1(n9183), .A2(n8329), .ZN(n5697) );
  AOI21_X1 U7407 ( .B1(n8097), .B2(n5822), .A(n5697), .ZN(n9013) );
  NOR2_X1 U7408 ( .A1(n9175), .A2(n9013), .ZN(n5698) );
  INV_X1 U7409 ( .A(n5700), .ZN(n9178) );
  AOI21_X1 U7410 ( .B1(n9013), .B2(n9175), .A(n9178), .ZN(n5701) );
  NAND3_X1 U7411 ( .A1(n9178), .A2(n9013), .A3(n9175), .ZN(n5702) );
  AND2_X1 U7412 ( .A1(n5703), .A2(n5702), .ZN(n5704) );
  INV_X1 U7413 ( .A(n5706), .ZN(n5707) );
  MUX2_X1 U7414 ( .A(n7438), .B(n7444), .S(n4409), .Z(n5753) );
  XNOR2_X1 U7415 ( .A(n5753), .B(SI_12_), .ZN(n5728) );
  NAND2_X1 U7416 ( .A1(n7437), .A2(n6953), .ZN(n5712) );
  NAND2_X1 U7417 ( .A1(n5456), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5708) );
  MUX2_X1 U7418 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5708), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n5710) );
  INV_X1 U7419 ( .A(n5733), .ZN(n5709) );
  NAND2_X1 U7420 ( .A1(n5710), .A2(n5709), .ZN(n8195) );
  INV_X1 U7421 ( .A(n8195), .ZN(n9513) );
  AOI22_X1 U7422 ( .A1(n5579), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5885), .B2(
        n9513), .ZN(n5711) );
  NAND2_X1 U7423 ( .A1(n6112), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5720) );
  NAND2_X1 U7424 ( .A1(n5713), .A2(n9087), .ZN(n5714) );
  AND2_X1 U7425 ( .A1(n5738), .A2(n5714), .ZN(n9088) );
  NAND2_X1 U7426 ( .A1(n4405), .A2(n9088), .ZN(n5719) );
  INV_X1 U7427 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5715) );
  OR2_X1 U7428 ( .A1(n4406), .A2(n5715), .ZN(n5718) );
  INV_X1 U7429 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n5716) );
  OR2_X1 U7430 ( .A1(n4408), .A2(n5716), .ZN(n5717) );
  AOI22_X1 U7431 ( .A1(n9093), .A2(n5822), .B1(n9036), .B2(n9479), .ZN(n5724)
         );
  NAND2_X1 U7432 ( .A1(n9093), .A2(n9041), .ZN(n5722) );
  NAND2_X1 U7433 ( .A1(n9479), .A2(n5822), .ZN(n5721) );
  NAND2_X1 U7434 ( .A1(n5722), .A2(n5721), .ZN(n5723) );
  XNOR2_X1 U7435 ( .A(n5723), .B(n8327), .ZN(n5725) );
  XOR2_X1 U7436 ( .A(n5724), .B(n5725), .Z(n9086) );
  NAND2_X1 U7437 ( .A1(n5725), .A2(n5724), .ZN(n5726) );
  NAND2_X1 U7438 ( .A1(n5727), .A2(n5726), .ZN(n9156) );
  INV_X1 U7439 ( .A(n5728), .ZN(n5730) );
  INV_X1 U7440 ( .A(n5753), .ZN(n5729) );
  NAND2_X1 U7441 ( .A1(n5729), .A2(SI_12_), .ZN(n5754) );
  MUX2_X1 U7442 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n4409), .Z(n5758) );
  XNOR2_X1 U7443 ( .A(n5758), .B(SI_13_), .ZN(n5751) );
  XNOR2_X1 U7444 ( .A(n5732), .B(n5751), .ZN(n7472) );
  NAND2_X1 U7445 ( .A1(n7472), .A2(n6953), .ZN(n5736) );
  OR2_X1 U7446 ( .A1(n5733), .A2(n10021), .ZN(n5734) );
  XNOR2_X1 U7447 ( .A(n5734), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9521) );
  AOI22_X1 U7448 ( .A1(n5579), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5885), .B2(
        n9521), .ZN(n5735) );
  NAND2_X1 U7449 ( .A1(n5738), .A2(n5737), .ZN(n5739) );
  AND2_X1 U7450 ( .A1(n5812), .A2(n5739), .ZN(n9826) );
  NAND2_X1 U7451 ( .A1(n4405), .A2(n9826), .ZN(n5744) );
  NAND2_X1 U7452 ( .A1(n6112), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5743) );
  INV_X1 U7453 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10009) );
  OR2_X1 U7454 ( .A1(n4406), .A2(n10009), .ZN(n5742) );
  INV_X1 U7455 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n5740) );
  OR2_X1 U7456 ( .A1(n4408), .A2(n5740), .ZN(n5741) );
  AOI22_X1 U7457 ( .A1(n9941), .A2(n5822), .B1(n9036), .B2(n9478), .ZN(n5748)
         );
  NAND2_X1 U7458 ( .A1(n9941), .A2(n9041), .ZN(n5746) );
  NAND2_X1 U7459 ( .A1(n9478), .A2(n5822), .ZN(n5745) );
  NAND2_X1 U7460 ( .A1(n5746), .A2(n5745), .ZN(n5747) );
  XNOR2_X1 U7461 ( .A(n5747), .B(n8327), .ZN(n5749) );
  XOR2_X1 U7462 ( .A(n5748), .B(n5749), .Z(n9157) );
  NAND2_X1 U7463 ( .A1(n5749), .A2(n5748), .ZN(n5750) );
  INV_X1 U7464 ( .A(n5751), .ZN(n5757) );
  INV_X1 U7465 ( .A(n5752), .ZN(n5755) );
  INV_X1 U7466 ( .A(SI_12_), .ZN(n10453) );
  AOI22_X1 U7467 ( .A1(n5755), .A2(n5754), .B1(n5753), .B2(n10453), .ZN(n5756)
         );
  MUX2_X1 U7468 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4409), .Z(n5760) );
  XNOR2_X1 U7469 ( .A(n5760), .B(SI_14_), .ZN(n5804) );
  INV_X1 U7470 ( .A(n5804), .ZN(n5759) );
  NAND2_X1 U7471 ( .A1(n5760), .A2(SI_14_), .ZN(n5761) );
  INV_X1 U7472 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n5763) );
  MUX2_X1 U7473 ( .A(n7516), .B(n5763), .S(n4409), .Z(n5765) );
  INV_X1 U7474 ( .A(SI_15_), .ZN(n5764) );
  NOR2_X1 U7475 ( .A1(n5765), .A2(n5764), .ZN(n5766) );
  INV_X1 U7476 ( .A(n5765), .ZN(n5787) );
  MUX2_X1 U7477 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n4409), .Z(n5834) );
  INV_X1 U7478 ( .A(n5834), .ZN(n5767) );
  XNOR2_X1 U7479 ( .A(n5767), .B(SI_16_), .ZN(n5768) );
  XNOR2_X1 U7480 ( .A(n5833), .B(n5768), .ZN(n7553) );
  NAND2_X1 U7481 ( .A1(n7553), .A2(n6953), .ZN(n5773) );
  NAND2_X1 U7482 ( .A1(n5769), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5770) );
  MUX2_X1 U7483 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5770), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n5771) );
  AOI22_X1 U7484 ( .A1(n5579), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5885), .B2(
        n10112), .ZN(n5772) );
  NAND2_X1 U7485 ( .A1(n9925), .A2(n9041), .ZN(n5783) );
  INV_X1 U7486 ( .A(n5814), .ZN(n5774) );
  NAND2_X1 U7487 ( .A1(n5796), .A2(n5775), .ZN(n5776) );
  AND2_X1 U7488 ( .A1(n5846), .A2(n5776), .ZN(n9761) );
  NAND2_X1 U7489 ( .A1(n9761), .A2(n4405), .ZN(n5781) );
  AOI22_X1 U7490 ( .A1(n5777), .A2(P1_REG0_REG_16__SCAN_IN), .B1(n6112), .B2(
        P1_REG1_REG_16__SCAN_IN), .ZN(n5780) );
  INV_X1 U7491 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n5778) );
  OR2_X1 U7492 ( .A1(n4408), .A2(n5778), .ZN(n5779) );
  OR2_X1 U7493 ( .A1(n9919), .A2(n6057), .ZN(n5782) );
  NAND2_X1 U7494 ( .A1(n5783), .A2(n5782), .ZN(n5784) );
  XNOR2_X1 U7495 ( .A(n5784), .B(n9039), .ZN(n9109) );
  NAND2_X1 U7496 ( .A1(n9925), .A2(n5822), .ZN(n5786) );
  OR2_X1 U7497 ( .A1(n9919), .A2(n6056), .ZN(n5785) );
  NAND2_X1 U7498 ( .A1(n5786), .A2(n5785), .ZN(n9108) );
  XNOR2_X1 U7499 ( .A(n5787), .B(SI_15_), .ZN(n5788) );
  NOR2_X1 U7500 ( .A1(n5789), .A2(n10021), .ZN(n5806) );
  INV_X1 U7501 ( .A(n5806), .ZN(n5791) );
  INV_X1 U7502 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U7503 ( .A1(n5791), .A2(n5790), .ZN(n5807) );
  NAND2_X1 U7504 ( .A1(n5807), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5792) );
  XNOR2_X1 U7505 ( .A(n5792), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9549) );
  AOI22_X1 U7506 ( .A1(n5579), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5885), .B2(
        n9549), .ZN(n5793) );
  INV_X1 U7507 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U7508 ( .A1(n5814), .A2(n5794), .ZN(n5795) );
  NAND2_X1 U7509 ( .A1(n5796), .A2(n5795), .ZN(n9786) );
  INV_X1 U7510 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9787) );
  OAI22_X1 U7511 ( .A1(n9786), .A2(n6985), .B1(n4408), .B2(n9787), .ZN(n5799)
         );
  INV_X1 U7512 ( .A(n6112), .ZN(n6989) );
  NAND2_X1 U7513 ( .A1(n5777), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5797) );
  OAI21_X1 U7514 ( .B1(n10572), .B2(n6989), .A(n5797), .ZN(n5798) );
  NAND2_X1 U7515 ( .A1(n9803), .A2(n5822), .ZN(n5800) );
  XNOR2_X1 U7516 ( .A(n5801), .B(n9039), .ZN(n9107) );
  NAND2_X1 U7517 ( .A1(n9789), .A2(n5822), .ZN(n5803) );
  NAND2_X1 U7518 ( .A1(n9803), .A2(n9036), .ZN(n5802) );
  NAND2_X1 U7519 ( .A1(n5803), .A2(n5802), .ZN(n9106) );
  AOI22_X1 U7520 ( .A1(n9109), .A2(n9108), .B1(n9107), .B2(n9106), .ZN(n5826)
         );
  XNOR2_X1 U7521 ( .A(n5805), .B(n5804), .ZN(n7439) );
  NAND2_X1 U7522 ( .A1(n7439), .A2(n6953), .ZN(n5810) );
  NAND2_X1 U7523 ( .A1(n5806), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5808) );
  AOI22_X1 U7524 ( .A1(n5579), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5885), .B2(
        n9535), .ZN(n5809) );
  NAND2_X1 U7525 ( .A1(n9937), .A2(n9041), .ZN(n5820) );
  NAND2_X1 U7526 ( .A1(n6112), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5818) );
  NAND2_X1 U7527 ( .A1(n5777), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5817) );
  INV_X1 U7528 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5811) );
  NAND2_X1 U7529 ( .A1(n5812), .A2(n5811), .ZN(n5813) );
  AND2_X1 U7530 ( .A1(n5814), .A2(n5813), .ZN(n9795) );
  NAND2_X1 U7531 ( .A1(n4405), .A2(n9795), .ZN(n5816) );
  NAND2_X1 U7532 ( .A1(n6986), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5815) );
  NAND4_X1 U7533 ( .A1(n5818), .A2(n5817), .A3(n5816), .A4(n5815), .ZN(n9779)
         );
  NAND2_X1 U7534 ( .A1(n9779), .A2(n5822), .ZN(n5819) );
  NAND2_X1 U7535 ( .A1(n5820), .A2(n5819), .ZN(n5821) );
  XNOR2_X1 U7536 ( .A(n5821), .B(n8327), .ZN(n9104) );
  NAND2_X1 U7537 ( .A1(n9937), .A2(n5822), .ZN(n5824) );
  NAND2_X1 U7538 ( .A1(n9036), .A2(n9779), .ZN(n5823) );
  NAND3_X1 U7539 ( .A1(n5826), .A2(n8994), .A3(n9104), .ZN(n5831) );
  INV_X1 U7540 ( .A(n9109), .ZN(n5829) );
  OAI21_X1 U7541 ( .B1(n9107), .B2(n9106), .A(n9108), .ZN(n5828) );
  NOR2_X1 U7542 ( .A1(n9108), .A2(n9106), .ZN(n5827) );
  INV_X1 U7543 ( .A(n9107), .ZN(n9105) );
  AOI22_X1 U7544 ( .A1(n5829), .A2(n5828), .B1(n5827), .B2(n9105), .ZN(n5830)
         );
  NAND2_X1 U7545 ( .A1(n5834), .A2(SI_16_), .ZN(n5835) );
  MUX2_X1 U7546 ( .A(n7691), .B(n5836), .S(n4409), .Z(n5837) );
  NAND2_X1 U7547 ( .A1(n5837), .A2(n10409), .ZN(n5858) );
  INV_X1 U7548 ( .A(n5837), .ZN(n5838) );
  NAND2_X1 U7549 ( .A1(n5838), .A2(SI_17_), .ZN(n5839) );
  NAND2_X1 U7550 ( .A1(n5858), .A2(n5839), .ZN(n5856) );
  NAND2_X1 U7551 ( .A1(n7641), .A2(n6953), .ZN(n5843) );
  NAND2_X1 U7552 ( .A1(n5840), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5841) );
  XNOR2_X1 U7553 ( .A(n5841), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10128) );
  AOI22_X1 U7554 ( .A1(n5579), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5885), .B2(
        n10128), .ZN(n5842) );
  INV_X1 U7555 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n5850) );
  INV_X1 U7556 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U7557 ( .A1(n5846), .A2(n5845), .ZN(n5847) );
  NAND2_X1 U7558 ( .A1(n5889), .A2(n5847), .ZN(n9748) );
  OR2_X1 U7559 ( .A1(n9748), .A2(n6985), .ZN(n5849) );
  AOI22_X1 U7560 ( .A1(n5777), .A2(P1_REG0_REG_17__SCAN_IN), .B1(n6112), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n5848) );
  OAI211_X1 U7561 ( .C1(n4408), .C2(n5850), .A(n5849), .B(n5848), .ZN(n9767)
         );
  AOI22_X1 U7562 ( .A1(n9755), .A2(n5468), .B1(n9036), .B2(n9767), .ZN(n5854)
         );
  NAND2_X1 U7563 ( .A1(n9755), .A2(n9041), .ZN(n5852) );
  NAND2_X1 U7564 ( .A1(n9767), .A2(n5822), .ZN(n5851) );
  NAND2_X1 U7565 ( .A1(n5852), .A2(n5851), .ZN(n5853) );
  XNOR2_X1 U7566 ( .A(n5853), .B(n8327), .ZN(n5855) );
  XOR2_X1 U7567 ( .A(n5854), .B(n5855), .Z(n9119) );
  NAND2_X1 U7568 ( .A1(n5859), .A2(n5858), .ZN(n5883) );
  MUX2_X1 U7569 ( .A(n10487), .B(n5860), .S(n4409), .Z(n5861) );
  XNOR2_X1 U7570 ( .A(n5861), .B(SI_18_), .ZN(n5882) );
  INV_X1 U7571 ( .A(n5882), .ZN(n5864) );
  INV_X1 U7572 ( .A(n5861), .ZN(n5862) );
  NAND2_X1 U7573 ( .A1(n5862), .A2(SI_18_), .ZN(n5863) );
  MUX2_X1 U7574 ( .A(n7858), .B(n8319), .S(n4403), .Z(n5866) );
  INV_X1 U7575 ( .A(SI_19_), .ZN(n5865) );
  NAND2_X1 U7576 ( .A1(n5866), .A2(n5865), .ZN(n5912) );
  INV_X1 U7577 ( .A(n5866), .ZN(n5867) );
  NAND2_X1 U7578 ( .A1(n5867), .A2(SI_19_), .ZN(n5868) );
  NAND2_X1 U7579 ( .A1(n5912), .A2(n5868), .ZN(n5910) );
  NAND2_X1 U7580 ( .A1(n7856), .A2(n6953), .ZN(n5871) );
  AOI22_X1 U7581 ( .A1(n9556), .A2(n5885), .B1(n5579), .B2(
        P2_DATAO_REG_19__SCAN_IN), .ZN(n5870) );
  INV_X1 U7582 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5872) );
  NAND2_X1 U7583 ( .A1(n5891), .A2(n5872), .ZN(n5873) );
  NAND2_X1 U7584 ( .A1(n5917), .A2(n5873), .ZN(n9722) );
  OR2_X1 U7585 ( .A1(n9722), .A2(n6985), .ZN(n5878) );
  INV_X1 U7586 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9721) );
  NAND2_X1 U7587 ( .A1(n6112), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U7588 ( .A1(n5777), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5874) );
  OAI211_X1 U7589 ( .C1(n9721), .C2(n4408), .A(n5875), .B(n5874), .ZN(n5876)
         );
  INV_X1 U7590 ( .A(n5876), .ZN(n5877) );
  NAND2_X1 U7591 ( .A1(n9720), .A2(n5468), .ZN(n5881) );
  NAND2_X1 U7592 ( .A1(n9477), .A2(n9036), .ZN(n5880) );
  NAND2_X1 U7593 ( .A1(n5881), .A2(n5880), .ZN(n5905) );
  XNOR2_X1 U7594 ( .A(n5883), .B(n5882), .ZN(n7741) );
  NAND2_X1 U7595 ( .A1(n7741), .A2(n6953), .ZN(n5887) );
  XNOR2_X1 U7596 ( .A(n5884), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10145) );
  AOI22_X1 U7597 ( .A1(n5579), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n10145), 
        .B2(n5885), .ZN(n5886) );
  NAND2_X1 U7598 ( .A1(n9914), .A2(n9041), .ZN(n5898) );
  NAND2_X1 U7599 ( .A1(n5889), .A2(n5888), .ZN(n5890) );
  AND2_X1 U7600 ( .A1(n5891), .A2(n5890), .ZN(n9736) );
  NAND2_X1 U7601 ( .A1(n9736), .A2(n4405), .ZN(n5896) );
  INV_X1 U7602 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10439) );
  NAND2_X1 U7603 ( .A1(n6112), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5893) );
  NAND2_X1 U7604 ( .A1(n6986), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5892) );
  OAI211_X1 U7605 ( .C1(n4406), .C2(n10439), .A(n5893), .B(n5892), .ZN(n5894)
         );
  INV_X1 U7606 ( .A(n5894), .ZN(n5895) );
  NAND2_X1 U7607 ( .A1(n5896), .A2(n5895), .ZN(n9744) );
  NAND2_X1 U7608 ( .A1(n9744), .A2(n5822), .ZN(n5897) );
  NAND2_X1 U7609 ( .A1(n5898), .A2(n5897), .ZN(n5899) );
  XNOR2_X1 U7610 ( .A(n5899), .B(n9039), .ZN(n9025) );
  NAND2_X1 U7611 ( .A1(n9914), .A2(n5822), .ZN(n5901) );
  NAND2_X1 U7612 ( .A1(n9744), .A2(n9036), .ZN(n5900) );
  NAND2_X1 U7613 ( .A1(n5901), .A2(n5900), .ZN(n9191) );
  OAI22_X1 U7614 ( .A1(n9028), .A2(n5905), .B1(n9025), .B2(n9191), .ZN(n5908)
         );
  NAND2_X1 U7615 ( .A1(n9025), .A2(n9191), .ZN(n5903) );
  INV_X1 U7616 ( .A(n5903), .ZN(n5906) );
  INV_X1 U7617 ( .A(n5905), .ZN(n9027) );
  INV_X1 U7618 ( .A(n9028), .ZN(n5902) );
  AOI21_X1 U7619 ( .B1(n9027), .B2(n5903), .A(n5902), .ZN(n5904) );
  AOI21_X1 U7620 ( .B1(n5906), .B2(n5905), .A(n5904), .ZN(n5907) );
  INV_X1 U7621 ( .A(n5909), .ZN(n5911) );
  MUX2_X1 U7622 ( .A(n6452), .B(n7962), .S(n4409), .Z(n5955) );
  XNOR2_X1 U7623 ( .A(n5955), .B(SI_20_), .ZN(n5913) );
  XNOR2_X1 U7624 ( .A(n5962), .B(n5913), .ZN(n6451) );
  NAND2_X1 U7625 ( .A1(n6451), .A2(n6953), .ZN(n5915) );
  OR2_X1 U7626 ( .A1(n9220), .A2(n7962), .ZN(n5914) );
  NAND2_X1 U7627 ( .A1(n9903), .A2(n9041), .ZN(n5926) );
  NAND2_X1 U7628 ( .A1(n5917), .A2(n5916), .ZN(n5918) );
  AND2_X1 U7629 ( .A1(n5941), .A2(n5918), .ZN(n9696) );
  NAND2_X1 U7630 ( .A1(n9696), .A2(n4405), .ZN(n5924) );
  INV_X1 U7631 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n5921) );
  NAND2_X1 U7632 ( .A1(n6112), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5920) );
  NAND2_X1 U7633 ( .A1(n5777), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5919) );
  OAI211_X1 U7634 ( .C1(n5921), .C2(n4408), .A(n5920), .B(n5919), .ZN(n5922)
         );
  INV_X1 U7635 ( .A(n5922), .ZN(n5923) );
  NAND2_X1 U7636 ( .A1(n9712), .A2(n5822), .ZN(n5925) );
  NAND2_X1 U7637 ( .A1(n5926), .A2(n5925), .ZN(n5927) );
  XNOR2_X1 U7638 ( .A(n5927), .B(n8327), .ZN(n5929) );
  AND2_X1 U7639 ( .A1(n9712), .A2(n9036), .ZN(n5928) );
  AOI21_X1 U7640 ( .B1(n9903), .B2(n5468), .A(n5928), .ZN(n5930) );
  NAND2_X1 U7641 ( .A1(n5929), .A2(n5930), .ZN(n9148) );
  INV_X1 U7642 ( .A(n5929), .ZN(n5932) );
  INV_X1 U7643 ( .A(n5930), .ZN(n5931) );
  NAND2_X1 U7644 ( .A1(n5932), .A2(n5931), .ZN(n9147) );
  NAND2_X1 U7645 ( .A1(n5962), .A2(n5954), .ZN(n5933) );
  NAND2_X1 U7646 ( .A1(n5934), .A2(n5933), .ZN(n5936) );
  MUX2_X1 U7647 ( .A(n8081), .B(n8090), .S(n4403), .Z(n5953) );
  XNOR2_X1 U7648 ( .A(n5953), .B(SI_21_), .ZN(n5935) );
  NAND2_X1 U7649 ( .A1(n8080), .A2(n6953), .ZN(n5938) );
  OR2_X1 U7650 ( .A1(n9220), .A2(n8090), .ZN(n5937) );
  NAND2_X2 U7651 ( .A1(n5938), .A2(n5937), .ZN(n9896) );
  INV_X1 U7652 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U7653 ( .A1(n5941), .A2(n5940), .ZN(n5942) );
  NAND2_X1 U7654 ( .A1(n5971), .A2(n5942), .ZN(n9679) );
  OR2_X1 U7655 ( .A1(n9679), .A2(n6985), .ZN(n5947) );
  INV_X1 U7656 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9678) );
  NAND2_X1 U7657 ( .A1(n6112), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5944) );
  NAND2_X1 U7658 ( .A1(n5777), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5943) );
  OAI211_X1 U7659 ( .C1(n9678), .C2(n4408), .A(n5944), .B(n5943), .ZN(n5945)
         );
  INV_X1 U7660 ( .A(n5945), .ZN(n5946) );
  AOI22_X1 U7661 ( .A1(n9896), .A2(n5468), .B1(n9036), .B2(n9702), .ZN(n5950)
         );
  AOI22_X1 U7662 ( .A1(n9896), .A2(n9041), .B1(n5468), .B2(n9702), .ZN(n5948)
         );
  INV_X1 U7663 ( .A(n5949), .ZN(n5951) );
  NAND2_X1 U7664 ( .A1(n5951), .A2(n5950), .ZN(n5952) );
  INV_X1 U7665 ( .A(n5955), .ZN(n5957) );
  INV_X1 U7666 ( .A(n5953), .ZN(n5958) );
  OAI22_X1 U7667 ( .A1(n5957), .A2(SI_20_), .B1(n5958), .B2(SI_21_), .ZN(n5961) );
  OAI21_X1 U7668 ( .B1(n5955), .B2(n5954), .A(n10399), .ZN(n5959) );
  AND2_X1 U7669 ( .A1(SI_20_), .A2(SI_21_), .ZN(n5956) );
  AOI22_X1 U7670 ( .A1(n5959), .A2(n5958), .B1(n5957), .B2(n5956), .ZN(n5960)
         );
  MUX2_X1 U7671 ( .A(n8087), .B(n8084), .S(n4409), .Z(n5964) );
  INV_X1 U7672 ( .A(SI_22_), .ZN(n5963) );
  NAND2_X1 U7673 ( .A1(n5964), .A2(n5963), .ZN(n5987) );
  INV_X1 U7674 ( .A(n5964), .ZN(n5965) );
  NAND2_X1 U7675 ( .A1(n5965), .A2(SI_22_), .ZN(n5966) );
  NAND2_X1 U7676 ( .A1(n5987), .A2(n5966), .ZN(n5985) );
  XNOR2_X1 U7677 ( .A(n5986), .B(n5985), .ZN(n8083) );
  NAND2_X1 U7678 ( .A1(n8083), .A2(n6953), .ZN(n5968) );
  OR2_X1 U7679 ( .A1(n9220), .A2(n8084), .ZN(n5967) );
  INV_X1 U7680 ( .A(n5971), .ZN(n5969) );
  INV_X1 U7681 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5970) );
  NAND2_X1 U7682 ( .A1(n5971), .A2(n5970), .ZN(n5972) );
  NAND2_X1 U7683 ( .A1(n5997), .A2(n5972), .ZN(n9668) );
  OR2_X1 U7684 ( .A1(n9668), .A2(n6985), .ZN(n5978) );
  INV_X1 U7685 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U7686 ( .A1(n6112), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5974) );
  NAND2_X1 U7687 ( .A1(n5777), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5973) );
  OAI211_X1 U7688 ( .C1(n5975), .C2(n4408), .A(n5974), .B(n5973), .ZN(n5976)
         );
  INV_X1 U7689 ( .A(n5976), .ZN(n5977) );
  OAI22_X1 U7690 ( .A1(n9990), .A2(n5979), .B1(n9300), .B2(n6057), .ZN(n5980)
         );
  XNOR2_X1 U7691 ( .A(n5980), .B(n8327), .ZN(n5982) );
  AOI22_X1 U7692 ( .A1(n9673), .A2(n5468), .B1(n9036), .B2(n9688), .ZN(n9166)
         );
  NAND2_X1 U7693 ( .A1(n9164), .A2(n9166), .ZN(n5984) );
  NAND2_X1 U7694 ( .A1(n5983), .A2(n5982), .ZN(n9165) );
  MUX2_X1 U7695 ( .A(n8163), .B(n5995), .S(n4403), .Z(n5988) );
  INV_X1 U7696 ( .A(SI_23_), .ZN(n10364) );
  NAND2_X1 U7697 ( .A1(n5988), .A2(n10364), .ZN(n6013) );
  INV_X1 U7698 ( .A(n5988), .ZN(n5989) );
  NAND2_X1 U7699 ( .A1(n5989), .A2(SI_23_), .ZN(n5990) );
  NAND2_X1 U7700 ( .A1(n6013), .A2(n5990), .ZN(n5992) );
  NAND2_X1 U7701 ( .A1(n5991), .A2(n5992), .ZN(n6487) );
  INV_X1 U7702 ( .A(n5992), .ZN(n5993) );
  NAND2_X1 U7703 ( .A1(n6487), .A2(n6489), .ZN(n8165) );
  OR2_X1 U7704 ( .A1(n9220), .A2(n5995), .ZN(n5996) );
  NAND2_X1 U7705 ( .A1(n9656), .A2(n9041), .ZN(n6005) );
  INV_X1 U7706 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9008) );
  NAND2_X1 U7707 ( .A1(n5997), .A2(n9008), .ZN(n5998) );
  NAND2_X1 U7708 ( .A1(n6021), .A2(n5998), .ZN(n9658) );
  OR2_X1 U7709 ( .A1(n9658), .A2(n6985), .ZN(n6003) );
  INV_X1 U7710 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9657) );
  NAND2_X1 U7711 ( .A1(n6112), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U7712 ( .A1(n5777), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5999) );
  OAI211_X1 U7713 ( .C1(n9657), .C2(n4408), .A(n6000), .B(n5999), .ZN(n6001)
         );
  INV_X1 U7714 ( .A(n6001), .ZN(n6002) );
  NAND2_X1 U7715 ( .A1(n9876), .A2(n5468), .ZN(n6004) );
  NAND2_X1 U7716 ( .A1(n6005), .A2(n6004), .ZN(n6006) );
  XNOR2_X1 U7717 ( .A(n6006), .B(n9039), .ZN(n6009) );
  NAND2_X1 U7718 ( .A1(n9656), .A2(n5468), .ZN(n6008) );
  NAND2_X1 U7719 ( .A1(n9876), .A2(n9036), .ZN(n6007) );
  NAND2_X1 U7720 ( .A1(n6008), .A2(n6007), .ZN(n6010) );
  NAND2_X1 U7721 ( .A1(n6009), .A2(n6010), .ZN(n9003) );
  INV_X1 U7722 ( .A(n6009), .ZN(n6012) );
  INV_X1 U7723 ( .A(n6010), .ZN(n6011) );
  NAND2_X1 U7724 ( .A1(n6012), .A2(n6011), .ZN(n9004) );
  MUX2_X1 U7725 ( .A(n10520), .B(n10038), .S(n4403), .Z(n6015) );
  INV_X1 U7726 ( .A(SI_24_), .ZN(n6014) );
  NAND2_X1 U7727 ( .A1(n6015), .A2(n6014), .ZN(n6731) );
  INV_X1 U7728 ( .A(n6015), .ZN(n6016) );
  NAND2_X1 U7729 ( .A1(n6016), .A2(SI_24_), .ZN(n6017) );
  NAND2_X1 U7730 ( .A1(n8990), .A2(n6953), .ZN(n6019) );
  OR2_X1 U7731 ( .A1(n9220), .A2(n10038), .ZN(n6018) );
  NAND2_X1 U7732 ( .A1(n6980), .A2(n9041), .ZN(n6029) );
  INV_X1 U7733 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6020) );
  NAND2_X1 U7734 ( .A1(n6021), .A2(n6020), .ZN(n6022) );
  NAND2_X1 U7735 ( .A1(n9637), .A2(n4405), .ZN(n6027) );
  INV_X1 U7736 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10526) );
  NAND2_X1 U7737 ( .A1(n6986), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6024) );
  NAND2_X1 U7738 ( .A1(n5777), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6023) );
  OAI211_X1 U7739 ( .C1(n6989), .C2(n10526), .A(n6024), .B(n6023), .ZN(n6025)
         );
  INV_X1 U7740 ( .A(n6025), .ZN(n6026) );
  NAND2_X2 U7741 ( .A1(n6027), .A2(n6026), .ZN(n9650) );
  NAND2_X1 U7742 ( .A1(n9650), .A2(n5468), .ZN(n6028) );
  NAND2_X1 U7743 ( .A1(n6029), .A2(n6028), .ZN(n6030) );
  XNOR2_X1 U7744 ( .A(n6030), .B(n9039), .ZN(n6034) );
  NAND2_X1 U7745 ( .A1(n6980), .A2(n5822), .ZN(n6032) );
  NAND2_X1 U7746 ( .A1(n9650), .A2(n9036), .ZN(n6031) );
  NAND2_X1 U7747 ( .A1(n6032), .A2(n6031), .ZN(n6033) );
  NOR2_X1 U7748 ( .A1(n6034), .A2(n6033), .ZN(n6035) );
  AOI21_X1 U7749 ( .B1(n6034), .B2(n6033), .A(n6035), .ZN(n9128) );
  INV_X1 U7750 ( .A(n6035), .ZN(n6036) );
  INV_X1 U7751 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8988) );
  INV_X1 U7752 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10034) );
  MUX2_X1 U7753 ( .A(n8988), .B(n10034), .S(n4403), .Z(n6040) );
  NAND2_X1 U7754 ( .A1(n6040), .A2(n6039), .ZN(n6544) );
  INV_X1 U7755 ( .A(n6040), .ZN(n6041) );
  NAND2_X1 U7756 ( .A1(n6041), .A2(SI_25_), .ZN(n6042) );
  NAND2_X1 U7757 ( .A1(n8987), .A2(n6953), .ZN(n6044) );
  OR2_X1 U7758 ( .A1(n9220), .A2(n10034), .ZN(n6043) );
  NAND2_X1 U7759 ( .A1(n9625), .A2(n9041), .ZN(n6054) );
  INV_X1 U7760 ( .A(n6046), .ZN(n6045) );
  INV_X1 U7761 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n10394) );
  NAND2_X1 U7762 ( .A1(n6046), .A2(n10394), .ZN(n6047) );
  NAND2_X1 U7763 ( .A1(n6071), .A2(n6047), .ZN(n9622) );
  INV_X1 U7764 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9621) );
  NAND2_X1 U7765 ( .A1(n6112), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U7766 ( .A1(n5777), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6048) );
  OAI211_X1 U7767 ( .C1(n9621), .C2(n4408), .A(n6049), .B(n6048), .ZN(n6050)
         );
  INV_X1 U7768 ( .A(n6050), .ZN(n6051) );
  NAND2_X1 U7769 ( .A1(n9633), .A2(n5468), .ZN(n6053) );
  NAND2_X1 U7770 ( .A1(n6054), .A2(n6053), .ZN(n6055) );
  XNOR2_X1 U7771 ( .A(n6055), .B(n8327), .ZN(n6058) );
  OAI22_X1 U7772 ( .A1(n9982), .A2(n6057), .B1(n9608), .B2(n6056), .ZN(n6059)
         );
  XNOR2_X1 U7773 ( .A(n6058), .B(n6059), .ZN(n9097) );
  INV_X1 U7774 ( .A(n6086), .ZN(n6082) );
  INV_X1 U7775 ( .A(n6058), .ZN(n6060) );
  NOR2_X1 U7776 ( .A1(n6060), .A2(n6059), .ZN(n6083) );
  NAND2_X1 U7777 ( .A1(n6541), .A2(n6540), .ZN(n6061) );
  NAND2_X1 U7778 ( .A1(n6061), .A2(n6544), .ZN(n6066) );
  INV_X1 U7779 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10031) );
  MUX2_X1 U7780 ( .A(n8985), .B(n10031), .S(n4409), .Z(n6063) );
  INV_X1 U7781 ( .A(SI_26_), .ZN(n6062) );
  NAND2_X1 U7782 ( .A1(n6063), .A2(n6062), .ZN(n6543) );
  INV_X1 U7783 ( .A(n6063), .ZN(n6064) );
  NAND2_X1 U7784 ( .A1(n6064), .A2(SI_26_), .ZN(n6542) );
  AND2_X1 U7785 ( .A1(n6543), .A2(n6542), .ZN(n6065) );
  NAND2_X1 U7786 ( .A1(n8984), .A2(n6953), .ZN(n6068) );
  OR2_X1 U7787 ( .A1(n9220), .A2(n10031), .ZN(n6067) );
  NAND2_X1 U7788 ( .A1(n9866), .A2(n9041), .ZN(n6079) );
  INV_X1 U7789 ( .A(n6071), .ZN(n6069) );
  NAND2_X1 U7790 ( .A1(n6069), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6110) );
  INV_X1 U7791 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7792 ( .A1(n6071), .A2(n6070), .ZN(n6072) );
  NAND2_X1 U7793 ( .A1(n6110), .A2(n6072), .ZN(n9601) );
  INV_X1 U7794 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10373) );
  INV_X1 U7795 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n10339) );
  OR2_X1 U7796 ( .A1(n4408), .A2(n10339), .ZN(n6074) );
  INV_X1 U7797 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10336) );
  OR2_X1 U7798 ( .A1(n4406), .A2(n10336), .ZN(n6073) );
  OAI211_X1 U7799 ( .C1(n6989), .C2(n10373), .A(n6074), .B(n6073), .ZN(n6075)
         );
  INV_X1 U7800 ( .A(n6075), .ZN(n6076) );
  NAND2_X1 U7801 ( .A1(n4412), .A2(n5468), .ZN(n6078) );
  NAND2_X1 U7802 ( .A1(n6079), .A2(n6078), .ZN(n6080) );
  XNOR2_X1 U7803 ( .A(n6080), .B(n8327), .ZN(n8321) );
  AND2_X1 U7804 ( .A1(n4412), .A2(n9036), .ZN(n6081) );
  AOI21_X1 U7805 ( .B1(n9866), .B2(n5468), .A(n6081), .ZN(n8322) );
  XNOR2_X1 U7806 ( .A(n8321), .B(n8322), .ZN(n6084) );
  OAI21_X1 U7807 ( .B1(n6082), .B2(n6083), .A(n6084), .ZN(n6132) );
  NOR2_X1 U7808 ( .A1(n6084), .A2(n6083), .ZN(n6085) );
  NAND2_X1 U7809 ( .A1(n10036), .A2(P1_B_REG_SCAN_IN), .ZN(n6088) );
  MUX2_X1 U7810 ( .A(P1_B_REG_SCAN_IN), .B(n6088), .S(n10041), .Z(n6089) );
  INV_X1 U7811 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U7812 ( .A1(n7002), .A2(n6090), .ZN(n6092) );
  NAND2_X1 U7813 ( .A1(n10041), .A2(n10033), .ZN(n10020) );
  NOR4_X1 U7814 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n10327) );
  NOR2_X1 U7815 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .ZN(
        n6095) );
  NOR4_X1 U7816 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n6094) );
  NOR4_X1 U7817 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n6093) );
  AND4_X1 U7818 ( .A1(n10327), .A2(n6095), .A3(n6094), .A4(n6093), .ZN(n6101)
         );
  NOR4_X1 U7819 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6099) );
  NOR4_X1 U7820 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6098) );
  NOR4_X1 U7821 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n6097) );
  NOR4_X1 U7822 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6096) );
  AND4_X1 U7823 ( .A1(n6099), .A2(n6098), .A3(n6097), .A4(n6096), .ZN(n6100)
         );
  NAND2_X1 U7824 ( .A1(n6101), .A2(n6100), .ZN(n7001) );
  INV_X1 U7825 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10482) );
  NOR2_X1 U7826 ( .A1(n7001), .A2(n10482), .ZN(n7612) );
  NAND2_X1 U7827 ( .A1(n10036), .A2(n10033), .ZN(n10019) );
  OAI21_X1 U7828 ( .B1(n7611), .B2(n7612), .A(n10019), .ZN(n6102) );
  NAND2_X1 U7829 ( .A1(n6103), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6105) );
  INV_X1 U7830 ( .A(n7620), .ZN(n7619) );
  NOR2_X1 U7831 ( .A1(n10154), .A2(n9421), .ZN(n6107) );
  NAND2_X1 U7832 ( .A1(n9402), .A2(n8088), .ZN(n6108) );
  AOI21_X2 U7833 ( .B1(n6118), .B2(n7618), .A(n9836), .ZN(n9213) );
  INV_X1 U7834 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6109) );
  OR2_X2 U7835 ( .A1(n6110), .A2(n6109), .ZN(n6960) );
  NAND2_X1 U7836 ( .A1(n6110), .A2(n6109), .ZN(n6111) );
  NAND2_X1 U7837 ( .A1(n9588), .A2(n4405), .ZN(n6117) );
  INV_X1 U7838 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10523) );
  NAND2_X1 U7839 ( .A1(n6986), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U7840 ( .A1(n6112), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6113) );
  OAI211_X1 U7841 ( .C1(n4406), .C2(n10523), .A(n6114), .B(n6113), .ZN(n6115)
         );
  INV_X1 U7842 ( .A(n6115), .ZN(n6116) );
  AND2_X2 U7843 ( .A1(n6117), .A2(n6116), .ZN(n9609) );
  INV_X1 U7844 ( .A(n6118), .ZN(n6119) );
  INV_X1 U7845 ( .A(n6126), .ZN(n6121) );
  NAND2_X1 U7846 ( .A1(n6121), .A2(n6120), .ZN(n9207) );
  INV_X1 U7847 ( .A(n7618), .ZN(n6122) );
  NAND2_X1 U7848 ( .A1(n10154), .A2(n6122), .ZN(n7005) );
  NAND2_X1 U7849 ( .A1(n6123), .A2(n7005), .ZN(n6124) );
  NAND2_X1 U7850 ( .A1(n9335), .A2(n9421), .ZN(n7615) );
  NAND2_X1 U7851 ( .A1(n6124), .A2(n7615), .ZN(n7693) );
  OAI21_X1 U7852 ( .B1(n7693), .B2(n4810), .A(P1_STATE_REG_SCAN_IN), .ZN(n6125) );
  AOI22_X1 U7853 ( .A1(n9633), .A2(n9210), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        n4401), .ZN(n6127) );
  OAI21_X1 U7854 ( .B1(n9206), .B2(n9601), .A(n6127), .ZN(n6128) );
  AOI21_X1 U7855 ( .B1(n9476), .B2(n9192), .A(n6128), .ZN(n6129) );
  OAI21_X1 U7856 ( .B1(n9600), .B2(n9213), .A(n6129), .ZN(n6130) );
  INV_X1 U7857 ( .A(n6133), .ZN(P1_U3240) );
  NOR2_X1 U7858 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n6137) );
  NAND4_X1 U7859 ( .A1(n6137), .A2(n6136), .A3(n6280), .A4(n6353), .ZN(n6140)
         );
  NAND4_X1 U7860 ( .A1(n10317), .A2(n6395), .A3(n6394), .A4(n6138), .ZN(n6139)
         );
  NOR2_X1 U7861 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n6143) );
  NOR2_X1 U7862 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n6142) );
  NOR2_X1 U7863 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n6141) );
  NAND2_X1 U7864 ( .A1(n6144), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6145) );
  XNOR2_X1 U7865 ( .A(n8992), .B(P2_B_REG_SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7866 ( .A1(n6147), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7867 ( .A1(n6153), .A2(n8989), .ZN(n6157) );
  NAND2_X1 U7868 ( .A1(n8992), .A2(n8986), .ZN(n7352) );
  INV_X1 U7869 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6159) );
  INV_X1 U7870 ( .A(n6579), .ZN(n6163) );
  NAND2_X1 U7871 ( .A1(n6165), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6167) );
  XNOR2_X2 U7872 ( .A(n6170), .B(n6173), .ZN(n7247) );
  XNOR2_X1 U7873 ( .A(n6172), .B(P2_IR_REG_1__SCAN_IN), .ZN(n10179) );
  XNOR2_X2 U7874 ( .A(n6174), .B(P2_IR_REG_30__SCAN_IN), .ZN(n6176) );
  INV_X1 U7875 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10169) );
  INV_X1 U7876 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7877 ( .A1(n4416), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6177) );
  INV_X1 U7878 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6836) );
  INV_X1 U7879 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6179) );
  NAND2_X1 U7880 ( .A1(n4416), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6180) );
  XNOR2_X1 U7881 ( .A(n6184), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8993) );
  NAND2_X1 U7882 ( .A1(n7604), .A2(n6653), .ZN(n7598) );
  NAND2_X1 U7883 ( .A1(n6528), .A2(n7532), .ZN(n6186) );
  INV_X1 U7884 ( .A(n6188), .ZN(n6189) );
  NAND2_X1 U7885 ( .A1(n6189), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6191) );
  XNOR2_X2 U7886 ( .A(n6191), .B(n6190), .ZN(n7508) );
  OR2_X1 U7887 ( .A1(n6225), .A2(n7317), .ZN(n6193) );
  OR2_X1 U7888 ( .A1(n7071), .A2(n4721), .ZN(n6192) );
  NAND2_X1 U7889 ( .A1(n6270), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6199) );
  NAND2_X1 U7890 ( .A1(n4414), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6198) );
  INV_X1 U7891 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6195) );
  OR2_X1 U7892 ( .A1(n6208), .A2(n6195), .ZN(n6197) );
  INV_X1 U7893 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10441) );
  OR2_X1 U7894 ( .A1(n6374), .A2(n10441), .ZN(n6196) );
  XNOR2_X1 U7895 ( .A(n6200), .B(n7605), .ZN(n7448) );
  INV_X1 U7896 ( .A(n6200), .ZN(n6201) );
  NAND2_X1 U7897 ( .A1(n7605), .A2(n6201), .ZN(n6202) );
  NAND2_X1 U7898 ( .A1(n6223), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6205) );
  XNOR2_X1 U7899 ( .A(n6204), .B(n6205), .ZN(n7306) );
  OR2_X1 U7900 ( .A1(n6225), .A2(n7318), .ZN(n6207) );
  OR2_X1 U7901 ( .A1(n7071), .A2(n7307), .ZN(n6206) );
  XNOR2_X1 U7902 ( .A(n6194), .B(n7666), .ZN(n6213) );
  NAND2_X1 U7903 ( .A1(n6265), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U7904 ( .A1(n6270), .A2(n6217), .ZN(n6211) );
  NAND2_X1 U7905 ( .A1(n4415), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6210) );
  INV_X1 U7906 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7665) );
  INV_X1 U7907 ( .A(n6213), .ZN(n6214) );
  NAND2_X1 U7908 ( .A1(n6214), .A2(n8497), .ZN(n6215) );
  NAND2_X1 U7909 ( .A1(n6265), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6222) );
  INV_X1 U7910 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U7911 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6218) );
  NAND2_X1 U7912 ( .A1(n6240), .A2(n6218), .ZN(n7674) );
  NAND2_X1 U7913 ( .A1(n6270), .A2(n7674), .ZN(n6221) );
  NAND2_X1 U7914 ( .A1(n4415), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6220) );
  OR2_X1 U7915 ( .A1(n7058), .A2(n10450), .ZN(n6219) );
  NAND4_X1 U7916 ( .A1(n6222), .A2(n6221), .A3(n6220), .A4(n6219), .ZN(n8496)
         );
  INV_X1 U7917 ( .A(n8496), .ZN(n7725) );
  NAND2_X1 U7918 ( .A1(n6232), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6224) );
  INV_X2 U7919 ( .A(n6225), .ZN(n6278) );
  NAND2_X1 U7920 ( .A1(n6278), .A2(n7308), .ZN(n6227) );
  OR2_X1 U7921 ( .A1(n7071), .A2(n4860), .ZN(n6226) );
  XNOR2_X1 U7922 ( .A(n7258), .B(n7673), .ZN(n6228) );
  NAND2_X1 U7923 ( .A1(n7725), .A2(n6228), .ZN(n7717) );
  INV_X1 U7924 ( .A(n6228), .ZN(n6229) );
  NAND2_X1 U7925 ( .A1(n6229), .A2(n8496), .ZN(n6230) );
  NAND2_X1 U7926 ( .A1(n7717), .A2(n6230), .ZN(n7670) );
  INV_X1 U7927 ( .A(n7670), .ZN(n6231) );
  NAND2_X1 U7928 ( .A1(n7311), .A2(n6278), .ZN(n6237) );
  INV_X1 U7929 ( .A(n6232), .ZN(n6234) );
  NAND2_X1 U7930 ( .A1(n6234), .A2(n6233), .ZN(n6248) );
  NAND2_X1 U7931 ( .A1(n6248), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6235) );
  XNOR2_X1 U7932 ( .A(n6235), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6847) );
  AOI22_X1 U7933 ( .A1(n6441), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6847), .B2(
        n5222), .ZN(n6236) );
  NAND2_X1 U7934 ( .A1(n6237), .A2(n6236), .ZN(n7824) );
  XNOR2_X1 U7935 ( .A(n7824), .B(n7258), .ZN(n6246) );
  NAND2_X1 U7936 ( .A1(n6265), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U7937 ( .A1(n4414), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6244) );
  INV_X1 U7938 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6239) );
  NAND2_X1 U7939 ( .A1(n6240), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6241) );
  NAND2_X1 U7940 ( .A1(n6252), .A2(n6241), .ZN(n7823) );
  NAND2_X1 U7941 ( .A1(n6270), .A2(n7823), .ZN(n6243) );
  OR2_X1 U7942 ( .A1(n7058), .A2(n5164), .ZN(n6242) );
  XNOR2_X1 U7943 ( .A(n6246), .B(n8495), .ZN(n7718) );
  INV_X1 U7944 ( .A(n8495), .ZN(n7793) );
  NAND2_X1 U7945 ( .A1(n6246), .A2(n7793), .ZN(n6247) );
  NAND2_X1 U7946 ( .A1(n7309), .A2(n6278), .ZN(n6251) );
  NAND2_X1 U7947 ( .A1(n6261), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6249) );
  XNOR2_X1 U7948 ( .A(n6249), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6851) );
  AOI22_X1 U7949 ( .A1(n6441), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6851), .B2(
        n5222), .ZN(n6250) );
  NAND2_X1 U7950 ( .A1(n6251), .A2(n6250), .ZN(n8064) );
  XNOR2_X1 U7951 ( .A(n8064), .B(n7258), .ZN(n6258) );
  NAND2_X1 U7952 ( .A1(n6252), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U7953 ( .A1(n6268), .A2(n6253), .ZN(n7923) );
  NAND2_X1 U7954 ( .A1(n6270), .A2(n7923), .ZN(n6257) );
  INV_X1 U7955 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7922) );
  OR2_X1 U7956 ( .A1(n7058), .A2(n7922), .ZN(n6256) );
  NAND2_X1 U7957 ( .A1(n6265), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U7958 ( .A1(n4414), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6254) );
  XNOR2_X1 U7959 ( .A(n6258), .B(n8494), .ZN(n7791) );
  INV_X1 U7960 ( .A(n6258), .ZN(n6259) );
  NAND2_X1 U7961 ( .A1(n6259), .A2(n8494), .ZN(n6260) );
  NAND2_X1 U7962 ( .A1(n7326), .A2(n6278), .ZN(n6264) );
  OAI21_X1 U7963 ( .B1(n6261), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6262) );
  XNOR2_X1 U7964 ( .A(n6262), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6855) );
  AOI22_X1 U7965 ( .A1(n6441), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6855), .B2(
        n5222), .ZN(n6263) );
  XNOR2_X1 U7966 ( .A(n7957), .B(n7258), .ZN(n6275) );
  NAND2_X1 U7967 ( .A1(n6265), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6274) );
  NAND2_X1 U7968 ( .A1(n4415), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6273) );
  INV_X1 U7969 ( .A(n6268), .ZN(n6267) );
  NAND2_X1 U7970 ( .A1(n6268), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U7971 ( .A1(n6317), .A2(n6269), .ZN(n8032) );
  NAND2_X1 U7972 ( .A1(n6270), .A2(n8032), .ZN(n6272) );
  INV_X1 U7973 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7649) );
  OR2_X1 U7974 ( .A1(n7058), .A2(n7649), .ZN(n6271) );
  NAND4_X1 U7975 ( .A1(n6274), .A2(n6273), .A3(n6272), .A4(n6271), .ZN(n8493)
         );
  XNOR2_X1 U7976 ( .A(n6275), .B(n8493), .ZN(n7929) );
  INV_X1 U7977 ( .A(n6275), .ZN(n6276) );
  NAND2_X1 U7978 ( .A1(n6276), .A2(n7792), .ZN(n6277) );
  NAND2_X1 U7979 ( .A1(n7392), .A2(n6278), .ZN(n6283) );
  NAND2_X1 U7980 ( .A1(n6279), .A2(n10317), .ZN(n6301) );
  INV_X1 U7981 ( .A(n6291), .ZN(n6281) );
  NAND2_X1 U7982 ( .A1(n6281), .A2(n6280), .ZN(n6391) );
  NAND2_X1 U7983 ( .A1(n6391), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6355) );
  XNOR2_X1 U7984 ( .A(n6355), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8507) );
  AOI22_X1 U7985 ( .A1(n6441), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8507), .B2(
        n5222), .ZN(n6282) );
  NAND2_X1 U7986 ( .A1(n6604), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6290) );
  NAND2_X1 U7987 ( .A1(n6296), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U7988 ( .A1(n6345), .A2(n6285), .ZN(n8446) );
  NAND2_X1 U7989 ( .A1(n6270), .A2(n8446), .ZN(n6289) );
  INV_X1 U7990 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n6286) );
  OR2_X1 U7991 ( .A1(n6208), .A2(n6286), .ZN(n6288) );
  INV_X1 U7992 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8503) );
  OR2_X1 U7993 ( .A1(n7058), .A2(n8503), .ZN(n6287) );
  NAND2_X1 U7994 ( .A1(n8447), .A2(n8357), .ZN(n7166) );
  XNOR2_X1 U7995 ( .A(n8234), .B(n7258), .ZN(n8440) );
  NAND2_X1 U7996 ( .A1(n7343), .A2(n6278), .ZN(n6294) );
  NAND2_X1 U7997 ( .A1(n6291), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6292) );
  XNOR2_X1 U7998 ( .A(n6292), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6867) );
  AOI22_X1 U7999 ( .A1(n6441), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6867), .B2(
        n5222), .ZN(n6293) );
  XNOR2_X1 U8000 ( .A(n8360), .B(n6528), .ZN(n8437) );
  NAND2_X1 U8001 ( .A1(n6265), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6300) );
  NAND2_X1 U8002 ( .A1(n4415), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6299) );
  NAND2_X1 U8003 ( .A1(n6306), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6295) );
  NAND2_X1 U8004 ( .A1(n6296), .A2(n6295), .ZN(n8359) );
  NAND2_X1 U8005 ( .A1(n6270), .A2(n8359), .ZN(n6298) );
  INV_X1 U8006 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6806) );
  OR2_X1 U8007 ( .A1(n6374), .A2(n6806), .ZN(n6297) );
  NAND4_X1 U8008 ( .A1(n6300), .A2(n6299), .A3(n6298), .A4(n6297), .ZN(n8490)
         );
  NAND2_X1 U8009 ( .A1(n7338), .A2(n6278), .ZN(n6304) );
  NAND2_X1 U8010 ( .A1(n6301), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6302) );
  XNOR2_X1 U8011 ( .A(n6302), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6863) );
  AOI22_X1 U8012 ( .A1(n6441), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6863), .B2(
        n5222), .ZN(n6303) );
  XNOR2_X1 U8013 ( .A(n8257), .B(n6528), .ZN(n6326) );
  NAND2_X1 U8014 ( .A1(n4414), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6311) );
  NAND2_X1 U8015 ( .A1(n6319), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6305) );
  NAND2_X1 U8016 ( .A1(n6306), .A2(n6305), .ZN(n8256) );
  NAND2_X1 U8017 ( .A1(n6270), .A2(n8256), .ZN(n6310) );
  INV_X1 U8018 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n6307) );
  OR2_X1 U8019 ( .A1(n6208), .A2(n6307), .ZN(n6309) );
  INV_X1 U8020 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7999) );
  OR2_X1 U8021 ( .A1(n6374), .A2(n7999), .ZN(n6308) );
  AND2_X1 U8022 ( .A1(n6326), .A2(n8491), .ZN(n8348) );
  AOI21_X1 U8023 ( .B1(n8437), .B2(n8490), .A(n8348), .ZN(n6312) );
  NAND2_X1 U8024 ( .A1(n7330), .A2(n6278), .ZN(n6316) );
  INV_X1 U8025 ( .A(n6279), .ZN(n6313) );
  NAND2_X1 U8026 ( .A1(n6313), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6314) );
  AOI22_X1 U8027 ( .A1(n6441), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7333), .B2(
        n5222), .ZN(n6315) );
  NAND2_X1 U8028 ( .A1(n6316), .A2(n6315), .ZN(n8269) );
  XNOR2_X1 U8029 ( .A(n8269), .B(n7258), .ZN(n8212) );
  NAND2_X1 U8030 ( .A1(n6265), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6323) );
  NAND2_X1 U8031 ( .A1(n4415), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6322) );
  NAND2_X1 U8032 ( .A1(n6317), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6318) );
  NAND2_X1 U8033 ( .A1(n6319), .A2(n6318), .ZN(n8268) );
  NAND2_X1 U8034 ( .A1(n6270), .A2(n8268), .ZN(n6321) );
  INV_X1 U8035 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6801) );
  OR2_X1 U8036 ( .A1(n6374), .A2(n6801), .ZN(n6320) );
  NAND2_X1 U8037 ( .A1(n8213), .A2(n6325), .ZN(n6338) );
  INV_X1 U8038 ( .A(n6326), .ZN(n6327) );
  XNOR2_X1 U8039 ( .A(n6327), .B(n8180), .ZN(n8216) );
  AOI21_X1 U8040 ( .B1(n8142), .B2(n8212), .A(n8216), .ZN(n6328) );
  INV_X1 U8041 ( .A(n6328), .ZN(n6335) );
  INV_X1 U8042 ( .A(n8490), .ZN(n8351) );
  NAND2_X1 U8043 ( .A1(n8351), .A2(n6528), .ZN(n6329) );
  OAI22_X1 U8044 ( .A1(n8360), .A2(n6329), .B1(n6528), .B2(n4718), .ZN(n6332)
         );
  NAND3_X1 U8045 ( .A1(n8360), .A2(n8351), .A3(n7258), .ZN(n6330) );
  OAI211_X1 U8046 ( .C1(n4718), .C2(n7258), .A(n8234), .B(n6330), .ZN(n6331)
         );
  OAI21_X1 U8047 ( .B1(n8234), .B2(n6332), .A(n6331), .ZN(n6333) );
  INV_X1 U8048 ( .A(n6333), .ZN(n6334) );
  NAND2_X1 U8049 ( .A1(n7437), .A2(n6278), .ZN(n6342) );
  NAND2_X1 U8050 ( .A1(n6355), .A2(n6353), .ZN(n6339) );
  NAND2_X1 U8051 ( .A1(n6339), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6340) );
  AOI22_X1 U8052 ( .A1(n6441), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6876), .B2(
        n5222), .ZN(n6341) );
  XNOR2_X1 U8053 ( .A(n8893), .B(n6528), .ZN(n6351) );
  NAND2_X1 U8054 ( .A1(n6265), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6350) );
  NAND2_X1 U8055 ( .A1(n6604), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6349) );
  NAND2_X1 U8056 ( .A1(n6345), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6346) );
  NAND2_X1 U8057 ( .A1(n6358), .A2(n6346), .ZN(n8120) );
  NAND2_X1 U8058 ( .A1(n6270), .A2(n8120), .ZN(n6348) );
  INV_X1 U8059 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8831) );
  OR2_X1 U8060 ( .A1(n7058), .A2(n8831), .ZN(n6347) );
  NAND4_X1 U8061 ( .A1(n6350), .A2(n6349), .A3(n6348), .A4(n6347), .ZN(n8815)
         );
  NAND2_X1 U8062 ( .A1(n6351), .A2(n8815), .ZN(n8117) );
  NAND2_X1 U8063 ( .A1(n7472), .A2(n6278), .ZN(n6357) );
  INV_X1 U8064 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6352) );
  NAND2_X1 U8065 ( .A1(n6353), .A2(n6352), .ZN(n6392) );
  NAND2_X1 U8066 ( .A1(n6392), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6354) );
  NAND2_X1 U8067 ( .A1(n6355), .A2(n6354), .ZN(n6366) );
  XNOR2_X1 U8068 ( .A(n6366), .B(n6394), .ZN(n6881) );
  AOI22_X1 U8069 ( .A1(n6441), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5222), .B2(
        n6881), .ZN(n6356) );
  XNOR2_X1 U8070 ( .A(n8964), .B(n7258), .ZN(n6364) );
  NAND2_X1 U8071 ( .A1(n6604), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6363) );
  NAND2_X1 U8072 ( .A1(n6265), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6362) );
  NAND2_X1 U8073 ( .A1(n6358), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6359) );
  NAND2_X1 U8074 ( .A1(n6372), .A2(n6359), .ZN(n8820) );
  NAND2_X1 U8075 ( .A1(n6270), .A2(n8820), .ZN(n6361) );
  INV_X1 U8076 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10468) );
  OR2_X1 U8077 ( .A1(n7058), .A2(n10468), .ZN(n6360) );
  NAND4_X1 U8078 ( .A1(n6363), .A2(n6362), .A3(n6361), .A4(n6360), .ZN(n8827)
         );
  XNOR2_X1 U8079 ( .A(n6364), .B(n8827), .ZN(n8168) );
  INV_X1 U8080 ( .A(n8827), .ZN(n6642) );
  NAND2_X1 U8081 ( .A1(n7439), .A2(n6278), .ZN(n6371) );
  NAND2_X1 U8082 ( .A1(n6367), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6368) );
  OR2_X1 U8083 ( .A1(n6368), .A2(n6393), .ZN(n6369) );
  NAND2_X1 U8084 ( .A1(n6368), .A2(n6393), .ZN(n6380) );
  AOI22_X1 U8085 ( .A1(n6441), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6886), .B2(
        n5222), .ZN(n6370) );
  NAND2_X1 U8086 ( .A1(n6371), .A2(n6370), .ZN(n8247) );
  XNOR2_X1 U8087 ( .A(n8247), .B(n7258), .ZN(n6379) );
  NAND2_X1 U8088 ( .A1(n6265), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6378) );
  NAND2_X1 U8089 ( .A1(n6372), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U8090 ( .A1(n6383), .A2(n6373), .ZN(n8801) );
  NAND2_X1 U8091 ( .A1(n6270), .A2(n8801), .ZN(n6377) );
  NAND2_X1 U8092 ( .A1(n6604), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6376) );
  INV_X1 U8093 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6812) );
  OR2_X1 U8094 ( .A1(n6374), .A2(n6812), .ZN(n6375) );
  NAND4_X1 U8095 ( .A1(n6378), .A2(n6377), .A3(n6376), .A4(n6375), .ZN(n8816)
         );
  XNOR2_X1 U8096 ( .A(n6379), .B(n8475), .ZN(n8245) );
  NAND2_X1 U8097 ( .A1(n6380), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6381) );
  XNOR2_X1 U8098 ( .A(n6381), .B(P2_IR_REG_15__SCAN_IN), .ZN(n6891) );
  AOI22_X1 U8099 ( .A1(n6891), .A2(n5222), .B1(n6441), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6382) );
  XNOR2_X1 U8100 ( .A(n8952), .B(n7258), .ZN(n6389) );
  INV_X1 U8101 ( .A(n6407), .ZN(n6408) );
  NAND2_X1 U8102 ( .A1(n6383), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6384) );
  NAND2_X1 U8103 ( .A1(n6408), .A2(n6384), .ZN(n8792) );
  NAND2_X1 U8104 ( .A1(n8792), .A2(n6270), .ZN(n6388) );
  NAND2_X1 U8105 ( .A1(n6604), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6387) );
  NAND2_X1 U8106 ( .A1(n6265), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6386) );
  INV_X1 U8107 ( .A(n7058), .ZN(n6766) );
  NAND2_X1 U8108 ( .A1(n6766), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6385) );
  NAND4_X1 U8109 ( .A1(n6388), .A2(n6387), .A3(n6386), .A4(n6385), .ZN(n8797)
         );
  XNOR2_X1 U8110 ( .A(n6389), .B(n8797), .ZN(n8472) );
  NAND2_X1 U8111 ( .A1(n7553), .A2(n6278), .ZN(n6405) );
  INV_X1 U8112 ( .A(n6391), .ZN(n6398) );
  INV_X1 U8113 ( .A(n6392), .ZN(n6396) );
  AND4_X1 U8114 ( .A1(n6396), .A2(n6395), .A3(n6394), .A4(n6393), .ZN(n6397)
         );
  INV_X1 U8115 ( .A(n6402), .ZN(n6399) );
  NAND2_X1 U8116 ( .A1(n6399), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6400) );
  MUX2_X1 U8117 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6400), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n6403) );
  INV_X1 U8118 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6401) );
  NAND2_X1 U8119 ( .A1(n6402), .A2(n6401), .ZN(n6416) );
  NAND2_X1 U8120 ( .A1(n6403), .A2(n6416), .ZN(n8578) );
  AOI22_X1 U8121 ( .A1(n6441), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6895), .B2(
        n5222), .ZN(n6404) );
  NAND2_X1 U8122 ( .A1(n6405), .A2(n6404), .ZN(n8779) );
  XNOR2_X1 U8123 ( .A(n8779), .B(n7258), .ZN(n6414) );
  INV_X1 U8124 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n6816) );
  INV_X1 U8125 ( .A(n6420), .ZN(n6421) );
  NAND2_X1 U8126 ( .A1(n6408), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6409) );
  NAND2_X1 U8127 ( .A1(n6421), .A2(n6409), .ZN(n8778) );
  NAND2_X1 U8128 ( .A1(n8778), .A2(n6270), .ZN(n6413) );
  NAND2_X1 U8129 ( .A1(n6604), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6411) );
  NAND2_X1 U8130 ( .A1(n6265), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6410) );
  AND2_X1 U8131 ( .A1(n6411), .A2(n6410), .ZN(n6412) );
  XNOR2_X1 U8132 ( .A(n6414), .B(n8789), .ZN(n8391) );
  INV_X1 U8133 ( .A(n8789), .ZN(n8402) );
  NAND2_X1 U8134 ( .A1(n6416), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6417) );
  XNOR2_X1 U8135 ( .A(n6417), .B(P2_IR_REG_17__SCAN_IN), .ZN(n6899) );
  AOI22_X1 U8136 ( .A1(n6441), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6899), .B2(
        n5222), .ZN(n6418) );
  XNOR2_X1 U8137 ( .A(n8941), .B(n6528), .ZN(n8397) );
  NAND2_X1 U8138 ( .A1(n6421), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6422) );
  NAND2_X1 U8139 ( .A1(n6432), .A2(n6422), .ZN(n8764) );
  NAND2_X1 U8140 ( .A1(n8764), .A2(n6270), .ZN(n6425) );
  AOI22_X1 U8141 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n6604), .B1(n6265), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n6424) );
  NAND2_X1 U8142 ( .A1(n6766), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6423) );
  INV_X1 U8143 ( .A(n8772), .ZN(n8489) );
  INV_X1 U8144 ( .A(n8397), .ZN(n6427) );
  NAND2_X1 U8145 ( .A1(n7741), .A2(n6278), .ZN(n6431) );
  NAND2_X1 U8146 ( .A1(n6149), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6429) );
  XNOR2_X1 U8147 ( .A(n6429), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8610) );
  AOI22_X1 U8148 ( .A1(n6441), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8610), .B2(
        n5222), .ZN(n6430) );
  XNOR2_X1 U8149 ( .A(n8938), .B(n7258), .ZN(n6440) );
  NAND2_X1 U8150 ( .A1(n6432), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6433) );
  NAND2_X1 U8151 ( .A1(n6446), .A2(n6433), .ZN(n8745) );
  NAND2_X1 U8152 ( .A1(n8745), .A2(n6270), .ZN(n6439) );
  INV_X1 U8153 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n6436) );
  NAND2_X1 U8154 ( .A1(n6766), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6435) );
  NAND2_X1 U8155 ( .A1(n6265), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6434) );
  OAI211_X1 U8156 ( .C1(n6769), .C2(n6436), .A(n6435), .B(n6434), .ZN(n6437)
         );
  INV_X1 U8157 ( .A(n6437), .ZN(n6438) );
  XNOR2_X1 U8158 ( .A(n6440), .B(n8732), .ZN(n8453) );
  NAND2_X1 U8159 ( .A1(n7856), .A2(n6278), .ZN(n6443) );
  AOI22_X1 U8160 ( .A1(n6441), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7080), .B2(
        n5222), .ZN(n6442) );
  XNOR2_X1 U8161 ( .A(n8933), .B(n7258), .ZN(n6463) );
  NAND2_X1 U8162 ( .A1(n6446), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6447) );
  NAND2_X1 U8163 ( .A1(n6455), .A2(n6447), .ZN(n8738) );
  INV_X1 U8164 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8869) );
  NAND2_X1 U8165 ( .A1(n6265), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6449) );
  NAND2_X1 U8166 ( .A1(n6766), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6448) );
  OAI211_X1 U8167 ( .C1(n6769), .C2(n8869), .A(n6449), .B(n6448), .ZN(n6450)
         );
  XNOR2_X1 U8168 ( .A(n6463), .B(n8722), .ZN(n8364) );
  NAND2_X1 U8169 ( .A1(n6451), .A2(n6278), .ZN(n6454) );
  OR2_X1 U8170 ( .A1(n7071), .A2(n6452), .ZN(n6453) );
  XNOR2_X1 U8171 ( .A(n8927), .B(n6528), .ZN(n6462) );
  NAND2_X1 U8172 ( .A1(n6455), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6456) );
  NAND2_X1 U8173 ( .A1(n6467), .A2(n6456), .ZN(n8726) );
  NAND2_X1 U8174 ( .A1(n8726), .A2(n6270), .ZN(n6461) );
  INV_X1 U8175 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8725) );
  NAND2_X1 U8176 ( .A1(n6604), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U8177 ( .A1(n6265), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6457) );
  OAI211_X1 U8178 ( .C1(n8725), .C2(n7058), .A(n6458), .B(n6457), .ZN(n6459)
         );
  INV_X1 U8179 ( .A(n6459), .ZN(n6460) );
  NOR2_X1 U8180 ( .A1(n6462), .A2(n8488), .ZN(n8372) );
  AOI21_X1 U8181 ( .B1(n6462), .B2(n8488), .A(n8372), .ZN(n8416) );
  INV_X1 U8182 ( .A(n6463), .ZN(n6464) );
  NAND2_X1 U8183 ( .A1(n6464), .A2(n8722), .ZN(n8417) );
  NAND2_X1 U8184 ( .A1(n8080), .A2(n6278), .ZN(n6466) );
  OR2_X1 U8185 ( .A1(n7071), .A2(n8081), .ZN(n6465) );
  XNOR2_X1 U8186 ( .A(n8863), .B(n7258), .ZN(n6473) );
  NAND2_X1 U8187 ( .A1(n6467), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6468) );
  NAND2_X1 U8188 ( .A1(n6477), .A2(n6468), .ZN(n8709) );
  INV_X1 U8189 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n6471) );
  NAND2_X1 U8190 ( .A1(n6604), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6470) );
  NAND2_X1 U8191 ( .A1(n6265), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6469) );
  OAI211_X1 U8192 ( .C1(n6471), .C2(n7058), .A(n6470), .B(n6469), .ZN(n6472)
         );
  AOI21_X1 U8193 ( .B1(n8709), .B2(n6270), .A(n6472), .ZN(n6644) );
  XNOR2_X1 U8194 ( .A(n6473), .B(n8723), .ZN(n8371) );
  NAND2_X1 U8195 ( .A1(n6473), .A2(n6644), .ZN(n6474) );
  NAND2_X1 U8196 ( .A1(n8083), .A2(n6278), .ZN(n6476) );
  OR2_X1 U8197 ( .A1(n7071), .A2(n8087), .ZN(n6475) );
  XNOR2_X1 U8198 ( .A(n8700), .B(n7258), .ZN(n6485) );
  NAND2_X1 U8199 ( .A1(n6477), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6478) );
  NAND2_X1 U8200 ( .A1(n6494), .A2(n6478), .ZN(n8429) );
  NAND2_X1 U8201 ( .A1(n8429), .A2(n6270), .ZN(n6483) );
  INV_X1 U8202 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8697) );
  NAND2_X1 U8203 ( .A1(n6265), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6480) );
  NAND2_X1 U8204 ( .A1(n6604), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6479) );
  OAI211_X1 U8205 ( .C1(n7058), .C2(n8697), .A(n6480), .B(n6479), .ZN(n6481)
         );
  INV_X1 U8206 ( .A(n6481), .ZN(n6482) );
  XNOR2_X1 U8207 ( .A(n6485), .B(n8708), .ZN(n8425) );
  OR2_X1 U8208 ( .A1(n7071), .A2(n8163), .ZN(n6490) );
  AND2_X1 U8209 ( .A1(n6487), .A2(n6490), .ZN(n6488) );
  NAND2_X1 U8210 ( .A1(n6489), .A2(n6488), .ZN(n6493) );
  INV_X1 U8211 ( .A(n6490), .ZN(n6491) );
  OR2_X1 U8212 ( .A1(n6491), .A2(n6278), .ZN(n6492) );
  XNOR2_X1 U8213 ( .A(n8313), .B(n6528), .ZN(n8297) );
  NAND2_X1 U8214 ( .A1(n6494), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6495) );
  NAND2_X1 U8215 ( .A1(n6505), .A2(n6495), .ZN(n8302) );
  NAND2_X1 U8216 ( .A1(n8302), .A2(n6270), .ZN(n6500) );
  INV_X1 U8217 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8294) );
  NAND2_X1 U8218 ( .A1(n6604), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6497) );
  NAND2_X1 U8219 ( .A1(n6265), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6496) );
  OAI211_X1 U8220 ( .C1(n8294), .C2(n7058), .A(n6497), .B(n6496), .ZN(n6498)
         );
  INV_X1 U8221 ( .A(n6498), .ZN(n6499) );
  OR2_X1 U8222 ( .A1(n7071), .A2(n10520), .ZN(n6502) );
  XNOR2_X1 U8223 ( .A(n6650), .B(n7258), .ZN(n6513) );
  NAND2_X1 U8224 ( .A1(n6505), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6506) );
  NAND2_X1 U8225 ( .A1(n6517), .A2(n6506), .ZN(n8683) );
  NAND2_X1 U8226 ( .A1(n8683), .A2(n6270), .ZN(n6512) );
  INV_X1 U8227 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6509) );
  NAND2_X1 U8228 ( .A1(n6604), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6508) );
  NAND2_X1 U8229 ( .A1(n6265), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6507) );
  OAI211_X1 U8230 ( .C1(n6509), .C2(n7058), .A(n6508), .B(n6507), .ZN(n6510)
         );
  INV_X1 U8231 ( .A(n6510), .ZN(n6511) );
  OAI21_X1 U8232 ( .B1(n6513), .B2(n8386), .A(n8380), .ZN(n8406) );
  AOI21_X1 U8233 ( .B1(n8297), .B2(n8695), .A(n8406), .ZN(n6514) );
  NAND2_X1 U8234 ( .A1(n8987), .A2(n6278), .ZN(n6516) );
  OR2_X1 U8235 ( .A1(n7071), .A2(n8988), .ZN(n6515) );
  XNOR2_X1 U8236 ( .A(n8912), .B(n7258), .ZN(n6524) );
  NAND2_X1 U8237 ( .A1(n6517), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6518) );
  NAND2_X1 U8238 ( .A1(n6529), .A2(n6518), .ZN(n8673) );
  NAND2_X1 U8239 ( .A1(n8673), .A2(n6270), .ZN(n6523) );
  INV_X1 U8240 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n10529) );
  NAND2_X1 U8241 ( .A1(n6604), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6520) );
  NAND2_X1 U8242 ( .A1(n6265), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6519) );
  OAI211_X1 U8243 ( .C1(n10529), .C2(n7058), .A(n6520), .B(n6519), .ZN(n6521)
         );
  INV_X1 U8244 ( .A(n6521), .ZN(n6522) );
  XNOR2_X1 U8245 ( .A(n6524), .B(n8486), .ZN(n8381) );
  NAND2_X1 U8246 ( .A1(n6524), .A2(n8680), .ZN(n6525) );
  NAND2_X1 U8247 ( .A1(n8984), .A2(n6278), .ZN(n6527) );
  OR2_X1 U8248 ( .A1(n7071), .A2(n8985), .ZN(n6526) );
  NAND2_X1 U8249 ( .A1(n6529), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6530) );
  NAND2_X1 U8250 ( .A1(n6558), .A2(n6530), .ZN(n8662) );
  NAND2_X1 U8251 ( .A1(n8662), .A2(n6270), .ZN(n6536) );
  INV_X1 U8252 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n6533) );
  NAND2_X1 U8253 ( .A1(n6604), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6532) );
  NAND2_X1 U8254 ( .A1(n6265), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6531) );
  OAI211_X1 U8255 ( .C1(n6533), .C2(n7058), .A(n6532), .B(n6531), .ZN(n6534)
         );
  INV_X1 U8256 ( .A(n6534), .ZN(n6535) );
  INV_X1 U8257 ( .A(n6537), .ZN(n6538) );
  NAND2_X1 U8258 ( .A1(n6539), .A2(n6538), .ZN(n6593) );
  NAND2_X1 U8259 ( .A1(n8463), .A2(n6593), .ZN(n6564) );
  AND2_X1 U8260 ( .A1(n6540), .A2(n6542), .ZN(n6736) );
  NAND2_X1 U8261 ( .A1(n6541), .A2(n6736), .ZN(n6547) );
  INV_X1 U8262 ( .A(n6542), .ZN(n6546) );
  AND2_X1 U8263 ( .A1(n6544), .A2(n6543), .ZN(n6545) );
  NAND2_X1 U8264 ( .A1(n6547), .A2(n6729), .ZN(n6552) );
  INV_X1 U8265 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6553) );
  MUX2_X1 U8266 ( .A(n6553), .B(n10030), .S(n4403), .Z(n6549) );
  INV_X1 U8267 ( .A(SI_27_), .ZN(n6548) );
  NAND2_X1 U8268 ( .A1(n6549), .A2(n6548), .ZN(n6733) );
  INV_X1 U8269 ( .A(n6549), .ZN(n6550) );
  NAND2_X1 U8270 ( .A1(n6550), .A2(SI_27_), .ZN(n6551) );
  NAND2_X1 U8271 ( .A1(n6733), .A2(n6551), .ZN(n6730) );
  INV_X1 U8272 ( .A(n6730), .ZN(n6735) );
  NAND2_X1 U8273 ( .A1(n8980), .A2(n6278), .ZN(n6555) );
  OR2_X1 U8274 ( .A1(n7071), .A2(n6553), .ZN(n6554) );
  XNOR2_X1 U8275 ( .A(n6725), .B(n7258), .ZN(n7267) );
  INV_X1 U8276 ( .A(n6558), .ZN(n6557) );
  INV_X1 U8277 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U8278 ( .A1(n6558), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6559) );
  NAND2_X1 U8279 ( .A1(n6602), .A2(n6559), .ZN(n8651) );
  INV_X1 U8280 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n10539) );
  NAND2_X1 U8281 ( .A1(n6766), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6561) );
  NAND2_X1 U8282 ( .A1(n6265), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6560) );
  OAI211_X1 U8283 ( .C1(n6769), .C2(n10539), .A(n6561), .B(n6560), .ZN(n6562)
         );
  INV_X1 U8284 ( .A(n6562), .ZN(n6563) );
  NAND2_X1 U8285 ( .A1(n6564), .A2(n6591), .ZN(n6595) );
  NOR2_X1 U8286 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .ZN(
        n10328) );
  NOR4_X1 U8287 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6569) );
  NOR4_X1 U8288 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6568) );
  NOR4_X1 U8289 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n6567) );
  NAND4_X1 U8290 ( .A1(n10328), .A2(n6569), .A3(n6568), .A4(n6567), .ZN(n6576)
         );
  NOR4_X1 U8291 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n6573) );
  NOR4_X1 U8292 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6572) );
  NOR4_X1 U8293 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n6571) );
  NOR4_X1 U8294 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6570) );
  NAND4_X1 U8295 ( .A1(n6573), .A2(n6572), .A3(n6571), .A4(n6570), .ZN(n6575)
         );
  INV_X1 U8296 ( .A(n6565), .ZN(n6574) );
  INV_X1 U8297 ( .A(n6700), .ZN(n6577) );
  NOR2_X1 U8298 ( .A1(n6702), .A2(n6577), .ZN(n6617) );
  NOR2_X1 U8299 ( .A1(n8992), .A2(n8986), .ZN(n6582) );
  NAND2_X1 U8300 ( .A1(n6617), .A2(n7332), .ZN(n6716) );
  AND2_X1 U8301 ( .A1(n7217), .A2(n10242), .ZN(n6588) );
  NAND2_X1 U8302 ( .A1(n7250), .A2(n7080), .ZN(n6694) );
  NAND2_X1 U8303 ( .A1(n6588), .A2(n6714), .ZN(n6612) );
  OR2_X1 U8304 ( .A1(n6716), .A2(n6612), .ZN(n6590) );
  NAND3_X1 U8305 ( .A1(n7522), .A2(n6705), .A3(n6700), .ZN(n6620) );
  INV_X1 U8306 ( .A(n6714), .ZN(n6615) );
  NAND2_X1 U8307 ( .A1(n6718), .A2(n6615), .ZN(n6589) );
  INV_X1 U8308 ( .A(n6591), .ZN(n6592) );
  AND2_X1 U8309 ( .A1(n6593), .A2(n6592), .ZN(n6594) );
  NAND3_X1 U8310 ( .A1(n6595), .A2(n8470), .A3(n7274), .ZN(n6630) );
  OR2_X1 U8311 ( .A1(n6716), .A2(n10242), .ZN(n6597) );
  NAND2_X1 U8312 ( .A1(n7936), .A2(n7080), .ZN(n7245) );
  INV_X1 U8313 ( .A(n7517), .ZN(n6621) );
  AND2_X1 U8314 ( .A1(n6718), .A2(n6621), .ZN(n6611) );
  INV_X1 U8315 ( .A(n6611), .ZN(n6601) );
  INV_X1 U8316 ( .A(n7247), .ZN(n6599) );
  INV_X1 U8317 ( .A(n6910), .ZN(n7248) );
  NAND2_X1 U8318 ( .A1(n6599), .A2(n7248), .ZN(n6600) );
  INV_X1 U8319 ( .A(n6695), .ZN(n6610) );
  NAND2_X1 U8320 ( .A1(n6602), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6603) );
  NAND2_X1 U8321 ( .A1(n8624), .A2(n6603), .ZN(n8645) );
  NAND2_X1 U8322 ( .A1(n8645), .A2(n6270), .ZN(n6609) );
  INV_X1 U8323 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n10303) );
  NAND2_X1 U8324 ( .A1(n6265), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6606) );
  NAND2_X1 U8325 ( .A1(n6604), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6605) );
  OAI211_X1 U8326 ( .C1(n10303), .C2(n7058), .A(n6606), .B(n6605), .ZN(n6607)
         );
  INV_X1 U8327 ( .A(n6607), .ZN(n6608) );
  INV_X1 U8328 ( .A(n7245), .ZN(n7595) );
  NAND2_X1 U8329 ( .A1(n6612), .A2(n10206), .ZN(n6717) );
  INV_X1 U8330 ( .A(n6717), .ZN(n6618) );
  AND2_X1 U8331 ( .A1(n7353), .A2(n6912), .ZN(n6614) );
  NAND2_X1 U8332 ( .A1(n6620), .A2(n6615), .ZN(n6616) );
  OAI211_X1 U8333 ( .C1(n6618), .C2(n6617), .A(n6701), .B(n6616), .ZN(n6619)
         );
  NAND2_X1 U8334 ( .A1(n6619), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6624) );
  INV_X1 U8335 ( .A(n6620), .ZN(n6622) );
  NAND2_X1 U8336 ( .A1(n6621), .A2(n7332), .ZN(n7249) );
  OR2_X1 U8337 ( .A1(n6622), .A2(n7249), .ZN(n6623) );
  AOI22_X1 U8338 ( .A1(n8651), .A2(n8478), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n6625) );
  OAI21_X1 U8339 ( .B1(n8465), .B2(n8476), .A(n6625), .ZN(n6626) );
  AOI21_X1 U8340 ( .B1(n8473), .B2(n8484), .A(n6626), .ZN(n6627) );
  OAI21_X1 U8341 ( .B1(n6726), .B2(n8481), .A(n6627), .ZN(n6628) );
  NAND2_X1 U8342 ( .A1(n6630), .A2(n6629), .ZN(P2_U3154) );
  NAND2_X1 U8343 ( .A1(n7250), .A2(n7857), .ZN(n6703) );
  NAND2_X1 U8344 ( .A1(n6703), .A2(n6631), .ZN(n6632) );
  NAND3_X1 U8345 ( .A1(n7517), .A2(n10242), .A3(n6632), .ZN(n8177) );
  INV_X1 U8346 ( .A(n7598), .ZN(n6634) );
  INV_X1 U8347 ( .A(n7605), .ZN(n8498) );
  NAND2_X1 U8348 ( .A1(n7605), .A2(n7450), .ZN(n7133) );
  INV_X1 U8349 ( .A(n7127), .ZN(n10210) );
  INV_X1 U8350 ( .A(n7666), .ZN(n10231) );
  NAND2_X1 U8351 ( .A1(n8497), .A2(n10231), .ZN(n7142) );
  INV_X1 U8352 ( .A(n7673), .ZN(n10235) );
  NAND2_X1 U8353 ( .A1(n7725), .A2(n7673), .ZN(n7145) );
  INV_X1 U8354 ( .A(n7819), .ZN(n6635) );
  NOR2_X1 U8355 ( .A1(n8495), .A2(n10243), .ZN(n7915) );
  INV_X1 U8356 ( .A(n8494), .ZN(n7724) );
  NAND2_X1 U8357 ( .A1(n7724), .A2(n8064), .ZN(n7141) );
  INV_X1 U8358 ( .A(n7141), .ZN(n7147) );
  NAND2_X1 U8359 ( .A1(n7957), .A2(n8493), .ZN(n8006) );
  NAND2_X1 U8360 ( .A1(n7792), .A2(n8033), .ZN(n7151) );
  INV_X1 U8361 ( .A(n8064), .ZN(n7940) );
  NAND2_X1 U8362 ( .A1(n8494), .A2(n7940), .ZN(n7140) );
  NAND2_X1 U8363 ( .A1(n8495), .A2(n10243), .ZN(n7916) );
  OR2_X1 U8364 ( .A1(n8269), .A2(n8142), .ZN(n7149) );
  AND2_X1 U8365 ( .A1(n7149), .A2(n8006), .ZN(n7156) );
  NAND2_X1 U8366 ( .A1(n7943), .A2(n7156), .ZN(n6636) );
  NAND2_X1 U8367 ( .A1(n8269), .A2(n8142), .ZN(n7152) );
  NAND2_X1 U8368 ( .A1(n6636), .A2(n7152), .ZN(n8128) );
  OR2_X1 U8369 ( .A1(n8257), .A2(n8180), .ZN(n8174) );
  AND2_X1 U8370 ( .A1(n8225), .A2(n8174), .ZN(n7155) );
  NAND2_X1 U8371 ( .A1(n8257), .A2(n8180), .ZN(n7153) );
  NAND2_X1 U8372 ( .A1(n7153), .A2(n8490), .ZN(n6638) );
  INV_X1 U8373 ( .A(n7153), .ZN(n6637) );
  AOI22_X1 U8374 ( .A1(n8360), .A2(n6638), .B1(n6637), .B2(n8351), .ZN(n6639)
         );
  NAND2_X1 U8375 ( .A1(n7166), .A2(n6639), .ZN(n6640) );
  INV_X1 U8376 ( .A(n8815), .ZN(n8444) );
  OR2_X1 U8377 ( .A1(n8893), .A2(n8444), .ZN(n7169) );
  NAND2_X1 U8378 ( .A1(n8964), .A2(n6642), .ZN(n7172) );
  OR2_X1 U8379 ( .A1(n8964), .A2(n6642), .ZN(n7173) );
  NAND2_X1 U8380 ( .A1(n8247), .A2(n8475), .ZN(n7175) );
  OR2_X1 U8381 ( .A1(n8247), .A2(n8475), .ZN(n7176) );
  NAND2_X1 U8382 ( .A1(n8952), .A2(n8771), .ZN(n6651) );
  OR2_X1 U8383 ( .A1(n8952), .A2(n8771), .ZN(n6652) );
  NAND2_X1 U8384 ( .A1(n8779), .A2(n8402), .ZN(n7182) );
  OR2_X1 U8385 ( .A1(n8779), .A2(n8402), .ZN(n7183) );
  OR2_X1 U8386 ( .A1(n8941), .A2(n8772), .ZN(n7180) );
  NAND2_X1 U8387 ( .A1(n8941), .A2(n8772), .ZN(n7190) );
  NAND2_X1 U8388 ( .A1(n8938), .A2(n8732), .ZN(n7189) );
  NAND2_X1 U8389 ( .A1(n7192), .A2(n7189), .ZN(n8741) );
  NAND2_X1 U8390 ( .A1(n8933), .A2(n8749), .ZN(n7193) );
  NAND2_X1 U8391 ( .A1(n8729), .A2(n8731), .ZN(n8716) );
  OR2_X1 U8392 ( .A1(n8927), .A2(n8733), .ZN(n7194) );
  AND2_X1 U8393 ( .A1(n7194), .A2(n8715), .ZN(n7187) );
  NAND2_X1 U8394 ( .A1(n8927), .A2(n8733), .ZN(n7195) );
  NAND2_X1 U8395 ( .A1(n8863), .A2(n6644), .ZN(n7200) );
  AND2_X1 U8396 ( .A1(n8700), .A2(n8708), .ZN(n8685) );
  NOR2_X1 U8397 ( .A1(n8685), .A2(n8288), .ZN(n6645) );
  OR2_X1 U8398 ( .A1(n8700), .A2(n8708), .ZN(n8289) );
  INV_X1 U8399 ( .A(n8685), .ZN(n7202) );
  NAND2_X1 U8400 ( .A1(n8313), .A2(n8681), .ZN(n8686) );
  NAND2_X1 U8401 ( .A1(n6650), .A2(n8386), .ZN(n7088) );
  OAI211_X1 U8402 ( .C1(n6646), .C2(n7202), .A(n8686), .B(n7088), .ZN(n6647)
         );
  OR2_X1 U8403 ( .A1(n6650), .A2(n8386), .ZN(n7212) );
  NAND2_X1 U8404 ( .A1(n8912), .A2(n8680), .ZN(n7113) );
  OR2_X1 U8405 ( .A1(n8462), .A2(n8465), .ZN(n7218) );
  NOR2_X1 U8406 ( .A1(n6725), .A2(n8659), .ZN(n7221) );
  XNOR2_X1 U8407 ( .A(n6765), .B(n4621), .ZN(n8654) );
  NAND2_X1 U8408 ( .A1(n8779), .A2(n8789), .ZN(n8758) );
  NAND2_X1 U8409 ( .A1(n6652), .A2(n6651), .ZN(n8787) );
  NAND2_X1 U8410 ( .A1(n8758), .A2(n8787), .ZN(n6677) );
  NAND2_X1 U8411 ( .A1(n7602), .A2(n7601), .ZN(n6655) );
  NAND2_X1 U8412 ( .A1(n6633), .A2(n7964), .ZN(n6654) );
  NAND2_X1 U8413 ( .A1(n6655), .A2(n6654), .ZN(n10209) );
  NAND2_X1 U8414 ( .A1(n7605), .A2(n10224), .ZN(n6656) );
  NAND2_X1 U8415 ( .A1(n8497), .A2(n7666), .ZN(n6658) );
  NAND2_X1 U8416 ( .A1(n7725), .A2(n10235), .ZN(n6659) );
  NOR2_X1 U8417 ( .A1(n8495), .A2(n7824), .ZN(n6660) );
  INV_X1 U8418 ( .A(n7920), .ZN(n6661) );
  NAND2_X1 U8419 ( .A1(n6661), .A2(n4486), .ZN(n6663) );
  NAND2_X1 U8420 ( .A1(n7724), .A2(n7940), .ZN(n6662) );
  NAND2_X1 U8421 ( .A1(n6663), .A2(n6662), .ZN(n7949) );
  NAND2_X1 U8422 ( .A1(n7957), .A2(n7792), .ZN(n6664) );
  NAND2_X1 U8423 ( .A1(n7149), .A2(n7152), .ZN(n7091) );
  OAI21_X1 U8424 ( .B1(n8257), .B2(n8491), .A(n7091), .ZN(n6669) );
  NAND2_X1 U8425 ( .A1(n8269), .A2(n8492), .ZN(n8130) );
  NAND2_X1 U8426 ( .A1(n8130), .A2(n8180), .ZN(n6667) );
  INV_X1 U8427 ( .A(n8130), .ZN(n6666) );
  AOI22_X1 U8428 ( .A1(n8257), .A2(n6667), .B1(n6666), .B2(n8491), .ZN(n6668)
         );
  OR2_X1 U8429 ( .A1(n8360), .A2(n8490), .ZN(n8233) );
  AND2_X1 U8430 ( .A1(n8229), .A2(n8233), .ZN(n6670) );
  NAND2_X1 U8431 ( .A1(n8893), .A2(n8815), .ZN(n8810) );
  NAND2_X1 U8432 ( .A1(n8447), .A2(n4718), .ZN(n8809) );
  OR2_X1 U8433 ( .A1(n8964), .A2(n8827), .ZN(n7090) );
  OR2_X1 U8434 ( .A1(n8893), .A2(n8815), .ZN(n8812) );
  AND2_X1 U8435 ( .A1(n7090), .A2(n8812), .ZN(n6671) );
  NAND2_X1 U8436 ( .A1(n8964), .A2(n8827), .ZN(n7089) );
  OR2_X1 U8437 ( .A1(n8247), .A2(n8816), .ZN(n6672) );
  NAND2_X1 U8438 ( .A1(n8247), .A2(n8816), .ZN(n6673) );
  NAND2_X1 U8439 ( .A1(n7180), .A2(n7190), .ZN(n7178) );
  OR2_X1 U8440 ( .A1(n8952), .A2(n8797), .ZN(n8767) );
  INV_X1 U8441 ( .A(n8767), .ZN(n8756) );
  OAI21_X1 U8442 ( .B1(n8767), .B2(n8789), .A(n8779), .ZN(n6675) );
  OAI21_X1 U8443 ( .B1(n8756), .B2(n8402), .A(n6675), .ZN(n6676) );
  NAND2_X1 U8444 ( .A1(n8941), .A2(n8489), .ZN(n6678) );
  OR2_X1 U8445 ( .A1(n8938), .A2(n8761), .ZN(n6679) );
  NAND2_X1 U8446 ( .A1(n8933), .A2(n8722), .ZN(n6681) );
  NAND2_X1 U8447 ( .A1(n7194), .A2(n7195), .ZN(n8720) );
  OR2_X1 U8448 ( .A1(n8927), .A2(n8488), .ZN(n6682) );
  NAND2_X1 U8449 ( .A1(n8288), .A2(n7200), .ZN(n8705) );
  NAND2_X1 U8450 ( .A1(n8706), .A2(n8705), .ZN(n6684) );
  OR2_X1 U8451 ( .A1(n8863), .A2(n8723), .ZN(n6683) );
  XNOR2_X1 U8452 ( .A(n8700), .B(n8708), .ZN(n8694) );
  OR2_X1 U8453 ( .A1(n8700), .A2(n8487), .ZN(n6685) );
  NOR2_X1 U8454 ( .A1(n8313), .A2(n8695), .ZN(n6688) );
  NAND2_X1 U8455 ( .A1(n8313), .A2(n8695), .ZN(n6687) );
  AND2_X1 U8456 ( .A1(n6650), .A2(n8669), .ZN(n6690) );
  OR2_X1 U8457 ( .A1(n8912), .A2(n8680), .ZN(n7213) );
  NAND2_X1 U8458 ( .A1(n7213), .A2(n7113), .ZN(n8675) );
  OR2_X1 U8459 ( .A1(n8912), .A2(n8486), .ZN(n6691) );
  NAND2_X1 U8460 ( .A1(n8462), .A2(n8670), .ZN(n6692) );
  INV_X1 U8461 ( .A(n7936), .ZN(n7081) );
  NAND2_X1 U8462 ( .A1(n7594), .A2(n7081), .ZN(n6693) );
  OR2_X1 U8463 ( .A1(n6703), .A2(n7936), .ZN(n6704) );
  NAND2_X1 U8464 ( .A1(n7524), .A2(n6706), .ZN(n6707) );
  NAND2_X1 U8465 ( .A1(n7525), .A2(n6707), .ZN(n6710) );
  INV_X1 U8466 ( .A(n7525), .ZN(n6708) );
  NAND2_X1 U8467 ( .A1(n6708), .A2(n7522), .ZN(n6709) );
  MUX2_X1 U8468 ( .A(n10539), .B(n6721), .S(n10254), .Z(n6713) );
  NAND2_X1 U8469 ( .A1(n6725), .A2(n8888), .ZN(n6712) );
  NAND2_X1 U8470 ( .A1(n6713), .A2(n6712), .ZN(P2_U3486) );
  INV_X1 U8471 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6722) );
  AND2_X1 U8472 ( .A1(n6714), .A2(n7517), .ZN(n6715) );
  OR2_X1 U8473 ( .A1(n6716), .A2(n6715), .ZN(n6720) );
  NAND2_X1 U8474 ( .A1(n6718), .A2(n6717), .ZN(n6719) );
  MUX2_X1 U8475 ( .A(n6722), .B(n6721), .S(n10247), .Z(n6724) );
  NAND2_X1 U8476 ( .A1(n6725), .A2(n6778), .ZN(n6723) );
  NAND2_X1 U8477 ( .A1(n6724), .A2(n6723), .ZN(P2_U3454) );
  AND2_X1 U8478 ( .A1(n6725), .A2(n8485), .ZN(n6727) );
  AND2_X1 U8479 ( .A1(n6731), .A2(n6734), .ZN(n6732) );
  AND2_X1 U8480 ( .A1(n6732), .A2(n6733), .ZN(n6741) );
  INV_X1 U8481 ( .A(n6733), .ZN(n6740) );
  INV_X1 U8482 ( .A(n6734), .ZN(n6738) );
  AND2_X1 U8483 ( .A1(n6736), .A2(n6735), .ZN(n6737) );
  INV_X1 U8484 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8979) );
  INV_X1 U8485 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10558) );
  MUX2_X1 U8486 ( .A(n8979), .B(n10558), .S(n4409), .Z(n6749) );
  XNOR2_X1 U8487 ( .A(n6749), .B(SI_28_), .ZN(n6746) );
  NAND2_X1 U8488 ( .A1(n8977), .A2(n6278), .ZN(n6744) );
  OR2_X1 U8489 ( .A1(n7071), .A2(n8979), .ZN(n6743) );
  NOR2_X1 U8490 ( .A1(n8844), .A2(n8484), .ZN(n6745) );
  INV_X1 U8491 ( .A(n8844), .ZN(n8647) );
  NAND2_X1 U8492 ( .A1(n6747), .A2(n6746), .ZN(n6751) );
  INV_X1 U8493 ( .A(SI_28_), .ZN(n6748) );
  NAND2_X1 U8494 ( .A1(n6749), .A2(n6748), .ZN(n6750) );
  INV_X1 U8495 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8975) );
  INV_X1 U8496 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10581) );
  MUX2_X1 U8497 ( .A(n8975), .B(n10581), .S(n4403), .Z(n7043) );
  XNOR2_X1 U8498 ( .A(n7043), .B(SI_29_), .ZN(n6752) );
  NAND2_X1 U8499 ( .A1(n8974), .A2(n6278), .ZN(n6754) );
  OR2_X1 U8500 ( .A1(n7071), .A2(n8975), .ZN(n6753) );
  NAND2_X1 U8501 ( .A1(n6754), .A2(n6753), .ZN(n6777) );
  INV_X1 U8502 ( .A(n8624), .ZN(n6755) );
  NAND2_X1 U8503 ( .A1(n6755), .A2(n6270), .ZN(n7062) );
  INV_X1 U8504 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n6758) );
  NAND2_X1 U8505 ( .A1(n6265), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6757) );
  NAND2_X1 U8506 ( .A1(n6604), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6756) );
  OAI211_X1 U8507 ( .C1(n7058), .C2(n6758), .A(n6757), .B(n6756), .ZN(n6759)
         );
  INV_X1 U8508 ( .A(n6759), .ZN(n6760) );
  OR2_X1 U8509 ( .A1(n6777), .A2(n8638), .ZN(n7086) );
  NAND2_X1 U8510 ( .A1(n6777), .A2(n8638), .ZN(n7074) );
  NAND2_X1 U8511 ( .A1(n7086), .A2(n7074), .ZN(n7237) );
  XNOR2_X1 U8512 ( .A(n6762), .B(n6761), .ZN(n6763) );
  NAND2_X1 U8513 ( .A1(n6763), .A2(n8829), .ZN(n6775) );
  INV_X1 U8514 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n10573) );
  NAND2_X1 U8515 ( .A1(n6766), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6768) );
  NAND2_X1 U8516 ( .A1(n6265), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6767) );
  OAI211_X1 U8517 ( .C1(n6769), .C2(n10573), .A(n6768), .B(n6767), .ZN(n6770)
         );
  INV_X1 U8518 ( .A(n6770), .ZN(n6771) );
  AND2_X1 U8519 ( .A1(n7062), .A2(n6771), .ZN(n7054) );
  NAND2_X1 U8520 ( .A1(n8826), .A2(n6772), .ZN(n8622) );
  OAI22_X1 U8521 ( .A1(n7223), .A2(n10211), .B1(n7054), .B2(n8622), .ZN(n6773)
         );
  INV_X1 U8522 ( .A(n6773), .ZN(n6774) );
  NOR2_X1 U8523 ( .A1(n8635), .A2(n8137), .ZN(n6776) );
  OR2_X1 U8524 ( .A1(n6782), .A2(n10249), .ZN(n6781) );
  NAND2_X1 U8525 ( .A1(n6777), .A2(n6778), .ZN(n6780) );
  NAND2_X1 U8526 ( .A1(n6781), .A2(n5363), .ZN(P2_U3456) );
  OR2_X1 U8527 ( .A1(n6782), .A2(n10257), .ZN(n6785) );
  NAND2_X1 U8528 ( .A1(n6777), .A2(n8888), .ZN(n6784) );
  NAND2_X1 U8529 ( .A1(n10257), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6783) );
  NAND2_X1 U8530 ( .A1(n6785), .A2(n5360), .ZN(P2_U3488) );
  NOR2_X1 U8531 ( .A1(n6912), .A2(P2_U3151), .ZN(n6786) );
  NAND2_X1 U8532 ( .A1(n7217), .A2(n6912), .ZN(n6787) );
  NAND2_X1 U8533 ( .A1(n6787), .A2(n7353), .ZN(n10286) );
  NAND2_X1 U8534 ( .A1(n6788), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NAND2_X1 U8535 ( .A1(n6188), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6790) );
  NAND2_X1 U8536 ( .A1(n6789), .A2(n6790), .ZN(n10168) );
  NOR2_X1 U8537 ( .A1(n10168), .A2(n10169), .ZN(n10167) );
  INV_X1 U8538 ( .A(n6790), .ZN(n6791) );
  XNOR2_X1 U8539 ( .A(n7508), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n7498) );
  NOR2_X1 U8540 ( .A1(n7497), .A2(n7498), .ZN(n7496) );
  INV_X1 U8541 ( .A(n6792), .ZN(n10188) );
  XNOR2_X1 U8542 ( .A(n10184), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n10189) );
  NOR2_X1 U8543 ( .A1(n6793), .A2(n10450), .ZN(n6794) );
  XOR2_X1 U8544 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6851), .Z(n7544) );
  INV_X1 U8545 ( .A(n6851), .ZN(n7545) );
  INV_X1 U8546 ( .A(n6799), .ZN(n7750) );
  XNOR2_X1 U8547 ( .A(n7333), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n7748) );
  NAND2_X1 U8548 ( .A1(n6802), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6803) );
  INV_X1 U8549 ( .A(n6863), .ZN(n7996) );
  OAI21_X1 U8550 ( .B1(n6804), .B2(n7996), .A(n6805), .ZN(n7998) );
  INV_X1 U8551 ( .A(n6805), .ZN(n7984) );
  XNOR2_X1 U8552 ( .A(n6867), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n7983) );
  INV_X1 U8553 ( .A(n6808), .ZN(n8522) );
  XNOR2_X1 U8554 ( .A(n6876), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n8521) );
  OR2_X1 U8555 ( .A1(n6876), .A2(n8831), .ZN(n6809) );
  INV_X1 U8556 ( .A(n6881), .ZN(n8535) );
  NAND2_X1 U8557 ( .A1(n6810), .A2(n8535), .ZN(n6811) );
  INV_X1 U8558 ( .A(n6811), .ZN(n8550) );
  XNOR2_X1 U8559 ( .A(n6886), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n8549) );
  NAND2_X1 U8560 ( .A1(n6813), .A2(n5242), .ZN(n8579) );
  NAND2_X1 U8561 ( .A1(n6814), .A2(n6891), .ZN(n6815) );
  INV_X1 U8562 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8791) );
  OAI21_X1 U8563 ( .B1(n6895), .B2(n6816), .A(n8581), .ZN(n6817) );
  INV_X1 U8564 ( .A(n6899), .ZN(n8594) );
  NAND2_X1 U8565 ( .A1(n6817), .A2(n8594), .ZN(n8603) );
  INV_X1 U8566 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8763) );
  INV_X1 U8567 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8747) );
  OR2_X1 U8568 ( .A1(n8610), .A2(n8747), .ZN(n6819) );
  NAND2_X1 U8569 ( .A1(n8610), .A2(n8747), .ZN(n6818) );
  NAND2_X1 U8570 ( .A1(n6819), .A2(n6818), .ZN(n8602) );
  XNOR2_X1 U8571 ( .A(n7080), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n6907) );
  XNOR2_X1 U8572 ( .A(n6820), .B(n6907), .ZN(n6822) );
  INV_X1 U8573 ( .A(n10286), .ZN(n6821) );
  OR2_X1 U8574 ( .A1(n7247), .A2(P2_U3151), .ZN(n10284) );
  INV_X1 U8575 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10308) );
  INV_X1 U8576 ( .A(n7508), .ZN(n6839) );
  INV_X1 U8577 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10250) );
  AND2_X1 U8578 ( .A1(n6188), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6824) );
  NAND2_X1 U8579 ( .A1(n10297), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6823) );
  OAI22_X1 U8580 ( .A1(n6824), .A2(n10179), .B1(n6188), .B2(n6823), .ZN(n10165) );
  NAND2_X1 U8581 ( .A1(n10165), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6826) );
  INV_X1 U8582 ( .A(n6824), .ZN(n6825) );
  NAND2_X1 U8583 ( .A1(n6826), .A2(n6825), .ZN(n7494) );
  INV_X1 U8584 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10255) );
  MUX2_X1 U8585 ( .A(n10255), .B(P2_REG1_REG_4__SCAN_IN), .S(n10184), .Z(
        n10187) );
  INV_X1 U8586 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6827) );
  MUX2_X1 U8587 ( .A(n10308), .B(P2_REG1_REG_6__SCAN_IN), .S(n6851), .Z(n7541)
         );
  XNOR2_X1 U8588 ( .A(n6828), .B(n6855), .ZN(n7644) );
  AOI22_X1 U8589 ( .A1(n7644), .A2(P2_REG1_REG_7__SCAN_IN), .B1(n6798), .B2(
        n6828), .ZN(n7743) );
  XOR2_X1 U8590 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n7333), .Z(n7744) );
  INV_X1 U8591 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10426) );
  INV_X1 U8592 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10438) );
  XNOR2_X1 U8593 ( .A(n6867), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n7978) );
  INV_X1 U8594 ( .A(n6867), .ZN(n7982) );
  INV_X1 U8595 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6831) );
  XNOR2_X1 U8596 ( .A(n6876), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n8515) );
  INV_X1 U8597 ( .A(n6876), .ZN(n8520) );
  XNOR2_X1 U8598 ( .A(n6832), .B(n6881), .ZN(n8530) );
  INV_X1 U8599 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8887) );
  XNOR2_X1 U8600 ( .A(n6886), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n8544) );
  INV_X1 U8601 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8881) );
  XNOR2_X1 U8602 ( .A(n6895), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8573) );
  INV_X1 U8603 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n10436) );
  XNOR2_X1 U8604 ( .A(n8610), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8601) );
  INV_X1 U8605 ( .A(n8610), .ZN(n8615) );
  XNOR2_X1 U8606 ( .A(n7857), .B(n8869), .ZN(n6906) );
  NOR2_X1 U8607 ( .A1(n10284), .A2(n7248), .ZN(n6834) );
  XNOR2_X1 U8608 ( .A(n6837), .B(n10179), .ZN(n10172) );
  INV_X1 U8609 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6835) );
  MUX2_X1 U8610 ( .A(n6836), .B(n6835), .S(n6910), .Z(n10290) );
  NAND2_X1 U8611 ( .A1(n10172), .A2(n10289), .ZN(n10171) );
  NAND2_X1 U8612 ( .A1(n6837), .A2(n5221), .ZN(n6838) );
  NAND2_X1 U8613 ( .A1(n10171), .A2(n6838), .ZN(n7505) );
  MUX2_X1 U8614 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n6910), .Z(n6840) );
  XNOR2_X1 U8615 ( .A(n6840), .B(n6839), .ZN(n7504) );
  NAND2_X1 U8616 ( .A1(n7505), .A2(n7504), .ZN(n7503) );
  NAND2_X1 U8617 ( .A1(n6840), .A2(n7508), .ZN(n6841) );
  MUX2_X1 U8618 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n6910), .Z(n6842) );
  XNOR2_X1 U8619 ( .A(n6842), .B(n7306), .ZN(n7427) );
  INV_X1 U8620 ( .A(n6842), .ZN(n6843) );
  NAND2_X1 U8621 ( .A1(n6843), .A2(n5247), .ZN(n6844) );
  MUX2_X1 U8622 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n6910), .Z(n6845) );
  XNOR2_X1 U8623 ( .A(n6845), .B(n10184), .ZN(n10183) );
  NAND2_X1 U8624 ( .A1(n6845), .A2(n10184), .ZN(n6846) );
  MUX2_X1 U8625 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n6910), .Z(n6848) );
  XNOR2_X1 U8626 ( .A(n6848), .B(n6847), .ZN(n7464) );
  NAND2_X1 U8627 ( .A1(n7465), .A2(n7464), .ZN(n7463) );
  NAND2_X1 U8628 ( .A1(n6848), .A2(n5233), .ZN(n6849) );
  NAND2_X1 U8629 ( .A1(n7463), .A2(n6849), .ZN(n7537) );
  MUX2_X1 U8630 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n6910), .Z(n6850) );
  XNOR2_X1 U8631 ( .A(n6850), .B(n7545), .ZN(n7538) );
  INV_X1 U8632 ( .A(n6850), .ZN(n6852) );
  NAND2_X1 U8633 ( .A1(n6852), .A2(n6851), .ZN(n6853) );
  MUX2_X1 U8634 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n6910), .Z(n6854) );
  XNOR2_X1 U8635 ( .A(n6854), .B(n6855), .ZN(n7646) );
  INV_X1 U8636 ( .A(n6854), .ZN(n6856) );
  NAND2_X1 U8637 ( .A1(n6856), .A2(n6855), .ZN(n6857) );
  MUX2_X1 U8638 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n6910), .Z(n6858) );
  XNOR2_X1 U8639 ( .A(n6858), .B(n7333), .ZN(n7745) );
  NAND2_X1 U8640 ( .A1(n7746), .A2(n7745), .ZN(n6861) );
  INV_X1 U8641 ( .A(n6858), .ZN(n6859) );
  NAND2_X1 U8642 ( .A1(n6859), .A2(n7333), .ZN(n6860) );
  MUX2_X1 U8643 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n6910), .Z(n6862) );
  XNOR2_X1 U8644 ( .A(n6862), .B(n6863), .ZN(n7993) );
  INV_X1 U8645 ( .A(n6862), .ZN(n6864) );
  NAND2_X1 U8646 ( .A1(n6864), .A2(n6863), .ZN(n6865) );
  MUX2_X1 U8647 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n6910), .Z(n6866) );
  XNOR2_X1 U8648 ( .A(n6866), .B(n6867), .ZN(n7979) );
  INV_X1 U8649 ( .A(n6866), .ZN(n6868) );
  NAND2_X1 U8650 ( .A1(n6868), .A2(n6867), .ZN(n6869) );
  NAND2_X1 U8651 ( .A1(n6870), .A2(n6869), .ZN(n8509) );
  MUX2_X1 U8652 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n6910), .Z(n6871) );
  XNOR2_X1 U8653 ( .A(n6871), .B(n8507), .ZN(n8508) );
  NAND2_X1 U8654 ( .A1(n8509), .A2(n8508), .ZN(n6874) );
  INV_X1 U8655 ( .A(n6871), .ZN(n6872) );
  NAND2_X1 U8656 ( .A1(n6872), .A2(n8507), .ZN(n6873) );
  NAND2_X1 U8657 ( .A1(n6874), .A2(n6873), .ZN(n8517) );
  MUX2_X1 U8658 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n6910), .Z(n6875) );
  XNOR2_X1 U8659 ( .A(n6875), .B(n6876), .ZN(n8516) );
  NAND2_X1 U8660 ( .A1(n8517), .A2(n8516), .ZN(n6879) );
  INV_X1 U8661 ( .A(n6875), .ZN(n6877) );
  NAND2_X1 U8662 ( .A1(n6877), .A2(n6876), .ZN(n6878) );
  NAND2_X1 U8663 ( .A1(n6879), .A2(n6878), .ZN(n8532) );
  MUX2_X1 U8664 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n6910), .Z(n6880) );
  XNOR2_X1 U8665 ( .A(n6880), .B(n6881), .ZN(n8531) );
  NAND2_X1 U8666 ( .A1(n8532), .A2(n8531), .ZN(n6884) );
  INV_X1 U8667 ( .A(n6880), .ZN(n6882) );
  NAND2_X1 U8668 ( .A1(n6882), .A2(n6881), .ZN(n6883) );
  MUX2_X1 U8669 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n6910), .Z(n6885) );
  XNOR2_X1 U8670 ( .A(n6885), .B(n6886), .ZN(n8545) );
  INV_X1 U8671 ( .A(n6885), .ZN(n6887) );
  NAND2_X1 U8672 ( .A1(n6887), .A2(n6886), .ZN(n6888) );
  MUX2_X1 U8673 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n6910), .Z(n6889) );
  XNOR2_X1 U8674 ( .A(n6891), .B(n6889), .ZN(n8560) );
  INV_X1 U8675 ( .A(n6889), .ZN(n6890) );
  NAND2_X1 U8676 ( .A1(n6891), .A2(n6890), .ZN(n6892) );
  NAND2_X1 U8677 ( .A1(n6893), .A2(n6892), .ZN(n8575) );
  MUX2_X1 U8678 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n6910), .Z(n6894) );
  XNOR2_X1 U8679 ( .A(n6894), .B(n6895), .ZN(n8574) );
  INV_X1 U8680 ( .A(n6894), .ZN(n6896) );
  NAND2_X1 U8681 ( .A1(n6896), .A2(n6895), .ZN(n6897) );
  MUX2_X1 U8682 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n6910), .Z(n6898) );
  XNOR2_X1 U8683 ( .A(n6898), .B(n6899), .ZN(n8590) );
  INV_X1 U8684 ( .A(n6898), .ZN(n6900) );
  AND2_X1 U8685 ( .A1(n6900), .A2(n6899), .ZN(n6901) );
  MUX2_X1 U8686 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n6910), .Z(n6903) );
  NAND2_X1 U8687 ( .A1(n8612), .A2(n8610), .ZN(n8608) );
  INV_X1 U8688 ( .A(n6902), .ZN(n6905) );
  INV_X1 U8689 ( .A(n6903), .ZN(n6904) );
  NAND2_X1 U8690 ( .A1(n6905), .A2(n6904), .ZN(n8611) );
  NAND2_X1 U8691 ( .A1(n8608), .A2(n8611), .ZN(n6909) );
  MUX2_X1 U8692 ( .A(n6907), .B(n6906), .S(n6910), .Z(n6908) );
  XNOR2_X1 U8693 ( .A(n6909), .B(n6908), .ZN(n6917) );
  NOR2_X1 U8694 ( .A1(n6910), .A2(P2_U3151), .ZN(n8981) );
  NAND2_X1 U8695 ( .A1(n10286), .A2(n8981), .ZN(n6911) );
  MUX2_X1 U8696 ( .A(n8606), .B(n6911), .S(n7247), .Z(n10298) );
  INV_X1 U8697 ( .A(n6912), .ZN(n6913) );
  AND2_X1 U8698 ( .A1(n7353), .A2(n6913), .ZN(n6914) );
  NAND2_X1 U8699 ( .A1(n10170), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n6915) );
  NAND2_X1 U8700 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8366) );
  OAI211_X1 U8701 ( .C1(n10298), .C2(n7857), .A(n6915), .B(n8366), .ZN(n6916)
         );
  NAND2_X1 U8702 ( .A1(n6970), .A2(n7572), .ZN(n7571) );
  INV_X1 U8703 ( .A(n7571), .ZN(n7585) );
  NAND2_X1 U8704 ( .A1(n9489), .A2(n7710), .ZN(n6919) );
  NAND2_X1 U8705 ( .A1(n7585), .A2(n6919), .ZN(n6921) );
  AOI22_X1 U8706 ( .A1(n7584), .A2(n6919), .B1(n7849), .B2(n7589), .ZN(n6920)
         );
  NAND2_X1 U8707 ( .A1(n6921), .A2(n6920), .ZN(n7678) );
  NOR2_X1 U8708 ( .A1(n9487), .A2(n9349), .ZN(n7731) );
  NAND2_X1 U8709 ( .A1(n7885), .A2(n10153), .ZN(n9226) );
  NOR2_X1 U8710 ( .A1(n9486), .A2(n10153), .ZN(n7763) );
  NOR2_X1 U8711 ( .A1(n9485), .A2(n7888), .ZN(n6924) );
  AOI21_X1 U8712 ( .B1(n9431), .B2(n7763), .A(n6924), .ZN(n6925) );
  NAND2_X1 U8713 ( .A1(n6926), .A2(n6925), .ZN(n7801) );
  NAND2_X1 U8714 ( .A1(n7897), .A2(n7912), .ZN(n9231) );
  NAND2_X1 U8715 ( .A1(n9484), .A2(n7909), .ZN(n9230) );
  NAND2_X1 U8716 ( .A1(n9231), .A2(n9230), .ZN(n7804) );
  NAND2_X1 U8717 ( .A1(n8058), .A2(n9483), .ZN(n6975) );
  INV_X1 U8718 ( .A(n9483), .ZN(n8101) );
  NAND2_X1 U8719 ( .A1(n6975), .A2(n8042), .ZN(n8043) );
  NAND2_X1 U8720 ( .A1(n7801), .A2(n5371), .ZN(n6929) );
  NOR2_X1 U8721 ( .A1(n9484), .A2(n7912), .ZN(n7893) );
  NOR2_X1 U8722 ( .A1(n7968), .A2(n9483), .ZN(n6927) );
  AOI21_X1 U8723 ( .B1(n8043), .B2(n7893), .A(n6927), .ZN(n6928) );
  NAND2_X1 U8724 ( .A1(n6929), .A2(n6928), .ZN(n8100) );
  NAND2_X1 U8725 ( .A1(n9965), .A2(n9142), .ZN(n9242) );
  NAND2_X1 U8726 ( .A1(n8045), .A2(n9242), .ZN(n8102) );
  OR2_X1 U8727 ( .A1(n9965), .A2(n5051), .ZN(n6930) );
  OR2_X1 U8728 ( .A1(n9838), .A2(n9063), .ZN(n9252) );
  NAND2_X1 U8729 ( .A1(n9838), .A2(n9063), .ZN(n9247) );
  NAND2_X1 U8730 ( .A1(n9252), .A2(n9247), .ZN(n8047) );
  NAND2_X1 U8731 ( .A1(n8039), .A2(n8047), .ZN(n8038) );
  OR2_X1 U8732 ( .A1(n9838), .A2(n9482), .ZN(n6931) );
  NAND2_X1 U8733 ( .A1(n8038), .A2(n6931), .ZN(n8021) );
  OR2_X1 U8734 ( .A1(n8097), .A2(n9183), .ZN(n9255) );
  NAND2_X1 U8735 ( .A1(n8097), .A2(n9183), .ZN(n9254) );
  NAND2_X1 U8736 ( .A1(n9255), .A2(n9254), .ZN(n8020) );
  OR2_X1 U8737 ( .A1(n8097), .A2(n9481), .ZN(n6932) );
  NAND2_X1 U8738 ( .A1(n8019), .A2(n6932), .ZN(n8071) );
  OR2_X1 U8739 ( .A1(n8074), .A2(n9091), .ZN(n9256) );
  NAND2_X1 U8740 ( .A1(n8074), .A2(n9091), .ZN(n9257) );
  NAND2_X1 U8741 ( .A1(n9256), .A2(n9257), .ZN(n8070) );
  NAND2_X1 U8742 ( .A1(n8071), .A2(n8070), .ZN(n8069) );
  OR2_X1 U8743 ( .A1(n8074), .A2(n9480), .ZN(n6933) );
  NAND2_X1 U8744 ( .A1(n8069), .A2(n6933), .ZN(n8153) );
  OR2_X1 U8745 ( .A1(n9093), .A2(n9944), .ZN(n9258) );
  NAND2_X1 U8746 ( .A1(n9093), .A2(n9944), .ZN(n9364) );
  NAND2_X1 U8747 ( .A1(n9258), .A2(n9364), .ZN(n9439) );
  OR2_X1 U8748 ( .A1(n9093), .A2(n9479), .ZN(n6934) );
  NAND2_X1 U8749 ( .A1(n9941), .A2(n9934), .ZN(n9799) );
  OR2_X1 U8750 ( .A1(n9941), .A2(n9478), .ZN(n6935) );
  NAND2_X1 U8751 ( .A1(n9937), .A2(n9779), .ZN(n6936) );
  OR2_X1 U8752 ( .A1(n9925), .A2(n9919), .ZN(n9274) );
  NAND2_X1 U8753 ( .A1(n9925), .A2(n9919), .ZN(n9742) );
  NAND2_X1 U8754 ( .A1(n9274), .A2(n9742), .ZN(n9759) );
  NAND2_X1 U8755 ( .A1(n9758), .A2(n9759), .ZN(n6938) );
  NAND2_X1 U8756 ( .A1(n9925), .A2(n9780), .ZN(n6937) );
  NAND2_X1 U8757 ( .A1(n6938), .A2(n6937), .ZN(n9746) );
  OR2_X1 U8758 ( .A1(n9755), .A2(n9767), .ZN(n6939) );
  NAND2_X1 U8759 ( .A1(n9746), .A2(n6939), .ZN(n6941) );
  NAND2_X1 U8760 ( .A1(n9755), .A2(n9767), .ZN(n6940) );
  AND2_X1 U8761 ( .A1(n9914), .A2(n9744), .ZN(n6943) );
  NAND2_X1 U8762 ( .A1(n9720), .A2(n9477), .ZN(n6944) );
  AND2_X1 U8763 ( .A1(n9903), .A2(n9712), .ZN(n6945) );
  OR2_X1 U8764 ( .A1(n9903), .A2(n9712), .ZN(n6946) );
  NAND2_X1 U8765 ( .A1(n9896), .A2(n9702), .ZN(n6947) );
  NOR2_X1 U8766 ( .A1(n9656), .A2(n9876), .ZN(n6949) );
  AND2_X1 U8767 ( .A1(n6980), .A2(n9650), .ZN(n6950) );
  OR2_X1 U8768 ( .A1(n6980), .A2(n9650), .ZN(n6951) );
  NOR2_X1 U8769 ( .A1(n9625), .A2(n9633), .ZN(n6952) );
  NAND2_X1 U8770 ( .A1(n8980), .A2(n6953), .ZN(n6955) );
  OR2_X1 U8771 ( .A1(n9220), .A2(n10030), .ZN(n6954) );
  OR2_X2 U8772 ( .A1(n9859), .A2(n9609), .ZN(n9342) );
  NAND2_X1 U8773 ( .A1(n9859), .A2(n9609), .ZN(n9308) );
  NAND2_X1 U8774 ( .A1(n9342), .A2(n9308), .ZN(n9586) );
  NAND2_X1 U8775 ( .A1(n8977), .A2(n6953), .ZN(n6957) );
  OR2_X1 U8776 ( .A1(n9220), .A2(n10558), .ZN(n6956) );
  INV_X1 U8777 ( .A(n6960), .ZN(n6958) );
  NAND2_X1 U8778 ( .A1(n6958), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8279) );
  INV_X1 U8779 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6959) );
  NAND2_X1 U8780 ( .A1(n6960), .A2(n6959), .ZN(n6961) );
  NAND2_X1 U8781 ( .A1(n8279), .A2(n6961), .ZN(n9045) );
  INV_X1 U8782 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n10496) );
  NAND2_X1 U8783 ( .A1(n6986), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6963) );
  NAND2_X1 U8784 ( .A1(n5777), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6962) );
  OAI211_X1 U8785 ( .C1(n6989), .C2(n10496), .A(n6963), .B(n6962), .ZN(n6964)
         );
  INV_X1 U8786 ( .A(n6964), .ZN(n6965) );
  XNOR2_X1 U8787 ( .A(n7017), .B(n4932), .ZN(n9572) );
  NAND2_X1 U8788 ( .A1(n9335), .A2(n6968), .ZN(n6969) );
  NAND3_X1 U8789 ( .A1(n9404), .A2(n7620), .A3(n6969), .ZN(n7705) );
  NAND2_X1 U8790 ( .A1(n7573), .A2(n7695), .ZN(n7574) );
  NAND2_X1 U8791 ( .A1(n9489), .A2(n7589), .ZN(n9353) );
  NAND2_X1 U8792 ( .A1(n7590), .A2(n9353), .ZN(n6972) );
  NAND2_X1 U8793 ( .A1(n7849), .A2(n7710), .ZN(n6971) );
  XNOR2_X1 U8794 ( .A(n9487), .B(n9349), .ZN(n9428) );
  NAND2_X1 U8795 ( .A1(n6922), .A2(n9349), .ZN(n6973) );
  INV_X1 U8796 ( .A(n9431), .ZN(n7765) );
  AND2_X1 U8797 ( .A1(n9223), .A2(n9231), .ZN(n9228) );
  NAND2_X1 U8798 ( .A1(n7760), .A2(n9228), .ZN(n7898) );
  NAND2_X1 U8799 ( .A1(n9242), .A2(n8042), .ZN(n9237) );
  INV_X1 U8800 ( .A(n9230), .ZN(n6976) );
  INV_X1 U8801 ( .A(n8020), .ZN(n9437) );
  AND2_X1 U8802 ( .A1(n9258), .A2(n9256), .ZN(n9250) );
  INV_X1 U8803 ( .A(n9779), .ZN(n9816) );
  OR2_X1 U8804 ( .A1(n9937), .A2(n9816), .ZN(n9365) );
  NAND2_X1 U8805 ( .A1(n9937), .A2(n9816), .ZN(n9270) );
  NAND2_X1 U8806 ( .A1(n9365), .A2(n9270), .ZN(n9440) );
  INV_X1 U8807 ( .A(n9799), .ZN(n9268) );
  NOR2_X1 U8808 ( .A1(n9440), .A2(n9268), .ZN(n9262) );
  INV_X1 U8809 ( .A(n9803), .ZN(n9113) );
  OR2_X1 U8810 ( .A1(n9789), .A2(n9113), .ZN(n9276) );
  NAND2_X1 U8811 ( .A1(n9789), .A2(n9113), .ZN(n9271) );
  NAND2_X1 U8812 ( .A1(n9276), .A2(n9271), .ZN(n9775) );
  INV_X1 U8813 ( .A(n9365), .ZN(n9776) );
  NOR2_X1 U8814 ( .A1(n9775), .A2(n9776), .ZN(n6977) );
  NAND2_X1 U8815 ( .A1(n9774), .A2(n6977), .ZN(n9777) );
  INV_X1 U8816 ( .A(n9759), .ZN(n9766) );
  INV_X1 U8817 ( .A(n9767), .ZN(n9734) );
  OR2_X1 U8818 ( .A1(n9755), .A2(n9734), .ZN(n9281) );
  NAND2_X1 U8819 ( .A1(n9755), .A2(n9734), .ZN(n9283) );
  NAND2_X1 U8820 ( .A1(n9281), .A2(n9283), .ZN(n9279) );
  INV_X1 U8821 ( .A(n9742), .ZN(n9277) );
  NOR2_X1 U8822 ( .A1(n9279), .A2(n9277), .ZN(n6978) );
  INV_X1 U8823 ( .A(n9744), .ZN(n9120) );
  OR2_X1 U8824 ( .A1(n9914), .A2(n9120), .ZN(n9282) );
  NAND2_X1 U8825 ( .A1(n9914), .A2(n9120), .ZN(n9284) );
  NAND2_X1 U8826 ( .A1(n9282), .A2(n9284), .ZN(n9731) );
  OR2_X1 U8827 ( .A1(n9720), .A2(n9900), .ZN(n9280) );
  NAND2_X1 U8828 ( .A1(n9720), .A2(n9900), .ZN(n9376) );
  INV_X1 U8829 ( .A(n9702), .ZN(n9888) );
  OR2_X1 U8830 ( .A1(n9896), .A2(n9888), .ZN(n9291) );
  INV_X1 U8831 ( .A(n9712), .ZN(n9893) );
  AND2_X1 U8832 ( .A1(n9291), .A2(n9685), .ZN(n9380) );
  NAND2_X1 U8833 ( .A1(n9896), .A2(n9888), .ZN(n9298) );
  NAND2_X1 U8834 ( .A1(n9903), .A2(n9893), .ZN(n9288) );
  NAND2_X1 U8835 ( .A1(n9298), .A2(n9288), .ZN(n9292) );
  NAND2_X1 U8836 ( .A1(n9292), .A2(n9291), .ZN(n9385) );
  XNOR2_X1 U8837 ( .A(n9673), .B(n9300), .ZN(n9297) );
  INV_X1 U8838 ( .A(n9876), .ZN(n9639) );
  OR2_X1 U8839 ( .A1(n9673), .A2(n9300), .ZN(n9630) );
  INV_X1 U8840 ( .A(n9650), .ZN(n9869) );
  OR2_X1 U8841 ( .A1(n6980), .A2(n9869), .ZN(n9343) );
  NAND2_X1 U8842 ( .A1(n6980), .A2(n9869), .ZN(n9387) );
  NAND2_X1 U8843 ( .A1(n9656), .A2(n9639), .ZN(n9423) );
  NAND2_X1 U8844 ( .A1(n9387), .A2(n9423), .ZN(n6981) );
  NAND2_X1 U8845 ( .A1(n9625), .A2(n9608), .ZN(n9388) );
  XNOR2_X1 U8846 ( .A(n9866), .B(n4402), .ZN(n9604) );
  INV_X1 U8847 ( .A(n9586), .ZN(n9582) );
  NAND2_X1 U8848 ( .A1(n9866), .A2(n4402), .ZN(n9581) );
  NAND3_X1 U8849 ( .A1(n9606), .A2(n9582), .A3(n9581), .ZN(n6982) );
  NAND2_X1 U8850 ( .A1(n9556), .A2(n9405), .ZN(n6983) );
  OAI211_X1 U8851 ( .C1(n9446), .C2(n6984), .A(n7024), .B(n9782), .ZN(n6994)
         );
  OR2_X1 U8852 ( .A1(n8279), .A2(n6985), .ZN(n6992) );
  INV_X1 U8853 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n10498) );
  NAND2_X1 U8854 ( .A1(n5777), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6988) );
  NAND2_X1 U8855 ( .A1(n6986), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6987) );
  OAI211_X1 U8856 ( .C1(n6989), .C2(n10498), .A(n6988), .B(n6987), .ZN(n6990)
         );
  INV_X1 U8857 ( .A(n6990), .ZN(n6991) );
  INV_X1 U8858 ( .A(n6120), .ZN(n7300) );
  NAND2_X1 U8859 ( .A1(n9475), .A2(n9804), .ZN(n6993) );
  INV_X1 U8860 ( .A(n7695), .ZN(n7625) );
  NAND2_X1 U8861 ( .A1(n7581), .A2(n7625), .ZN(n7587) );
  NOR2_X2 U8862 ( .A1(n7805), .A2(n7912), .ZN(n7896) );
  INV_X1 U8863 ( .A(n8097), .ZN(n9018) );
  AND2_X2 U8864 ( .A1(n8023), .A2(n9018), .ZN(n8022) );
  NOR2_X4 U8865 ( .A1(n8072), .A2(n9093), .ZN(n8154) );
  INV_X1 U8866 ( .A(n9941), .ZN(n6996) );
  NOR2_X2 U8867 ( .A1(n9751), .A2(n9755), .ZN(n9735) );
  INV_X1 U8868 ( .A(n9914), .ZN(n9739) );
  NAND2_X1 U8869 ( .A1(n9717), .A2(n9996), .ZN(n9694) );
  INV_X1 U8870 ( .A(n9592), .ZN(n6997) );
  OAI211_X1 U8871 ( .C1(n5174), .C2(n6997), .A(n4450), .B(n9784), .ZN(n9575)
         );
  OAI21_X1 U8872 ( .B1(n9609), .B2(n9943), .A(n9575), .ZN(n6998) );
  AND2_X1 U8873 ( .A1(n7615), .A2(n9402), .ZN(n7006) );
  OAI21_X1 U8874 ( .B1(n7611), .B2(P1_D_REG_1__SCAN_IN), .A(n10019), .ZN(n7004) );
  NAND2_X1 U8875 ( .A1(n7002), .A2(n7001), .ZN(n7003) );
  NAND4_X1 U8876 ( .A1(n7006), .A2(n7005), .A3(n7004), .A4(n7003), .ZN(n7010)
         );
  INV_X1 U8877 ( .A(n7007), .ZN(n7008) );
  OAI21_X1 U8878 ( .B1(n7015), .B2(n10162), .A(n7008), .ZN(P1_U3550) );
  INV_X1 U8879 ( .A(n7616), .ZN(n7009) );
  INV_X1 U8880 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n7012) );
  NOR2_X1 U8881 ( .A1(n7011), .A2(n7013), .ZN(n7014) );
  OAI21_X1 U8882 ( .B1(n7015), .B2(n10160), .A(n7014), .ZN(P1_U3518) );
  NOR2_X1 U8883 ( .A1(n9578), .A2(n9584), .ZN(n7016) );
  INV_X1 U8884 ( .A(n8275), .ZN(n7021) );
  NAND2_X1 U8885 ( .A1(n8974), .A2(n6953), .ZN(n7019) );
  OR2_X1 U8886 ( .A1(n9220), .A2(n10581), .ZN(n7018) );
  OR2_X1 U8887 ( .A1(n8283), .A2(n7020), .ZN(n9447) );
  NAND2_X1 U8888 ( .A1(n8283), .A2(n7020), .ZN(n9339) );
  NAND2_X1 U8889 ( .A1(n9447), .A2(n9339), .ZN(n9321) );
  NAND3_X1 U8890 ( .A1(n7021), .A2(n9959), .A3(n5132), .ZN(n7036) );
  NAND2_X1 U8891 ( .A1(n9578), .A2(n9584), .ZN(n8274) );
  NAND4_X1 U8892 ( .A1(n8275), .A2(n9959), .A3(n9321), .A4(n8274), .ZN(n7035)
         );
  OR3_X1 U8893 ( .A1(n9321), .A2(n10157), .A3(n8274), .ZN(n7023) );
  AOI21_X1 U8894 ( .B1(n8283), .B2(n4450), .A(n9822), .ZN(n7022) );
  NAND2_X1 U8895 ( .A1(n9566), .A2(n7022), .ZN(n8280) );
  AND2_X1 U8896 ( .A1(n7023), .A2(n8280), .ZN(n7034) );
  NAND2_X1 U8897 ( .A1(n6112), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7028) );
  INV_X1 U8898 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9568) );
  OR2_X1 U8899 ( .A1(n4408), .A2(n9568), .ZN(n7027) );
  INV_X1 U8900 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n7025) );
  OR2_X1 U8901 ( .A1(n4406), .A2(n7025), .ZN(n7026) );
  AND3_X1 U8902 ( .A1(n7028), .A2(n7027), .A3(n7026), .ZN(n9338) );
  INV_X1 U8903 ( .A(n4413), .ZN(n7294) );
  NAND2_X1 U8904 ( .A1(n7294), .A2(P1_B_REG_SCAN_IN), .ZN(n7030) );
  NAND2_X1 U8905 ( .A1(n9804), .A2(n7030), .ZN(n9562) );
  NAND2_X1 U8906 ( .A1(n9584), .A2(n9877), .ZN(n7031) );
  OAI21_X1 U8907 ( .B1(n9338), .B2(n9562), .A(n7031), .ZN(n7032) );
  NAND4_X1 U8908 ( .A1(n7036), .A2(n7035), .A3(n7034), .A4(n8286), .ZN(n7255)
         );
  NAND2_X1 U8909 ( .A1(n7255), .A2(n10161), .ZN(n7041) );
  INV_X1 U8910 ( .A(n7039), .ZN(n7040) );
  NAND2_X1 U8911 ( .A1(n7041), .A2(n7040), .ZN(P1_U3519) );
  INV_X1 U8912 ( .A(SI_29_), .ZN(n7042) );
  AND2_X1 U8913 ( .A1(n7043), .A2(n7042), .ZN(n7046) );
  INV_X1 U8914 ( .A(n7043), .ZN(n7044) );
  NAND2_X1 U8915 ( .A1(n7044), .A2(SI_29_), .ZN(n7045) );
  INV_X1 U8916 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n10346) );
  INV_X1 U8917 ( .A(SI_30_), .ZN(n7048) );
  NAND2_X1 U8918 ( .A1(n7049), .A2(n7048), .ZN(n7064) );
  INV_X1 U8919 ( .A(n7049), .ZN(n7050) );
  NAND2_X1 U8920 ( .A1(n7050), .A2(SI_30_), .ZN(n7051) );
  NAND2_X1 U8921 ( .A1(n7064), .A2(n7051), .ZN(n7065) );
  NAND2_X1 U8922 ( .A1(n9218), .A2(n6278), .ZN(n7053) );
  OR2_X1 U8923 ( .A1(n7071), .A2(n10346), .ZN(n7052) );
  NAND2_X1 U8924 ( .A1(n7053), .A2(n7052), .ZN(n8841) );
  NAND2_X1 U8925 ( .A1(n8841), .A2(n7054), .ZN(n7226) );
  NAND2_X1 U8926 ( .A1(n7226), .A2(n7074), .ZN(n7229) );
  INV_X1 U8927 ( .A(n8841), .ZN(n8904) );
  INV_X1 U8928 ( .A(n7054), .ZN(n8483) );
  AND2_X1 U8929 ( .A1(n8904), .A2(n8483), .ZN(n7227) );
  INV_X1 U8930 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n7059) );
  NAND2_X1 U8931 ( .A1(n6604), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n7057) );
  INV_X1 U8932 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n7055) );
  OR2_X1 U8933 ( .A1(n6208), .A2(n7055), .ZN(n7056) );
  OAI211_X1 U8934 ( .C1(n7059), .C2(n7058), .A(n7057), .B(n7056), .ZN(n7060)
         );
  INV_X1 U8935 ( .A(n7060), .ZN(n7061) );
  AOI21_X1 U8936 ( .B1(n7063), .B2(n4701), .A(n5367), .ZN(n7079) );
  OAI21_X1 U8937 ( .B1(n7066), .B2(n7065), .A(n7064), .ZN(n7069) );
  INV_X1 U8938 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9215) );
  INV_X1 U8939 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n7070) );
  XNOR2_X1 U8940 ( .A(n7067), .B(SI_31_), .ZN(n7068) );
  XNOR2_X1 U8941 ( .A(n7069), .B(n7068), .ZN(n9214) );
  NAND2_X1 U8942 ( .A1(n9214), .A2(n6278), .ZN(n7073) );
  OR2_X1 U8943 ( .A1(n7071), .A2(n7070), .ZN(n7072) );
  INV_X1 U8944 ( .A(n7074), .ZN(n7075) );
  NAND3_X1 U8945 ( .A1(n7077), .A2(n8623), .A3(n8904), .ZN(n7078) );
  OAI21_X1 U8946 ( .B1(n7079), .B2(n8901), .A(n7078), .ZN(n7084) );
  NAND2_X1 U8947 ( .A1(n7081), .A2(n7080), .ZN(n7105) );
  NAND2_X1 U8948 ( .A1(n7081), .A2(n7857), .ZN(n7107) );
  NOR2_X1 U8949 ( .A1(n8082), .A2(n7107), .ZN(n7082) );
  NAND2_X1 U8950 ( .A1(n7084), .A2(n7082), .ZN(n7083) );
  OAI21_X1 U8951 ( .B1(n7084), .B2(n5362), .A(n7083), .ZN(n7085) );
  INV_X1 U8952 ( .A(n7227), .ZN(n7087) );
  INV_X1 U8953 ( .A(n7236), .ZN(n7104) );
  NAND2_X1 U8954 ( .A1(n7208), .A2(n8686), .ZN(n8292) );
  INV_X1 U8955 ( .A(n8720), .ZN(n8717) );
  NAND2_X1 U8956 ( .A1(n7090), .A2(n7089), .ZN(n8814) );
  NAND2_X1 U8957 ( .A1(n7598), .A2(n7125), .ZN(n7518) );
  NOR2_X1 U8958 ( .A1(n7602), .A2(n7518), .ZN(n7092) );
  NAND2_X1 U8959 ( .A1(n7145), .A2(n7138), .ZN(n7135) );
  INV_X1 U8960 ( .A(n7135), .ZN(n7635) );
  NAND4_X1 U8961 ( .A1(n7092), .A2(n7635), .A3(n10210), .A4(n7663), .ZN(n7094)
         );
  INV_X1 U8962 ( .A(n7916), .ZN(n7093) );
  OR2_X1 U8963 ( .A1(n7093), .A2(n7915), .ZN(n7820) );
  NAND2_X1 U8964 ( .A1(n7141), .A2(n7140), .ZN(n7919) );
  NOR4_X1 U8965 ( .A1(n7094), .A2(n7950), .A3(n7820), .A4(n7919), .ZN(n7095)
         );
  AND4_X1 U8966 ( .A1(n8234), .A2(n8132), .A3(n8008), .A4(n7095), .ZN(n7096)
         );
  XNOR2_X1 U8967 ( .A(n8360), .B(n8490), .ZN(n8179) );
  AND3_X1 U8968 ( .A1(n8814), .A2(n7096), .A3(n8179), .ZN(n7099) );
  INV_X1 U8969 ( .A(n8802), .ZN(n7097) );
  INV_X1 U8970 ( .A(n8833), .ZN(n7171) );
  NOR2_X1 U8971 ( .A1(n7097), .A2(n7171), .ZN(n7098) );
  NAND4_X1 U8972 ( .A1(n8776), .A2(n8783), .A3(n7099), .A4(n7098), .ZN(n7100)
         );
  NOR2_X1 U8973 ( .A1(n7178), .A2(n7100), .ZN(n7101) );
  NAND4_X1 U8974 ( .A1(n8717), .A2(n8731), .A3(n6643), .A4(n7101), .ZN(n7102)
         );
  NOR3_X1 U8975 ( .A1(n8292), .A2(n8705), .A3(n7102), .ZN(n7103) );
  INV_X1 U8976 ( .A(n7105), .ZN(n7106) );
  NAND2_X1 U8977 ( .A1(n7106), .A2(n8082), .ZN(n7111) );
  INV_X1 U8978 ( .A(n7107), .ZN(n7108) );
  NAND3_X1 U8979 ( .A1(n7112), .A2(n7108), .A3(n8082), .ZN(n7110) );
  OR2_X1 U8980 ( .A1(n7353), .A2(P2_U3151), .ZN(n8161) );
  INV_X1 U8981 ( .A(n8161), .ZN(n7109) );
  OAI211_X1 U8982 ( .C1(n7112), .C2(n7111), .A(n7110), .B(n7109), .ZN(n7244)
         );
  OAI21_X1 U8983 ( .B1(n7217), .B2(n7212), .A(n7113), .ZN(n7114) );
  NAND2_X1 U8984 ( .A1(n7215), .A2(n7114), .ZN(n7116) );
  NAND4_X1 U8985 ( .A1(n7213), .A2(n8386), .A3(n7217), .A4(n6650), .ZN(n7115)
         );
  OAI211_X1 U8986 ( .C1(n7213), .C2(n7217), .A(n7116), .B(n7115), .ZN(n7117)
         );
  INV_X1 U8987 ( .A(n7117), .ZN(n7216) );
  AND2_X1 U8988 ( .A1(n8797), .A2(n7217), .ZN(n7119) );
  OAI21_X1 U8989 ( .B1(n8797), .B2(n7217), .A(n8952), .ZN(n7118) );
  OAI21_X1 U8990 ( .B1(n7119), .B2(n8952), .A(n7118), .ZN(n7120) );
  AND3_X1 U8991 ( .A1(n7183), .A2(n7182), .A3(n7120), .ZN(n7179) );
  INV_X1 U8992 ( .A(n7121), .ZN(n7122) );
  OAI21_X1 U8993 ( .B1(n7128), .B2(n7122), .A(n7123), .ZN(n7124) );
  INV_X1 U8994 ( .A(n7125), .ZN(n7126) );
  NOR2_X1 U8995 ( .A1(n7602), .A2(n7126), .ZN(n7129) );
  AOI21_X1 U8996 ( .B1(n7129), .B2(n7128), .A(n7127), .ZN(n7130) );
  NAND2_X1 U8997 ( .A1(n7131), .A2(n7130), .ZN(n7136) );
  NAND2_X1 U8998 ( .A1(n7143), .A2(n7137), .ZN(n7139) );
  NAND2_X1 U8999 ( .A1(n7143), .A2(n7142), .ZN(n7146) );
  INV_X1 U9000 ( .A(n7915), .ZN(n7144) );
  AND2_X1 U9001 ( .A1(n7152), .A2(n7151), .ZN(n7154) );
  NAND2_X1 U9002 ( .A1(n8360), .A2(n8351), .ZN(n8226) );
  OAI211_X1 U9003 ( .C1(n7157), .C2(n7154), .A(n7153), .B(n8226), .ZN(n7159)
         );
  OAI21_X1 U9004 ( .B1(n7157), .B2(n7156), .A(n7155), .ZN(n7158) );
  INV_X1 U9005 ( .A(n7160), .ZN(n7161) );
  NAND2_X1 U9006 ( .A1(n7162), .A2(n7161), .ZN(n7164) );
  NAND3_X1 U9007 ( .A1(n7164), .A2(n7166), .A3(n8226), .ZN(n7163) );
  NAND2_X1 U9008 ( .A1(n7164), .A2(n8225), .ZN(n7167) );
  NAND2_X1 U9009 ( .A1(n8893), .A2(n8444), .ZN(n7168) );
  MUX2_X1 U9010 ( .A(n7169), .B(n7168), .S(n7217), .Z(n7170) );
  MUX2_X1 U9011 ( .A(n7173), .B(n7172), .S(n4420), .Z(n7174) );
  MUX2_X1 U9012 ( .A(n7176), .B(n7175), .S(n7217), .Z(n7177) );
  NAND2_X1 U9013 ( .A1(n7192), .A2(n7180), .ZN(n7181) );
  NAND2_X1 U9014 ( .A1(n7184), .A2(n7183), .ZN(n7185) );
  NAND2_X1 U9015 ( .A1(n7193), .A2(n7189), .ZN(n7188) );
  NAND2_X1 U9016 ( .A1(n8288), .A2(n7194), .ZN(n7197) );
  NAND2_X1 U9017 ( .A1(n7200), .A2(n7195), .ZN(n7196) );
  MUX2_X1 U9018 ( .A(n7197), .B(n7196), .S(n7217), .Z(n7198) );
  INV_X1 U9019 ( .A(n7198), .ZN(n7199) );
  MUX2_X1 U9020 ( .A(n8288), .B(n7200), .S(n4420), .Z(n7201) );
  AND2_X1 U9021 ( .A1(n7201), .A2(n5103), .ZN(n7206) );
  NAND2_X1 U9022 ( .A1(n7208), .A2(n8289), .ZN(n7204) );
  NAND2_X1 U9023 ( .A1(n7202), .A2(n8686), .ZN(n7203) );
  MUX2_X1 U9024 ( .A(n7204), .B(n7203), .S(n7217), .Z(n7205) );
  INV_X1 U9025 ( .A(n7208), .ZN(n7209) );
  NAND2_X1 U9026 ( .A1(n7209), .A2(n7217), .ZN(n7210) );
  OAI211_X1 U9027 ( .C1(n8686), .C2(n7217), .A(n7088), .B(n7210), .ZN(n7211)
         );
  INV_X1 U9028 ( .A(n7211), .ZN(n7214) );
  MUX2_X1 U9029 ( .A(n7218), .B(n4527), .S(n7217), .Z(n7219) );
  MUX2_X1 U9030 ( .A(n7223), .B(n8647), .S(n7217), .Z(n7232) );
  MUX2_X1 U9031 ( .A(n7221), .B(n4793), .S(n4420), .Z(n7231) );
  AOI21_X1 U9032 ( .B1(n7232), .B2(n8484), .A(n7231), .ZN(n7222) );
  INV_X1 U9033 ( .A(n7232), .ZN(n7233) );
  OAI21_X1 U9034 ( .B1(n7227), .B2(n4420), .A(n7226), .ZN(n7228) );
  AOI21_X1 U9035 ( .B1(n7232), .B2(n8844), .A(n7231), .ZN(n7235) );
  AOI22_X1 U9036 ( .A1(n7235), .A2(n7234), .B1(n8647), .B2(n7233), .ZN(n7238)
         );
  NOR3_X1 U9037 ( .A1(n7249), .A2(n7248), .A3(n7247), .ZN(n7252) );
  OAI21_X1 U9038 ( .B1(n8161), .B2(n7250), .A(P2_B_REG_SCAN_IN), .ZN(n7251) );
  OR2_X1 U9039 ( .A1(n7252), .A2(n7251), .ZN(n7253) );
  NAND2_X1 U9040 ( .A1(n10162), .A2(n10498), .ZN(n7254) );
  OAI21_X1 U9041 ( .B1(n7255), .B2(n10162), .A(n7254), .ZN(n7257) );
  NAND2_X1 U9042 ( .A1(n8283), .A2(n9856), .ZN(n7256) );
  NAND2_X1 U9043 ( .A1(n7257), .A2(n7256), .ZN(P1_U3551) );
  XNOR2_X1 U9044 ( .A(n8484), .B(n7258), .ZN(n7259) );
  XNOR2_X1 U9045 ( .A(n8844), .B(n7259), .ZN(n7268) );
  INV_X1 U9046 ( .A(n7268), .ZN(n7260) );
  NAND2_X1 U9047 ( .A1(n7260), .A2(n8470), .ZN(n7273) );
  INV_X1 U9048 ( .A(n7267), .ZN(n7261) );
  NAND2_X1 U9049 ( .A1(n7261), .A2(n8485), .ZN(n7263) );
  NAND2_X1 U9050 ( .A1(n7274), .A2(n7264), .ZN(n7272) );
  AOI22_X1 U9051 ( .A1(n8645), .A2(n8478), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n7266) );
  NAND2_X1 U9052 ( .A1(n8485), .A2(n8441), .ZN(n7265) );
  OAI211_X1 U9053 ( .C1(n8638), .C2(n8454), .A(n7266), .B(n7265), .ZN(n7270)
         );
  NOR4_X1 U9054 ( .A1(n7268), .A2(n7267), .A3(n8659), .A4(n8460), .ZN(n7269)
         );
  AOI211_X1 U9055 ( .C1(n8844), .C2(n8457), .A(n7270), .B(n7269), .ZN(n7271)
         );
  OAI211_X1 U9056 ( .C1(n7274), .C2(n7273), .A(n7272), .B(n7271), .ZN(P2_U3160) );
  NAND2_X1 U9057 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n7284) );
  NOR2_X1 U9058 ( .A1(n7277), .A2(n7276), .ZN(n7278) );
  NOR2_X1 U9059 ( .A1(n7279), .A2(n7278), .ZN(n7694) );
  MUX2_X1 U9060 ( .A(n7284), .B(n7694), .S(n4413), .Z(n7280) );
  OR2_X1 U9061 ( .A1(n7280), .A2(n6120), .ZN(n7283) );
  NOR2_X1 U9062 ( .A1(n4413), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7281) );
  OR2_X1 U9063 ( .A1(n6120), .A2(n7281), .ZN(n10082) );
  NAND2_X1 U9064 ( .A1(n10082), .A2(n4764), .ZN(n10087) );
  AND2_X1 U9065 ( .A1(P1_U3973), .A2(n10087), .ZN(n7282) );
  AND2_X1 U9066 ( .A1(n7283), .A2(n7282), .ZN(n10104) );
  XNOR2_X1 U9067 ( .A(n7321), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9493) );
  INV_X1 U9068 ( .A(n7284), .ZN(n9492) );
  NAND2_X1 U9069 ( .A1(n9493), .A2(n9492), .ZN(n9491) );
  INV_X1 U9070 ( .A(n7321), .ZN(n9497) );
  NAND2_X1 U9071 ( .A1(n9497), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7285) );
  NAND2_X1 U9072 ( .A1(n9491), .A2(n7285), .ZN(n7291) );
  NAND2_X1 U9073 ( .A1(n7692), .A2(n9456), .ZN(n7299) );
  NAND2_X1 U9074 ( .A1(n9421), .A2(n7286), .ZN(n7288) );
  AND2_X1 U9075 ( .A1(n7288), .A2(n7287), .ZN(n7297) );
  NAND2_X1 U9076 ( .A1(n7299), .A2(n7297), .ZN(n10092) );
  NOR2_X1 U9077 ( .A1(n6120), .A2(n4413), .ZN(n9401) );
  INV_X1 U9078 ( .A(n9401), .ZN(n7289) );
  INV_X1 U9079 ( .A(n7360), .ZN(n7290) );
  OAI211_X1 U9080 ( .C1(n7292), .C2(n7291), .A(n10127), .B(n7290), .ZN(n7304)
         );
  XNOR2_X1 U9081 ( .A(n7321), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n9496) );
  AND2_X1 U9082 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9495) );
  NAND2_X1 U9083 ( .A1(n9496), .A2(n9495), .ZN(n9494) );
  NAND2_X1 U9084 ( .A1(n9497), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7293) );
  OAI211_X1 U9085 ( .C1(n7296), .C2(n7295), .A(n10131), .B(n5068), .ZN(n7303)
         );
  INV_X1 U9086 ( .A(n7297), .ZN(n7298) );
  AOI22_X1 U9087 ( .A1(n10089), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n7302) );
  OR2_X1 U9088 ( .A1(n10092), .A2(n7300), .ZN(n10100) );
  INV_X1 U9089 ( .A(n7316), .ZN(n7361) );
  NAND2_X1 U9090 ( .A1(n10146), .A2(n7361), .ZN(n7301) );
  NAND4_X1 U9091 ( .A1(n7304), .A2(n7303), .A3(n7302), .A4(n7301), .ZN(n7305)
         );
  OR2_X1 U9092 ( .A1(n10104), .A2(n7305), .ZN(P1_U3245) );
  INV_X2 U9093 ( .A(n8982), .ZN(n8991) );
  OAI222_X1 U9094 ( .A1(n8991), .A2(n4997), .B1(P2_U3151), .B2(n5221), .C1(
        n4411), .C2(n7322), .ZN(P2_U3294) );
  OAI222_X1 U9095 ( .A1(n8991), .A2(n7307), .B1(n4411), .B2(n7318), .C1(n7306), 
        .C2(P2_U3151), .ZN(P2_U3292) );
  OAI222_X1 U9096 ( .A1(n8991), .A2(n4721), .B1(n4411), .B2(n7317), .C1(n7508), 
        .C2(P2_U3151), .ZN(P2_U3293) );
  INV_X1 U9097 ( .A(n7308), .ZN(n7319) );
  OAI222_X1 U9098 ( .A1(n8991), .A2(n4860), .B1(n4411), .B2(n7319), .C1(n10184), .C2(P2_U3151), .ZN(P2_U3291) );
  INV_X1 U9099 ( .A(n7309), .ZN(n7324) );
  INV_X1 U9100 ( .A(n10037), .ZN(n10024) );
  AOI22_X1 U9101 ( .A1(n7400), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n10024), .ZN(n7310) );
  OAI21_X1 U9102 ( .B1(n7324), .B2(n10040), .A(n7310), .ZN(P1_U3349) );
  INV_X1 U9103 ( .A(n7311), .ZN(n7313) );
  INV_X1 U9104 ( .A(n10040), .ZN(n8164) );
  INV_X1 U9105 ( .A(n8164), .ZN(n10026) );
  AOI22_X1 U9106 ( .A1(n7384), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n10024), .ZN(n7312) );
  OAI21_X1 U9107 ( .B1(n7313), .B2(n10026), .A(n7312), .ZN(P1_U3350) );
  OAI222_X1 U9108 ( .A1(n8991), .A2(n4851), .B1(n4411), .B2(n7313), .C1(n5233), 
        .C2(P2_U3151), .ZN(P2_U3290) );
  NAND2_X1 U9109 ( .A1(n7315), .A2(P2_D_REG_1__SCAN_IN), .ZN(n7314) );
  OAI21_X1 U9110 ( .B1(n7315), .B2(n7522), .A(n7314), .ZN(P2_U3377) );
  OAI222_X1 U9111 ( .A1(n10037), .A2(n10306), .B1(n10026), .B2(n7317), .C1(
        n4401), .C2(n7316), .ZN(P1_U3353) );
  OAI222_X1 U9112 ( .A1(n10037), .A2(n10329), .B1(n10026), .B2(n7318), .C1(
        P1_U3086), .C2(n7357), .ZN(P1_U3352) );
  OAI222_X1 U9113 ( .A1(n10037), .A2(n7320), .B1(n10026), .B2(n7319), .C1(
        P1_U3086), .C2(n10099), .ZN(P1_U3351) );
  OAI222_X1 U9114 ( .A1(n10037), .A2(n7323), .B1(n10026), .B2(n7322), .C1(
        n7321), .C2(P1_U3086), .ZN(P1_U3354) );
  INV_X1 U9115 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7325) );
  OAI222_X1 U9116 ( .A1(n8991), .A2(n7325), .B1(n4411), .B2(n7324), .C1(n7545), 
        .C2(P2_U3151), .ZN(P2_U3289) );
  INV_X1 U9117 ( .A(n7326), .ZN(n7328) );
  AOI22_X1 U9118 ( .A1(n7479), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10024), .ZN(n7327) );
  OAI21_X1 U9119 ( .B1(n7328), .B2(n10040), .A(n7327), .ZN(P1_U3348) );
  INV_X1 U9120 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7329) );
  OAI222_X1 U9121 ( .A1(n8991), .A2(n7329), .B1(n4411), .B2(n7328), .C1(n6798), 
        .C2(P2_U3151), .ZN(P2_U3288) );
  INV_X1 U9122 ( .A(n7330), .ZN(n7334) );
  AOI22_X1 U9123 ( .A1(n7562), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10024), .ZN(n7331) );
  OAI21_X1 U9124 ( .B1(n7334), .B2(n10040), .A(n7331), .ZN(P1_U3347) );
  INV_X1 U9125 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n10508) );
  NOR2_X1 U9126 ( .A1(n7351), .A2(n10508), .ZN(P2_U3251) );
  INV_X1 U9127 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n10372) );
  NOR2_X1 U9128 ( .A1(n7351), .A2(n10372), .ZN(P2_U3252) );
  INV_X1 U9129 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n10507) );
  NOR2_X1 U9130 ( .A1(n7351), .A2(n10507), .ZN(P2_U3254) );
  INV_X1 U9131 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10541) );
  NOR2_X1 U9132 ( .A1(n7351), .A2(n10541), .ZN(P2_U3255) );
  INV_X1 U9133 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n10424) );
  NOR2_X1 U9134 ( .A1(n7351), .A2(n10424), .ZN(P2_U3260) );
  INV_X1 U9135 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10556) );
  NOR2_X1 U9136 ( .A1(n7351), .A2(n10556), .ZN(P2_U3256) );
  OAI222_X1 U9137 ( .A1(n8991), .A2(n7335), .B1(n4411), .B2(n7334), .C1(n6802), 
        .C2(P2_U3151), .ZN(P2_U3287) );
  NOR2_X1 U9138 ( .A1(n10089), .A2(P1_U3973), .ZN(P1_U3085) );
  NAND2_X1 U9139 ( .A1(n7336), .A2(P2_U3893), .ZN(n7337) );
  OAI21_X1 U9140 ( .B1(P2_U3893), .B2(n5488), .A(n7337), .ZN(P2_U3491) );
  INV_X1 U9141 ( .A(n7338), .ZN(n7342) );
  AOI22_X1 U9142 ( .A1(n7776), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n10024), .ZN(n7339) );
  OAI21_X1 U9143 ( .B1(n7342), .B2(n10026), .A(n7339), .ZN(P1_U3346) );
  AND2_X1 U9144 ( .A1(n7340), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U9145 ( .A1(n7340), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U9146 ( .A1(n7340), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U9147 ( .A1(n7340), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U9148 ( .A1(n7340), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U9149 ( .A1(n7340), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U9150 ( .A1(n7340), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  OAI222_X1 U9151 ( .A1(n4411), .A2(n7342), .B1(P2_U3151), .B2(n7996), .C1(
        n7341), .C2(n8991), .ZN(P2_U3286) );
  INV_X1 U9152 ( .A(n7343), .ZN(n7345) );
  AOI22_X1 U9153 ( .A1(n7863), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10024), .ZN(n7344) );
  OAI21_X1 U9154 ( .B1(n7345), .B2(n10040), .A(n7344), .ZN(P1_U3345) );
  OAI222_X1 U9155 ( .A1(n4411), .A2(n7345), .B1(P2_U3151), .B2(n7982), .C1(
        n10330), .C2(n8991), .ZN(P2_U3285) );
  NAND2_X1 U9156 ( .A1(n6112), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n7349) );
  INV_X1 U9157 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n7346) );
  OR2_X1 U9158 ( .A1(n4408), .A2(n7346), .ZN(n7348) );
  INV_X1 U9159 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10410) );
  OR2_X1 U9160 ( .A1(n4406), .A2(n10410), .ZN(n7347) );
  AND3_X1 U9161 ( .A1(n7349), .A2(n7348), .A3(n7347), .ZN(n9563) );
  INV_X1 U9162 ( .A(n9563), .ZN(n9419) );
  NAND2_X1 U9163 ( .A1(n9419), .A2(P1_U3973), .ZN(n7350) );
  OAI21_X1 U9164 ( .B1(P1_U3973), .B2(n7070), .A(n7350), .ZN(P1_U3585) );
  AND2_X1 U9165 ( .A1(n7340), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U9166 ( .A1(n7340), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U9167 ( .A1(n7340), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U9168 ( .A1(n7340), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U9169 ( .A1(n7340), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U9170 ( .A1(n7340), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U9171 ( .A1(n7340), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U9172 ( .A1(n7340), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U9173 ( .A1(n7340), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U9174 ( .A1(n7340), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U9175 ( .A1(n7340), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U9176 ( .A1(n7340), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U9177 ( .A1(n7340), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U9178 ( .A1(n7340), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U9179 ( .A1(n7340), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U9180 ( .A1(n7340), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U9181 ( .A1(n7340), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  INV_X1 U9182 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n7355) );
  NOR2_X1 U9183 ( .A1(n7352), .A2(P2_U3151), .ZN(n7354) );
  AOI22_X1 U9184 ( .A1(n7340), .A2(n7355), .B1(n7354), .B2(n7353), .ZN(
        P2_U3376) );
  INV_X1 U9185 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n10395) );
  INV_X1 U9186 ( .A(n10089), .ZN(n10148) );
  NAND2_X1 U9187 ( .A1(n10146), .A2(n7372), .ZN(n7356) );
  NAND2_X1 U9188 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(n4401), .ZN(n7785) );
  OAI211_X1 U9189 ( .C1(n10395), .C2(n10148), .A(n7356), .B(n7785), .ZN(n7366)
         );
  AOI211_X1 U9190 ( .C1(n7359), .C2(n7358), .A(n7367), .B(n10137), .ZN(n7365)
         );
  AOI211_X1 U9191 ( .C1(n7363), .C2(n7362), .A(n7371), .B(n10141), .ZN(n7364)
         );
  OR3_X1 U9192 ( .A1(n7366), .A2(n7365), .A3(n7364), .ZN(P1_U3246) );
  INV_X1 U9193 ( .A(n10099), .ZN(n7373) );
  INV_X1 U9194 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7368) );
  MUX2_X1 U9195 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n7368), .S(n10099), .Z(n10094) );
  NOR2_X1 U9196 ( .A1(n10095), .A2(n10094), .ZN(n10093) );
  XNOR2_X1 U9197 ( .A(n7384), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n7369) );
  AOI211_X1 U9198 ( .C1(n7370), .C2(n7369), .A(n10137), .B(n7383), .ZN(n7379)
         );
  MUX2_X1 U9199 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7736), .S(n10099), .Z(n10097) );
  XNOR2_X1 U9200 ( .A(n7384), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n7374) );
  AOI211_X1 U9201 ( .C1(n7375), .C2(n7374), .A(n10141), .B(n7380), .ZN(n7378)
         );
  INV_X1 U9202 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10511) );
  NAND2_X1 U9203 ( .A1(n10146), .A2(n7384), .ZN(n7376) );
  NAND2_X1 U9204 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7884) );
  OAI211_X1 U9205 ( .C1(n10511), .C2(n10148), .A(n7376), .B(n7884), .ZN(n7377)
         );
  OR3_X1 U9206 ( .A1(n7379), .A2(n7378), .A3(n7377), .ZN(P1_U3248) );
  XNOR2_X1 U9207 ( .A(n7400), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n7381) );
  AOI211_X1 U9208 ( .C1(n7382), .C2(n7381), .A(n10141), .B(n7399), .ZN(n7391)
         );
  XNOR2_X1 U9209 ( .A(n7400), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n7385) );
  AOI211_X1 U9210 ( .C1(n7386), .C2(n7385), .A(n10137), .B(n7396), .ZN(n7390)
         );
  INV_X1 U9211 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n7388) );
  NAND2_X1 U9212 ( .A1(n10146), .A2(n7400), .ZN(n7387) );
  NAND2_X1 U9213 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(n4401), .ZN(n7875) );
  OAI211_X1 U9214 ( .C1(n7388), .C2(n10148), .A(n7387), .B(n7875), .ZN(n7389)
         );
  OR3_X1 U9215 ( .A1(n7391), .A2(n7390), .A3(n7389), .ZN(P1_U3249) );
  INV_X1 U9216 ( .A(n7392), .ZN(n7394) );
  AOI22_X1 U9217 ( .A1(n8194), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10024), .ZN(n7393) );
  OAI21_X1 U9218 ( .B1(n7394), .B2(n10026), .A(n7393), .ZN(P1_U3344) );
  OAI222_X1 U9219 ( .A1(n8991), .A2(n7395), .B1(n4411), .B2(n7394), .C1(n4675), 
        .C2(P2_U3151), .ZN(P2_U3284) );
  XNOR2_X1 U9220 ( .A(n7479), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n7397) );
  AOI211_X1 U9221 ( .C1(n7398), .C2(n7397), .A(n10137), .B(n7475), .ZN(n7408)
         );
  INV_X1 U9222 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7401) );
  MUX2_X1 U9223 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n7401), .S(n7479), .Z(n7402)
         );
  INV_X1 U9224 ( .A(n7402), .ZN(n7403) );
  AOI211_X1 U9225 ( .C1(n7404), .C2(n7403), .A(n10141), .B(n7478), .ZN(n7407)
         );
  INV_X1 U9226 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10521) );
  NAND2_X1 U9227 ( .A1(n10146), .A2(n7479), .ZN(n7405) );
  NAND2_X1 U9228 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8056) );
  OAI211_X1 U9229 ( .C1(n10521), .C2(n10148), .A(n7405), .B(n8056), .ZN(n7406)
         );
  OR3_X1 U9230 ( .A1(n7408), .A2(n7407), .A3(n7406), .ZN(P1_U3250) );
  AOI22_X1 U9231 ( .A1(n8473), .A2(n5112), .B1(n7518), .B2(n8470), .ZN(n7410)
         );
  OR2_X1 U9232 ( .A1(n8478), .A2(P2_U3151), .ZN(n7449) );
  NAND2_X1 U9233 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(n7449), .ZN(n7409) );
  OAI211_X1 U9234 ( .C1(n8481), .C2(n7532), .A(n7410), .B(n7409), .ZN(P2_U3172) );
  INV_X1 U9235 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7414) );
  NAND2_X1 U9236 ( .A1(n7574), .A2(n9350), .ZN(n9426) );
  OAI21_X1 U9237 ( .B1(n9782), .B2(n9959), .A(n9426), .ZN(n7412) );
  NOR2_X1 U9238 ( .A1(n6918), .A2(n9815), .ZN(n7622) );
  INV_X1 U9239 ( .A(n7622), .ZN(n7411) );
  OAI211_X1 U9240 ( .C1(n7625), .C2(n7620), .A(n7412), .B(n7411), .ZN(n7491)
         );
  NAND2_X1 U9241 ( .A1(n7491), .A2(n10161), .ZN(n7413) );
  OAI21_X1 U9242 ( .B1(n10161), .B2(n7414), .A(n7413), .ZN(P1_U3453) );
  INV_X1 U9243 ( .A(n7415), .ZN(n7419) );
  INV_X1 U9244 ( .A(n7416), .ZN(n7417) );
  AOI21_X1 U9245 ( .B1(n7419), .B2(n7418), .A(n7417), .ZN(n7423) );
  AOI22_X1 U9246 ( .A1(n8473), .A2(n8498), .B1(n8457), .B2(n7607), .ZN(n7420)
         );
  OAI21_X1 U9247 ( .B1(n7604), .B2(n8476), .A(n7420), .ZN(n7421) );
  AOI21_X1 U9248 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7449), .A(n7421), .ZN(
        n7422) );
  OAI21_X1 U9249 ( .B1(n7423), .B2(n8460), .A(n7422), .ZN(P2_U3162) );
  INV_X1 U9250 ( .A(n7424), .ZN(n7425) );
  AOI21_X1 U9251 ( .B1(n7427), .B2(n7426), .A(n7425), .ZN(n7436) );
  INV_X1 U9252 ( .A(n10288), .ZN(n8609) );
  INV_X1 U9253 ( .A(n10298), .ZN(n10178) );
  XOR2_X1 U9254 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n7428), .Z(n7433) );
  OAI21_X1 U9255 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n7429), .A(n10190), .ZN(
        n7430) );
  NOR2_X1 U9256 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6217), .ZN(n7512) );
  AOI21_X1 U9257 ( .B1(n10191), .B2(n7430), .A(n7512), .ZN(n7432) );
  NAND2_X1 U9258 ( .A1(n10170), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n7431) );
  OAI211_X1 U9259 ( .C1(n7433), .C2(n10197), .A(n7432), .B(n7431), .ZN(n7434)
         );
  AOI21_X1 U9260 ( .B1(n5247), .B2(n10178), .A(n7434), .ZN(n7435) );
  OAI21_X1 U9261 ( .B1(n7436), .B2(n8609), .A(n7435), .ZN(P2_U3185) );
  INV_X1 U9262 ( .A(n7437), .ZN(n7443) );
  OAI222_X1 U9263 ( .A1(n4411), .A2(n7443), .B1(P2_U3151), .B2(n8520), .C1(
        n7438), .C2(n8991), .ZN(P2_U3283) );
  INV_X1 U9264 ( .A(n7439), .ZN(n7469) );
  AOI22_X1 U9265 ( .A1(n9535), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n10024), .ZN(n7440) );
  OAI21_X1 U9266 ( .B1(n7469), .B2(n10026), .A(n7440), .ZN(P1_U3341) );
  OAI21_X1 U9267 ( .B1(n8829), .B2(n10245), .A(n7518), .ZN(n7441) );
  NAND2_X1 U9268 ( .A1(n5112), .A2(n8826), .ZN(n7519) );
  OAI211_X1 U9269 ( .C1(n10242), .C2(n7532), .A(n7441), .B(n7519), .ZN(n8898)
         );
  NAND2_X1 U9270 ( .A1(n8898), .A2(n10247), .ZN(n7442) );
  OAI21_X1 U9271 ( .B1(n6179), .B2(n10247), .A(n7442), .ZN(P2_U3390) );
  OAI222_X1 U9272 ( .A1(n10037), .A2(n7444), .B1(n10026), .B2(n7443), .C1(
        n8195), .C2(n4401), .ZN(P1_U3343) );
  NAND2_X1 U9273 ( .A1(n9712), .A2(P1_U3973), .ZN(n7445) );
  OAI21_X1 U9274 ( .B1(n6452), .B2(P1_U3973), .A(n7445), .ZN(P1_U3574) );
  OAI21_X1 U9275 ( .B1(n7448), .B2(n7447), .A(n7446), .ZN(n7454) );
  NAND2_X1 U9276 ( .A1(n7449), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7452) );
  AOI22_X1 U9277 ( .A1(n8473), .A2(n8497), .B1(n8457), .B2(n7450), .ZN(n7451)
         );
  OAI211_X1 U9278 ( .C1(n6633), .C2(n8476), .A(n7452), .B(n7451), .ZN(n7453)
         );
  AOI21_X1 U9279 ( .B1(n7454), .B2(n8470), .A(n7453), .ZN(n7455) );
  INV_X1 U9280 ( .A(n7455), .ZN(P2_U3177) );
  XNOR2_X1 U9281 ( .A(n7456), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n7468) );
  XNOR2_X1 U9282 ( .A(n7457), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n7462) );
  NOR2_X1 U9283 ( .A1(n10298), .A2(n5233), .ZN(n7461) );
  INV_X1 U9284 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7459) );
  AND2_X1 U9285 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7727) );
  INV_X1 U9286 ( .A(n7727), .ZN(n7458) );
  OAI21_X1 U9287 ( .B1(n10294), .B2(n7459), .A(n7458), .ZN(n7460) );
  AOI211_X1 U9288 ( .C1(n7462), .C2(n10191), .A(n7461), .B(n7460), .ZN(n7467)
         );
  OAI211_X1 U9289 ( .C1(n7465), .C2(n7464), .A(n7463), .B(n10288), .ZN(n7466)
         );
  OAI211_X1 U9290 ( .C1(n7468), .C2(n10197), .A(n7467), .B(n7466), .ZN(
        P2_U3187) );
  INV_X1 U9291 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7470) );
  OAI222_X1 U9292 ( .A1(n8991), .A2(n7470), .B1(n4411), .B2(n7469), .C1(n5154), 
        .C2(P2_U3151), .ZN(P2_U3281) );
  OAI21_X1 U9293 ( .B1(P1_U3973), .B2(n5274), .A(n7471), .ZN(P1_U3554) );
  INV_X1 U9294 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10338) );
  INV_X1 U9295 ( .A(n7472), .ZN(n7474) );
  OAI222_X1 U9296 ( .A1(n10338), .A2(n8991), .B1(n4411), .B2(n7474), .C1(
        P2_U3151), .C2(n8535), .ZN(P2_U3282) );
  INV_X1 U9297 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10300) );
  INV_X1 U9298 ( .A(n9521), .ZN(n7473) );
  OAI222_X1 U9299 ( .A1(n10037), .A2(n10300), .B1(n10040), .B2(n7474), .C1(
        n4401), .C2(n7473), .ZN(P1_U3342) );
  XNOR2_X1 U9300 ( .A(n7562), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n7476) );
  AOI211_X1 U9301 ( .C1(n7477), .C2(n7476), .A(n10137), .B(n7554), .ZN(n7488)
         );
  XNOR2_X1 U9302 ( .A(n7562), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n7480) );
  AOI211_X1 U9303 ( .C1(n7481), .C2(n7480), .A(n10141), .B(n7561), .ZN(n7487)
         );
  INV_X1 U9304 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n7485) );
  NAND2_X1 U9305 ( .A1(n10146), .A2(n7562), .ZN(n7484) );
  NOR2_X1 U9306 ( .A1(n7482), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9060) );
  INV_X1 U9307 ( .A(n9060), .ZN(n7483) );
  OAI211_X1 U9308 ( .C1(n7485), .C2(n10148), .A(n7484), .B(n7483), .ZN(n7486)
         );
  OR3_X1 U9309 ( .A1(n7488), .A2(n7487), .A3(n7486), .ZN(P1_U3251) );
  INV_X1 U9310 ( .A(n7489), .ZN(n7515) );
  AOI22_X1 U9311 ( .A1(n9549), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n10024), .ZN(n7490) );
  OAI21_X1 U9312 ( .B1(n7515), .B2(n10026), .A(n7490), .ZN(P1_U3340) );
  INV_X1 U9313 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10083) );
  NAND2_X1 U9314 ( .A1(n7491), .A2(n10164), .ZN(n7492) );
  OAI21_X1 U9315 ( .B1(n10164), .B2(n10083), .A(n7492), .ZN(P1_U3522) );
  OAI21_X1 U9316 ( .B1(n7495), .B2(n7494), .A(n7493), .ZN(n7502) );
  INV_X1 U9317 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10452) );
  NOR2_X1 U9318 ( .A1(n10294), .A2(n10452), .ZN(n7501) );
  AOI21_X1 U9319 ( .B1(n7498), .B2(n7497), .A(n7496), .ZN(n7499) );
  INV_X1 U9320 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10208) );
  OAI22_X1 U9321 ( .A1(n10176), .A2(n7499), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10208), .ZN(n7500) );
  AOI211_X1 U9322 ( .C1(n5231), .C2(n7502), .A(n7501), .B(n7500), .ZN(n7507)
         );
  OAI211_X1 U9323 ( .C1(n7505), .C2(n7504), .A(n7503), .B(n10288), .ZN(n7506)
         );
  OAI211_X1 U9324 ( .C1(n10298), .C2(n7508), .A(n7507), .B(n7506), .ZN(
        P2_U3184) );
  INV_X1 U9325 ( .A(n8478), .ZN(n8431) );
  OAI211_X1 U9326 ( .C1(n4561), .C2(n7510), .A(n7509), .B(n8470), .ZN(n7514)
         );
  OAI22_X1 U9327 ( .A1(n8476), .A2(n7605), .B1(n7725), .B2(n8454), .ZN(n7511)
         );
  AOI211_X1 U9328 ( .C1(n7666), .C2(n8457), .A(n7512), .B(n7511), .ZN(n7513)
         );
  OAI211_X1 U9329 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8431), .A(n7514), .B(
        n7513), .ZN(P2_U3158) );
  OAI222_X1 U9330 ( .A1(n8991), .A2(n7516), .B1(n4411), .B2(n7515), .C1(n5242), 
        .C2(P2_U3151), .ZN(P2_U3280) );
  NAND3_X1 U9331 ( .A1(n7518), .A2(n10242), .A3(n7517), .ZN(n7520) );
  NAND2_X1 U9332 ( .A1(n7520), .A2(n7519), .ZN(n7529) );
  INV_X1 U9333 ( .A(n7521), .ZN(n7528) );
  NAND2_X1 U9334 ( .A1(n7525), .A2(n7522), .ZN(n7523) );
  OAI21_X1 U9335 ( .B1(n7525), .B2(n7524), .A(n7523), .ZN(n7526) );
  INV_X1 U9336 ( .A(n7526), .ZN(n7527) );
  MUX2_X1 U9337 ( .A(n7529), .B(P2_REG2_REG_0__SCAN_IN), .S(n10223), .Z(n7534)
         );
  INV_X1 U9338 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7531) );
  OAI22_X1 U9339 ( .A1(n8711), .A2(n7532), .B1(n7531), .B2(n10207), .ZN(n7533)
         );
  OR2_X1 U9340 ( .A1(n7534), .A2(n7533), .ZN(P2_U3233) );
  INV_X1 U9341 ( .A(n7535), .ZN(n7536) );
  AOI21_X1 U9342 ( .B1(n7538), .B2(n7537), .A(n7536), .ZN(n7552) );
  OAI21_X1 U9343 ( .B1(n7541), .B2(n7540), .A(n7539), .ZN(n7550) );
  AOI21_X1 U9344 ( .B1(n7544), .B2(n7543), .A(n7542), .ZN(n7548) );
  AND2_X1 U9345 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7795) );
  NOR2_X1 U9346 ( .A1(n10298), .A2(n7545), .ZN(n7546) );
  AOI211_X1 U9347 ( .C1(n10170), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n7795), .B(
        n7546), .ZN(n7547) );
  OAI21_X1 U9348 ( .B1(n7548), .B2(n10176), .A(n7547), .ZN(n7549) );
  AOI21_X1 U9349 ( .B1(n5231), .B2(n7550), .A(n7549), .ZN(n7551) );
  OAI21_X1 U9350 ( .B1(n7552), .B2(n8609), .A(n7551), .ZN(P2_U3188) );
  INV_X1 U9351 ( .A(n7553), .ZN(n7569) );
  INV_X1 U9352 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10467) );
  OAI222_X1 U9353 ( .A1(n4411), .A2(n7569), .B1(P2_U3151), .B2(n8578), .C1(
        n10467), .C2(n8991), .ZN(P2_U3279) );
  XOR2_X1 U9354 ( .A(n7776), .B(P1_REG1_REG_9__SCAN_IN), .Z(n7556) );
  NAND2_X1 U9355 ( .A1(n7555), .A2(n7556), .ZN(n7772) );
  OAI21_X1 U9356 ( .B1(n7556), .B2(n7555), .A(n7772), .ZN(n7560) );
  INV_X1 U9357 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7558) );
  NAND2_X1 U9358 ( .A1(n10146), .A2(n7776), .ZN(n7557) );
  NAND2_X1 U9359 ( .A1(n4401), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9140) );
  OAI211_X1 U9360 ( .C1(n7558), .C2(n10148), .A(n7557), .B(n9140), .ZN(n7559)
         );
  AOI21_X1 U9361 ( .B1(n7560), .B2(n10131), .A(n7559), .ZN(n7568) );
  MUX2_X1 U9362 ( .A(n5621), .B(P1_REG2_REG_9__SCAN_IN), .S(n7776), .Z(n7563)
         );
  INV_X1 U9363 ( .A(n7563), .ZN(n7564) );
  OAI21_X1 U9364 ( .B1(n7565), .B2(n7564), .A(n7775), .ZN(n7566) );
  NAND2_X1 U9365 ( .A1(n7566), .A2(n10127), .ZN(n7567) );
  NAND2_X1 U9366 ( .A1(n7568), .A2(n7567), .ZN(P1_U3252) );
  INV_X1 U9367 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7570) );
  INV_X1 U9368 ( .A(n10112), .ZN(n9550) );
  OAI222_X1 U9369 ( .A1(n10037), .A2(n7570), .B1(n10040), .B2(n7569), .C1(
        n9550), .C2(P1_U3086), .ZN(P1_U3339) );
  OAI21_X1 U9370 ( .B1(n6970), .B2(n7572), .A(n7571), .ZN(n7830) );
  INV_X1 U9371 ( .A(n7830), .ZN(n7580) );
  INV_X1 U9372 ( .A(n7705), .ZN(n8107) );
  OAI22_X1 U9373 ( .A1(n7573), .A2(n9943), .B1(n7849), .B2(n9815), .ZN(n7578)
         );
  NAND2_X1 U9374 ( .A1(n6970), .A2(n7574), .ZN(n7575) );
  AOI21_X1 U9375 ( .B1(n7576), .B2(n7575), .A(n9817), .ZN(n7577) );
  AOI211_X1 U9376 ( .C1(n8107), .C2(n7830), .A(n7578), .B(n7577), .ZN(n7828)
         );
  AOI21_X1 U9377 ( .B1(n9072), .B2(n7695), .A(n9822), .ZN(n7579) );
  NAND2_X1 U9378 ( .A1(n7579), .A2(n7587), .ZN(n7832) );
  OAI211_X1 U9379 ( .C1(n7580), .C2(n9968), .A(n7828), .B(n7832), .ZN(n7657)
         );
  OAI22_X1 U9380 ( .A1(n10016), .A2(n7581), .B1(n10161), .B2(n5471), .ZN(n7582) );
  AOI21_X1 U9381 ( .B1(n7657), .B2(n10161), .A(n7582), .ZN(n7583) );
  INV_X1 U9382 ( .A(n7583), .ZN(P1_U3456) );
  XNOR2_X1 U9383 ( .A(n9489), .B(n7589), .ZN(n9432) );
  NOR2_X1 U9384 ( .A1(n7585), .A2(n7584), .ZN(n7586) );
  XOR2_X1 U9385 ( .A(n9432), .B(n7586), .Z(n7714) );
  INV_X1 U9386 ( .A(n10154), .ZN(n9950) );
  INV_X1 U9387 ( .A(n7587), .ZN(n7588) );
  OAI211_X1 U9388 ( .C1(n7589), .C2(n7588), .A(n5190), .B(n9784), .ZN(n7712)
         );
  OAI21_X1 U9389 ( .B1(n7589), .B2(n9950), .A(n7712), .ZN(n7592) );
  XNOR2_X1 U9390 ( .A(n7590), .B(n9432), .ZN(n7591) );
  OAI222_X1 U9391 ( .A1(n9815), .A2(n6922), .B1(n9943), .B2(n6918), .C1(n9817), 
        .C2(n7591), .ZN(n7703) );
  AOI211_X1 U9392 ( .C1(n7714), .C2(n9959), .A(n7592), .B(n7703), .ZN(n10151)
         );
  NAND2_X1 U9393 ( .A1(n10162), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7593) );
  OAI21_X1 U9394 ( .B1(n10151), .B2(n10162), .A(n7593), .ZN(P1_U3524) );
  AND2_X1 U9395 ( .A1(n7595), .A2(n7594), .ZN(n10220) );
  INV_X1 U9396 ( .A(n10220), .ZN(n7596) );
  NAND2_X1 U9397 ( .A1(n8177), .A2(n7596), .ZN(n7597) );
  OAI21_X1 U9398 ( .B1(n7600), .B2(n6634), .A(n7599), .ZN(n7628) );
  INV_X1 U9399 ( .A(n7628), .ZN(n7610) );
  XOR2_X1 U9400 ( .A(n7602), .B(n7601), .Z(n7603) );
  OAI222_X1 U9401 ( .A1(n10212), .A2(n7605), .B1(n10211), .B2(n7604), .C1(
        n10218), .C2(n7603), .ZN(n7627) );
  INV_X1 U9402 ( .A(n7627), .ZN(n7606) );
  MUX2_X1 U9403 ( .A(n10169), .B(n7606), .S(n10221), .Z(n7609) );
  AOI22_X1 U9404 ( .A1(n8838), .A2(n7607), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8821), .ZN(n7608) );
  OAI211_X1 U9405 ( .C1(n8835), .C2(n7610), .A(n7609), .B(n7608), .ZN(P2_U3232) );
  NAND2_X1 U9406 ( .A1(n9402), .A2(n7612), .ZN(n7613) );
  NAND2_X1 U9407 ( .A1(n10150), .A2(n7613), .ZN(n7614) );
  NAND4_X1 U9408 ( .A1(n7616), .A2(n10019), .A3(n7615), .A4(n7614), .ZN(n7617)
         );
  AOI21_X1 U9409 ( .B1(n9807), .B2(n7619), .A(n9837), .ZN(n7626) );
  AND3_X1 U9410 ( .A1(n9426), .A2(n9404), .A3(n7620), .ZN(n7621) );
  AOI211_X1 U9411 ( .C1(n9836), .C2(P1_REG3_REG_0__SCAN_IN), .A(n7622), .B(
        n7621), .ZN(n7623) );
  MUX2_X1 U9412 ( .A(n5483), .B(n7623), .S(n9842), .Z(n7624) );
  OAI21_X1 U9413 ( .B1(n7626), .B2(n7625), .A(n7624), .ZN(P1_U3293) );
  AOI21_X1 U9414 ( .B1(n10245), .B2(n7628), .A(n7627), .ZN(n7967) );
  OAI22_X1 U9415 ( .A1(n8957), .A2(n7964), .B1(n6175), .B2(n10247), .ZN(n7629)
         );
  INV_X1 U9416 ( .A(n7629), .ZN(n7630) );
  OAI21_X1 U9417 ( .B1(n7967), .B2(n10249), .A(n7630), .ZN(P2_U3393) );
  XNOR2_X1 U9418 ( .A(n7631), .B(n7635), .ZN(n7632) );
  NAND2_X1 U9419 ( .A1(n7632), .A2(n8829), .ZN(n7634) );
  AOI22_X1 U9420 ( .A1(n8825), .A2(n8497), .B1(n8495), .B2(n8826), .ZN(n7633)
         );
  NAND2_X1 U9421 ( .A1(n7634), .A2(n7633), .ZN(n10236) );
  INV_X1 U9422 ( .A(n10236), .ZN(n7640) );
  XNOR2_X1 U9423 ( .A(n7636), .B(n7635), .ZN(n10238) );
  INV_X1 U9424 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10450) );
  AOI22_X1 U9425 ( .A1(n8838), .A2(n7673), .B1(n8821), .B2(n7674), .ZN(n7637)
         );
  OAI21_X1 U9426 ( .B1(n10450), .B2(n10221), .A(n7637), .ZN(n7638) );
  AOI21_X1 U9427 ( .B1(n10238), .B2(n8804), .A(n7638), .ZN(n7639) );
  OAI21_X1 U9428 ( .B1(n7640), .B2(n10223), .A(n7639), .ZN(P2_U3229) );
  INV_X1 U9429 ( .A(n7641), .ZN(n7690) );
  AOI22_X1 U9430 ( .A1(n10128), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10024), .ZN(n7642) );
  OAI21_X1 U9431 ( .B1(n7690), .B2(n10026), .A(n7642), .ZN(P1_U3338) );
  NAND2_X1 U9432 ( .A1(n9876), .A2(P1_U3973), .ZN(n7643) );
  OAI21_X1 U9433 ( .B1(P1_U3973), .B2(n8163), .A(n7643), .ZN(P1_U3577) );
  XOR2_X1 U9434 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n7644), .Z(n7656) );
  OAI21_X1 U9435 ( .B1(n7647), .B2(n7646), .A(n7645), .ZN(n7654) );
  AOI21_X1 U9436 ( .B1(n7649), .B2(n7648), .A(n7749), .ZN(n7652) );
  NOR2_X1 U9437 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6266), .ZN(n7926) );
  NOR2_X1 U9438 ( .A1(n10298), .A2(n6798), .ZN(n7650) );
  AOI211_X1 U9439 ( .C1(n10170), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n7926), .B(
        n7650), .ZN(n7651) );
  OAI21_X1 U9440 ( .B1(n7652), .B2(n10176), .A(n7651), .ZN(n7653) );
  AOI21_X1 U9441 ( .B1(n10288), .B2(n7654), .A(n7653), .ZN(n7655) );
  OAI21_X1 U9442 ( .B1(n7656), .B2(n10197), .A(n7655), .ZN(P2_U3189) );
  INV_X1 U9443 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7660) );
  NAND2_X1 U9444 ( .A1(n7657), .A2(n10164), .ZN(n7659) );
  NAND2_X1 U9445 ( .A1(n9856), .A2(n9072), .ZN(n7658) );
  OAI211_X1 U9446 ( .C1(n10164), .C2(n7660), .A(n7659), .B(n7658), .ZN(
        P1_U3523) );
  XOR2_X1 U9447 ( .A(n7661), .B(n7663), .Z(n10229) );
  XOR2_X1 U9448 ( .A(n7663), .B(n7662), .Z(n7664) );
  AOI222_X1 U9449 ( .A1(n8829), .A2(n7664), .B1(n8496), .B2(n8826), .C1(n8498), 
        .C2(n8825), .ZN(n10230) );
  MUX2_X1 U9450 ( .A(n7665), .B(n10230), .S(n10221), .Z(n7668) );
  AOI22_X1 U9451 ( .A1(n8838), .A2(n7666), .B1(n6217), .B2(n8821), .ZN(n7667)
         );
  OAI211_X1 U9452 ( .C1(n8835), .C2(n10229), .A(n7668), .B(n7667), .ZN(
        P2_U3230) );
  INV_X1 U9453 ( .A(n7669), .ZN(n7720) );
  AOI21_X1 U9454 ( .B1(n7671), .B2(n7670), .A(n7720), .ZN(n7677) );
  AND2_X1 U9455 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n10194) );
  OAI22_X1 U9456 ( .A1(n8476), .A2(n10213), .B1(n7793), .B2(n8454), .ZN(n7672)
         );
  AOI211_X1 U9457 ( .C1(n7673), .C2(n8457), .A(n10194), .B(n7672), .ZN(n7676)
         );
  NAND2_X1 U9458 ( .A1(n8478), .A2(n7674), .ZN(n7675) );
  OAI211_X1 U9459 ( .C1(n7677), .C2(n8460), .A(n7676), .B(n7675), .ZN(P2_U3170) );
  INV_X1 U9460 ( .A(n7678), .ZN(n7679) );
  NOR2_X1 U9461 ( .A1(n7679), .A2(n9428), .ZN(n7732) );
  INV_X1 U9462 ( .A(n7732), .ZN(n7680) );
  OAI21_X1 U9463 ( .B1(n4734), .B2(n7678), .A(n7680), .ZN(n7853) );
  OAI211_X1 U9464 ( .C1(n7682), .C2(n7848), .A(n9784), .B(n7681), .ZN(n7850)
         );
  OAI21_X1 U9465 ( .B1(n7849), .B2(n9943), .A(n7850), .ZN(n7685) );
  XOR2_X1 U9466 ( .A(n9428), .B(n7683), .Z(n7684) );
  OAI22_X1 U9467 ( .A1(n7684), .A2(n9817), .B1(n7885), .B2(n9815), .ZN(n7845)
         );
  AOI211_X1 U9468 ( .C1(n9959), .C2(n7853), .A(n7685), .B(n7845), .ZN(n7689)
         );
  OAI22_X1 U9469 ( .A1(n10016), .A2(n7848), .B1(n10161), .B2(n5523), .ZN(n7686) );
  INV_X1 U9470 ( .A(n7686), .ZN(n7687) );
  OAI21_X1 U9471 ( .B1(n7689), .B2(n10160), .A(n7687), .ZN(P1_U3462) );
  AOI22_X1 U9472 ( .A1(n9856), .A2(n9349), .B1(n10162), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n7688) );
  OAI21_X1 U9473 ( .B1(n7689), .B2(n10162), .A(n7688), .ZN(P1_U3525) );
  OAI222_X1 U9474 ( .A1(n8991), .A2(n7691), .B1(n4411), .B2(n7690), .C1(n8594), 
        .C2(P2_U3151), .ZN(P2_U3278) );
  OR2_X1 U9475 ( .A1(n7693), .A2(n7692), .ZN(n9071) );
  AOI22_X1 U9476 ( .A1(n7694), .A2(n9204), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n9071), .ZN(n7697) );
  AOI22_X1 U9477 ( .A1(n9171), .A2(n7695), .B1(n9192), .B2(n9490), .ZN(n7696)
         );
  NAND2_X1 U9478 ( .A1(n7697), .A2(n7696), .ZN(P1_U3232) );
  XOR2_X1 U9479 ( .A(n7699), .B(n7698), .Z(n7702) );
  AOI22_X1 U9480 ( .A1(n9171), .A2(n7710), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n9071), .ZN(n7701) );
  AOI22_X1 U9481 ( .A1(n9210), .A2(n9490), .B1(n9192), .B2(n9487), .ZN(n7700)
         );
  OAI211_X1 U9482 ( .C1(n7702), .C2(n9199), .A(n7701), .B(n7700), .ZN(P1_U3237) );
  INV_X1 U9483 ( .A(n7703), .ZN(n7716) );
  OR2_X1 U9484 ( .A1(n5869), .A2(n7704), .ZN(n7827) );
  NAND2_X1 U9485 ( .A1(n7705), .A2(n7827), .ZN(n7706) );
  INV_X1 U9486 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7708) );
  INV_X1 U9487 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7707) );
  OAI22_X1 U9488 ( .A1(n9842), .A2(n7708), .B1(n7707), .B2(n9785), .ZN(n7709)
         );
  AOI21_X1 U9489 ( .B1(n9837), .B2(n7710), .A(n7709), .ZN(n7711) );
  OAI21_X1 U9490 ( .B1(n9840), .B2(n7712), .A(n7711), .ZN(n7713) );
  AOI21_X1 U9491 ( .B1(n7714), .B2(n9847), .A(n7713), .ZN(n7715) );
  OAI21_X1 U9492 ( .B1(n7716), .B2(n9827), .A(n7715), .ZN(P1_U3291) );
  INV_X1 U9493 ( .A(n7823), .ZN(n7730) );
  INV_X1 U9494 ( .A(n7717), .ZN(n7719) );
  NOR3_X1 U9495 ( .A1(n7720), .A2(n7719), .A3(n7718), .ZN(n7723) );
  INV_X1 U9496 ( .A(n7721), .ZN(n7722) );
  OAI21_X1 U9497 ( .B1(n7723), .B2(n7722), .A(n8470), .ZN(n7729) );
  OAI22_X1 U9498 ( .A1(n8476), .A2(n7725), .B1(n7724), .B2(n8454), .ZN(n7726)
         );
  AOI211_X1 U9499 ( .C1(n7824), .C2(n8457), .A(n7727), .B(n7726), .ZN(n7728)
         );
  OAI211_X1 U9500 ( .C1(n7730), .C2(n8431), .A(n7729), .B(n7728), .ZN(P2_U3167) );
  NOR2_X1 U9501 ( .A1(n7732), .A2(n7731), .ZN(n7733) );
  INV_X1 U9502 ( .A(n9427), .ZN(n7734) );
  NOR2_X1 U9503 ( .A1(n7733), .A2(n7734), .ZN(n7764) );
  AOI21_X1 U9504 ( .B1(n7733), .B2(n7734), .A(n7764), .ZN(n10158) );
  XNOR2_X1 U9505 ( .A(n9227), .B(n7734), .ZN(n7735) );
  AOI222_X1 U9506 ( .A1(n9782), .A2(n7735), .B1(n9487), .B2(n9877), .C1(n9485), 
        .C2(n9804), .ZN(n10156) );
  MUX2_X1 U9507 ( .A(n7736), .B(n10156), .S(n9842), .Z(n7740) );
  AOI211_X1 U9508 ( .C1(n10153), .C2(n7681), .A(n9822), .B(n4549), .ZN(n10152)
         );
  OAI22_X1 U9509 ( .A1(n9763), .A2(n7812), .B1(n9785), .B2(n7737), .ZN(n7738)
         );
  AOI21_X1 U9510 ( .B1(n10152), .B2(n9807), .A(n7738), .ZN(n7739) );
  OAI211_X1 U9511 ( .C1(n10158), .C2(n9809), .A(n7740), .B(n7739), .ZN(
        P1_U3289) );
  INV_X1 U9512 ( .A(n7741), .ZN(n7759) );
  AOI22_X1 U9513 ( .A1(n10145), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10024), .ZN(n7742) );
  OAI21_X1 U9514 ( .B1(n7759), .B2(n10026), .A(n7742), .ZN(P1_U3337) );
  XOR2_X1 U9515 ( .A(n7744), .B(n7743), .Z(n7757) );
  XNOR2_X1 U9516 ( .A(n7746), .B(n7745), .ZN(n7755) );
  NAND2_X1 U9517 ( .A1(n10170), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7747) );
  NAND2_X1 U9518 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8144) );
  OAI211_X1 U9519 ( .C1(n10298), .C2(n6802), .A(n7747), .B(n8144), .ZN(n7754)
         );
  OR3_X1 U9520 ( .A1(n7750), .A2(n7749), .A3(n7748), .ZN(n7751) );
  AOI21_X1 U9521 ( .B1(n7752), .B2(n7751), .A(n10176), .ZN(n7753) );
  AOI211_X1 U9522 ( .C1(n10288), .C2(n7755), .A(n7754), .B(n7753), .ZN(n7756)
         );
  OAI21_X1 U9523 ( .B1(n7757), .B2(n10197), .A(n7756), .ZN(P2_U3190) );
  NAND2_X1 U9524 ( .A1(n8695), .A2(P2_U3893), .ZN(n7758) );
  OAI21_X1 U9525 ( .B1(P2_U3893), .B2(n5995), .A(n7758), .ZN(P2_U3514) );
  OAI222_X1 U9526 ( .A1(n4411), .A2(n7759), .B1(P2_U3151), .B2(n8615), .C1(
        n10487), .C2(n8991), .ZN(P2_U3277) );
  NAND3_X1 U9527 ( .A1(n9225), .A2(n9431), .A3(n9226), .ZN(n7761) );
  AOI21_X1 U9528 ( .B1(n7760), .B2(n7761), .A(n9817), .ZN(n7762) );
  AOI21_X1 U9529 ( .B1(n9804), .B2(n9484), .A(n7762), .ZN(n7837) );
  NOR2_X1 U9530 ( .A1(n7764), .A2(n7763), .ZN(n7766) );
  XNOR2_X1 U9531 ( .A(n7766), .B(n7765), .ZN(n7839) );
  OAI211_X1 U9532 ( .C1(n4549), .C2(n7840), .A(n7805), .B(n9784), .ZN(n7836)
         );
  NAND2_X1 U9533 ( .A1(n9842), .A2(n9877), .ZN(n9829) );
  INV_X1 U9534 ( .A(n9829), .ZN(n9681) );
  AOI22_X1 U9535 ( .A1(n9827), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7889), .B2(
        n9836), .ZN(n7767) );
  OAI21_X1 U9536 ( .B1(n9763), .B2(n7840), .A(n7767), .ZN(n7768) );
  AOI21_X1 U9537 ( .B1(n9681), .B2(n9486), .A(n7768), .ZN(n7769) );
  OAI21_X1 U9538 ( .B1(n9840), .B2(n7836), .A(n7769), .ZN(n7770) );
  AOI21_X1 U9539 ( .B1(n7839), .B2(n9847), .A(n7770), .ZN(n7771) );
  OAI21_X1 U9540 ( .B1(n9827), .B2(n7837), .A(n7771), .ZN(P1_U3288) );
  XNOR2_X1 U9541 ( .A(n7863), .B(P1_REG1_REG_10__SCAN_IN), .ZN(n7774) );
  OAI21_X1 U9542 ( .B1(n7776), .B2(P1_REG1_REG_9__SCAN_IN), .A(n7772), .ZN(
        n7773) );
  AOI211_X1 U9543 ( .C1(n7774), .C2(n7773), .A(n10137), .B(n7859), .ZN(n7782)
         );
  XNOR2_X1 U9544 ( .A(n7863), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n7778) );
  AOI211_X1 U9545 ( .C1(n7778), .C2(n7777), .A(n10141), .B(n7862), .ZN(n7781)
         );
  INV_X1 U9546 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10382) );
  NAND2_X1 U9547 ( .A1(n10146), .A2(n7863), .ZN(n7779) );
  NAND2_X1 U9548 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9016) );
  OAI211_X1 U9549 ( .C1(n10382), .C2(n10148), .A(n7779), .B(n9016), .ZN(n7780)
         );
  OR3_X1 U9550 ( .A1(n7782), .A2(n7781), .A3(n7780), .ZN(P1_U3253) );
  XOR2_X1 U9551 ( .A(n7784), .B(n7783), .Z(n7789) );
  AOI22_X1 U9552 ( .A1(n9210), .A2(n9489), .B1(n9192), .B2(n9486), .ZN(n7786)
         );
  OAI211_X1 U9553 ( .C1(n7848), .C2(n9213), .A(n7786), .B(n7785), .ZN(n7787)
         );
  AOI21_X1 U9554 ( .B1(n7846), .B2(n9197), .A(n7787), .ZN(n7788) );
  OAI21_X1 U9555 ( .B1(n7789), .B2(n9199), .A(n7788), .ZN(P1_U3218) );
  INV_X1 U9556 ( .A(n7923), .ZN(n7798) );
  OAI211_X1 U9557 ( .C1(n4547), .C2(n7791), .A(n7790), .B(n8470), .ZN(n7797)
         );
  OAI22_X1 U9558 ( .A1(n8476), .A2(n7793), .B1(n7792), .B2(n8454), .ZN(n7794)
         );
  AOI211_X1 U9559 ( .C1(n8064), .C2(n8457), .A(n7795), .B(n7794), .ZN(n7796)
         );
  OAI211_X1 U9560 ( .C1(n7798), .C2(n8431), .A(n7797), .B(n7796), .ZN(P2_U3179) );
  NAND2_X1 U9561 ( .A1(n7760), .A2(n9223), .ZN(n7799) );
  XNOR2_X1 U9562 ( .A(n7799), .B(n7804), .ZN(n7800) );
  OAI222_X1 U9563 ( .A1(n9943), .A2(n4645), .B1(n9815), .B2(n8101), .C1(n7800), 
        .C2(n9817), .ZN(n7906) );
  INV_X1 U9564 ( .A(n7906), .ZN(n7810) );
  INV_X1 U9565 ( .A(n7801), .ZN(n7802) );
  INV_X1 U9566 ( .A(n7804), .ZN(n9429) );
  NOR2_X1 U9567 ( .A1(n7802), .A2(n9429), .ZN(n7894) );
  INV_X1 U9568 ( .A(n7894), .ZN(n7803) );
  OAI21_X1 U9569 ( .B1(n7804), .B2(n7801), .A(n7803), .ZN(n7908) );
  AOI211_X1 U9570 ( .C1(n7912), .C2(n7805), .A(n9822), .B(n7896), .ZN(n7907)
         );
  NAND2_X1 U9571 ( .A1(n7907), .A2(n9807), .ZN(n7807) );
  AOI22_X1 U9572 ( .A1(n9827), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n7878), .B2(
        n9836), .ZN(n7806) );
  OAI211_X1 U9573 ( .C1(n7909), .C2(n9763), .A(n7807), .B(n7806), .ZN(n7808)
         );
  AOI21_X1 U9574 ( .B1(n9847), .B2(n7908), .A(n7808), .ZN(n7809) );
  OAI21_X1 U9575 ( .B1(n7810), .B2(n9827), .A(n7809), .ZN(P1_U3287) );
  AOI22_X1 U9576 ( .A1(n9210), .A2(n9487), .B1(n9192), .B2(n9485), .ZN(n7811)
         );
  NAND2_X1 U9577 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n10105) );
  OAI211_X1 U9578 ( .C1(n7812), .C2(n9213), .A(n7811), .B(n10105), .ZN(n7816)
         );
  AOI211_X1 U9579 ( .C1(n7814), .C2(n7813), .A(n9199), .B(n4545), .ZN(n7815)
         );
  AOI211_X1 U9580 ( .C1(n7817), .C2(n9197), .A(n7816), .B(n7815), .ZN(n7818)
         );
  INV_X1 U9581 ( .A(n7818), .ZN(P1_U3230) );
  XNOR2_X1 U9582 ( .A(n7819), .B(n7820), .ZN(n10240) );
  XNOR2_X1 U9583 ( .A(n7821), .B(n7820), .ZN(n7822) );
  AOI222_X1 U9584 ( .A1(n8829), .A2(n7822), .B1(n8494), .B2(n8826), .C1(n8496), 
        .C2(n8825), .ZN(n10241) );
  MUX2_X1 U9585 ( .A(n5164), .B(n10241), .S(n10221), .Z(n7826) );
  AOI22_X1 U9586 ( .A1(n8838), .A2(n7824), .B1(n8821), .B2(n7823), .ZN(n7825)
         );
  OAI211_X1 U9587 ( .C1(n8835), .C2(n10240), .A(n7826), .B(n7825), .ZN(
        P2_U3228) );
  INV_X1 U9588 ( .A(n7827), .ZN(n8109) );
  INV_X1 U9589 ( .A(n7828), .ZN(n7829) );
  AOI21_X1 U9590 ( .B1(n8109), .B2(n7830), .A(n7829), .ZN(n7835) );
  AOI22_X1 U9591 ( .A1(n9827), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n9836), .ZN(n7831) );
  OAI21_X1 U9592 ( .B1(n9840), .B2(n7832), .A(n7831), .ZN(n7833) );
  AOI21_X1 U9593 ( .B1(n9837), .B2(n9072), .A(n7833), .ZN(n7834) );
  OAI21_X1 U9594 ( .B1(n7835), .B2(n9827), .A(n7834), .ZN(P1_U3292) );
  OAI211_X1 U9595 ( .C1(n7885), .C2(n9943), .A(n7837), .B(n7836), .ZN(n7838)
         );
  AOI21_X1 U9596 ( .B1(n9959), .B2(n7839), .A(n7838), .ZN(n7844) );
  OAI22_X1 U9597 ( .A1(n10016), .A2(n7840), .B1(n10161), .B2(n5559), .ZN(n7841) );
  INV_X1 U9598 ( .A(n7841), .ZN(n7842) );
  OAI21_X1 U9599 ( .B1(n7844), .B2(n10160), .A(n7842), .ZN(P1_U3468) );
  AOI22_X1 U9600 ( .A1(n9856), .A2(n7888), .B1(n10162), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n7843) );
  OAI21_X1 U9601 ( .B1(n7844), .B2(n10162), .A(n7843), .ZN(P1_U3527) );
  INV_X1 U9602 ( .A(n7845), .ZN(n7855) );
  AOI22_X1 U9603 ( .A1(n9827), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9836), .B2(
        n7846), .ZN(n7847) );
  OAI21_X1 U9604 ( .B1(n9763), .B2(n7848), .A(n7847), .ZN(n7852) );
  OAI22_X1 U9605 ( .A1(n7850), .A2(n9840), .B1(n7849), .B2(n9829), .ZN(n7851)
         );
  AOI211_X1 U9606 ( .C1(n7853), .C2(n9847), .A(n7852), .B(n7851), .ZN(n7854)
         );
  OAI21_X1 U9607 ( .B1(n7855), .B2(n9827), .A(n7854), .ZN(P1_U3290) );
  INV_X1 U9608 ( .A(n7856), .ZN(n8318) );
  OAI222_X1 U9609 ( .A1(n8991), .A2(n7858), .B1(n4411), .B2(n8318), .C1(n7857), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  XNOR2_X1 U9610 ( .A(n8194), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n7860) );
  AOI211_X1 U9611 ( .C1(n7861), .C2(n7860), .A(n10137), .B(n8190), .ZN(n7870)
         );
  XNOR2_X1 U9612 ( .A(n8194), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n7864) );
  AOI211_X1 U9613 ( .C1(n7865), .C2(n7864), .A(n10141), .B(n8193), .ZN(n7869)
         );
  INV_X1 U9614 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7867) );
  NAND2_X1 U9615 ( .A1(n10146), .A2(n8194), .ZN(n7866) );
  NAND2_X1 U9616 ( .A1(n4401), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9181) );
  OAI211_X1 U9617 ( .C1(n7867), .C2(n10148), .A(n7866), .B(n9181), .ZN(n7868)
         );
  OR3_X1 U9618 ( .A1(n7870), .A2(n7869), .A3(n7868), .ZN(P1_U3254) );
  XNOR2_X1 U9619 ( .A(n7872), .B(n7871), .ZN(n7873) );
  XNOR2_X1 U9620 ( .A(n7874), .B(n7873), .ZN(n7880) );
  AOI22_X1 U9621 ( .A1(n9210), .A2(n9485), .B1(n9192), .B2(n9483), .ZN(n7876)
         );
  OAI211_X1 U9622 ( .C1(n7909), .C2(n9213), .A(n7876), .B(n7875), .ZN(n7877)
         );
  AOI21_X1 U9623 ( .B1(n7878), .B2(n9197), .A(n7877), .ZN(n7879) );
  OAI21_X1 U9624 ( .B1(n7880), .B2(n9199), .A(n7879), .ZN(P1_U3239) );
  NOR2_X1 U9625 ( .A1(n7881), .A2(n4542), .ZN(n7883) );
  XNOR2_X1 U9626 ( .A(n7883), .B(n7882), .ZN(n7892) );
  INV_X1 U9627 ( .A(n7884), .ZN(n7887) );
  OAI22_X1 U9628 ( .A1(n9207), .A2(n7897), .B1(n7885), .B2(n9194), .ZN(n7886)
         );
  AOI211_X1 U9629 ( .C1(n7888), .C2(n9171), .A(n7887), .B(n7886), .ZN(n7891)
         );
  NAND2_X1 U9630 ( .A1(n9197), .A2(n7889), .ZN(n7890) );
  OAI211_X1 U9631 ( .C1(n7892), .C2(n9199), .A(n7891), .B(n7890), .ZN(P1_U3227) );
  NOR2_X1 U9632 ( .A1(n7894), .A2(n7893), .ZN(n7895) );
  INV_X1 U9633 ( .A(n8043), .ZN(n9235) );
  XNOR2_X1 U9634 ( .A(n7895), .B(n9235), .ZN(n7975) );
  OAI211_X1 U9635 ( .C1(n7896), .C2(n8058), .A(n8112), .B(n9784), .ZN(n7971)
         );
  OAI21_X1 U9636 ( .B1(n7897), .B2(n9943), .A(n7971), .ZN(n7900) );
  NAND2_X1 U9637 ( .A1(n7898), .A2(n9230), .ZN(n8044) );
  XNOR2_X1 U9638 ( .A(n8044), .B(n9235), .ZN(n7899) );
  OAI22_X1 U9639 ( .A1(n7899), .A2(n9817), .B1(n9142), .B2(n9815), .ZN(n7972)
         );
  AOI211_X1 U9640 ( .C1(n9959), .C2(n7975), .A(n7900), .B(n7972), .ZN(n7905)
         );
  INV_X1 U9641 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7901) );
  OAI22_X1 U9642 ( .A1(n10016), .A2(n8058), .B1(n10161), .B2(n7901), .ZN(n7902) );
  INV_X1 U9643 ( .A(n7902), .ZN(n7903) );
  OAI21_X1 U9644 ( .B1(n7905), .B2(n10160), .A(n7903), .ZN(P1_U3474) );
  AOI22_X1 U9645 ( .A1(n9856), .A2(n7968), .B1(n10162), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7904) );
  OAI21_X1 U9646 ( .B1(n7905), .B2(n10162), .A(n7904), .ZN(P1_U3529) );
  AOI211_X1 U9647 ( .C1(n9959), .C2(n7908), .A(n7907), .B(n7906), .ZN(n7914)
         );
  OAI22_X1 U9648 ( .A1(n10016), .A2(n7909), .B1(n10161), .B2(n5411), .ZN(n7910) );
  INV_X1 U9649 ( .A(n7910), .ZN(n7911) );
  OAI21_X1 U9650 ( .B1(n7914), .B2(n10160), .A(n7911), .ZN(P1_U3471) );
  AOI22_X1 U9651 ( .A1(n9856), .A2(n7912), .B1(n10162), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n7913) );
  OAI21_X1 U9652 ( .B1(n7914), .B2(n10162), .A(n7913), .ZN(P1_U3528) );
  OR2_X1 U9653 ( .A1(n7819), .A2(n7915), .ZN(n7917) );
  NAND2_X1 U9654 ( .A1(n7917), .A2(n7916), .ZN(n7918) );
  XOR2_X1 U9655 ( .A(n7919), .B(n7918), .Z(n7938) );
  XOR2_X1 U9656 ( .A(n7920), .B(n7919), .Z(n7921) );
  AOI222_X1 U9657 ( .A1(n8829), .A2(n7921), .B1(n8493), .B2(n8826), .C1(n8495), 
        .C2(n8825), .ZN(n7937) );
  MUX2_X1 U9658 ( .A(n7922), .B(n7937), .S(n10221), .Z(n7925) );
  AOI22_X1 U9659 ( .A1(n8838), .A2(n8064), .B1(n8821), .B2(n7923), .ZN(n7924)
         );
  OAI211_X1 U9660 ( .C1(n7938), .C2(n8835), .A(n7925), .B(n7924), .ZN(P2_U3227) );
  AOI21_X1 U9661 ( .B1(n8441), .B2(n8494), .A(n7926), .ZN(n7928) );
  NAND2_X1 U9662 ( .A1(n8478), .A2(n8032), .ZN(n7927) );
  OAI211_X1 U9663 ( .C1(n8142), .C2(n8454), .A(n7928), .B(n7927), .ZN(n7934)
         );
  NAND2_X1 U9664 ( .A1(n7930), .A2(n7929), .ZN(n7931) );
  AOI21_X1 U9665 ( .B1(n7932), .B2(n7931), .A(n8460), .ZN(n7933) );
  AOI211_X1 U9666 ( .C1(n8033), .C2(n8457), .A(n7934), .B(n7933), .ZN(n7935)
         );
  INV_X1 U9667 ( .A(n7935), .ZN(P2_U3153) );
  INV_X1 U9668 ( .A(n6451), .ZN(n7961) );
  OAI222_X1 U9669 ( .A1(n4411), .A2(n7961), .B1(n8991), .B2(n6452), .C1(
        P2_U3151), .C2(n7936), .ZN(P2_U3275) );
  INV_X1 U9670 ( .A(n10245), .ZN(n8897) );
  OAI21_X1 U9671 ( .B1(n8897), .B2(n7938), .A(n7937), .ZN(n8063) );
  INV_X1 U9672 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7939) );
  OAI22_X1 U9673 ( .A1(n8957), .A2(n7940), .B1(n7939), .B2(n10247), .ZN(n7941)
         );
  AOI21_X1 U9674 ( .B1(n8063), .B2(n10247), .A(n7941), .ZN(n7942) );
  INV_X1 U9675 ( .A(n7942), .ZN(P2_U3408) );
  OR2_X1 U9676 ( .A1(n7819), .A2(n7944), .ZN(n7946) );
  AND2_X1 U9677 ( .A1(n7946), .A2(n7945), .ZN(n7947) );
  NAND2_X1 U9678 ( .A1(n7947), .A2(n7950), .ZN(n7948) );
  NAND2_X1 U9679 ( .A1(n7943), .A2(n7948), .ZN(n8036) );
  INV_X1 U9680 ( .A(n8036), .ZN(n7954) );
  XNOR2_X1 U9681 ( .A(n7949), .B(n7950), .ZN(n7951) );
  NAND2_X1 U9682 ( .A1(n7951), .A2(n8829), .ZN(n7953) );
  AOI22_X1 U9683 ( .A1(n8826), .A2(n8492), .B1(n8494), .B2(n8825), .ZN(n7952)
         );
  OAI211_X1 U9684 ( .C1(n8036), .C2(n8177), .A(n7953), .B(n7952), .ZN(n8030)
         );
  AOI21_X1 U9685 ( .B1(n10228), .B2(n7954), .A(n8030), .ZN(n7960) );
  AOI22_X1 U9686 ( .A1(n6778), .A2(n8033), .B1(P2_REG0_REG_7__SCAN_IN), .B2(
        n10249), .ZN(n7955) );
  OAI21_X1 U9687 ( .B1(n7960), .B2(n10249), .A(n7955), .ZN(P2_U3411) );
  INV_X1 U9688 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7956) );
  OAI22_X1 U9689 ( .A1(n8884), .A2(n7957), .B1(n10259), .B2(n7956), .ZN(n7958)
         );
  INV_X1 U9690 ( .A(n7958), .ZN(n7959) );
  OAI21_X1 U9691 ( .B1(n7960), .B2(n10257), .A(n7959), .ZN(P2_U3466) );
  OAI222_X1 U9692 ( .A1(n10037), .A2(n7962), .B1(n10040), .B2(n7961), .C1(
        n9455), .C2(n4401), .ZN(P1_U3335) );
  INV_X1 U9693 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7963) );
  OAI22_X1 U9694 ( .A1(n8884), .A2(n7964), .B1(n10259), .B2(n7963), .ZN(n7965)
         );
  INV_X1 U9695 ( .A(n7965), .ZN(n7966) );
  OAI21_X1 U9696 ( .B1(n7967), .B2(n10257), .A(n7966), .ZN(P2_U3460) );
  AOI22_X1 U9697 ( .A1(n9837), .A2(n7968), .B1(n9836), .B2(n8060), .ZN(n7970)
         );
  NAND2_X1 U9698 ( .A1(n9681), .A2(n9484), .ZN(n7969) );
  OAI211_X1 U9699 ( .C1(n7971), .C2(n9840), .A(n7970), .B(n7969), .ZN(n7974)
         );
  MUX2_X1 U9700 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n7972), .S(n9842), .Z(n7973)
         );
  AOI211_X1 U9701 ( .C1(n9847), .C2(n7975), .A(n7974), .B(n7973), .ZN(n7976)
         );
  INV_X1 U9702 ( .A(n7976), .ZN(P1_U3286) );
  XOR2_X1 U9703 ( .A(n7977), .B(n7978), .Z(n7991) );
  XNOR2_X1 U9704 ( .A(n7980), .B(n7979), .ZN(n7989) );
  NAND2_X1 U9705 ( .A1(n10170), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7981) );
  NAND2_X1 U9706 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8355) );
  OAI211_X1 U9707 ( .C1(n10298), .C2(n7982), .A(n7981), .B(n8355), .ZN(n7988)
         );
  OR3_X1 U9708 ( .A1(n7997), .A2(n7984), .A3(n7983), .ZN(n7985) );
  AOI21_X1 U9709 ( .B1(n7986), .B2(n7985), .A(n10176), .ZN(n7987) );
  AOI211_X1 U9710 ( .C1(n10288), .C2(n7989), .A(n7988), .B(n7987), .ZN(n7990)
         );
  OAI21_X1 U9711 ( .B1(n7991), .B2(n10197), .A(n7990), .ZN(P2_U3192) );
  XNOR2_X1 U9712 ( .A(n7992), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n8005) );
  XNOR2_X1 U9713 ( .A(n7994), .B(n7993), .ZN(n8003) );
  NAND2_X1 U9714 ( .A1(n10170), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7995) );
  NAND2_X1 U9715 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8219) );
  OAI211_X1 U9716 ( .C1(n10298), .C2(n7996), .A(n7995), .B(n8219), .ZN(n8002)
         );
  AOI21_X1 U9717 ( .B1(n7999), .B2(n7998), .A(n7997), .ZN(n8000) );
  NOR2_X1 U9718 ( .A1(n8000), .A2(n10176), .ZN(n8001) );
  AOI211_X1 U9719 ( .C1(n10288), .C2(n8003), .A(n8002), .B(n8001), .ZN(n8004)
         );
  OAI21_X1 U9720 ( .B1(n8005), .B2(n10197), .A(n8004), .ZN(P2_U3191) );
  NAND2_X1 U9721 ( .A1(n7943), .A2(n8006), .ZN(n8007) );
  XNOR2_X1 U9722 ( .A(n8007), .B(n8008), .ZN(n8271) );
  AOI21_X1 U9723 ( .B1(n8009), .B2(n8008), .A(n10218), .ZN(n8010) );
  OR2_X1 U9724 ( .A1(n8009), .A2(n8008), .ZN(n8131) );
  NAND2_X1 U9725 ( .A1(n8010), .A2(n8131), .ZN(n8012) );
  AOI22_X1 U9726 ( .A1(n8491), .A2(n8826), .B1(n8825), .B2(n8493), .ZN(n8011)
         );
  NAND2_X1 U9727 ( .A1(n8012), .A2(n8011), .ZN(n8267) );
  NAND2_X1 U9728 ( .A1(n8267), .A2(n10247), .ZN(n8014) );
  AOI22_X1 U9729 ( .A1(n6778), .A2(n8269), .B1(P2_REG0_REG_8__SCAN_IN), .B2(
        n10249), .ZN(n8013) );
  OAI211_X1 U9730 ( .C1(n8271), .C2(n8967), .A(n8014), .B(n8013), .ZN(P2_U3414) );
  INV_X1 U9731 ( .A(n8015), .ZN(n8017) );
  AOI21_X1 U9732 ( .B1(n9359), .B2(n9357), .A(n9437), .ZN(n8016) );
  OAI21_X1 U9733 ( .B1(n8017), .B2(n8016), .A(n9782), .ZN(n8018) );
  OAI21_X1 U9734 ( .B1(n9091), .B2(n9815), .A(n8018), .ZN(n8092) );
  INV_X1 U9735 ( .A(n8092), .ZN(n8029) );
  OAI21_X1 U9736 ( .B1(n8021), .B2(n8020), .A(n8019), .ZN(n8094) );
  INV_X1 U9737 ( .A(n8022), .ZN(n8073) );
  OAI211_X1 U9738 ( .C1(n9018), .C2(n8023), .A(n8073), .B(n9784), .ZN(n8091)
         );
  AOI22_X1 U9739 ( .A1(n9827), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n9021), .B2(
        n9836), .ZN(n8024) );
  OAI21_X1 U9740 ( .B1(n9063), .B2(n9829), .A(n8024), .ZN(n8025) );
  AOI21_X1 U9741 ( .B1(n9837), .B2(n8097), .A(n8025), .ZN(n8026) );
  OAI21_X1 U9742 ( .B1(n8091), .B2(n9840), .A(n8026), .ZN(n8027) );
  AOI21_X1 U9743 ( .B1(n9847), .B2(n8094), .A(n8027), .ZN(n8028) );
  OAI21_X1 U9744 ( .B1(n8029), .B2(n9827), .A(n8028), .ZN(P1_U3283) );
  NAND2_X1 U9745 ( .A1(n10221), .A2(n10220), .ZN(n8634) );
  MUX2_X1 U9746 ( .A(n8030), .B(P2_REG2_REG_7__SCAN_IN), .S(n10223), .Z(n8031)
         );
  INV_X1 U9747 ( .A(n8031), .ZN(n8035) );
  AOI22_X1 U9748 ( .A1(n8838), .A2(n8033), .B1(n8821), .B2(n8032), .ZN(n8034)
         );
  OAI211_X1 U9749 ( .C1(n8036), .C2(n8634), .A(n8035), .B(n8034), .ZN(P2_U3226) );
  NAND2_X1 U9750 ( .A1(n8606), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8037) );
  OAI21_X1 U9751 ( .B1(n8638), .B2(n8606), .A(n8037), .ZN(P2_U3520) );
  OAI21_X1 U9752 ( .B1(n8039), .B2(n8047), .A(n8038), .ZN(n9846) );
  INV_X1 U9753 ( .A(n9838), .ZN(n8041) );
  XOR2_X1 U9754 ( .A(n8110), .B(n9838), .Z(n8040) );
  AOI22_X1 U9755 ( .A1(n8040), .A2(n9784), .B1(n9804), .B2(n9481), .ZN(n9841)
         );
  OAI21_X1 U9756 ( .B1(n8041), .B2(n9950), .A(n9841), .ZN(n8049) );
  OAI21_X1 U9757 ( .B1(n8044), .B2(n8043), .A(n8042), .ZN(n8103) );
  OAI21_X1 U9758 ( .B1(n8103), .B2(n8102), .A(n8045), .ZN(n8046) );
  XOR2_X1 U9759 ( .A(n8047), .B(n8046), .Z(n8048) );
  OAI22_X1 U9760 ( .A1(n8048), .A2(n9817), .B1(n9142), .B2(n9943), .ZN(n9843)
         );
  AOI211_X1 U9761 ( .C1(n9959), .C2(n9846), .A(n8049), .B(n9843), .ZN(n8052)
         );
  NAND2_X1 U9762 ( .A1(n10160), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8050) );
  OAI21_X1 U9763 ( .B1(n8052), .B2(n10160), .A(n8050), .ZN(P1_U3480) );
  NAND2_X1 U9764 ( .A1(n10162), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n8051) );
  OAI21_X1 U9765 ( .B1(n8052), .B2(n10162), .A(n8051), .ZN(P1_U3531) );
  NAND2_X1 U9766 ( .A1(n4555), .A2(n8053), .ZN(n8054) );
  XNOR2_X1 U9767 ( .A(n8055), .B(n8054), .ZN(n8062) );
  AOI22_X1 U9768 ( .A1(n9210), .A2(n9484), .B1(n9192), .B2(n5051), .ZN(n8057)
         );
  OAI211_X1 U9769 ( .C1(n8058), .C2(n9213), .A(n8057), .B(n8056), .ZN(n8059)
         );
  AOI21_X1 U9770 ( .B1(n8060), .B2(n9197), .A(n8059), .ZN(n8061) );
  OAI21_X1 U9771 ( .B1(n8062), .B2(n9199), .A(n8061), .ZN(P1_U3213) );
  INV_X1 U9772 ( .A(n8063), .ZN(n8066) );
  AOI22_X1 U9773 ( .A1(n8888), .A2(n8064), .B1(n10257), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n8065) );
  OAI21_X1 U9774 ( .B1(n8066), .B2(n10257), .A(n8065), .ZN(P2_U3465) );
  OAI211_X1 U9775 ( .C1(n4540), .C2(n4940), .A(n9782), .B(n8149), .ZN(n8068)
         );
  AOI22_X1 U9776 ( .A1(n9877), .A2(n9481), .B1(n9479), .B2(n9804), .ZN(n8067)
         );
  NAND2_X1 U9777 ( .A1(n8068), .A2(n8067), .ZN(n9957) );
  INV_X1 U9778 ( .A(n9957), .ZN(n8079) );
  OAI21_X1 U9779 ( .B1(n8071), .B2(n8070), .A(n8069), .ZN(n9958) );
  INV_X1 U9780 ( .A(n8072), .ZN(n8155) );
  AOI211_X1 U9781 ( .C1(n8074), .C2(n8073), .A(n9822), .B(n8155), .ZN(n9956)
         );
  NAND2_X1 U9782 ( .A1(n9956), .A2(n9807), .ZN(n8076) );
  AOI22_X1 U9783 ( .A1(n9827), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9186), .B2(
        n9836), .ZN(n8075) );
  OAI211_X1 U9784 ( .C1(n10017), .C2(n9763), .A(n8076), .B(n8075), .ZN(n8077)
         );
  AOI21_X1 U9785 ( .B1(n9847), .B2(n9958), .A(n8077), .ZN(n8078) );
  OAI21_X1 U9786 ( .B1(n9827), .B2(n8079), .A(n8078), .ZN(P1_U3282) );
  INV_X1 U9787 ( .A(n8080), .ZN(n8089) );
  OAI222_X1 U9788 ( .A1(n4411), .A2(n8089), .B1(P2_U3151), .B2(n8082), .C1(
        n8081), .C2(n8991), .ZN(P2_U3274) );
  INV_X1 U9789 ( .A(n8083), .ZN(n8086) );
  OAI222_X1 U9790 ( .A1(n10037), .A2(n8084), .B1(n10040), .B2(n8086), .C1(
        P1_U3086), .C2(n9465), .ZN(P1_U3333) );
  OAI222_X1 U9791 ( .A1(n8991), .A2(n8087), .B1(n4411), .B2(n8086), .C1(n8085), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  OAI222_X1 U9792 ( .A1(n10037), .A2(n8090), .B1(n10040), .B2(n8089), .C1(
        n8088), .C2(P1_U3086), .ZN(P1_U3334) );
  OAI21_X1 U9793 ( .B1(n9063), .B2(n9943), .A(n8091), .ZN(n8093) );
  AOI211_X1 U9794 ( .C1(n9959), .C2(n8094), .A(n8093), .B(n8092), .ZN(n8099)
         );
  AOI22_X1 U9795 ( .A1(n8097), .A2(n9856), .B1(P1_REG1_REG_10__SCAN_IN), .B2(
        n10162), .ZN(n8095) );
  OAI21_X1 U9796 ( .B1(n8099), .B2(n10162), .A(n8095), .ZN(P1_U3532) );
  INV_X1 U9797 ( .A(n10016), .ZN(n8096) );
  AOI22_X1 U9798 ( .A1(n8097), .A2(n8096), .B1(P1_REG0_REG_10__SCAN_IN), .B2(
        n10160), .ZN(n8098) );
  OAI21_X1 U9799 ( .B1(n8099), .B2(n10160), .A(n8098), .ZN(P1_U3483) );
  OAI22_X1 U9800 ( .A1(n8101), .A2(n9943), .B1(n9063), .B2(n9815), .ZN(n8106)
         );
  XNOR2_X1 U9801 ( .A(n8103), .B(n8102), .ZN(n8104) );
  NOR2_X1 U9802 ( .A1(n8104), .A2(n9817), .ZN(n8105) );
  AOI211_X1 U9803 ( .C1(n8107), .C2(n9963), .A(n8106), .B(n8105), .ZN(n9967)
         );
  INV_X1 U9804 ( .A(n9967), .ZN(n8108) );
  AOI21_X1 U9805 ( .B1(n8109), .B2(n9963), .A(n8108), .ZN(n8116) );
  INV_X1 U9806 ( .A(n8110), .ZN(n8111) );
  AOI211_X1 U9807 ( .C1(n9965), .C2(n8112), .A(n9822), .B(n8111), .ZN(n9964)
         );
  AOI22_X1 U9808 ( .A1(n9827), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n9059), .B2(
        n9836), .ZN(n8113) );
  OAI21_X1 U9809 ( .B1(n9763), .B2(n5052), .A(n8113), .ZN(n8114) );
  AOI21_X1 U9810 ( .B1(n9964), .B2(n9807), .A(n8114), .ZN(n8115) );
  OAI21_X1 U9811 ( .B1(n8116), .B2(n9827), .A(n8115), .ZN(P1_U3285) );
  NAND2_X1 U9812 ( .A1(n4553), .A2(n8117), .ZN(n8118) );
  XNOR2_X1 U9813 ( .A(n8119), .B(n8118), .ZN(n8125) );
  INV_X1 U9814 ( .A(n8120), .ZN(n8830) );
  NAND2_X1 U9815 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8518) );
  OAI21_X1 U9816 ( .B1(n8476), .B2(n8357), .A(n8518), .ZN(n8121) );
  AOI21_X1 U9817 ( .B1(n8473), .B2(n8827), .A(n8121), .ZN(n8122) );
  OAI21_X1 U9818 ( .B1(n8830), .B2(n8431), .A(n8122), .ZN(n8123) );
  AOI21_X1 U9819 ( .B1(n8893), .B2(n8457), .A(n8123), .ZN(n8124) );
  OAI21_X1 U9820 ( .B1(n8125), .B2(n8460), .A(n8124), .ZN(P2_U3164) );
  INV_X1 U9821 ( .A(n8128), .ZN(n8126) );
  NAND2_X1 U9822 ( .A1(n8126), .A2(n8132), .ZN(n8175) );
  INV_X1 U9823 ( .A(n8132), .ZN(n8127) );
  NAND2_X1 U9824 ( .A1(n8128), .A2(n8127), .ZN(n8129) );
  NAND2_X1 U9825 ( .A1(n8175), .A2(n8129), .ZN(n8259) );
  NAND2_X1 U9826 ( .A1(n8131), .A2(n8130), .ZN(n8133) );
  XNOR2_X1 U9827 ( .A(n8133), .B(n8132), .ZN(n8134) );
  NAND2_X1 U9828 ( .A1(n8134), .A2(n8829), .ZN(n8136) );
  AOI22_X1 U9829 ( .A1(n8826), .A2(n8490), .B1(n8492), .B2(n8825), .ZN(n8135)
         );
  OAI211_X1 U9830 ( .C1(n8259), .C2(n8177), .A(n8136), .B(n8135), .ZN(n8255)
         );
  INV_X1 U9831 ( .A(n8257), .ZN(n8224) );
  OAI22_X1 U9832 ( .A1(n8259), .A2(n8137), .B1(n8224), .B2(n10242), .ZN(n8138)
         );
  NOR2_X1 U9833 ( .A1(n8255), .A2(n8138), .ZN(n8210) );
  NAND2_X1 U9834 ( .A1(n10249), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8139) );
  OAI21_X1 U9835 ( .B1(n8210), .B2(n10249), .A(n8139), .ZN(P2_U3417) );
  INV_X1 U9836 ( .A(n8269), .ZN(n8252) );
  INV_X1 U9837 ( .A(n8212), .ZN(n8140) );
  XNOR2_X1 U9838 ( .A(n8213), .B(n8140), .ZN(n8141) );
  NAND2_X1 U9839 ( .A1(n8141), .A2(n8142), .ZN(n8215) );
  OAI21_X1 U9840 ( .B1(n8142), .B2(n8141), .A(n8215), .ZN(n8143) );
  NAND2_X1 U9841 ( .A1(n8143), .A2(n8470), .ZN(n8148) );
  NAND2_X1 U9842 ( .A1(n8441), .A2(n8493), .ZN(n8145) );
  OAI211_X1 U9843 ( .C1(n8180), .C2(n8454), .A(n8145), .B(n8144), .ZN(n8146)
         );
  AOI21_X1 U9844 ( .B1(n8268), .B2(n8478), .A(n8146), .ZN(n8147) );
  OAI211_X1 U9845 ( .C1(n8252), .C2(n8481), .A(n8148), .B(n8147), .ZN(P2_U3161) );
  NAND2_X1 U9846 ( .A1(n8149), .A2(n9256), .ZN(n8150) );
  XOR2_X1 U9847 ( .A(n9439), .B(n8150), .Z(n8151) );
  OAI222_X1 U9848 ( .A1(n9815), .A2(n9934), .B1(n9943), .B2(n9091), .C1(n9817), 
        .C2(n8151), .ZN(n9952) );
  INV_X1 U9849 ( .A(n9952), .ZN(n8160) );
  OAI21_X1 U9850 ( .B1(n8153), .B2(n9439), .A(n8152), .ZN(n9954) );
  INV_X1 U9851 ( .A(n9093), .ZN(n9951) );
  OAI211_X1 U9852 ( .C1(n8155), .C2(n9951), .A(n9784), .B(n9823), .ZN(n9949)
         );
  AOI22_X1 U9853 ( .A1(n9827), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n9088), .B2(
        n9836), .ZN(n8157) );
  NAND2_X1 U9854 ( .A1(n9093), .A2(n9837), .ZN(n8156) );
  OAI211_X1 U9855 ( .C1(n9949), .C2(n9840), .A(n8157), .B(n8156), .ZN(n8158)
         );
  AOI21_X1 U9856 ( .B1(n9954), .B2(n9847), .A(n8158), .ZN(n8159) );
  OAI21_X1 U9857 ( .B1(n8160), .B2(n9827), .A(n8159), .ZN(P1_U3281) );
  NAND2_X1 U9858 ( .A1(n8165), .A2(n8976), .ZN(n8162) );
  OAI211_X1 U9859 ( .C1(n8163), .C2(n8991), .A(n8162), .B(n8161), .ZN(P2_U3272) );
  NAND2_X1 U9860 ( .A1(n8165), .A2(n8164), .ZN(n8166) );
  OAI211_X1 U9861 ( .C1(n5995), .C2(n10037), .A(n8166), .B(n9456), .ZN(
        P1_U3332) );
  INV_X1 U9862 ( .A(n8964), .ZN(n8818) );
  OAI211_X1 U9863 ( .C1(n8169), .C2(n8168), .A(n8167), .B(n8470), .ZN(n8173)
         );
  NOR2_X1 U9864 ( .A1(n10583), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8533) );
  AOI21_X1 U9865 ( .B1(n8473), .B2(n8816), .A(n8533), .ZN(n8170) );
  OAI21_X1 U9866 ( .B1(n8476), .B2(n8444), .A(n8170), .ZN(n8171) );
  AOI21_X1 U9867 ( .B1(n8820), .B2(n8478), .A(n8171), .ZN(n8172) );
  OAI211_X1 U9868 ( .C1(n8818), .C2(n8481), .A(n8173), .B(n8172), .ZN(P2_U3174) );
  INV_X1 U9869 ( .A(n8360), .ZN(n8189) );
  INV_X1 U9870 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n8185) );
  NAND2_X1 U9871 ( .A1(n8175), .A2(n8174), .ZN(n8228) );
  INV_X1 U9872 ( .A(n8179), .ZN(n8176) );
  XNOR2_X1 U9873 ( .A(n8228), .B(n8176), .ZN(n8204) );
  INV_X1 U9874 ( .A(n8177), .ZN(n10215) );
  NAND2_X1 U9875 ( .A1(n8204), .A2(n10215), .ZN(n8184) );
  XNOR2_X1 U9876 ( .A(n8178), .B(n8179), .ZN(n8182) );
  OAI22_X1 U9877 ( .A1(n8180), .A2(n10211), .B1(n8357), .B2(n10212), .ZN(n8181) );
  AOI21_X1 U9878 ( .B1(n8182), .B2(n8829), .A(n8181), .ZN(n8183) );
  NAND2_X1 U9879 ( .A1(n8184), .A2(n8183), .ZN(n8205) );
  AOI21_X1 U9880 ( .B1(n10228), .B2(n8204), .A(n8205), .ZN(n8187) );
  MUX2_X1 U9881 ( .A(n8185), .B(n8187), .S(n10247), .Z(n8186) );
  OAI21_X1 U9882 ( .B1(n8189), .B2(n8957), .A(n8186), .ZN(P2_U3420) );
  MUX2_X1 U9883 ( .A(n5228), .B(n8187), .S(n10259), .Z(n8188) );
  OAI21_X1 U9884 ( .B1(n8189), .B2(n8884), .A(n8188), .ZN(P2_U3469) );
  XNOR2_X1 U9885 ( .A(n9521), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n8192) );
  XNOR2_X1 U9886 ( .A(n8195), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n9508) );
  AOI211_X1 U9887 ( .C1(n8192), .C2(n8191), .A(n10137), .B(n9517), .ZN(n8203)
         );
  XNOR2_X1 U9888 ( .A(n9521), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n8198) );
  MUX2_X1 U9889 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n5716), .S(n8195), .Z(n8196)
         );
  INV_X1 U9890 ( .A(n8196), .ZN(n9503) );
  AOI211_X1 U9891 ( .C1(n8198), .C2(n8197), .A(n10141), .B(n9520), .ZN(n8202)
         );
  INV_X1 U9892 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n8200) );
  NAND2_X1 U9893 ( .A1(n10146), .A2(n9521), .ZN(n8199) );
  NAND2_X1 U9894 ( .A1(n4401), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9158) );
  OAI211_X1 U9895 ( .C1(n8200), .C2(n10148), .A(n8199), .B(n9158), .ZN(n8201)
         );
  OR3_X1 U9896 ( .A1(n8203), .A2(n8202), .A3(n8201), .ZN(P1_U3256) );
  INV_X1 U9897 ( .A(n8204), .ZN(n8209) );
  MUX2_X1 U9898 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n8205), .S(n10221), .Z(n8206) );
  INV_X1 U9899 ( .A(n8206), .ZN(n8208) );
  AOI22_X1 U9900 ( .A1(n8360), .A2(n8838), .B1(n8821), .B2(n8359), .ZN(n8207)
         );
  OAI211_X1 U9901 ( .C1(n8209), .C2(n8634), .A(n8208), .B(n8207), .ZN(P2_U3223) );
  MUX2_X1 U9902 ( .A(n8210), .B(n10438), .S(n10257), .Z(n8211) );
  INV_X1 U9903 ( .A(n8211), .ZN(P2_U3468) );
  NAND2_X1 U9904 ( .A1(n8213), .A2(n8212), .ZN(n8214) );
  AND2_X1 U9905 ( .A1(n8215), .A2(n8214), .ZN(n8218) );
  INV_X1 U9906 ( .A(n8216), .ZN(n8217) );
  NAND2_X1 U9907 ( .A1(n8218), .A2(n8217), .ZN(n8350) );
  OAI211_X1 U9908 ( .C1(n8218), .C2(n8217), .A(n8350), .B(n8470), .ZN(n8223)
         );
  NAND2_X1 U9909 ( .A1(n8441), .A2(n8492), .ZN(n8220) );
  OAI211_X1 U9910 ( .C1(n8351), .C2(n8454), .A(n8220), .B(n8219), .ZN(n8221)
         );
  AOI21_X1 U9911 ( .B1(n8256), .B2(n8478), .A(n8221), .ZN(n8222) );
  OAI211_X1 U9912 ( .C1(n8224), .C2(n8481), .A(n8223), .B(n8222), .ZN(P2_U3171) );
  INV_X1 U9913 ( .A(n8225), .ZN(n8227) );
  OAI21_X1 U9914 ( .B1(n8228), .B2(n8227), .A(n8226), .ZN(n8230) );
  XNOR2_X1 U9915 ( .A(n8230), .B(n8229), .ZN(n8264) );
  OAI22_X1 U9916 ( .A1(n8264), .A2(n8967), .B1(n4719), .B2(n8957), .ZN(n8240)
         );
  NAND2_X1 U9917 ( .A1(n8232), .A2(n8233), .ZN(n8235) );
  NAND2_X1 U9918 ( .A1(n8235), .A2(n8234), .ZN(n8236) );
  NAND3_X1 U9919 ( .A1(n8231), .A2(n8829), .A3(n8236), .ZN(n8238) );
  AOI22_X1 U9920 ( .A1(n8825), .A2(n8490), .B1(n8815), .B2(n8826), .ZN(n8237)
         );
  NAND2_X1 U9921 ( .A1(n8238), .A2(n8237), .ZN(n8262) );
  MUX2_X1 U9922 ( .A(n8262), .B(P2_REG0_REG_11__SCAN_IN), .S(n10249), .Z(n8239) );
  OR2_X1 U9923 ( .A1(n8240), .A2(n8239), .ZN(P2_U3423) );
  OAI22_X1 U9924 ( .A1(n8264), .A2(n8891), .B1(n4719), .B2(n8884), .ZN(n8242)
         );
  MUX2_X1 U9925 ( .A(n8262), .B(P2_REG1_REG_11__SCAN_IN), .S(n10257), .Z(n8241) );
  OR2_X1 U9926 ( .A1(n8242), .A2(n8241), .ZN(P2_U3470) );
  AOI21_X1 U9927 ( .B1(n8245), .B2(n8244), .A(n8243), .ZN(n8251) );
  NAND2_X1 U9928 ( .A1(n8441), .A2(n8827), .ZN(n8246) );
  NAND2_X1 U9929 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8547) );
  OAI211_X1 U9930 ( .C1(n8771), .C2(n8454), .A(n8246), .B(n8547), .ZN(n8249)
         );
  INV_X1 U9931 ( .A(n8247), .ZN(n8958) );
  NOR2_X1 U9932 ( .A1(n8958), .A2(n8481), .ZN(n8248) );
  AOI211_X1 U9933 ( .C1(n8801), .C2(n8478), .A(n8249), .B(n8248), .ZN(n8250)
         );
  OAI21_X1 U9934 ( .B1(n8251), .B2(n8460), .A(n8250), .ZN(P2_U3155) );
  MUX2_X1 U9935 ( .A(n8267), .B(P2_REG1_REG_8__SCAN_IN), .S(n10257), .Z(n8254)
         );
  OAI22_X1 U9936 ( .A1(n8271), .A2(n8891), .B1(n8252), .B2(n8884), .ZN(n8253)
         );
  OR2_X1 U9937 ( .A1(n8254), .A2(n8253), .ZN(P2_U3467) );
  MUX2_X1 U9938 ( .A(n8255), .B(P2_REG2_REG_9__SCAN_IN), .S(n10223), .Z(n8261)
         );
  AOI22_X1 U9939 ( .A1(n8257), .A2(n8838), .B1(n8821), .B2(n8256), .ZN(n8258)
         );
  OAI21_X1 U9940 ( .B1(n8259), .B2(n8634), .A(n8258), .ZN(n8260) );
  OR2_X1 U9941 ( .A1(n8261), .A2(n8260), .ZN(P2_U3224) );
  MUX2_X1 U9942 ( .A(n8262), .B(P2_REG2_REG_11__SCAN_IN), .S(n10223), .Z(n8266) );
  AOI22_X1 U9943 ( .A1(n8447), .A2(n8838), .B1(n8821), .B2(n8446), .ZN(n8263)
         );
  OAI21_X1 U9944 ( .B1(n8264), .B2(n8835), .A(n8263), .ZN(n8265) );
  OR2_X1 U9945 ( .A1(n8266), .A2(n8265), .ZN(P2_U3222) );
  MUX2_X1 U9946 ( .A(n8267), .B(P2_REG2_REG_8__SCAN_IN), .S(n10223), .Z(n8273)
         );
  AOI22_X1 U9947 ( .A1(n8838), .A2(n8269), .B1(n8821), .B2(n8268), .ZN(n8270)
         );
  OAI21_X1 U9948 ( .B1(n8271), .B2(n8835), .A(n8270), .ZN(n8272) );
  OR2_X1 U9949 ( .A1(n8273), .A2(n8272), .ZN(P2_U3225) );
  NAND2_X1 U9950 ( .A1(n8275), .A2(n8274), .ZN(n8276) );
  XNOR2_X1 U9951 ( .A(n8276), .B(n5132), .ZN(n8277) );
  NAND2_X1 U9952 ( .A1(n8277), .A2(n9847), .ZN(n8285) );
  INV_X1 U9953 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8278) );
  OAI22_X1 U9954 ( .A1(n8279), .A2(n9785), .B1(n8278), .B2(n9842), .ZN(n8282)
         );
  NOR2_X1 U9955 ( .A1(n8280), .A2(n9840), .ZN(n8281) );
  AOI211_X1 U9956 ( .C1(n9837), .C2(n8283), .A(n8282), .B(n8281), .ZN(n8284)
         );
  OAI211_X1 U9957 ( .C1(n8286), .C2(n9827), .A(n8285), .B(n8284), .ZN(P1_U3356) );
  NAND2_X1 U9958 ( .A1(n8287), .A2(n8288), .ZN(n8701) );
  NAND2_X1 U9959 ( .A1(n8701), .A2(n5103), .ZN(n8857) );
  NAND2_X1 U9960 ( .A1(n8857), .A2(n8289), .ZN(n8290) );
  XOR2_X1 U9961 ( .A(n8292), .B(n8290), .Z(n8316) );
  XNOR2_X1 U9962 ( .A(n8291), .B(n8292), .ZN(n8293) );
  AOI222_X1 U9963 ( .A1(n8829), .A2(n8293), .B1(n8669), .B2(n8826), .C1(n8487), 
        .C2(n8825), .ZN(n8311) );
  MUX2_X1 U9964 ( .A(n8294), .B(n8311), .S(n10221), .Z(n8296) );
  AOI22_X1 U9965 ( .A1(n8313), .A2(n8838), .B1(n8821), .B2(n8302), .ZN(n8295)
         );
  OAI211_X1 U9966 ( .C1(n8316), .C2(n8835), .A(n8296), .B(n8295), .ZN(P2_U3210) );
  INV_X1 U9967 ( .A(n8298), .ZN(n8300) );
  INV_X1 U9968 ( .A(n8297), .ZN(n8299) );
  OR2_X1 U9969 ( .A1(n8298), .A2(n8297), .ZN(n8407) );
  OAI21_X1 U9970 ( .B1(n8300), .B2(n8299), .A(n8407), .ZN(n8301) );
  NOR2_X1 U9971 ( .A1(n8301), .A2(n8695), .ZN(n8410) );
  AOI21_X1 U9972 ( .B1(n8695), .B2(n8301), .A(n8410), .ZN(n8307) );
  AOI22_X1 U9973 ( .A1(n8487), .A2(n8441), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8304) );
  NAND2_X1 U9974 ( .A1(n8302), .A2(n8478), .ZN(n8303) );
  OAI211_X1 U9975 ( .C1(n8386), .C2(n8454), .A(n8304), .B(n8303), .ZN(n8305)
         );
  AOI21_X1 U9976 ( .B1(n8313), .B2(n8457), .A(n8305), .ZN(n8306) );
  OAI21_X1 U9977 ( .B1(n8307), .B2(n8460), .A(n8306), .ZN(P2_U3156) );
  INV_X1 U9978 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8308) );
  MUX2_X1 U9979 ( .A(n8308), .B(n8311), .S(n10247), .Z(n8310) );
  NAND2_X1 U9980 ( .A1(n8313), .A2(n6778), .ZN(n8309) );
  OAI211_X1 U9981 ( .C1(n8316), .C2(n8967), .A(n8310), .B(n8309), .ZN(P2_U3450) );
  INV_X1 U9982 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8312) );
  MUX2_X1 U9983 ( .A(n8312), .B(n8311), .S(n10254), .Z(n8315) );
  NAND2_X1 U9984 ( .A1(n8313), .A2(n8888), .ZN(n8314) );
  OAI211_X1 U9985 ( .C1(n8316), .C2(n8891), .A(n8315), .B(n8314), .ZN(P2_U3482) );
  INV_X1 U9986 ( .A(n9218), .ZN(n8320) );
  OAI222_X1 U9987 ( .A1(n8991), .A2(n10346), .B1(n4411), .B2(n8320), .C1(
        P2_U3151), .C2(n8317), .ZN(P2_U3265) );
  OAI222_X1 U9988 ( .A1(n10037), .A2(n8319), .B1(n10040), .B2(n8318), .C1(
        n4401), .C2(n5869), .ZN(P1_U3336) );
  OAI222_X1 U9989 ( .A1(P1_U3086), .A2(n5410), .B1(n10026), .B2(n8320), .C1(
        n9219), .C2(n10037), .ZN(P1_U3325) );
  INV_X1 U9990 ( .A(n9859), .ZN(n8346) );
  INV_X1 U9991 ( .A(n8321), .ZN(n8324) );
  INV_X1 U9992 ( .A(n8322), .ZN(n8323) );
  NAND2_X1 U9993 ( .A1(n8324), .A2(n8323), .ZN(n8336) );
  NAND2_X1 U9994 ( .A1(n9859), .A2(n9041), .ZN(n8326) );
  NAND2_X1 U9995 ( .A1(n9476), .A2(n5468), .ZN(n8325) );
  NAND2_X1 U9996 ( .A1(n8326), .A2(n8325), .ZN(n8328) );
  XNOR2_X1 U9997 ( .A(n8328), .B(n8327), .ZN(n8332) );
  INV_X1 U9998 ( .A(n8332), .ZN(n8334) );
  NOR2_X1 U9999 ( .A1(n9609), .A2(n8329), .ZN(n8330) );
  AOI21_X1 U10000 ( .B1(n9859), .B2(n5468), .A(n8330), .ZN(n8331) );
  INV_X1 U10001 ( .A(n8331), .ZN(n8333) );
  AOI21_X1 U10002 ( .B1(n8340), .B2(n8336), .A(n8335), .ZN(n8341) );
  INV_X1 U10003 ( .A(n8335), .ZN(n8338) );
  INV_X1 U10004 ( .A(n8336), .ZN(n8337) );
  NOR2_X1 U10005 ( .A1(n8338), .A2(n8337), .ZN(n8339) );
  OAI21_X1 U10006 ( .B1(n8341), .B2(n9044), .A(n9204), .ZN(n8345) );
  AOI22_X1 U10007 ( .A1(n9588), .A2(n9197), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n8342) );
  OAI21_X1 U10008 ( .B1(n4402), .B2(n9194), .A(n8342), .ZN(n8343) );
  AOI21_X1 U10009 ( .B1(n9192), .B2(n9584), .A(n8343), .ZN(n8344) );
  OAI211_X1 U10010 ( .C1(n8346), .C2(n9213), .A(n8345), .B(n8344), .ZN(
        P1_U3214) );
  INV_X1 U10011 ( .A(n8977), .ZN(n8347) );
  OAI222_X1 U10012 ( .A1(n10037), .A2(n10558), .B1(n10040), .B2(n8347), .C1(
        n6120), .C2(n4401), .ZN(P1_U3327) );
  INV_X1 U10013 ( .A(n8348), .ZN(n8349) );
  NAND2_X1 U10014 ( .A1(n8352), .A2(n8351), .ZN(n8436) );
  INV_X1 U10015 ( .A(n8352), .ZN(n8353) );
  NAND2_X1 U10016 ( .A1(n8353), .A2(n8490), .ZN(n8435) );
  NAND2_X1 U10017 ( .A1(n8436), .A2(n8435), .ZN(n8354) );
  XOR2_X1 U10018 ( .A(n8437), .B(n8354), .Z(n8363) );
  NAND2_X1 U10019 ( .A1(n8441), .A2(n8491), .ZN(n8356) );
  OAI211_X1 U10020 ( .C1(n8357), .C2(n8454), .A(n8356), .B(n8355), .ZN(n8358)
         );
  AOI21_X1 U10021 ( .B1(n8359), .B2(n8478), .A(n8358), .ZN(n8362) );
  NAND2_X1 U10022 ( .A1(n8360), .A2(n8457), .ZN(n8361) );
  OAI211_X1 U10023 ( .C1(n8363), .C2(n8460), .A(n8362), .B(n8361), .ZN(
        P2_U3157) );
  INV_X1 U10024 ( .A(n8933), .ZN(n8370) );
  OAI211_X1 U10025 ( .C1(n4530), .C2(n8364), .A(n8418), .B(n8470), .ZN(n8369)
         );
  NAND2_X1 U10026 ( .A1(n8761), .A2(n8441), .ZN(n8365) );
  OAI211_X1 U10027 ( .C1(n8733), .C2(n8454), .A(n8366), .B(n8365), .ZN(n8367)
         );
  AOI21_X1 U10028 ( .B1(n8738), .B2(n8478), .A(n8367), .ZN(n8368) );
  OAI211_X1 U10029 ( .C1(n8370), .C2(n8481), .A(n8369), .B(n8368), .ZN(
        P2_U3159) );
  INV_X1 U10030 ( .A(n8863), .ZN(n8712) );
  NOR3_X1 U10031 ( .A1(n4447), .A2(n8372), .A3(n8371), .ZN(n8375) );
  INV_X1 U10032 ( .A(n8373), .ZN(n8374) );
  OAI21_X1 U10033 ( .B1(n8375), .B2(n8374), .A(n8470), .ZN(n8379) );
  AOI22_X1 U10034 ( .A1(n8488), .A2(n8441), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8376) );
  OAI21_X1 U10035 ( .B1(n8708), .B2(n8454), .A(n8376), .ZN(n8377) );
  AOI21_X1 U10036 ( .B1(n8709), .B2(n8478), .A(n8377), .ZN(n8378) );
  OAI211_X1 U10037 ( .C1(n8712), .C2(n8481), .A(n8379), .B(n8378), .ZN(
        P2_U3163) );
  INV_X1 U10038 ( .A(n8912), .ZN(n8667) );
  NOR3_X1 U10039 ( .A1(n4448), .A2(n4828), .A3(n8381), .ZN(n8384) );
  INV_X1 U10040 ( .A(n8382), .ZN(n8383) );
  OAI21_X1 U10041 ( .B1(n8384), .B2(n8383), .A(n8470), .ZN(n8389) );
  AOI22_X1 U10042 ( .A1(n8673), .A2(n8478), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8385) );
  OAI21_X1 U10043 ( .B1(n8386), .B2(n8476), .A(n8385), .ZN(n8387) );
  AOI21_X1 U10044 ( .B1(n8473), .B2(n8670), .A(n8387), .ZN(n8388) );
  OAI211_X1 U10045 ( .C1(n8667), .C2(n8481), .A(n8389), .B(n8388), .ZN(
        P2_U3165) );
  INV_X1 U10046 ( .A(n8779), .ZN(n8946) );
  OAI211_X1 U10047 ( .C1(n8392), .C2(n8391), .A(n8390), .B(n8470), .ZN(n8396)
         );
  NAND2_X1 U10048 ( .A1(n8441), .A2(n8797), .ZN(n8393) );
  NAND2_X1 U10049 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8576) );
  OAI211_X1 U10050 ( .C1(n8772), .C2(n8454), .A(n8393), .B(n8576), .ZN(n8394)
         );
  AOI21_X1 U10051 ( .B1(n8778), .B2(n8478), .A(n8394), .ZN(n8395) );
  OAI211_X1 U10052 ( .C1(n8946), .C2(n8481), .A(n8396), .B(n8395), .ZN(
        P2_U3166) );
  XNOR2_X1 U10053 ( .A(n8397), .B(n8772), .ZN(n8398) );
  XNOR2_X1 U10054 ( .A(n8399), .B(n8398), .ZN(n8405) );
  NOR2_X1 U10055 ( .A1(n10528), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8592) );
  AOI21_X1 U10056 ( .B1(n8761), .B2(n8473), .A(n8592), .ZN(n8401) );
  NAND2_X1 U10057 ( .A1(n8478), .A2(n8764), .ZN(n8400) );
  OAI211_X1 U10058 ( .C1(n8402), .C2(n8476), .A(n8401), .B(n8400), .ZN(n8403)
         );
  AOI21_X1 U10059 ( .B1(n8941), .B2(n8457), .A(n8403), .ZN(n8404) );
  OAI21_X1 U10060 ( .B1(n8405), .B2(n8460), .A(n8404), .ZN(P2_U3168) );
  INV_X1 U10061 ( .A(n8406), .ZN(n8409) );
  INV_X1 U10062 ( .A(n8407), .ZN(n8408) );
  NOR3_X1 U10063 ( .A1(n8410), .A2(n8409), .A3(n8408), .ZN(n8411) );
  OAI21_X1 U10064 ( .B1(n8411), .B2(n4448), .A(n8470), .ZN(n8415) );
  AOI22_X1 U10065 ( .A1(n8683), .A2(n8478), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8412) );
  OAI21_X1 U10066 ( .B1(n8681), .B2(n8476), .A(n8412), .ZN(n8413) );
  AOI21_X1 U10067 ( .B1(n8486), .B2(n8473), .A(n8413), .ZN(n8414) );
  OAI211_X1 U10068 ( .C1(n8917), .C2(n8481), .A(n8415), .B(n8414), .ZN(
        P2_U3169) );
  INV_X1 U10069 ( .A(n8927), .ZN(n8424) );
  AOI21_X1 U10070 ( .B1(n8418), .B2(n8417), .A(n8416), .ZN(n8419) );
  OAI21_X1 U10071 ( .B1(n4447), .B2(n8419), .A(n8470), .ZN(n8423) );
  AOI22_X1 U10072 ( .A1(n8723), .A2(n8473), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8420) );
  OAI21_X1 U10073 ( .B1(n8749), .B2(n8476), .A(n8420), .ZN(n8421) );
  AOI21_X1 U10074 ( .B1(n8726), .B2(n8478), .A(n8421), .ZN(n8422) );
  OAI211_X1 U10075 ( .C1(n8424), .C2(n8481), .A(n8423), .B(n8422), .ZN(
        P2_U3173) );
  INV_X1 U10076 ( .A(n8700), .ZN(n8861) );
  AOI21_X1 U10077 ( .B1(n8426), .B2(n8425), .A(n8460), .ZN(n8428) );
  NAND2_X1 U10078 ( .A1(n8428), .A2(n8427), .ZN(n8434) );
  INV_X1 U10079 ( .A(n8429), .ZN(n8698) );
  AOI22_X1 U10080 ( .A1(n8723), .A2(n8441), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8430) );
  OAI21_X1 U10081 ( .B1(n8698), .B2(n8431), .A(n8430), .ZN(n8432) );
  AOI21_X1 U10082 ( .B1(n8473), .B2(n8695), .A(n8432), .ZN(n8433) );
  OAI211_X1 U10083 ( .C1(n8861), .C2(n8481), .A(n8434), .B(n8433), .ZN(
        P2_U3175) );
  INV_X1 U10084 ( .A(n8435), .ZN(n8438) );
  OAI21_X1 U10085 ( .B1(n8438), .B2(n8437), .A(n8436), .ZN(n8439) );
  XOR2_X1 U10086 ( .A(n8440), .B(n8439), .Z(n8450) );
  NAND2_X1 U10087 ( .A1(n8441), .A2(n8490), .ZN(n8443) );
  NAND2_X1 U10088 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8500) );
  OAI211_X1 U10089 ( .C1(n8444), .C2(n8454), .A(n8443), .B(n8500), .ZN(n8445)
         );
  AOI21_X1 U10090 ( .B1(n8446), .B2(n8478), .A(n8445), .ZN(n8449) );
  NAND2_X1 U10091 ( .A1(n8447), .A2(n8457), .ZN(n8448) );
  OAI211_X1 U10092 ( .C1(n8450), .C2(n8460), .A(n8449), .B(n8448), .ZN(
        P2_U3176) );
  AOI21_X1 U10093 ( .B1(n8453), .B2(n8452), .A(n8451), .ZN(n8461) );
  NOR2_X1 U10094 ( .A1(n8476), .A2(n8772), .ZN(n8456) );
  NAND2_X1 U10095 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8613) );
  OAI21_X1 U10096 ( .B1(n8749), .B2(n8454), .A(n8613), .ZN(n8455) );
  AOI211_X1 U10097 ( .C1(n8745), .C2(n8478), .A(n8456), .B(n8455), .ZN(n8459)
         );
  NAND2_X1 U10098 ( .A1(n8938), .A2(n8457), .ZN(n8458) );
  OAI211_X1 U10099 ( .C1(n8461), .C2(n8460), .A(n8459), .B(n8458), .ZN(
        P2_U3178) );
  OAI21_X1 U10100 ( .B1(n8465), .B2(n8464), .A(n8463), .ZN(n8466) );
  AOI22_X1 U10101 ( .A1(n8662), .A2(n8478), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8467) );
  OAI21_X1 U10102 ( .B1(n8680), .B2(n8476), .A(n8467), .ZN(n8468) );
  AOI21_X1 U10103 ( .B1(n8485), .B2(n8473), .A(n8468), .ZN(n8469) );
  INV_X1 U10104 ( .A(n8952), .ZN(n8482) );
  OAI211_X1 U10105 ( .C1(n4548), .C2(n8472), .A(n8471), .B(n8470), .ZN(n8480)
         );
  INV_X1 U10106 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10465) );
  NOR2_X1 U10107 ( .A1(n10465), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8562) );
  AOI21_X1 U10108 ( .B1(n8473), .B2(n8789), .A(n8562), .ZN(n8474) );
  OAI21_X1 U10109 ( .B1(n8476), .B2(n8475), .A(n8474), .ZN(n8477) );
  AOI21_X1 U10110 ( .B1(n8792), .B2(n8478), .A(n8477), .ZN(n8479) );
  OAI211_X1 U10111 ( .C1(n8482), .C2(n8481), .A(n8480), .B(n8479), .ZN(
        P2_U3181) );
  MUX2_X1 U10112 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n7239), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10113 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8483), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10114 ( .A(n8484), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8606), .Z(
        P2_U3519) );
  MUX2_X1 U10115 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8485), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10116 ( .A(n8670), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8606), .Z(
        P2_U3517) );
  MUX2_X1 U10117 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8486), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10118 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8669), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10119 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8487), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10120 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8723), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10121 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8488), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10122 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8722), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10123 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8761), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10124 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8489), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10125 ( .A(n8789), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8606), .Z(
        P2_U3507) );
  MUX2_X1 U10126 ( .A(n8797), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8606), .Z(
        P2_U3506) );
  MUX2_X1 U10127 ( .A(n8816), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8606), .Z(
        P2_U3505) );
  MUX2_X1 U10128 ( .A(n8827), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8606), .Z(
        P2_U3504) );
  MUX2_X1 U10129 ( .A(n8815), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8606), .Z(
        P2_U3503) );
  MUX2_X1 U10130 ( .A(n4718), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8606), .Z(
        P2_U3502) );
  MUX2_X1 U10131 ( .A(n8490), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8606), .Z(
        P2_U3501) );
  MUX2_X1 U10132 ( .A(n8491), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8606), .Z(
        P2_U3500) );
  MUX2_X1 U10133 ( .A(n8492), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8606), .Z(
        P2_U3499) );
  MUX2_X1 U10134 ( .A(n8493), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8606), .Z(
        P2_U3498) );
  MUX2_X1 U10135 ( .A(n8494), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8606), .Z(
        P2_U3497) );
  MUX2_X1 U10136 ( .A(n8495), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8606), .Z(
        P2_U3496) );
  MUX2_X1 U10137 ( .A(n8496), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8606), .Z(
        P2_U3495) );
  MUX2_X1 U10138 ( .A(n8497), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8606), .Z(
        P2_U3494) );
  MUX2_X1 U10139 ( .A(n8498), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8606), .Z(
        P2_U3493) );
  MUX2_X1 U10140 ( .A(n5112), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8606), .Z(
        P2_U3492) );
  XNOR2_X1 U10141 ( .A(n8499), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n8513) );
  INV_X1 U10142 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n8501) );
  OAI21_X1 U10143 ( .B1(n10294), .B2(n8501), .A(n8500), .ZN(n8506) );
  AOI21_X1 U10144 ( .B1(n8503), .B2(n8502), .A(n8523), .ZN(n8504) );
  NOR2_X1 U10145 ( .A1(n8504), .A2(n10176), .ZN(n8505) );
  AOI211_X1 U10146 ( .C1(n10178), .C2(n8507), .A(n8506), .B(n8505), .ZN(n8512)
         );
  XNOR2_X1 U10147 ( .A(n8509), .B(n8508), .ZN(n8510) );
  NAND2_X1 U10148 ( .A1(n8510), .A2(n10288), .ZN(n8511) );
  OAI211_X1 U10149 ( .C1(n8513), .C2(n10197), .A(n8512), .B(n8511), .ZN(
        P2_U3193) );
  XOR2_X1 U10150 ( .A(n8515), .B(n8514), .Z(n8529) );
  XNOR2_X1 U10151 ( .A(n8517), .B(n8516), .ZN(n8527) );
  NAND2_X1 U10152 ( .A1(n10170), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n8519) );
  OAI211_X1 U10153 ( .C1(n10298), .C2(n8520), .A(n8519), .B(n8518), .ZN(n8526)
         );
  OR3_X1 U10154 ( .A1(n8523), .A2(n8522), .A3(n8521), .ZN(n8524) );
  AOI21_X1 U10155 ( .B1(n4546), .B2(n8524), .A(n10176), .ZN(n8525) );
  AOI211_X1 U10156 ( .C1(n10288), .C2(n8527), .A(n8526), .B(n8525), .ZN(n8528)
         );
  OAI21_X1 U10157 ( .B1(n8529), .B2(n10197), .A(n8528), .ZN(P2_U3194) );
  XNOR2_X1 U10158 ( .A(n8530), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n8542) );
  XNOR2_X1 U10159 ( .A(n8532), .B(n8531), .ZN(n8540) );
  AOI21_X1 U10160 ( .B1(n10170), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n8533), .ZN(
        n8534) );
  OAI21_X1 U10161 ( .B1(n8535), .B2(n10298), .A(n8534), .ZN(n8539) );
  AOI21_X1 U10162 ( .B1(n10468), .B2(n8536), .A(n8551), .ZN(n8537) );
  NOR2_X1 U10163 ( .A1(n8537), .A2(n10176), .ZN(n8538) );
  AOI211_X1 U10164 ( .C1(n10288), .C2(n8540), .A(n8539), .B(n8538), .ZN(n8541)
         );
  OAI21_X1 U10165 ( .B1(n10197), .B2(n8542), .A(n8541), .ZN(P2_U3195) );
  XOR2_X1 U10166 ( .A(n8544), .B(n8543), .Z(n8558) );
  XNOR2_X1 U10167 ( .A(n8546), .B(n8545), .ZN(n8556) );
  NAND2_X1 U10168 ( .A1(n10170), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n8548) );
  OAI211_X1 U10169 ( .C1(n10298), .C2(n5154), .A(n8548), .B(n8547), .ZN(n8555)
         );
  OR3_X1 U10170 ( .A1(n8551), .A2(n8550), .A3(n8549), .ZN(n8552) );
  AOI21_X1 U10171 ( .B1(n8553), .B2(n8552), .A(n10176), .ZN(n8554) );
  AOI211_X1 U10172 ( .C1(n10288), .C2(n8556), .A(n8555), .B(n8554), .ZN(n8557)
         );
  OAI21_X1 U10173 ( .B1(n8558), .B2(n10197), .A(n8557), .ZN(P2_U3196) );
  XNOR2_X1 U10174 ( .A(n8559), .B(P2_REG1_REG_15__SCAN_IN), .ZN(n8571) );
  XNOR2_X1 U10175 ( .A(n8561), .B(n8560), .ZN(n8569) );
  AOI21_X1 U10176 ( .B1(n10170), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8562), .ZN(
        n8563) );
  OAI21_X1 U10177 ( .B1(n5242), .B2(n10298), .A(n8563), .ZN(n8568) );
  NAND2_X1 U10178 ( .A1(n8565), .A2(n8791), .ZN(n8566) );
  AOI21_X1 U10179 ( .B1(n8564), .B2(n8566), .A(n10176), .ZN(n8567) );
  AOI211_X1 U10180 ( .C1(n10288), .C2(n8569), .A(n8568), .B(n8567), .ZN(n8570)
         );
  OAI21_X1 U10181 ( .B1(n8571), .B2(n10197), .A(n8570), .ZN(P2_U3197) );
  XOR2_X1 U10182 ( .A(n8573), .B(n8572), .Z(n8586) );
  XNOR2_X1 U10183 ( .A(n8575), .B(n8574), .ZN(n8584) );
  NAND2_X1 U10184 ( .A1(n10170), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n8577) );
  OAI211_X1 U10185 ( .C1(n10298), .C2(n8578), .A(n8577), .B(n8576), .ZN(n8583)
         );
  NAND3_X1 U10186 ( .A1(n8564), .A2(n4552), .A3(n8579), .ZN(n8580) );
  AOI21_X1 U10187 ( .B1(n8581), .B2(n8580), .A(n10176), .ZN(n8582) );
  AOI211_X1 U10188 ( .C1(n10288), .C2(n8584), .A(n8583), .B(n8582), .ZN(n8585)
         );
  OAI21_X1 U10189 ( .B1(n8586), .B2(n10197), .A(n8585), .ZN(P2_U3198) );
  XNOR2_X1 U10190 ( .A(n8587), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8599) );
  OAI21_X1 U10191 ( .B1(n4482), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8588), .ZN(
        n8589) );
  NAND2_X1 U10192 ( .A1(n8589), .A2(n10191), .ZN(n8598) );
  XNOR2_X1 U10193 ( .A(n8591), .B(n8590), .ZN(n8596) );
  AOI21_X1 U10194 ( .B1(n10170), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8592), .ZN(
        n8593) );
  OAI21_X1 U10195 ( .B1(n8594), .B2(n10298), .A(n8593), .ZN(n8595) );
  AOI21_X1 U10196 ( .B1(n8596), .B2(n10288), .A(n8595), .ZN(n8597) );
  OAI211_X1 U10197 ( .C1(n8599), .C2(n10197), .A(n8598), .B(n8597), .ZN(
        P2_U3199) );
  XOR2_X1 U10198 ( .A(n8601), .B(n8600), .Z(n8621) );
  AND3_X1 U10199 ( .A1(n8588), .A2(n8603), .A3(n8602), .ZN(n8604) );
  OAI21_X1 U10200 ( .B1(n8605), .B2(n8604), .A(n10191), .ZN(n8620) );
  INV_X1 U10201 ( .A(n8611), .ZN(n8607) );
  NOR3_X1 U10202 ( .A1(n8608), .A2(n8607), .A3(n8606), .ZN(n8618) );
  AOI211_X1 U10203 ( .C1(n8612), .C2(n8611), .A(n8610), .B(n8609), .ZN(n8617)
         );
  NAND2_X1 U10204 ( .A1(n10170), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n8614) );
  OAI211_X1 U10205 ( .C1(n10298), .C2(n8615), .A(n8614), .B(n8613), .ZN(n8616)
         );
  NOR3_X1 U10206 ( .A1(n8618), .A2(n8617), .A3(n8616), .ZN(n8619) );
  OAI211_X1 U10207 ( .C1(n8621), .C2(n10197), .A(n8620), .B(n8619), .ZN(
        P2_U3200) );
  NOR2_X1 U10208 ( .A1(n8624), .A2(n10207), .ZN(n8631) );
  AOI21_X1 U10209 ( .B1(n8899), .B2(n10221), .A(n8631), .ZN(n8627) );
  NAND2_X1 U10210 ( .A1(n10223), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8625) );
  OAI211_X1 U10211 ( .C1(n8901), .C2(n8711), .A(n8627), .B(n8625), .ZN(
        P2_U3202) );
  NAND2_X1 U10212 ( .A1(n10223), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8626) );
  OAI211_X1 U10213 ( .C1(n8904), .C2(n8711), .A(n8627), .B(n8626), .ZN(
        P2_U3203) );
  NAND2_X1 U10214 ( .A1(n8628), .A2(n10221), .ZN(n8633) );
  NOR2_X1 U10215 ( .A1(n8629), .A2(n8711), .ZN(n8630) );
  AOI211_X1 U10216 ( .C1(n10223), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8631), .B(
        n8630), .ZN(n8632) );
  OAI211_X1 U10217 ( .C1(n8635), .C2(n8634), .A(n8633), .B(n8632), .ZN(
        P2_U3204) );
  INV_X1 U10218 ( .A(n8641), .ZN(n8637) );
  XNOR2_X1 U10219 ( .A(n8636), .B(n8637), .ZN(n8640) );
  OAI22_X1 U10220 ( .A1(n8638), .A2(n10212), .B1(n8659), .B2(n10211), .ZN(
        n8639) );
  AOI21_X1 U10221 ( .B1(n8640), .B2(n8829), .A(n8639), .ZN(n8847) );
  OR2_X1 U10222 ( .A1(n8642), .A2(n8641), .ZN(n8643) );
  NAND2_X1 U10223 ( .A1(n8644), .A2(n8643), .ZN(n8845) );
  AOI22_X1 U10224 ( .A1(n8645), .A2(n8821), .B1(n10223), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n8646) );
  OAI21_X1 U10225 ( .B1(n8647), .B2(n8711), .A(n8646), .ZN(n8648) );
  AOI21_X1 U10226 ( .B1(n8845), .B2(n8804), .A(n8648), .ZN(n8649) );
  OAI21_X1 U10227 ( .B1(n8847), .B2(n10223), .A(n8649), .ZN(P2_U3205) );
  INV_X1 U10228 ( .A(n8650), .ZN(n8656) );
  AOI22_X1 U10229 ( .A1(n8651), .A2(n8821), .B1(n10223), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8652) );
  OAI21_X1 U10230 ( .B1(n6726), .B2(n8711), .A(n8652), .ZN(n8653) );
  AOI21_X1 U10231 ( .B1(n8654), .B2(n8804), .A(n8653), .ZN(n8655) );
  OAI21_X1 U10232 ( .B1(n8656), .B2(n10223), .A(n8655), .ZN(P2_U3206) );
  XNOR2_X1 U10233 ( .A(n8657), .B(n8661), .ZN(n8658) );
  OAI222_X1 U10234 ( .A1(n10211), .A2(n8680), .B1(n10212), .B2(n8659), .C1(
        n10218), .C2(n8658), .ZN(n8848) );
  INV_X1 U10235 ( .A(n8848), .ZN(n8666) );
  XNOR2_X1 U10236 ( .A(n8660), .B(n8661), .ZN(n8849) );
  AOI22_X1 U10237 ( .A1(n8662), .A2(n8821), .B1(n10223), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8663) );
  OAI21_X1 U10238 ( .B1(n8909), .B2(n8711), .A(n8663), .ZN(n8664) );
  AOI21_X1 U10239 ( .B1(n8849), .B2(n8804), .A(n8664), .ZN(n8665) );
  OAI21_X1 U10240 ( .B1(n8666), .B2(n10223), .A(n8665), .ZN(P2_U3207) );
  NOR2_X1 U10241 ( .A1(n8667), .A2(n10206), .ZN(n8672) );
  XNOR2_X1 U10242 ( .A(n8668), .B(n8675), .ZN(n8671) );
  AOI222_X1 U10243 ( .A1(n8829), .A2(n8671), .B1(n8670), .B2(n8826), .C1(n8669), .C2(n8825), .ZN(n8910) );
  XOR2_X1 U10244 ( .A(n8675), .B(n8674), .Z(n8915) );
  INV_X1 U10245 ( .A(n8915), .ZN(n8676) );
  AOI22_X1 U10246 ( .A1(n8676), .A2(n8804), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n10223), .ZN(n8677) );
  OAI21_X1 U10247 ( .B1(n8678), .B2(n10223), .A(n8677), .ZN(P2_U3208) );
  NOR2_X1 U10248 ( .A1(n8917), .A2(n10206), .ZN(n8682) );
  AOI211_X1 U10249 ( .C1(n8821), .C2(n8683), .A(n8682), .B(n8916), .ZN(n8692)
         );
  OAI21_X1 U10250 ( .B1(n8287), .B2(n8685), .A(n8684), .ZN(n8687) );
  NAND2_X1 U10251 ( .A1(n8687), .A2(n8686), .ZN(n8688) );
  XOR2_X1 U10252 ( .A(n8689), .B(n8688), .Z(n8918) );
  INV_X1 U10253 ( .A(n8918), .ZN(n8690) );
  AOI22_X1 U10254 ( .A1(n8690), .A2(n8804), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n10223), .ZN(n8691) );
  OAI21_X1 U10255 ( .B1(n8692), .B2(n10223), .A(n8691), .ZN(P2_U3209) );
  XNOR2_X1 U10256 ( .A(n8693), .B(n8694), .ZN(n8696) );
  AOI222_X1 U10257 ( .A1(n8829), .A2(n8696), .B1(n8723), .B2(n8825), .C1(n8695), .C2(n8826), .ZN(n8860) );
  OAI22_X1 U10258 ( .A1(n8698), .A2(n10207), .B1(n10221), .B2(n8697), .ZN(
        n8699) );
  AOI21_X1 U10259 ( .B1(n8700), .B2(n8838), .A(n8699), .ZN(n8703) );
  OR2_X1 U10260 ( .A1(n8701), .A2(n5103), .ZN(n8858) );
  NAND3_X1 U10261 ( .A1(n8858), .A2(n8857), .A3(n8804), .ZN(n8702) );
  OAI211_X1 U10262 ( .C1(n8860), .C2(n10223), .A(n8703), .B(n8702), .ZN(
        P2_U3211) );
  XNOR2_X1 U10263 ( .A(n8704), .B(n8705), .ZN(n8924) );
  XOR2_X1 U10264 ( .A(n8706), .B(n8705), .Z(n8707) );
  OAI222_X1 U10265 ( .A1(n10212), .A2(n8708), .B1(n10211), .B2(n8733), .C1(
        n10218), .C2(n8707), .ZN(n8862) );
  AOI22_X1 U10266 ( .A1(n8709), .A2(n8821), .B1(n10223), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n8710) );
  OAI21_X1 U10267 ( .B1(n8712), .B2(n8711), .A(n8710), .ZN(n8713) );
  AOI21_X1 U10268 ( .B1(n8862), .B2(n10221), .A(n8713), .ZN(n8714) );
  OAI21_X1 U10269 ( .B1(n8835), .B2(n8924), .A(n8714), .ZN(P2_U3212) );
  NAND2_X1 U10270 ( .A1(n8716), .A2(n8715), .ZN(n8718) );
  XNOR2_X1 U10271 ( .A(n8718), .B(n8717), .ZN(n8929) );
  OAI21_X1 U10272 ( .B1(n8721), .B2(n8720), .A(n8719), .ZN(n8724) );
  AOI222_X1 U10273 ( .A1(n8829), .A2(n8724), .B1(n8723), .B2(n8826), .C1(n8722), .C2(n8825), .ZN(n8866) );
  MUX2_X1 U10274 ( .A(n8725), .B(n8866), .S(n10221), .Z(n8728) );
  AOI22_X1 U10275 ( .A1(n8927), .A2(n8838), .B1(n8821), .B2(n8726), .ZN(n8727)
         );
  OAI211_X1 U10276 ( .C1(n8929), .C2(n8835), .A(n8728), .B(n8727), .ZN(
        P2_U3213) );
  XNOR2_X1 U10277 ( .A(n8729), .B(n8731), .ZN(n8935) );
  AOI21_X1 U10278 ( .B1(n8730), .B2(n8731), .A(n10218), .ZN(n8736) );
  OAI22_X1 U10279 ( .A1(n8733), .A2(n10212), .B1(n8732), .B2(n10211), .ZN(
        n8734) );
  AOI21_X1 U10280 ( .B1(n8736), .B2(n8735), .A(n8734), .ZN(n8930) );
  INV_X1 U10281 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8737) );
  MUX2_X1 U10282 ( .A(n8930), .B(n8737), .S(n10223), .Z(n8740) );
  AOI22_X1 U10283 ( .A1(n8933), .A2(n8838), .B1(n8821), .B2(n8738), .ZN(n8739)
         );
  OAI211_X1 U10284 ( .C1(n8935), .C2(n8835), .A(n8740), .B(n8739), .ZN(
        P2_U3214) );
  NAND2_X1 U10285 ( .A1(n8742), .A2(n8741), .ZN(n8743) );
  NAND2_X1 U10286 ( .A1(n8744), .A2(n8743), .ZN(n8872) );
  INV_X1 U10287 ( .A(n8745), .ZN(n8746) );
  OAI22_X1 U10288 ( .A1(n8747), .A2(n10221), .B1(n8746), .B2(n10207), .ZN(
        n8753) );
  XNOR2_X1 U10289 ( .A(n8748), .B(n6643), .ZN(n8751) );
  OAI22_X1 U10290 ( .A1(n8749), .A2(n10212), .B1(n8772), .B2(n10211), .ZN(
        n8750) );
  AOI21_X1 U10291 ( .B1(n8751), .B2(n8829), .A(n8750), .ZN(n8873) );
  NOR2_X1 U10292 ( .A1(n8873), .A2(n10223), .ZN(n8752) );
  AOI211_X1 U10293 ( .C1(n8838), .C2(n8938), .A(n8753), .B(n8752), .ZN(n8754)
         );
  OAI21_X1 U10294 ( .B1(n8835), .B2(n8872), .A(n8754), .ZN(P2_U3215) );
  XNOR2_X1 U10295 ( .A(n8755), .B(n8759), .ZN(n8944) );
  NOR2_X1 U10296 ( .A1(n8776), .A2(n8756), .ZN(n8757) );
  NAND2_X1 U10297 ( .A1(n8786), .A2(n8757), .ZN(n8769) );
  NAND2_X1 U10298 ( .A1(n8769), .A2(n8758), .ZN(n8760) );
  XNOR2_X1 U10299 ( .A(n8760), .B(n8759), .ZN(n8762) );
  AOI222_X1 U10300 ( .A1(n8829), .A2(n8762), .B1(n8761), .B2(n8826), .C1(n8789), .C2(n8825), .ZN(n8940) );
  MUX2_X1 U10301 ( .A(n8763), .B(n8940), .S(n10221), .Z(n8766) );
  AOI22_X1 U10302 ( .A1(n8941), .A2(n8838), .B1(n8821), .B2(n8764), .ZN(n8765)
         );
  OAI211_X1 U10303 ( .C1(n8944), .C2(n8835), .A(n8766), .B(n8765), .ZN(
        P2_U3216) );
  NAND2_X1 U10304 ( .A1(n8786), .A2(n8767), .ZN(n8768) );
  NAND2_X1 U10305 ( .A1(n8768), .A2(n8776), .ZN(n8770) );
  NAND3_X1 U10306 ( .A1(n8770), .A2(n8829), .A3(n8769), .ZN(n8775) );
  OAI22_X1 U10307 ( .A1(n8772), .A2(n10212), .B1(n8771), .B2(n10211), .ZN(
        n8773) );
  INV_X1 U10308 ( .A(n8773), .ZN(n8774) );
  NAND2_X1 U10309 ( .A1(n8775), .A2(n8774), .ZN(n8945) );
  MUX2_X1 U10310 ( .A(n8945), .B(P2_REG2_REG_16__SCAN_IN), .S(n10223), .Z(
        n8782) );
  XNOR2_X1 U10311 ( .A(n8777), .B(n8776), .ZN(n8947) );
  AOI22_X1 U10312 ( .A1(n8779), .A2(n8838), .B1(n8821), .B2(n8778), .ZN(n8780)
         );
  OAI21_X1 U10313 ( .B1(n8947), .B2(n8835), .A(n8780), .ZN(n8781) );
  XNOR2_X1 U10314 ( .A(n8784), .B(n8783), .ZN(n8955) );
  INV_X1 U10315 ( .A(n8785), .ZN(n8788) );
  OAI21_X1 U10316 ( .B1(n8788), .B2(n8787), .A(n8786), .ZN(n8790) );
  AOI222_X1 U10317 ( .A1(n8829), .A2(n8790), .B1(n8816), .B2(n8825), .C1(n8789), .C2(n8826), .ZN(n8950) );
  MUX2_X1 U10318 ( .A(n8791), .B(n8950), .S(n10221), .Z(n8794) );
  AOI22_X1 U10319 ( .A1(n8952), .A2(n8838), .B1(n8821), .B2(n8792), .ZN(n8793)
         );
  OAI211_X1 U10320 ( .C1(n8955), .C2(n8835), .A(n8794), .B(n8793), .ZN(
        P2_U3218) );
  NOR2_X1 U10321 ( .A1(n8958), .A2(n10206), .ZN(n8800) );
  XNOR2_X1 U10322 ( .A(n8795), .B(n8802), .ZN(n8796) );
  NAND2_X1 U10323 ( .A1(n8796), .A2(n8829), .ZN(n8799) );
  AOI22_X1 U10324 ( .A1(n8797), .A2(n8826), .B1(n8827), .B2(n8825), .ZN(n8798)
         );
  NAND2_X1 U10325 ( .A1(n8799), .A2(n8798), .ZN(n8956) );
  AOI211_X1 U10326 ( .C1(n8821), .C2(n8801), .A(n8800), .B(n8956), .ZN(n8807)
         );
  XNOR2_X1 U10327 ( .A(n8803), .B(n8802), .ZN(n8959) );
  INV_X1 U10328 ( .A(n8959), .ZN(n8805) );
  AOI22_X1 U10329 ( .A1(n8805), .A2(n8804), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n10223), .ZN(n8806) );
  OAI21_X1 U10330 ( .B1(n8807), .B2(n10223), .A(n8806), .ZN(P2_U3219) );
  XNOR2_X1 U10331 ( .A(n8808), .B(n8814), .ZN(n8968) );
  NAND2_X1 U10332 ( .A1(n8231), .A2(n8809), .ZN(n8824) );
  INV_X1 U10333 ( .A(n8810), .ZN(n8811) );
  AOI21_X1 U10334 ( .B1(n8824), .B2(n8812), .A(n8811), .ZN(n8813) );
  XOR2_X1 U10335 ( .A(n8814), .B(n8813), .Z(n8817) );
  AOI222_X1 U10336 ( .A1(n8829), .A2(n8817), .B1(n8816), .B2(n8826), .C1(n8815), .C2(n8825), .ZN(n8962) );
  OAI21_X1 U10337 ( .B1(n8818), .B2(n10206), .A(n8962), .ZN(n8819) );
  NAND2_X1 U10338 ( .A1(n8819), .A2(n10221), .ZN(n8823) );
  AOI22_X1 U10339 ( .A1(n10223), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8821), 
        .B2(n8820), .ZN(n8822) );
  OAI211_X1 U10340 ( .C1(n8968), .C2(n8835), .A(n8823), .B(n8822), .ZN(
        P2_U3220) );
  XNOR2_X1 U10341 ( .A(n8824), .B(n8833), .ZN(n8828) );
  AOI222_X1 U10342 ( .A1(n8829), .A2(n8828), .B1(n8827), .B2(n8826), .C1(n4718), .C2(n8825), .ZN(n8895) );
  OAI22_X1 U10343 ( .A1(n10221), .A2(n8831), .B1(n8830), .B2(n10207), .ZN(
        n8837) );
  OAI21_X1 U10344 ( .B1(n8834), .B2(n8833), .A(n8832), .ZN(n8896) );
  NOR2_X1 U10345 ( .A1(n8896), .A2(n8835), .ZN(n8836) );
  AOI211_X1 U10346 ( .C1(n8838), .C2(n8893), .A(n8837), .B(n8836), .ZN(n8839)
         );
  OAI21_X1 U10347 ( .B1(n8895), .B2(n10223), .A(n8839), .ZN(P2_U3221) );
  NAND2_X1 U10348 ( .A1(n8899), .A2(n10259), .ZN(n8842) );
  NAND2_X1 U10349 ( .A1(n10257), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8840) );
  OAI211_X1 U10350 ( .C1(n8901), .C2(n8884), .A(n8842), .B(n8840), .ZN(
        P2_U3490) );
  NAND2_X1 U10351 ( .A1(n8841), .A2(n8888), .ZN(n8843) );
  OAI211_X1 U10352 ( .C1(n10259), .C2(n10573), .A(n8843), .B(n8842), .ZN(
        P2_U3489) );
  AOI22_X1 U10353 ( .A1(n8845), .A2(n10245), .B1(n8892), .B2(n8844), .ZN(n8846) );
  NAND2_X1 U10354 ( .A1(n8847), .A2(n8846), .ZN(n8905) );
  MUX2_X1 U10355 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8905), .S(n10254), .Z(
        P2_U3487) );
  INV_X1 U10356 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8850) );
  AOI21_X1 U10357 ( .B1(n8849), .B2(n10245), .A(n8848), .ZN(n8906) );
  MUX2_X1 U10358 ( .A(n8850), .B(n8906), .S(n10259), .Z(n8851) );
  OAI21_X1 U10359 ( .B1(n8909), .B2(n8884), .A(n8851), .ZN(P2_U3485) );
  INV_X1 U10360 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8852) );
  MUX2_X1 U10361 ( .A(n8852), .B(n8910), .S(n10254), .Z(n8854) );
  NAND2_X1 U10362 ( .A1(n8912), .A2(n8888), .ZN(n8853) );
  OAI211_X1 U10363 ( .C1(n8915), .C2(n8891), .A(n8854), .B(n8853), .ZN(
        P2_U3484) );
  MUX2_X1 U10364 ( .A(n8916), .B(P2_REG1_REG_24__SCAN_IN), .S(n10257), .Z(
        n8856) );
  OAI22_X1 U10365 ( .A1(n8918), .A2(n8891), .B1(n8917), .B2(n8884), .ZN(n8855)
         );
  OR2_X1 U10366 ( .A1(n8856), .A2(n8855), .ZN(P2_U3483) );
  NAND3_X1 U10367 ( .A1(n8858), .A2(n10245), .A3(n8857), .ZN(n8859) );
  OAI211_X1 U10368 ( .C1(n8861), .C2(n10242), .A(n8860), .B(n8859), .ZN(n8920)
         );
  MUX2_X1 U10369 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8920), .S(n10254), .Z(
        P2_U3481) );
  INV_X1 U10370 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8864) );
  AOI21_X1 U10371 ( .B1(n8892), .B2(n8863), .A(n8862), .ZN(n8921) );
  MUX2_X1 U10372 ( .A(n8864), .B(n8921), .S(n10254), .Z(n8865) );
  OAI21_X1 U10373 ( .B1(n8891), .B2(n8924), .A(n8865), .ZN(P2_U3480) );
  INV_X1 U10374 ( .A(n8866), .ZN(n8925) );
  MUX2_X1 U10375 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8925), .S(n10259), .Z(
        n8867) );
  AOI21_X1 U10376 ( .B1(n8888), .B2(n8927), .A(n8867), .ZN(n8868) );
  OAI21_X1 U10377 ( .B1(n8929), .B2(n8891), .A(n8868), .ZN(P2_U3479) );
  MUX2_X1 U10378 ( .A(n8930), .B(n8869), .S(n10257), .Z(n8871) );
  NAND2_X1 U10379 ( .A1(n8933), .A2(n8888), .ZN(n8870) );
  OAI211_X1 U10380 ( .C1(n8935), .C2(n8891), .A(n8871), .B(n8870), .ZN(
        P2_U3478) );
  OR2_X1 U10381 ( .A1(n8872), .A2(n8897), .ZN(n8874) );
  NAND2_X1 U10382 ( .A1(n8874), .A2(n8873), .ZN(n8936) );
  MUX2_X1 U10383 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8936), .S(n10254), .Z(
        n8875) );
  AOI21_X1 U10384 ( .B1(n8888), .B2(n8938), .A(n8875), .ZN(n8876) );
  INV_X1 U10385 ( .A(n8876), .ZN(P2_U3477) );
  MUX2_X1 U10386 ( .A(n10436), .B(n8940), .S(n10259), .Z(n8878) );
  NAND2_X1 U10387 ( .A1(n8941), .A2(n8888), .ZN(n8877) );
  OAI211_X1 U10388 ( .C1(n8944), .C2(n8891), .A(n8878), .B(n8877), .ZN(
        P2_U3476) );
  MUX2_X1 U10389 ( .A(n8945), .B(P2_REG1_REG_16__SCAN_IN), .S(n10257), .Z(
        n8880) );
  OAI22_X1 U10390 ( .A1(n8947), .A2(n8891), .B1(n8946), .B2(n8884), .ZN(n8879)
         );
  MUX2_X1 U10391 ( .A(n8881), .B(n8950), .S(n10259), .Z(n8883) );
  NAND2_X1 U10392 ( .A1(n8952), .A2(n8888), .ZN(n8882) );
  OAI211_X1 U10393 ( .C1(n8955), .C2(n8891), .A(n8883), .B(n8882), .ZN(
        P2_U3474) );
  MUX2_X1 U10394 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8956), .S(n10259), .Z(
        n8886) );
  OAI22_X1 U10395 ( .A1(n8959), .A2(n8891), .B1(n8958), .B2(n8884), .ZN(n8885)
         );
  OR2_X1 U10396 ( .A1(n8886), .A2(n8885), .ZN(P2_U3473) );
  MUX2_X1 U10397 ( .A(n8887), .B(n8962), .S(n10259), .Z(n8890) );
  NAND2_X1 U10398 ( .A1(n8964), .A2(n8888), .ZN(n8889) );
  OAI211_X1 U10399 ( .C1(n8891), .C2(n8968), .A(n8890), .B(n8889), .ZN(
        P2_U3472) );
  NAND2_X1 U10400 ( .A1(n8893), .A2(n8892), .ZN(n8894) );
  OAI211_X1 U10401 ( .C1(n8897), .C2(n8896), .A(n8895), .B(n8894), .ZN(n8969)
         );
  MUX2_X1 U10402 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n8969), .S(n10259), .Z(
        P2_U3471) );
  MUX2_X1 U10403 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n8898), .S(n10259), .Z(
        P2_U3459) );
  NAND2_X1 U10404 ( .A1(n8899), .A2(n10247), .ZN(n8902) );
  NAND2_X1 U10405 ( .A1(n10249), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8900) );
  OAI211_X1 U10406 ( .C1(n8901), .C2(n8957), .A(n8902), .B(n8900), .ZN(
        P2_U3458) );
  NAND2_X1 U10407 ( .A1(n10249), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8903) );
  OAI211_X1 U10408 ( .C1(n8904), .C2(n8957), .A(n8903), .B(n8902), .ZN(
        P2_U3457) );
  MUX2_X1 U10409 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8905), .S(n10247), .Z(
        P2_U3455) );
  INV_X1 U10410 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8907) );
  MUX2_X1 U10411 ( .A(n8907), .B(n8906), .S(n10247), .Z(n8908) );
  OAI21_X1 U10412 ( .B1(n8909), .B2(n8957), .A(n8908), .ZN(P2_U3453) );
  INV_X1 U10413 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8911) );
  MUX2_X1 U10414 ( .A(n8911), .B(n8910), .S(n10247), .Z(n8914) );
  NAND2_X1 U10415 ( .A1(n8912), .A2(n6778), .ZN(n8913) );
  OAI211_X1 U10416 ( .C1(n8915), .C2(n8967), .A(n8914), .B(n8913), .ZN(
        P2_U3452) );
  OAI22_X1 U10417 ( .A1(n8918), .A2(n8967), .B1(n8917), .B2(n8957), .ZN(n8919)
         );
  MUX2_X1 U10418 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8920), .S(n10247), .Z(
        P2_U3449) );
  INV_X1 U10419 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8922) );
  MUX2_X1 U10420 ( .A(n8922), .B(n8921), .S(n10247), .Z(n8923) );
  OAI21_X1 U10421 ( .B1(n8924), .B2(n8967), .A(n8923), .ZN(P2_U3448) );
  MUX2_X1 U10422 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8925), .S(n10247), .Z(
        n8926) );
  AOI21_X1 U10423 ( .B1(n6778), .B2(n8927), .A(n8926), .ZN(n8928) );
  OAI21_X1 U10424 ( .B1(n8929), .B2(n8967), .A(n8928), .ZN(P2_U3447) );
  INV_X1 U10425 ( .A(n8930), .ZN(n8931) );
  MUX2_X1 U10426 ( .A(n8931), .B(P2_REG0_REG_19__SCAN_IN), .S(n10249), .Z(
        n8932) );
  AOI21_X1 U10427 ( .B1(n6778), .B2(n8933), .A(n8932), .ZN(n8934) );
  OAI21_X1 U10428 ( .B1(n8935), .B2(n8967), .A(n8934), .ZN(P2_U3446) );
  MUX2_X1 U10429 ( .A(n8936), .B(P2_REG0_REG_18__SCAN_IN), .S(n10249), .Z(
        n8937) );
  AOI21_X1 U10430 ( .B1(n6778), .B2(n8938), .A(n8937), .ZN(n8939) );
  INV_X1 U10431 ( .A(n8939), .ZN(P2_U3444) );
  INV_X1 U10432 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n10570) );
  MUX2_X1 U10433 ( .A(n10570), .B(n8940), .S(n10247), .Z(n8943) );
  NAND2_X1 U10434 ( .A1(n8941), .A2(n6778), .ZN(n8942) );
  OAI211_X1 U10435 ( .C1(n8944), .C2(n8967), .A(n8943), .B(n8942), .ZN(
        P2_U3441) );
  MUX2_X1 U10436 ( .A(n8945), .B(P2_REG0_REG_16__SCAN_IN), .S(n10249), .Z(
        n8949) );
  OAI22_X1 U10437 ( .A1(n8947), .A2(n8967), .B1(n8946), .B2(n8957), .ZN(n8948)
         );
  INV_X1 U10438 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8951) );
  MUX2_X1 U10439 ( .A(n8951), .B(n8950), .S(n10247), .Z(n8954) );
  NAND2_X1 U10440 ( .A1(n8952), .A2(n6778), .ZN(n8953) );
  OAI211_X1 U10441 ( .C1(n8955), .C2(n8967), .A(n8954), .B(n8953), .ZN(
        P2_U3435) );
  MUX2_X1 U10442 ( .A(n8956), .B(P2_REG0_REG_14__SCAN_IN), .S(n10249), .Z(
        n8961) );
  OAI22_X1 U10443 ( .A1(n8959), .A2(n8967), .B1(n8958), .B2(n8957), .ZN(n8960)
         );
  OR2_X1 U10444 ( .A1(n8961), .A2(n8960), .ZN(P2_U3432) );
  INV_X1 U10445 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8963) );
  MUX2_X1 U10446 ( .A(n8963), .B(n8962), .S(n10247), .Z(n8966) );
  NAND2_X1 U10447 ( .A1(n8964), .A2(n6778), .ZN(n8965) );
  OAI211_X1 U10448 ( .C1(n8968), .C2(n8967), .A(n8966), .B(n8965), .ZN(
        P2_U3429) );
  MUX2_X1 U10449 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n8969), .S(n10247), .Z(
        P2_U3426) );
  INV_X1 U10450 ( .A(n9214), .ZN(n10027) );
  NAND2_X1 U10451 ( .A1(n8982), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8973) );
  INV_X1 U10452 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8971) );
  NAND4_X1 U10453 ( .A1(n5090), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .A4(n8971), .ZN(n8972) );
  OAI211_X1 U10454 ( .C1(n10027), .C2(n4411), .A(n8973), .B(n8972), .ZN(
        P2_U3264) );
  INV_X1 U10455 ( .A(n8974), .ZN(n10028) );
  OAI222_X1 U10456 ( .A1(n4411), .A2(n10028), .B1(n5307), .B2(P2_U3151), .C1(
        n8975), .C2(n8991), .ZN(P2_U3266) );
  NAND2_X1 U10457 ( .A1(n8977), .A2(n8976), .ZN(n8978) );
  OAI211_X1 U10458 ( .C1(n8979), .C2(n8991), .A(n8978), .B(n10284), .ZN(
        P2_U3267) );
  INV_X1 U10459 ( .A(n8980), .ZN(n10029) );
  AOI21_X1 U10460 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n8982), .A(n8981), .ZN(
        n8983) );
  OAI21_X1 U10461 ( .B1(n10029), .B2(n4411), .A(n8983), .ZN(P2_U3268) );
  INV_X1 U10462 ( .A(n8984), .ZN(n10032) );
  OAI222_X1 U10463 ( .A1(n4411), .A2(n10032), .B1(P2_U3151), .B2(n8986), .C1(
        n8985), .C2(n8991), .ZN(P2_U3269) );
  INV_X1 U10464 ( .A(n8987), .ZN(n10035) );
  OAI222_X1 U10465 ( .A1(n4411), .A2(n10035), .B1(P2_U3151), .B2(n8989), .C1(
        n8988), .C2(n8991), .ZN(P2_U3270) );
  INV_X1 U10466 ( .A(n8990), .ZN(n10039) );
  OAI222_X1 U10467 ( .A1(n4411), .A2(n10039), .B1(P2_U3151), .B2(n8992), .C1(
        n10520), .C2(n8991), .ZN(P2_U3271) );
  INV_X1 U10468 ( .A(n8994), .ZN(n8997) );
  XNOR2_X1 U10469 ( .A(n8995), .B(n9104), .ZN(n8996) );
  NOR2_X1 U10470 ( .A1(n8996), .A2(n8997), .ZN(n9103) );
  AOI21_X1 U10471 ( .B1(n8997), .B2(n8996), .A(n9103), .ZN(n9002) );
  NAND2_X1 U10472 ( .A1(n9192), .A2(n9803), .ZN(n8998) );
  NAND2_X1 U10473 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9526) );
  OAI211_X1 U10474 ( .C1(n9934), .C2(n9194), .A(n8998), .B(n9526), .ZN(n8999)
         );
  AOI21_X1 U10475 ( .B1(n9795), .B2(n9197), .A(n8999), .ZN(n9001) );
  NAND2_X1 U10476 ( .A1(n9937), .A2(n9171), .ZN(n9000) );
  OAI211_X1 U10477 ( .C1(n9002), .C2(n9199), .A(n9001), .B(n9000), .ZN(
        P1_U3215) );
  NAND2_X1 U10478 ( .A1(n9004), .A2(n9003), .ZN(n9006) );
  XOR2_X1 U10479 ( .A(n9006), .B(n9005), .Z(n9007) );
  NAND2_X1 U10480 ( .A1(n9007), .A2(n9204), .ZN(n9012) );
  NOR2_X1 U10481 ( .A1(n9658), .A2(n9206), .ZN(n9010) );
  OAI22_X1 U10482 ( .A1(n9300), .A2(n9194), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9008), .ZN(n9009) );
  AOI211_X1 U10483 ( .C1(n9192), .C2(n9650), .A(n9010), .B(n9009), .ZN(n9011)
         );
  OAI211_X1 U10484 ( .C1(n5012), .C2(n9213), .A(n9012), .B(n9011), .ZN(
        P1_U3216) );
  INV_X1 U10485 ( .A(n9013), .ZN(n9015) );
  XNOR2_X1 U10486 ( .A(n9176), .B(n9175), .ZN(n9014) );
  NOR2_X1 U10487 ( .A1(n9014), .A2(n9015), .ZN(n9174) );
  AOI21_X1 U10488 ( .B1(n9015), .B2(n9014), .A(n9174), .ZN(n9023) );
  NAND2_X1 U10489 ( .A1(n9192), .A2(n9480), .ZN(n9017) );
  OAI211_X1 U10490 ( .C1(n9063), .C2(n9194), .A(n9017), .B(n9016), .ZN(n9020)
         );
  NOR2_X1 U10491 ( .A1(n9018), .A2(n9213), .ZN(n9019) );
  AOI211_X1 U10492 ( .C1(n9021), .C2(n9197), .A(n9020), .B(n9019), .ZN(n9022)
         );
  OAI21_X1 U10493 ( .B1(n9023), .B2(n9199), .A(n9022), .ZN(P1_U3217) );
  INV_X1 U10494 ( .A(n9025), .ZN(n9026) );
  XOR2_X1 U10495 ( .A(n9024), .B(n9025), .Z(n9190) );
  NOR2_X1 U10496 ( .A1(n9190), .A2(n9191), .ZN(n9189) );
  AOI21_X1 U10497 ( .B1(n9024), .B2(n9026), .A(n9189), .ZN(n9030) );
  XNOR2_X1 U10498 ( .A(n9028), .B(n9027), .ZN(n9029) );
  XNOR2_X1 U10499 ( .A(n9030), .B(n9029), .ZN(n9035) );
  NAND2_X1 U10500 ( .A1(n4401), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9560) );
  OAI21_X1 U10501 ( .B1(n9194), .B2(n9120), .A(n9560), .ZN(n9031) );
  AOI21_X1 U10502 ( .B1(n9192), .B2(n9712), .A(n9031), .ZN(n9032) );
  OAI21_X1 U10503 ( .B1(n9206), .B2(n9722), .A(n9032), .ZN(n9033) );
  AOI21_X1 U10504 ( .B1(n9720), .B2(n9171), .A(n9033), .ZN(n9034) );
  OAI21_X1 U10505 ( .B1(n9035), .B2(n9199), .A(n9034), .ZN(P1_U3219) );
  NAND2_X1 U10506 ( .A1(n9578), .A2(n5822), .ZN(n9038) );
  NAND2_X1 U10507 ( .A1(n9584), .A2(n9036), .ZN(n9037) );
  NAND2_X1 U10508 ( .A1(n9038), .A2(n9037), .ZN(n9040) );
  XNOR2_X1 U10509 ( .A(n9040), .B(n9039), .ZN(n9043) );
  AOI22_X1 U10510 ( .A1(n9578), .A2(n9041), .B1(n5822), .B2(n9584), .ZN(n9042)
         );
  XNOR2_X1 U10511 ( .A(n9043), .B(n9042), .ZN(n9050) );
  OR4_X2 U10512 ( .A1(n9044), .A2(n9050), .A3(n9199), .A4(n9049), .ZN(n9054)
         );
  NAND3_X1 U10513 ( .A1(n9044), .A2(n9204), .A3(n9050), .ZN(n9053) );
  INV_X1 U10514 ( .A(n9045), .ZN(n9573) );
  AOI22_X1 U10515 ( .A1(n9573), .A2(n9197), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n9046) );
  OAI21_X1 U10516 ( .B1(n9609), .B2(n9194), .A(n9046), .ZN(n9048) );
  NOR2_X1 U10517 ( .A1(n5174), .A2(n9213), .ZN(n9047) );
  AOI211_X1 U10518 ( .C1(n9192), .C2(n9475), .A(n9048), .B(n9047), .ZN(n9052)
         );
  NAND3_X1 U10519 ( .A1(n9050), .A2(n9204), .A3(n9049), .ZN(n9051) );
  NAND4_X1 U10520 ( .A1(n9054), .A2(n9053), .A3(n9052), .A4(n9051), .ZN(
        P1_U3220) );
  XNOR2_X1 U10521 ( .A(n9055), .B(n9056), .ZN(n9057) );
  NAND2_X1 U10522 ( .A1(n9057), .A2(n9058), .ZN(n9134) );
  OAI21_X1 U10523 ( .B1(n9058), .B2(n9057), .A(n9134), .ZN(n9065) );
  AOI22_X1 U10524 ( .A1(n9171), .A2(n9965), .B1(n9059), .B2(n9197), .ZN(n9062)
         );
  AOI21_X1 U10525 ( .B1(n9210), .B2(n9483), .A(n9060), .ZN(n9061) );
  OAI211_X1 U10526 ( .C1(n9063), .C2(n9207), .A(n9062), .B(n9061), .ZN(n9064)
         );
  AOI21_X1 U10527 ( .B1(n9065), .B2(n9204), .A(n9064), .ZN(n9066) );
  INV_X1 U10528 ( .A(n9066), .ZN(P1_U3221) );
  OAI21_X1 U10529 ( .B1(n9069), .B2(n9068), .A(n9067), .ZN(n9070) );
  NAND2_X1 U10530 ( .A1(n9070), .A2(n9204), .ZN(n9075) );
  AOI22_X1 U10531 ( .A1(n9171), .A2(n9072), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n9071), .ZN(n9074) );
  NAND3_X1 U10532 ( .A1(n9075), .A2(n9074), .A3(n9073), .ZN(P1_U3222) );
  INV_X1 U10533 ( .A(n9076), .ZN(n9077) );
  AOI21_X1 U10534 ( .B1(n9079), .B2(n9078), .A(n9077), .ZN(n9084) );
  AOI22_X1 U10535 ( .A1(n9688), .A2(n9192), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        n4401), .ZN(n9081) );
  NAND2_X1 U10536 ( .A1(n9712), .A2(n9210), .ZN(n9080) );
  OAI211_X1 U10537 ( .C1(n9206), .C2(n9679), .A(n9081), .B(n9080), .ZN(n9082)
         );
  AOI21_X1 U10538 ( .B1(n9896), .B2(n9171), .A(n9082), .ZN(n9083) );
  OAI21_X1 U10539 ( .B1(n9084), .B2(n9199), .A(n9083), .ZN(P1_U3223) );
  XOR2_X1 U10540 ( .A(n9085), .B(n9086), .Z(n9095) );
  NOR2_X1 U10541 ( .A1(n9087), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9512) );
  AOI21_X1 U10542 ( .B1(n9192), .B2(n9478), .A(n9512), .ZN(n9090) );
  NAND2_X1 U10543 ( .A1(n9197), .A2(n9088), .ZN(n9089) );
  OAI211_X1 U10544 ( .C1(n9091), .C2(n9194), .A(n9090), .B(n9089), .ZN(n9092)
         );
  AOI21_X1 U10545 ( .B1(n9093), .B2(n9171), .A(n9092), .ZN(n9094) );
  OAI21_X1 U10546 ( .B1(n9095), .B2(n9199), .A(n9094), .ZN(P1_U3224) );
  OAI21_X1 U10547 ( .B1(n9097), .B2(n9096), .A(n6086), .ZN(n9098) );
  NAND2_X1 U10548 ( .A1(n9098), .A2(n9204), .ZN(n9102) );
  AOI22_X1 U10549 ( .A1(n9650), .A2(n9210), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        n4401), .ZN(n9099) );
  OAI21_X1 U10550 ( .B1(n9206), .B2(n9622), .A(n9099), .ZN(n9100) );
  AOI21_X1 U10551 ( .B1(n9192), .B2(n4412), .A(n9100), .ZN(n9101) );
  OAI211_X1 U10552 ( .C1(n9982), .C2(n9213), .A(n9102), .B(n9101), .ZN(
        P1_U3225) );
  INV_X1 U10553 ( .A(n9106), .ZN(n9203) );
  XNOR2_X1 U10554 ( .A(n9109), .B(n9108), .ZN(n9110) );
  XNOR2_X1 U10555 ( .A(n9111), .B(n9110), .ZN(n9117) );
  NAND2_X1 U10556 ( .A1(n9192), .A2(n9767), .ZN(n9112) );
  NAND2_X1 U10557 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10118)
         );
  OAI211_X1 U10558 ( .C1(n9113), .C2(n9194), .A(n9112), .B(n10118), .ZN(n9114)
         );
  AOI21_X1 U10559 ( .B1(n9761), .B2(n9197), .A(n9114), .ZN(n9116) );
  NAND2_X1 U10560 ( .A1(n9925), .A2(n9171), .ZN(n9115) );
  OAI211_X1 U10561 ( .C1(n9117), .C2(n9199), .A(n9116), .B(n9115), .ZN(
        P1_U3226) );
  XOR2_X1 U10562 ( .A(n9118), .B(n9119), .Z(n9125) );
  NAND2_X1 U10563 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10133)
         );
  OAI21_X1 U10564 ( .B1(n9207), .B2(n9120), .A(n10133), .ZN(n9121) );
  AOI21_X1 U10565 ( .B1(n9210), .B2(n9780), .A(n9121), .ZN(n9122) );
  OAI21_X1 U10566 ( .B1(n9206), .B2(n9748), .A(n9122), .ZN(n9123) );
  AOI21_X1 U10567 ( .B1(n9755), .B2(n9171), .A(n9123), .ZN(n9124) );
  OAI21_X1 U10568 ( .B1(n9125), .B2(n9199), .A(n9124), .ZN(P1_U3228) );
  OAI21_X1 U10569 ( .B1(n9128), .B2(n9127), .A(n9126), .ZN(n9129) );
  NAND2_X1 U10570 ( .A1(n9129), .A2(n9204), .ZN(n9133) );
  AOI22_X1 U10571 ( .A1(n9876), .A2(n9210), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n9130) );
  OAI21_X1 U10572 ( .B1(n9608), .B2(n9207), .A(n9130), .ZN(n9131) );
  AOI21_X1 U10573 ( .B1(n9637), .B2(n9197), .A(n9131), .ZN(n9132) );
  OAI211_X1 U10574 ( .C1(n5192), .C2(n9213), .A(n9133), .B(n9132), .ZN(
        P1_U3229) );
  OAI21_X1 U10575 ( .B1(n9135), .B2(n9055), .A(n9134), .ZN(n9139) );
  XNOR2_X1 U10576 ( .A(n9137), .B(n9136), .ZN(n9138) );
  XNOR2_X1 U10577 ( .A(n9139), .B(n9138), .ZN(n9146) );
  NAND2_X1 U10578 ( .A1(n9192), .A2(n9481), .ZN(n9141) );
  OAI211_X1 U10579 ( .C1(n9142), .C2(n9194), .A(n9141), .B(n9140), .ZN(n9143)
         );
  AOI21_X1 U10580 ( .B1(n9835), .B2(n9197), .A(n9143), .ZN(n9145) );
  NAND2_X1 U10581 ( .A1(n9171), .A2(n9838), .ZN(n9144) );
  OAI211_X1 U10582 ( .C1(n9146), .C2(n9199), .A(n9145), .B(n9144), .ZN(
        P1_U3231) );
  NAND2_X1 U10583 ( .A1(n9148), .A2(n9147), .ZN(n9150) );
  XOR2_X1 U10584 ( .A(n9150), .B(n9149), .Z(n9155) );
  AOI22_X1 U10585 ( .A1(n9210), .A2(n9477), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        n4401), .ZN(n9152) );
  NAND2_X1 U10586 ( .A1(n9197), .A2(n9696), .ZN(n9151) );
  OAI211_X1 U10587 ( .C1(n9888), .C2(n9207), .A(n9152), .B(n9151), .ZN(n9153)
         );
  AOI21_X1 U10588 ( .B1(n9903), .B2(n9171), .A(n9153), .ZN(n9154) );
  OAI21_X1 U10589 ( .B1(n9155), .B2(n9199), .A(n9154), .ZN(P1_U3233) );
  XOR2_X1 U10590 ( .A(n9156), .B(n9157), .Z(n9163) );
  NAND2_X1 U10591 ( .A1(n9192), .A2(n9779), .ZN(n9159) );
  OAI211_X1 U10592 ( .C1(n9944), .C2(n9194), .A(n9159), .B(n9158), .ZN(n9160)
         );
  AOI21_X1 U10593 ( .B1(n9826), .B2(n9197), .A(n9160), .ZN(n9162) );
  NAND2_X1 U10594 ( .A1(n9941), .A2(n9171), .ZN(n9161) );
  OAI211_X1 U10595 ( .C1(n9163), .C2(n9199), .A(n9162), .B(n9161), .ZN(
        P1_U3234) );
  NAND2_X1 U10596 ( .A1(n9164), .A2(n9165), .ZN(n9167) );
  XNOR2_X1 U10597 ( .A(n9167), .B(n9166), .ZN(n9173) );
  AOI22_X1 U10598 ( .A1(n9876), .A2(n9192), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9169) );
  NAND2_X1 U10599 ( .A1(n9702), .A2(n9210), .ZN(n9168) );
  OAI211_X1 U10600 ( .C1(n9206), .C2(n9668), .A(n9169), .B(n9168), .ZN(n9170)
         );
  AOI21_X1 U10601 ( .B1(n9673), .B2(n9171), .A(n9170), .ZN(n9172) );
  OAI21_X1 U10602 ( .B1(n9173), .B2(n9199), .A(n9172), .ZN(P1_U3235) );
  AOI21_X1 U10603 ( .B1(n9176), .B2(n9175), .A(n9174), .ZN(n9180) );
  XNOR2_X1 U10604 ( .A(n9178), .B(n9177), .ZN(n9179) );
  XNOR2_X1 U10605 ( .A(n9180), .B(n9179), .ZN(n9188) );
  NAND2_X1 U10606 ( .A1(n9192), .A2(n9479), .ZN(n9182) );
  OAI211_X1 U10607 ( .C1(n9183), .C2(n9194), .A(n9182), .B(n9181), .ZN(n9185)
         );
  NOR2_X1 U10608 ( .A1(n10017), .A2(n9213), .ZN(n9184) );
  AOI211_X1 U10609 ( .C1(n9186), .C2(n9197), .A(n9185), .B(n9184), .ZN(n9187)
         );
  OAI21_X1 U10610 ( .B1(n9188), .B2(n9199), .A(n9187), .ZN(P1_U3236) );
  AOI21_X1 U10611 ( .B1(n9191), .B2(n9190), .A(n9189), .ZN(n9200) );
  NAND2_X1 U10612 ( .A1(n9192), .A2(n9477), .ZN(n9193) );
  NAND2_X1 U10613 ( .A1(n4401), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10147) );
  OAI211_X1 U10614 ( .C1(n9734), .C2(n9194), .A(n9193), .B(n10147), .ZN(n9196)
         );
  NOR2_X1 U10615 ( .A1(n9739), .A2(n9213), .ZN(n9195) );
  AOI211_X1 U10616 ( .C1(n9736), .C2(n9197), .A(n9196), .B(n9195), .ZN(n9198)
         );
  OAI21_X1 U10617 ( .B1(n9200), .B2(n9199), .A(n9198), .ZN(P1_U3238) );
  OAI21_X1 U10618 ( .B1(n9203), .B2(n9202), .A(n9201), .ZN(n9205) );
  NAND2_X1 U10619 ( .A1(n9205), .A2(n9204), .ZN(n9212) );
  NOR2_X1 U10620 ( .A1(n9206), .A2(n9786), .ZN(n9209) );
  NAND2_X1 U10621 ( .A1(n4401), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9537) );
  OAI21_X1 U10622 ( .B1(n9207), .B2(n9919), .A(n9537), .ZN(n9208) );
  AOI211_X1 U10623 ( .C1(n9210), .C2(n9779), .A(n9209), .B(n9208), .ZN(n9211)
         );
  OAI211_X1 U10624 ( .C1(n10006), .C2(n9213), .A(n9212), .B(n9211), .ZN(
        P1_U3241) );
  INV_X1 U10625 ( .A(n9323), .ZN(n9330) );
  NAND2_X1 U10626 ( .A1(n9214), .A2(n6953), .ZN(n9217) );
  OR2_X1 U10627 ( .A1(n9220), .A2(n9215), .ZN(n9216) );
  NAND2_X1 U10628 ( .A1(n9331), .A2(n9563), .ZN(n9420) );
  INV_X1 U10629 ( .A(n9420), .ZN(n9329) );
  NAND2_X1 U10630 ( .A1(n9218), .A2(n6953), .ZN(n9222) );
  OR2_X1 U10631 ( .A1(n9220), .A2(n9219), .ZN(n9221) );
  AOI21_X1 U10632 ( .B1(n9855), .B2(n9323), .A(n9419), .ZN(n9328) );
  INV_X1 U10633 ( .A(n9423), .ZN(n9631) );
  NAND2_X1 U10634 ( .A1(n9343), .A2(n9387), .ZN(n9636) );
  AND4_X1 U10635 ( .A1(n9223), .A2(n9226), .A3(n9231), .A4(n9323), .ZN(n9224)
         );
  NAND2_X1 U10636 ( .A1(n9225), .A2(n9224), .ZN(n9236) );
  NAND3_X1 U10637 ( .A1(n9229), .A2(n9330), .A3(n9230), .ZN(n9234) );
  NAND2_X1 U10638 ( .A1(n9355), .A2(n9230), .ZN(n9232) );
  NAND3_X1 U10639 ( .A1(n9232), .A2(n9231), .A3(n9323), .ZN(n9233) );
  NAND4_X1 U10640 ( .A1(n9234), .A2(n9235), .A3(n9236), .A4(n9233), .ZN(n9241)
         );
  INV_X1 U10641 ( .A(n9237), .ZN(n9238) );
  MUX2_X1 U10642 ( .A(n9239), .B(n9238), .S(n9323), .Z(n9240) );
  NAND2_X1 U10643 ( .A1(n9241), .A2(n9240), .ZN(n9246) );
  AND2_X1 U10644 ( .A1(n9247), .A2(n9242), .ZN(n9244) );
  MUX2_X1 U10645 ( .A(n9244), .B(n9243), .S(n9323), .Z(n9245) );
  NAND2_X1 U10646 ( .A1(n9246), .A2(n9245), .ZN(n9253) );
  AND2_X1 U10647 ( .A1(n9257), .A2(n9254), .ZN(n9362) );
  NAND3_X1 U10648 ( .A1(n9253), .A2(n9362), .A3(n9247), .ZN(n9251) );
  INV_X1 U10649 ( .A(n9362), .ZN(n9248) );
  OR2_X1 U10650 ( .A1(n9248), .A2(n9255), .ZN(n9249) );
  AND2_X1 U10651 ( .A1(n9250), .A2(n9249), .ZN(n9360) );
  AOI21_X1 U10652 ( .B1(n9251), .B2(n9360), .A(n5048), .ZN(n9261) );
  AND2_X1 U10653 ( .A1(n9364), .A2(n9257), .ZN(n9259) );
  INV_X1 U10654 ( .A(n9366), .ZN(n9263) );
  OAI21_X1 U10655 ( .B1(n9269), .B2(n9263), .A(n9262), .ZN(n9264) );
  AND2_X1 U10656 ( .A1(n9274), .A2(n9276), .ZN(n9369) );
  NAND3_X1 U10657 ( .A1(n9264), .A2(n9369), .A3(n9365), .ZN(n9267) );
  INV_X1 U10658 ( .A(n9271), .ZN(n9265) );
  NAND2_X1 U10659 ( .A1(n9274), .A2(n9265), .ZN(n9266) );
  INV_X1 U10660 ( .A(n9440), .ZN(n9798) );
  OAI211_X1 U10661 ( .C1(n9269), .C2(n9268), .A(n9798), .B(n9366), .ZN(n9273)
         );
  AND2_X1 U10662 ( .A1(n9271), .A2(n9270), .ZN(n9272) );
  AND2_X1 U10663 ( .A1(n9742), .A2(n9272), .ZN(n9372) );
  NAND2_X1 U10664 ( .A1(n9273), .A2(n9372), .ZN(n9275) );
  OAI211_X1 U10665 ( .C1(n9277), .C2(n9276), .A(n9275), .B(n9274), .ZN(n9278)
         );
  NAND2_X1 U10666 ( .A1(n9280), .A2(n9282), .ZN(n9377) );
  AND2_X1 U10667 ( .A1(n9282), .A2(n9281), .ZN(n9375) );
  AOI21_X1 U10668 ( .B1(n9900), .B2(n9323), .A(n9996), .ZN(n9287) );
  AOI21_X1 U10669 ( .B1(n9330), .B2(n9477), .A(n9720), .ZN(n9286) );
  NAND2_X1 U10670 ( .A1(n9284), .A2(n9283), .ZN(n9373) );
  NAND2_X1 U10671 ( .A1(n9373), .A2(n9323), .ZN(n9285) );
  OAI22_X1 U10672 ( .A1(n9287), .A2(n9286), .B1(n9377), .B2(n9285), .ZN(n9290)
         );
  NAND2_X1 U10673 ( .A1(n9685), .A2(n9288), .ZN(n9289) );
  OAI21_X1 U10674 ( .B1(n9295), .B2(n9292), .A(n9291), .ZN(n9294) );
  INV_X1 U10675 ( .A(n9344), .ZN(n9293) );
  NAND2_X1 U10676 ( .A1(n9296), .A2(n9380), .ZN(n9299) );
  NAND2_X1 U10677 ( .A1(n9673), .A2(n9300), .ZN(n9301) );
  NAND2_X1 U10678 ( .A1(n9423), .A2(n9301), .ZN(n9384) );
  INV_X1 U10679 ( .A(n9343), .ZN(n9304) );
  INV_X1 U10680 ( .A(n9387), .ZN(n9303) );
  MUX2_X1 U10681 ( .A(n9304), .B(n9303), .S(n9323), .Z(n9305) );
  NAND2_X1 U10682 ( .A1(n9307), .A2(n9388), .ZN(n9306) );
  OR2_X1 U10683 ( .A1(n9866), .A2(n4402), .ZN(n9341) );
  NAND3_X1 U10684 ( .A1(n9581), .A2(n9330), .A3(n9388), .ZN(n9310) );
  NAND2_X1 U10685 ( .A1(n9309), .A2(n9308), .ZN(n9393) );
  OAI21_X1 U10686 ( .B1(n9323), .B2(n9341), .A(n9342), .ZN(n9311) );
  NAND2_X1 U10687 ( .A1(n9393), .A2(n9323), .ZN(n9312) );
  OAI211_X1 U10688 ( .C1(n9330), .C2(n9581), .A(n9312), .B(n9394), .ZN(n9313)
         );
  OAI21_X1 U10689 ( .B1(n9393), .B2(n9342), .A(n9394), .ZN(n9315) );
  INV_X1 U10690 ( .A(n9339), .ZN(n9318) );
  INV_X1 U10691 ( .A(n9338), .ZN(n9474) );
  NAND3_X1 U10692 ( .A1(n9474), .A2(n9330), .A3(n9419), .ZN(n9322) );
  INV_X1 U10693 ( .A(n9855), .ZN(n9976) );
  NAND3_X1 U10694 ( .A1(n9976), .A2(n9330), .A3(n9339), .ZN(n9317) );
  NAND2_X1 U10695 ( .A1(n9447), .A2(n9323), .ZN(n9316) );
  OAI211_X1 U10696 ( .C1(n9318), .C2(n9322), .A(n9317), .B(n9316), .ZN(n9320)
         );
  NOR2_X1 U10697 ( .A1(n9855), .A2(n9338), .ZN(n9336) );
  OAI21_X1 U10698 ( .B1(n9336), .B2(n9563), .A(n9331), .ZN(n9319) );
  INV_X1 U10699 ( .A(n9322), .ZN(n9326) );
  NAND3_X1 U10700 ( .A1(n9338), .A2(n9323), .A3(n9419), .ZN(n9324) );
  NAND2_X1 U10701 ( .A1(n9855), .A2(n9324), .ZN(n9325) );
  OAI21_X1 U10702 ( .B1(n9855), .B2(n9326), .A(n9325), .ZN(n9327) );
  AOI21_X1 U10703 ( .B1(n9330), .B2(n9329), .A(n9466), .ZN(n9473) );
  INV_X1 U10704 ( .A(n9456), .ZN(n9334) );
  NOR2_X1 U10705 ( .A1(n9405), .A2(n9332), .ZN(n9333) );
  OAI211_X1 U10706 ( .C1(n4512), .C2(n5869), .A(n9334), .B(n9333), .ZN(n9472)
         );
  INV_X1 U10707 ( .A(n9336), .ZN(n9337) );
  NAND2_X1 U10708 ( .A1(n9420), .A2(n9337), .ZN(n9451) );
  NAND2_X1 U10709 ( .A1(n9855), .A2(n9338), .ZN(n9340) );
  NAND2_X1 U10710 ( .A1(n9340), .A2(n9339), .ZN(n9450) );
  INV_X1 U10711 ( .A(n9450), .ZN(n9397) );
  NAND2_X1 U10712 ( .A1(n9342), .A2(n9341), .ZN(n9411) );
  INV_X1 U10713 ( .A(n9411), .ZN(n9383) );
  OAI21_X1 U10714 ( .B1(n9344), .B2(n9631), .A(n9343), .ZN(n9345) );
  NAND2_X1 U10715 ( .A1(n9345), .A2(n9387), .ZN(n9346) );
  AND2_X1 U10716 ( .A1(n9347), .A2(n9346), .ZN(n9391) );
  INV_X1 U10717 ( .A(n9391), .ZN(n9413) );
  OAI21_X1 U10718 ( .B1(n6922), .B2(n9349), .A(n9348), .ZN(n9352) );
  NAND2_X1 U10719 ( .A1(n9350), .A2(n9464), .ZN(n9351) );
  NOR2_X1 U10720 ( .A1(n9352), .A2(n9351), .ZN(n9356) );
  AND4_X1 U10721 ( .A1(n9356), .A2(n9355), .A3(n9354), .A4(n9353), .ZN(n9358)
         );
  OAI21_X1 U10722 ( .B1(n9359), .B2(n9358), .A(n9357), .ZN(n9363) );
  INV_X1 U10723 ( .A(n9360), .ZN(n9361) );
  AOI21_X1 U10724 ( .B1(n9363), .B2(n9362), .A(n9361), .ZN(n9368) );
  NAND2_X1 U10725 ( .A1(n9799), .A2(n9364), .ZN(n9367) );
  OAI211_X1 U10726 ( .C1(n9368), .C2(n9367), .A(n9366), .B(n9365), .ZN(n9371)
         );
  INV_X1 U10727 ( .A(n9369), .ZN(n9370) );
  AOI22_X1 U10728 ( .A1(n9372), .A2(n9371), .B1(n9370), .B2(n9742), .ZN(n9374)
         );
  AOI21_X1 U10729 ( .B1(n9375), .B2(n9374), .A(n9373), .ZN(n9378) );
  OAI21_X1 U10730 ( .B1(n9378), .B2(n9377), .A(n9376), .ZN(n9379) );
  NAND2_X1 U10731 ( .A1(n9380), .A2(n9379), .ZN(n9381) );
  OAI21_X1 U10732 ( .B1(n9413), .B2(n9381), .A(n9581), .ZN(n9382) );
  INV_X1 U10733 ( .A(n9384), .ZN(n9386) );
  NAND3_X1 U10734 ( .A1(n9387), .A2(n9386), .A3(n9385), .ZN(n9390) );
  INV_X1 U10735 ( .A(n9388), .ZN(n9389) );
  AOI21_X1 U10736 ( .B1(n9391), .B2(n9390), .A(n9389), .ZN(n9392) );
  OAI21_X1 U10737 ( .B1(n9395), .B2(n9414), .A(n4483), .ZN(n9396) );
  AND2_X1 U10738 ( .A1(n9397), .A2(n9396), .ZN(n9398) );
  NAND2_X1 U10739 ( .A1(n9399), .A2(n4512), .ZN(n9409) );
  INV_X1 U10740 ( .A(n9409), .ZN(n9462) );
  OR3_X1 U10741 ( .A1(n9456), .A2(n5869), .A3(n9400), .ZN(n9408) );
  NAND2_X1 U10742 ( .A1(n9402), .A2(n9401), .ZN(n9403) );
  NOR2_X1 U10743 ( .A1(n9404), .A2(n9403), .ZN(n9407) );
  OAI21_X1 U10744 ( .B1(n9456), .B2(n9405), .A(P1_B_REG_SCAN_IN), .ZN(n9406)
         );
  OAI22_X1 U10745 ( .A1(n9409), .A2(n9408), .B1(n9407), .B2(n9406), .ZN(n9410)
         );
  INV_X1 U10746 ( .A(n9410), .ZN(n9461) );
  OAI21_X1 U10747 ( .B1(n9413), .B2(n9412), .A(n9581), .ZN(n9415) );
  NAND2_X1 U10748 ( .A1(n9474), .A2(n9419), .ZN(n9416) );
  OAI22_X1 U10749 ( .A1(n9417), .A2(n9450), .B1(n9855), .B2(n9416), .ZN(n9418)
         );
  OAI211_X1 U10750 ( .C1(n9976), .C2(n9419), .A(n9418), .B(n4512), .ZN(n9422)
         );
  NAND3_X1 U10751 ( .A1(n9422), .A2(n9421), .A3(n9420), .ZN(n9458) );
  NAND2_X1 U10752 ( .A1(n9424), .A2(n9423), .ZN(n9653) );
  INV_X1 U10753 ( .A(n9710), .ZN(n9715) );
  INV_X1 U10754 ( .A(n9775), .ZN(n9773) );
  INV_X1 U10755 ( .A(n9425), .ZN(n9436) );
  NOR4_X1 U10756 ( .A1(n6970), .A2(n9427), .A3(n9426), .A4(n9464), .ZN(n9430)
         );
  NAND3_X1 U10757 ( .A1(n9430), .A2(n9429), .A3(n9428), .ZN(n9434) );
  NOR4_X1 U10758 ( .A1(n9434), .A2(n9433), .A3(n9432), .A4(n9431), .ZN(n9435)
         );
  NAND4_X1 U10759 ( .A1(n4940), .A2(n9437), .A3(n9436), .A4(n9435), .ZN(n9438)
         );
  NOR4_X1 U10760 ( .A1(n9440), .A2(n9820), .A3(n9439), .A4(n9438), .ZN(n9441)
         );
  NAND4_X1 U10761 ( .A1(n9747), .A2(n9766), .A3(n9773), .A4(n9441), .ZN(n9442)
         );
  NOR4_X1 U10762 ( .A1(n9653), .A2(n9731), .A3(n9715), .A4(n9442), .ZN(n9443)
         );
  XNOR2_X1 U10763 ( .A(n9896), .B(n9702), .ZN(n9687) );
  XNOR2_X1 U10764 ( .A(n9903), .B(n9712), .ZN(n9699) );
  NAND4_X1 U10765 ( .A1(n9443), .A2(n9667), .A3(n9687), .A4(n9699), .ZN(n9444)
         );
  NOR4_X1 U10766 ( .A1(n9586), .A2(n9445), .A3(n9636), .A4(n9444), .ZN(n9454)
         );
  INV_X1 U10767 ( .A(n9604), .ZN(n9448) );
  NAND3_X1 U10768 ( .A1(n9448), .A2(n9447), .A3(n9446), .ZN(n9449) );
  NOR2_X1 U10769 ( .A1(n9450), .A2(n9449), .ZN(n9453) );
  INV_X1 U10770 ( .A(n9451), .ZN(n9452) );
  NAND4_X1 U10771 ( .A1(n4512), .A2(n9454), .A3(n9453), .A4(n9452), .ZN(n9467)
         );
  NOR2_X1 U10772 ( .A1(n9456), .A2(n9455), .ZN(n9468) );
  INV_X1 U10773 ( .A(n9468), .ZN(n9457) );
  AOI211_X1 U10774 ( .C1(n9458), .C2(n9467), .A(n9556), .B(n9457), .ZN(n9459)
         );
  INV_X1 U10775 ( .A(n9459), .ZN(n9460) );
  INV_X1 U10776 ( .A(n9463), .ZN(n9471) );
  OAI21_X1 U10777 ( .B1(n9466), .B2(n9465), .A(n9464), .ZN(n9469) );
  NAND4_X1 U10778 ( .A1(n9469), .A2(n9556), .A3(n9468), .A4(n9467), .ZN(n9470)
         );
  OAI211_X1 U10779 ( .C1(n9473), .C2(n9472), .A(n9471), .B(n9470), .ZN(
        P1_U3242) );
  MUX2_X1 U10780 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9474), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10781 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9475), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10782 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9584), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10783 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9476), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10784 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n4412), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10785 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9633), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10786 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9650), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10787 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9688), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10788 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9702), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10789 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9477), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10790 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9744), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10791 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9767), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10792 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9780), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10793 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9803), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10794 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9779), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10795 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9478), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10796 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9479), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10797 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9480), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10798 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9481), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10799 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9482), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10800 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n5051), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10801 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9483), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10802 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9484), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10803 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9485), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10804 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9486), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10805 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9487), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10806 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9489), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10807 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9490), .S(P1_U3973), .Z(
        P1_U3555) );
  OAI211_X1 U10808 ( .C1(n9493), .C2(n9492), .A(n10127), .B(n9491), .ZN(n9501)
         );
  OAI211_X1 U10809 ( .C1(n9496), .C2(n9495), .A(n10131), .B(n9494), .ZN(n9500)
         );
  AOI22_X1 U10810 ( .A1(n10089), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9499) );
  NAND2_X1 U10811 ( .A1(n10146), .A2(n9497), .ZN(n9498) );
  NAND4_X1 U10812 ( .A1(n9501), .A2(n9500), .A3(n9499), .A4(n9498), .ZN(
        P1_U3244) );
  OAI21_X1 U10813 ( .B1(n9504), .B2(n9503), .A(n9502), .ZN(n9505) );
  NAND2_X1 U10814 ( .A1(n9505), .A2(n10127), .ZN(n9516) );
  OAI21_X1 U10815 ( .B1(n9508), .B2(n9507), .A(n9506), .ZN(n9509) );
  NAND2_X1 U10816 ( .A1(n9509), .A2(n10131), .ZN(n9515) );
  INV_X1 U10817 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9510) );
  NOR2_X1 U10818 ( .A1(n10148), .A2(n9510), .ZN(n9511) );
  AOI211_X1 U10819 ( .C1(n9513), .C2(n10146), .A(n9512), .B(n9511), .ZN(n9514)
         );
  NAND3_X1 U10820 ( .A1(n9516), .A2(n9515), .A3(n9514), .ZN(P1_U3255) );
  XNOR2_X1 U10821 ( .A(n9535), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9518) );
  AOI211_X1 U10822 ( .C1(n9519), .C2(n9518), .A(n10137), .B(n9532), .ZN(n9531)
         );
  INV_X1 U10823 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9522) );
  MUX2_X1 U10824 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n9522), .S(n9535), .Z(n9523) );
  INV_X1 U10825 ( .A(n9523), .ZN(n9524) );
  AOI211_X1 U10826 ( .C1(n9525), .C2(n9524), .A(n10141), .B(n9534), .ZN(n9530)
         );
  INV_X1 U10827 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9528) );
  NAND2_X1 U10828 ( .A1(n10146), .A2(n9535), .ZN(n9527) );
  OAI211_X1 U10829 ( .C1(n9528), .C2(n10148), .A(n9527), .B(n9526), .ZN(n9529)
         );
  OR3_X1 U10830 ( .A1(n9531), .A2(n9530), .A3(n9529), .ZN(P1_U3257) );
  AOI211_X1 U10831 ( .C1(n9533), .C2(n10572), .A(n10137), .B(n9544), .ZN(n9542) );
  AOI211_X1 U10832 ( .C1(n9787), .C2(n9536), .A(n10141), .B(n9548), .ZN(n9541)
         );
  INV_X1 U10833 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9539) );
  NAND2_X1 U10834 ( .A1(n10146), .A2(n9549), .ZN(n9538) );
  OAI211_X1 U10835 ( .C1(n9539), .C2(n10148), .A(n9538), .B(n9537), .ZN(n9540)
         );
  OR3_X1 U10836 ( .A1(n9542), .A2(n9541), .A3(n9540), .ZN(P1_U3258) );
  NAND2_X1 U10837 ( .A1(n10145), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9545) );
  OAI21_X1 U10838 ( .B1(n10145), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9545), .ZN(
        n10139) );
  INV_X1 U10839 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9922) );
  XNOR2_X1 U10840 ( .A(n10128), .B(n9922), .ZN(n10121) );
  XNOR2_X1 U10841 ( .A(n9550), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n10114) );
  NAND2_X1 U10842 ( .A1(n10136), .A2(n9545), .ZN(n9546) );
  NOR2_X1 U10843 ( .A1(n10128), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9551) );
  AOI21_X1 U10844 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n10128), .A(n9551), .ZN(
        n10125) );
  AOI22_X1 U10845 ( .A1(n10112), .A2(n5778), .B1(P1_REG2_REG_16__SCAN_IN), 
        .B2(n9550), .ZN(n10109) );
  INV_X1 U10846 ( .A(n9551), .ZN(n9552) );
  INV_X1 U10847 ( .A(n10143), .ZN(n9554) );
  NAND2_X1 U10848 ( .A1(n10145), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9555) );
  OAI21_X1 U10849 ( .B1(n10145), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9555), .ZN(
        n10142) );
  INV_X1 U10850 ( .A(n10142), .ZN(n9553) );
  OAI21_X1 U10851 ( .B1(n9557), .B2(n10141), .A(n10100), .ZN(n9558) );
  NOR2_X2 U10852 ( .A1(n9855), .A2(n9566), .ZN(n9567) );
  XNOR2_X1 U10853 ( .A(n9972), .B(n9567), .ZN(n9561) );
  NAND2_X1 U10854 ( .A1(n9850), .A2(n9807), .ZN(n9565) );
  NOR2_X1 U10855 ( .A1(n9563), .A2(n9562), .ZN(n9849) );
  INV_X1 U10856 ( .A(n9849), .ZN(n9853) );
  NOR2_X1 U10857 ( .A1(n9853), .A2(n9827), .ZN(n9569) );
  AOI21_X1 U10858 ( .B1(n9827), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9569), .ZN(
        n9564) );
  OAI211_X1 U10859 ( .C1(n9972), .C2(n9763), .A(n9565), .B(n9564), .ZN(
        P1_U3263) );
  NOR2_X1 U10860 ( .A1(n9842), .A2(n9568), .ZN(n9570) );
  AOI211_X1 U10861 ( .C1(n9855), .C2(n9837), .A(n9570), .B(n9569), .ZN(n9571)
         );
  OAI21_X1 U10862 ( .B1(n9854), .B2(n9840), .A(n9571), .ZN(P1_U3264) );
  NAND2_X1 U10863 ( .A1(n9572), .A2(n9847), .ZN(n9580) );
  AOI22_X1 U10864 ( .A1(n9573), .A2(n9836), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9827), .ZN(n9574) );
  OAI21_X1 U10865 ( .B1(n9609), .B2(n9829), .A(n9574), .ZN(n9577) );
  NOR2_X1 U10866 ( .A1(n9575), .A2(n9840), .ZN(n9576) );
  AOI211_X1 U10867 ( .C1(n9837), .C2(n9578), .A(n9577), .B(n9576), .ZN(n9579)
         );
  OAI211_X1 U10868 ( .C1(n5380), .C2(n9827), .A(n9580), .B(n9579), .ZN(
        P1_U3265) );
  NAND2_X1 U10869 ( .A1(n9606), .A2(n9581), .ZN(n9583) );
  XNOR2_X1 U10870 ( .A(n9583), .B(n9582), .ZN(n9585) );
  AOI22_X1 U10871 ( .A1(n9585), .A2(n9782), .B1(n9804), .B2(n9584), .ZN(n9862)
         );
  XNOR2_X1 U10872 ( .A(n9587), .B(n9586), .ZN(n9858) );
  NAND2_X1 U10873 ( .A1(n9858), .A2(n9847), .ZN(n9596) );
  AOI22_X1 U10874 ( .A1(n9588), .A2(n9836), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9827), .ZN(n9589) );
  OAI21_X1 U10875 ( .B1(n4402), .B2(n9829), .A(n9589), .ZN(n9594) );
  NAND2_X1 U10876 ( .A1(n9590), .A2(n9859), .ZN(n9591) );
  NAND3_X1 U10877 ( .A1(n9592), .A2(n9784), .A3(n9591), .ZN(n9860) );
  NOR2_X1 U10878 ( .A1(n9860), .A2(n9840), .ZN(n9593) );
  AOI211_X1 U10879 ( .C1(n9837), .C2(n9859), .A(n9594), .B(n9593), .ZN(n9595)
         );
  OAI211_X1 U10880 ( .C1(n9862), .C2(n9827), .A(n9596), .B(n9595), .ZN(
        P1_U3266) );
  XNOR2_X1 U10881 ( .A(n9597), .B(n9604), .ZN(n9867) );
  INV_X1 U10882 ( .A(n9598), .ZN(n9619) );
  INV_X1 U10883 ( .A(n9590), .ZN(n9599) );
  AOI211_X1 U10884 ( .C1(n9866), .C2(n9619), .A(n9822), .B(n9599), .ZN(n9865)
         );
  NOR2_X1 U10885 ( .A1(n9600), .A2(n9763), .ZN(n9603) );
  OAI22_X1 U10886 ( .A1(n9601), .A2(n9785), .B1(n10339), .B2(n9842), .ZN(n9602) );
  AOI211_X1 U10887 ( .C1(n9865), .C2(n9807), .A(n9603), .B(n9602), .ZN(n9613)
         );
  OAI22_X1 U10888 ( .A1(n9609), .A2(n9815), .B1(n9943), .B2(n9608), .ZN(n9610)
         );
  NAND2_X1 U10889 ( .A1(n9864), .A2(n9842), .ZN(n9612) );
  OAI211_X1 U10890 ( .C1(n9867), .C2(n9809), .A(n9613), .B(n9612), .ZN(
        P1_U3267) );
  XOR2_X1 U10891 ( .A(n9616), .B(n9614), .Z(n9872) );
  INV_X1 U10892 ( .A(n9872), .ZN(n9629) );
  OAI211_X1 U10893 ( .C1(n9617), .C2(n9616), .A(n9615), .B(n9782), .ZN(n9618)
         );
  OAI21_X1 U10894 ( .B1(n4402), .B2(n9815), .A(n9618), .ZN(n9871) );
  INV_X1 U10895 ( .A(n9641), .ZN(n9620) );
  OAI211_X1 U10896 ( .C1(n9982), .C2(n9620), .A(n9619), .B(n9784), .ZN(n9868)
         );
  NOR2_X1 U10897 ( .A1(n9869), .A2(n9829), .ZN(n9624) );
  OAI22_X1 U10898 ( .A1(n9622), .A2(n9785), .B1(n9621), .B2(n9842), .ZN(n9623)
         );
  AOI211_X1 U10899 ( .C1(n9625), .C2(n9837), .A(n9624), .B(n9623), .ZN(n9626)
         );
  OAI21_X1 U10900 ( .B1(n9868), .B2(n9840), .A(n9626), .ZN(n9627) );
  AOI21_X1 U10901 ( .B1(n9842), .B2(n9871), .A(n9627), .ZN(n9628) );
  OAI21_X1 U10902 ( .B1(n9629), .B2(n9809), .A(n9628), .ZN(P1_U3268) );
  NAND2_X1 U10903 ( .A1(n5382), .A2(n9630), .ZN(n9647) );
  NOR2_X1 U10904 ( .A1(n9647), .A2(n9653), .ZN(n9649) );
  NOR2_X1 U10905 ( .A1(n9649), .A2(n9631), .ZN(n9632) );
  XNOR2_X1 U10906 ( .A(n9632), .B(n9636), .ZN(n9634) );
  AOI22_X1 U10907 ( .A1(n9634), .A2(n9782), .B1(n9804), .B2(n9633), .ZN(n9880)
         );
  XOR2_X1 U10908 ( .A(n9635), .B(n9636), .Z(n9875) );
  NAND2_X1 U10909 ( .A1(n9875), .A2(n9847), .ZN(n9646) );
  AOI22_X1 U10910 ( .A1(n9637), .A2(n9836), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9827), .ZN(n9638) );
  OAI21_X1 U10911 ( .B1(n9639), .B2(n9829), .A(n9638), .ZN(n9644) );
  AOI21_X1 U10912 ( .B1(n9640), .B2(n6980), .A(n9822), .ZN(n9642) );
  NAND2_X1 U10913 ( .A1(n9642), .A2(n9641), .ZN(n9878) );
  NOR2_X1 U10914 ( .A1(n9878), .A2(n9840), .ZN(n9643) );
  AOI211_X1 U10915 ( .C1(n9837), .C2(n6980), .A(n9644), .B(n9643), .ZN(n9645)
         );
  OAI211_X1 U10916 ( .C1(n9827), .C2(n9880), .A(n9646), .B(n9645), .ZN(
        P1_U3269) );
  AND2_X1 U10917 ( .A1(n9647), .A2(n9653), .ZN(n9648) );
  OAI21_X1 U10918 ( .B1(n9649), .B2(n9648), .A(n9782), .ZN(n9652) );
  AOI22_X1 U10919 ( .A1(n9650), .A2(n9804), .B1(n9877), .B2(n9688), .ZN(n9651)
         );
  NAND2_X1 U10920 ( .A1(n9652), .A2(n9651), .ZN(n9882) );
  INV_X1 U10921 ( .A(n9882), .ZN(n9663) );
  XNOR2_X1 U10922 ( .A(n9654), .B(n9653), .ZN(n9884) );
  NAND2_X1 U10923 ( .A1(n9884), .A2(n9847), .ZN(n9662) );
  INV_X1 U10924 ( .A(n9640), .ZN(n9655) );
  AOI211_X1 U10925 ( .C1(n9656), .C2(n4449), .A(n9822), .B(n9655), .ZN(n9883)
         );
  NOR2_X1 U10926 ( .A1(n5012), .A2(n9763), .ZN(n9660) );
  OAI22_X1 U10927 ( .A1(n9658), .A2(n9785), .B1(n9657), .B2(n9842), .ZN(n9659)
         );
  AOI211_X1 U10928 ( .C1(n9883), .C2(n9807), .A(n9660), .B(n9659), .ZN(n9661)
         );
  OAI211_X1 U10929 ( .C1(n9827), .C2(n9663), .A(n9662), .B(n9661), .ZN(
        P1_U3270) );
  XNOR2_X1 U10930 ( .A(n9664), .B(n9667), .ZN(n9665) );
  AOI22_X1 U10931 ( .A1(n9665), .A2(n9782), .B1(n9804), .B2(n9876), .ZN(n9887)
         );
  XNOR2_X1 U10932 ( .A(n9666), .B(n9667), .ZN(n9890) );
  NAND2_X1 U10933 ( .A1(n9890), .A2(n9847), .ZN(n9675) );
  INV_X1 U10934 ( .A(n9668), .ZN(n9669) );
  AOI22_X1 U10935 ( .A1(n9669), .A2(n9836), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9827), .ZN(n9670) );
  OAI21_X1 U10936 ( .B1(n9888), .B2(n9829), .A(n9670), .ZN(n9672) );
  OAI211_X1 U10937 ( .C1(n9990), .C2(n9677), .A(n4449), .B(n9784), .ZN(n9886)
         );
  NOR2_X1 U10938 ( .A1(n9886), .A2(n9840), .ZN(n9671) );
  AOI211_X1 U10939 ( .C1(n9837), .C2(n9673), .A(n9672), .B(n9671), .ZN(n9674)
         );
  OAI211_X1 U10940 ( .C1(n9827), .C2(n9887), .A(n9675), .B(n9674), .ZN(
        P1_U3271) );
  XNOR2_X1 U10941 ( .A(n9676), .B(n9687), .ZN(n9899) );
  AOI211_X1 U10942 ( .C1(n9896), .C2(n9695), .A(n9822), .B(n9677), .ZN(n9894)
         );
  INV_X1 U10943 ( .A(n9896), .ZN(n9683) );
  OAI22_X1 U10944 ( .A1(n9679), .A2(n9785), .B1(n9678), .B2(n9842), .ZN(n9680)
         );
  AOI21_X1 U10945 ( .B1(n9681), .B2(n9712), .A(n9680), .ZN(n9682) );
  OAI21_X1 U10946 ( .B1(n9683), .B2(n9763), .A(n9682), .ZN(n9691) );
  INV_X1 U10947 ( .A(n9701), .ZN(n9684) );
  NAND2_X1 U10948 ( .A1(n9684), .A2(n9699), .ZN(n9704) );
  NAND2_X1 U10949 ( .A1(n9704), .A2(n9685), .ZN(n9686) );
  XOR2_X1 U10950 ( .A(n9687), .B(n9686), .Z(n9689) );
  AOI22_X1 U10951 ( .A1(n9689), .A2(n9782), .B1(n9804), .B2(n9688), .ZN(n9898)
         );
  NOR2_X1 U10952 ( .A1(n9898), .A2(n9827), .ZN(n9690) );
  AOI211_X1 U10953 ( .C1(n9894), .C2(n9807), .A(n9691), .B(n9690), .ZN(n9692)
         );
  OAI21_X1 U10954 ( .B1(n9809), .B2(n9899), .A(n9692), .ZN(P1_U3272) );
  XOR2_X1 U10955 ( .A(n9693), .B(n9699), .Z(n9906) );
  AOI211_X1 U10956 ( .C1(n9903), .C2(n9694), .A(n9822), .B(n5193), .ZN(n9901)
         );
  NAND2_X1 U10957 ( .A1(n9903), .A2(n9837), .ZN(n9698) );
  AOI22_X1 U10958 ( .A1(n9696), .A2(n9836), .B1(P1_REG2_REG_20__SCAN_IN), .B2(
        n9827), .ZN(n9697) );
  OAI211_X1 U10959 ( .C1(n9900), .C2(n9829), .A(n9698), .B(n9697), .ZN(n9706)
         );
  INV_X1 U10960 ( .A(n9699), .ZN(n9700) );
  AOI21_X1 U10961 ( .B1(n9701), .B2(n9700), .A(n9817), .ZN(n9703) );
  AOI22_X1 U10962 ( .A1(n9704), .A2(n9703), .B1(n9804), .B2(n9702), .ZN(n9905)
         );
  NOR2_X1 U10963 ( .A1(n9905), .A2(n9827), .ZN(n9705) );
  AOI211_X1 U10964 ( .C1(n9901), .C2(n9807), .A(n9706), .B(n9705), .ZN(n9707)
         );
  OAI21_X1 U10965 ( .B1(n9906), .B2(n9809), .A(n9707), .ZN(P1_U3273) );
  OAI21_X1 U10966 ( .B1(n9710), .B2(n9709), .A(n9708), .ZN(n9711) );
  NAND2_X1 U10967 ( .A1(n9711), .A2(n9782), .ZN(n9714) );
  AOI22_X1 U10968 ( .A1(n9712), .A2(n9804), .B1(n9877), .B2(n9744), .ZN(n9713)
         );
  NAND2_X1 U10969 ( .A1(n9714), .A2(n9713), .ZN(n9907) );
  INV_X1 U10970 ( .A(n9907), .ZN(n9727) );
  XNOR2_X1 U10971 ( .A(n9716), .B(n9715), .ZN(n9909) );
  NAND2_X1 U10972 ( .A1(n9909), .A2(n9847), .ZN(n9726) );
  INV_X1 U10973 ( .A(n9717), .ZN(n9719) );
  INV_X1 U10974 ( .A(n9694), .ZN(n9718) );
  AOI211_X1 U10975 ( .C1(n9720), .C2(n9719), .A(n9822), .B(n9718), .ZN(n9908)
         );
  NOR2_X1 U10976 ( .A1(n9996), .A2(n9763), .ZN(n9724) );
  OAI22_X1 U10977 ( .A1(n9722), .A2(n9785), .B1(n9721), .B2(n9842), .ZN(n9723)
         );
  AOI211_X1 U10978 ( .C1(n9908), .C2(n9807), .A(n9724), .B(n9723), .ZN(n9725)
         );
  OAI211_X1 U10979 ( .C1(n9827), .C2(n9727), .A(n9726), .B(n9725), .ZN(
        P1_U3274) );
  XNOR2_X1 U10980 ( .A(n9728), .B(n9731), .ZN(n9916) );
  INV_X1 U10981 ( .A(n9729), .ZN(n9730) );
  AOI21_X1 U10982 ( .B1(n9732), .B2(n9731), .A(n9730), .ZN(n9733) );
  OAI222_X1 U10983 ( .A1(n9815), .A2(n9900), .B1(n9943), .B2(n9734), .C1(n9817), .C2(n9733), .ZN(n9912) );
  INV_X1 U10984 ( .A(n9735), .ZN(n9752) );
  AOI211_X1 U10985 ( .C1(n9914), .C2(n9752), .A(n9822), .B(n9717), .ZN(n9913)
         );
  NAND2_X1 U10986 ( .A1(n9913), .A2(n9807), .ZN(n9738) );
  AOI22_X1 U10987 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n9827), .B1(n9736), .B2(
        n9836), .ZN(n9737) );
  OAI211_X1 U10988 ( .C1(n9739), .C2(n9763), .A(n9738), .B(n9737), .ZN(n9740)
         );
  AOI21_X1 U10989 ( .B1(n9912), .B2(n9842), .A(n9740), .ZN(n9741) );
  OAI21_X1 U10990 ( .B1(n9809), .B2(n9916), .A(n9741), .ZN(P1_U3275) );
  NAND2_X1 U10991 ( .A1(n9764), .A2(n9742), .ZN(n9743) );
  XNOR2_X1 U10992 ( .A(n9743), .B(n9747), .ZN(n9745) );
  AOI22_X1 U10993 ( .A1(n9745), .A2(n9782), .B1(n9804), .B2(n9744), .ZN(n9918)
         );
  XNOR2_X1 U10994 ( .A(n9746), .B(n9747), .ZN(n9921) );
  NAND2_X1 U10995 ( .A1(n9921), .A2(n9847), .ZN(n9757) );
  INV_X1 U10996 ( .A(n9748), .ZN(n9749) );
  AOI22_X1 U10997 ( .A1(n9827), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9749), .B2(
        n9836), .ZN(n9750) );
  OAI21_X1 U10998 ( .B1(n9919), .B2(n9829), .A(n9750), .ZN(n9754) );
  INV_X1 U10999 ( .A(n9755), .ZN(n10001) );
  INV_X1 U11000 ( .A(n9751), .ZN(n9760) );
  OAI211_X1 U11001 ( .C1(n10001), .C2(n9760), .A(n9752), .B(n9784), .ZN(n9917)
         );
  NOR2_X1 U11002 ( .A1(n9917), .A2(n9840), .ZN(n9753) );
  AOI211_X1 U11003 ( .C1(n9837), .C2(n9755), .A(n9754), .B(n9753), .ZN(n9756)
         );
  OAI211_X1 U11004 ( .C1(n9827), .C2(n9918), .A(n9757), .B(n9756), .ZN(
        P1_U3276) );
  XNOR2_X1 U11005 ( .A(n9758), .B(n9759), .ZN(n9928) );
  AOI211_X1 U11006 ( .C1(n9925), .C2(n9783), .A(n9822), .B(n9760), .ZN(n9924)
         );
  AOI22_X1 U11007 ( .A1(n9827), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9761), .B2(
        n9836), .ZN(n9762) );
  OAI21_X1 U11008 ( .B1(n5187), .B2(n9763), .A(n9762), .ZN(n9770) );
  OAI21_X1 U11009 ( .B1(n9766), .B2(n9765), .A(n9764), .ZN(n9768) );
  AOI222_X1 U11010 ( .A1(n9782), .A2(n9768), .B1(n9803), .B2(n9877), .C1(n9767), .C2(n9804), .ZN(n9927) );
  NOR2_X1 U11011 ( .A1(n9927), .A2(n9827), .ZN(n9769) );
  AOI211_X1 U11012 ( .C1(n9924), .C2(n9807), .A(n9770), .B(n9769), .ZN(n9771)
         );
  OAI21_X1 U11013 ( .B1(n9809), .B2(n9928), .A(n9771), .ZN(P1_U3277) );
  XNOR2_X1 U11014 ( .A(n9772), .B(n9773), .ZN(n9931) );
  INV_X1 U11015 ( .A(n9774), .ZN(n9801) );
  OAI21_X1 U11016 ( .B1(n9801), .B2(n9776), .A(n9775), .ZN(n9778) );
  NAND2_X1 U11017 ( .A1(n9778), .A2(n9777), .ZN(n9781) );
  AOI222_X1 U11018 ( .A1(n9782), .A2(n9781), .B1(n9780), .B2(n9804), .C1(n9779), .C2(n9877), .ZN(n9930) );
  INV_X1 U11019 ( .A(n9930), .ZN(n9792) );
  OAI211_X1 U11020 ( .C1(n4537), .C2(n10006), .A(n9784), .B(n9783), .ZN(n9929)
         );
  OAI22_X1 U11021 ( .A1(n9842), .A2(n9787), .B1(n9786), .B2(n9785), .ZN(n9788)
         );
  AOI21_X1 U11022 ( .B1(n9789), .B2(n9837), .A(n9788), .ZN(n9790) );
  OAI21_X1 U11023 ( .B1(n9929), .B2(n9840), .A(n9790), .ZN(n9791) );
  AOI21_X1 U11024 ( .B1(n9792), .B2(n9842), .A(n9791), .ZN(n9793) );
  OAI21_X1 U11025 ( .B1(n9931), .B2(n9809), .A(n9793), .ZN(P1_U3278) );
  XNOR2_X1 U11026 ( .A(n9794), .B(n9798), .ZN(n9940) );
  AOI211_X1 U11027 ( .C1(n9937), .C2(n9824), .A(n9822), .B(n4537), .ZN(n9935)
         );
  NAND2_X1 U11028 ( .A1(n9937), .A2(n9837), .ZN(n9797) );
  AOI22_X1 U11029 ( .A1(n9827), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9795), .B2(
        n9836), .ZN(n9796) );
  OAI211_X1 U11030 ( .C1(n9934), .C2(n9829), .A(n9797), .B(n9796), .ZN(n9806)
         );
  AOI21_X1 U11031 ( .B1(n9811), .B2(n9799), .A(n9798), .ZN(n9800) );
  NOR3_X1 U11032 ( .A1(n9801), .A2(n9800), .A3(n9817), .ZN(n9802) );
  AOI21_X1 U11033 ( .B1(n9804), .B2(n9803), .A(n9802), .ZN(n9938) );
  NOR2_X1 U11034 ( .A1(n9938), .A2(n9827), .ZN(n9805) );
  AOI211_X1 U11035 ( .C1(n9935), .C2(n9807), .A(n9806), .B(n9805), .ZN(n9808)
         );
  OAI21_X1 U11036 ( .B1(n9940), .B2(n9809), .A(n9808), .ZN(P1_U3279) );
  NOR2_X1 U11037 ( .A1(n9810), .A2(n5048), .ZN(n9814) );
  INV_X1 U11038 ( .A(n9811), .ZN(n9812) );
  AOI21_X1 U11039 ( .B1(n9814), .B2(n9813), .A(n9812), .ZN(n9818) );
  OAI22_X1 U11040 ( .A1(n9818), .A2(n9817), .B1(n9816), .B2(n9815), .ZN(n9945)
         );
  INV_X1 U11041 ( .A(n9945), .ZN(n9834) );
  OAI21_X1 U11042 ( .B1(n9821), .B2(n9820), .A(n9819), .ZN(n9947) );
  AOI21_X1 U11043 ( .B1(n9823), .B2(n9941), .A(n9822), .ZN(n9825) );
  NAND2_X1 U11044 ( .A1(n9825), .A2(n9824), .ZN(n9942) );
  AOI22_X1 U11045 ( .A1(n9827), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9826), .B2(
        n9836), .ZN(n9828) );
  OAI21_X1 U11046 ( .B1(n9944), .B2(n9829), .A(n9828), .ZN(n9830) );
  AOI21_X1 U11047 ( .B1(n9941), .B2(n9837), .A(n9830), .ZN(n9831) );
  OAI21_X1 U11048 ( .B1(n9942), .B2(n9840), .A(n9831), .ZN(n9832) );
  AOI21_X1 U11049 ( .B1(n9947), .B2(n9847), .A(n9832), .ZN(n9833) );
  OAI21_X1 U11050 ( .B1(n9834), .B2(n9827), .A(n9833), .ZN(P1_U3280) );
  AOI22_X1 U11051 ( .A1(n9838), .A2(n9837), .B1(n9836), .B2(n9835), .ZN(n9839)
         );
  OAI21_X1 U11052 ( .B1(n9841), .B2(n9840), .A(n9839), .ZN(n9845) );
  MUX2_X1 U11053 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n9843), .S(n9842), .Z(n9844)
         );
  AOI211_X1 U11054 ( .C1(n9847), .C2(n9846), .A(n9845), .B(n9844), .ZN(n9848)
         );
  INV_X1 U11055 ( .A(n9848), .ZN(P1_U3284) );
  INV_X1 U11056 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9851) );
  NOR2_X1 U11057 ( .A1(n9850), .A2(n9849), .ZN(n9970) );
  MUX2_X1 U11058 ( .A(n9851), .B(n9970), .S(n10164), .Z(n9852) );
  OAI21_X1 U11059 ( .B1(n9972), .B2(n9962), .A(n9852), .ZN(P1_U3553) );
  INV_X1 U11060 ( .A(n9857), .ZN(P1_U3552) );
  NAND2_X1 U11061 ( .A1(n9858), .A2(n9959), .ZN(n9863) );
  AOI22_X1 U11062 ( .A1(n9859), .A2(n10154), .B1(n9877), .B2(n4412), .ZN(n9861) );
  NAND4_X1 U11063 ( .A1(n9863), .A2(n9862), .A3(n9861), .A4(n9860), .ZN(n9977)
         );
  MUX2_X1 U11064 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9977), .S(n10164), .Z(
        P1_U3549) );
  MUX2_X1 U11065 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9978), .S(n10164), .Z(
        P1_U3548) );
  INV_X1 U11066 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9873) );
  OAI21_X1 U11067 ( .B1(n9869), .B2(n9943), .A(n9868), .ZN(n9870) );
  AOI211_X1 U11068 ( .C1(n9872), .C2(n9959), .A(n9871), .B(n9870), .ZN(n9979)
         );
  MUX2_X1 U11069 ( .A(n9873), .B(n9979), .S(n10164), .Z(n9874) );
  OAI21_X1 U11070 ( .B1(n9982), .B2(n9962), .A(n9874), .ZN(P1_U3547) );
  NAND2_X1 U11071 ( .A1(n9875), .A2(n9959), .ZN(n9881) );
  AOI22_X1 U11072 ( .A1(n6980), .A2(n10154), .B1(n9877), .B2(n9876), .ZN(n9879) );
  NAND4_X1 U11073 ( .A1(n9881), .A2(n9880), .A3(n9879), .A4(n9878), .ZN(n9983)
         );
  MUX2_X1 U11074 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9983), .S(n10164), .Z(
        P1_U3546) );
  INV_X1 U11075 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10544) );
  AOI211_X1 U11076 ( .C1(n9884), .C2(n9959), .A(n9883), .B(n9882), .ZN(n9984)
         );
  MUX2_X1 U11077 ( .A(n10544), .B(n9984), .S(n10164), .Z(n9885) );
  OAI21_X1 U11078 ( .B1(n5012), .B2(n9962), .A(n9885), .ZN(P1_U3545) );
  INV_X1 U11079 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9891) );
  OAI211_X1 U11080 ( .C1(n9888), .C2(n9943), .A(n9887), .B(n9886), .ZN(n9889)
         );
  AOI21_X1 U11081 ( .B1(n9890), .B2(n9959), .A(n9889), .ZN(n9987) );
  MUX2_X1 U11082 ( .A(n9891), .B(n9987), .S(n10164), .Z(n9892) );
  OAI21_X1 U11083 ( .B1(n9990), .B2(n9962), .A(n9892), .ZN(P1_U3544) );
  NOR2_X1 U11084 ( .A1(n9893), .A2(n9943), .ZN(n9895) );
  AOI211_X1 U11085 ( .C1(n10154), .C2(n9896), .A(n9895), .B(n9894), .ZN(n9897)
         );
  OAI211_X1 U11086 ( .C1(n9899), .C2(n10157), .A(n9898), .B(n9897), .ZN(n9991)
         );
  MUX2_X1 U11087 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9991), .S(n10164), .Z(
        P1_U3543) );
  NOR2_X1 U11088 ( .A1(n9900), .A2(n9943), .ZN(n9902) );
  AOI211_X1 U11089 ( .C1(n10154), .C2(n9903), .A(n9902), .B(n9901), .ZN(n9904)
         );
  OAI211_X1 U11090 ( .C1(n9906), .C2(n10157), .A(n9905), .B(n9904), .ZN(n9992)
         );
  MUX2_X1 U11091 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9992), .S(n10164), .Z(
        P1_U3542) );
  INV_X1 U11092 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9910) );
  AOI211_X1 U11093 ( .C1(n9909), .C2(n9959), .A(n9908), .B(n9907), .ZN(n9993)
         );
  MUX2_X1 U11094 ( .A(n9910), .B(n9993), .S(n10164), .Z(n9911) );
  OAI21_X1 U11095 ( .B1(n9996), .B2(n9962), .A(n9911), .ZN(P1_U3541) );
  AOI211_X1 U11096 ( .C1(n10154), .C2(n9914), .A(n9913), .B(n9912), .ZN(n9915)
         );
  OAI21_X1 U11097 ( .B1(n10157), .B2(n9916), .A(n9915), .ZN(n9997) );
  MUX2_X1 U11098 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9997), .S(n10164), .Z(
        P1_U3540) );
  OAI211_X1 U11099 ( .C1(n9919), .C2(n9943), .A(n9918), .B(n9917), .ZN(n9920)
         );
  AOI21_X1 U11100 ( .B1(n9921), .B2(n9959), .A(n9920), .ZN(n9998) );
  MUX2_X1 U11101 ( .A(n9922), .B(n9998), .S(n10164), .Z(n9923) );
  OAI21_X1 U11102 ( .B1(n10001), .B2(n9962), .A(n9923), .ZN(P1_U3539) );
  AOI21_X1 U11103 ( .B1(n10154), .B2(n9925), .A(n9924), .ZN(n9926) );
  OAI211_X1 U11104 ( .C1(n10157), .C2(n9928), .A(n9927), .B(n9926), .ZN(n10002) );
  MUX2_X1 U11105 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10002), .S(n10164), .Z(
        P1_U3538) );
  OAI211_X1 U11106 ( .C1(n10157), .C2(n9931), .A(n9930), .B(n9929), .ZN(n9932)
         );
  INV_X1 U11107 ( .A(n9932), .ZN(n10003) );
  MUX2_X1 U11108 ( .A(n10572), .B(n10003), .S(n10164), .Z(n9933) );
  OAI21_X1 U11109 ( .B1(n10006), .B2(n9962), .A(n9933), .ZN(P1_U3537) );
  NOR2_X1 U11110 ( .A1(n9934), .A2(n9943), .ZN(n9936) );
  AOI211_X1 U11111 ( .C1(n10154), .C2(n9937), .A(n9936), .B(n9935), .ZN(n9939)
         );
  OAI211_X1 U11112 ( .C1(n10157), .C2(n9940), .A(n9939), .B(n9938), .ZN(n10007) );
  MUX2_X1 U11113 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10007), .S(n10164), .Z(
        P1_U3536) );
  INV_X1 U11114 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10481) );
  OAI21_X1 U11115 ( .B1(n9944), .B2(n9943), .A(n9942), .ZN(n9946) );
  AOI211_X1 U11116 ( .C1(n9959), .C2(n9947), .A(n9946), .B(n9945), .ZN(n10008)
         );
  MUX2_X1 U11117 ( .A(n10481), .B(n10008), .S(n10164), .Z(n9948) );
  OAI21_X1 U11118 ( .B1(n6996), .B2(n9962), .A(n9948), .ZN(P1_U3535) );
  OAI21_X1 U11119 ( .B1(n9951), .B2(n9950), .A(n9949), .ZN(n9953) );
  AOI211_X1 U11120 ( .C1(n9959), .C2(n9954), .A(n9953), .B(n9952), .ZN(n10012)
         );
  NAND2_X1 U11121 ( .A1(n10162), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9955) );
  OAI21_X1 U11122 ( .B1(n10012), .B2(n10162), .A(n9955), .ZN(P1_U3534) );
  INV_X1 U11123 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9960) );
  AOI211_X1 U11124 ( .C1(n9959), .C2(n9958), .A(n9957), .B(n9956), .ZN(n10013)
         );
  MUX2_X1 U11125 ( .A(n9960), .B(n10013), .S(n10164), .Z(n9961) );
  OAI21_X1 U11126 ( .B1(n10017), .B2(n9962), .A(n9961), .ZN(P1_U3533) );
  INV_X1 U11127 ( .A(n9963), .ZN(n9969) );
  AOI21_X1 U11128 ( .B1(n10154), .B2(n9965), .A(n9964), .ZN(n9966) );
  OAI211_X1 U11129 ( .C1(n9969), .C2(n9968), .A(n9967), .B(n9966), .ZN(n10018)
         );
  MUX2_X1 U11130 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10018), .S(n10164), .Z(
        P1_U3530) );
  MUX2_X1 U11131 ( .A(n10410), .B(n9970), .S(n10161), .Z(n9971) );
  OAI21_X1 U11132 ( .B1(n9972), .B2(n10016), .A(n9971), .ZN(P1_U3521) );
  MUX2_X1 U11133 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9973), .S(n10161), .Z(
        n9974) );
  INV_X1 U11134 ( .A(n9974), .ZN(n9975) );
  OAI21_X1 U11135 ( .B1(n9976), .B2(n10016), .A(n9975), .ZN(P1_U3520) );
  MUX2_X1 U11136 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9977), .S(n10161), .Z(
        P1_U3517) );
  MUX2_X1 U11137 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9978), .S(n10161), .Z(
        P1_U3516) );
  INV_X1 U11138 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9980) );
  MUX2_X1 U11139 ( .A(n9980), .B(n9979), .S(n10161), .Z(n9981) );
  OAI21_X1 U11140 ( .B1(n9982), .B2(n10016), .A(n9981), .ZN(P1_U3515) );
  MUX2_X1 U11141 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9983), .S(n10161), .Z(
        P1_U3514) );
  INV_X1 U11142 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9985) );
  MUX2_X1 U11143 ( .A(n9985), .B(n9984), .S(n10161), .Z(n9986) );
  OAI21_X1 U11144 ( .B1(n5012), .B2(n10016), .A(n9986), .ZN(P1_U3513) );
  INV_X1 U11145 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9988) );
  MUX2_X1 U11146 ( .A(n9988), .B(n9987), .S(n10161), .Z(n9989) );
  OAI21_X1 U11147 ( .B1(n9990), .B2(n10016), .A(n9989), .ZN(P1_U3512) );
  MUX2_X1 U11148 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9991), .S(n10161), .Z(
        P1_U3511) );
  MUX2_X1 U11149 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9992), .S(n10161), .Z(
        P1_U3510) );
  INV_X1 U11150 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9994) );
  MUX2_X1 U11151 ( .A(n9994), .B(n9993), .S(n10161), .Z(n9995) );
  OAI21_X1 U11152 ( .B1(n9996), .B2(n10016), .A(n9995), .ZN(P1_U3509) );
  MUX2_X1 U11153 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9997), .S(n10161), .Z(
        P1_U3507) );
  INV_X1 U11154 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9999) );
  MUX2_X1 U11155 ( .A(n9999), .B(n9998), .S(n10161), .Z(n10000) );
  OAI21_X1 U11156 ( .B1(n10001), .B2(n10016), .A(n10000), .ZN(P1_U3504) );
  MUX2_X1 U11157 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10002), .S(n10161), .Z(
        P1_U3501) );
  INV_X1 U11158 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10004) );
  MUX2_X1 U11159 ( .A(n10004), .B(n10003), .S(n10161), .Z(n10005) );
  OAI21_X1 U11160 ( .B1(n10006), .B2(n10016), .A(n10005), .ZN(P1_U3498) );
  MUX2_X1 U11161 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10007), .S(n10161), .Z(
        P1_U3495) );
  MUX2_X1 U11162 ( .A(n10009), .B(n10008), .S(n10161), .Z(n10010) );
  OAI21_X1 U11163 ( .B1(n6996), .B2(n10016), .A(n10010), .ZN(P1_U3492) );
  NAND2_X1 U11164 ( .A1(n10160), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10011) );
  OAI21_X1 U11165 ( .B1(n10012), .B2(n10160), .A(n10011), .ZN(P1_U3489) );
  MUX2_X1 U11166 ( .A(n10014), .B(n10013), .S(n10161), .Z(n10015) );
  OAI21_X1 U11167 ( .B1(n10017), .B2(n10016), .A(n10015), .ZN(P1_U3486) );
  MUX2_X1 U11168 ( .A(P1_REG0_REG_8__SCAN_IN), .B(n10018), .S(n10161), .Z(
        P1_U3477) );
  MUX2_X1 U11169 ( .A(n10019), .B(P1_D_REG_1__SCAN_IN), .S(n10150), .Z(
        P1_U3440) );
  MUX2_X1 U11170 ( .A(n10020), .B(P1_D_REG_0__SCAN_IN), .S(n10150), .Z(
        P1_U3439) );
  NOR4_X1 U11171 ( .A1(n10022), .A2(P1_IR_REG_30__SCAN_IN), .A3(n10021), .A4(
        n4401), .ZN(n10023) );
  AOI21_X1 U11172 ( .B1(n10024), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10023), 
        .ZN(n10025) );
  OAI21_X1 U11173 ( .B1(n10027), .B2(n10026), .A(n10025), .ZN(P1_U3324) );
  OAI222_X1 U11174 ( .A1(n5409), .A2(n4401), .B1(n10040), .B2(n10028), .C1(
        n10581), .C2(n10037), .ZN(P1_U3326) );
  OAI222_X1 U11175 ( .A1(n10037), .A2(n10030), .B1(n10040), .B2(n10029), .C1(
        n4413), .C2(P1_U3086), .ZN(P1_U3328) );
  OAI222_X1 U11176 ( .A1(n4401), .A2(n10033), .B1(n10040), .B2(n10032), .C1(
        n10031), .C2(n10037), .ZN(P1_U3329) );
  OAI222_X1 U11177 ( .A1(P1_U3086), .A2(n10036), .B1(n10040), .B2(n10035), 
        .C1(n10034), .C2(n10037), .ZN(P1_U3330) );
  OAI222_X1 U11178 ( .A1(n4401), .A2(n10041), .B1(n10040), .B2(n10039), .C1(
        n10038), .C2(n10037), .ZN(P1_U3331) );
  MUX2_X1 U11179 ( .A(n10042), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  NOR2_X1 U11180 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10077) );
  NOR2_X1 U11181 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10074) );
  NOR2_X1 U11182 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10071) );
  NOR2_X1 U11183 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10069) );
  NOR2_X1 U11184 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10067) );
  NOR2_X1 U11185 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10065) );
  NOR2_X1 U11186 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10063) );
  NOR2_X1 U11187 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10061) );
  NOR2_X1 U11188 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10059) );
  NOR2_X1 U11189 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10057) );
  NOR2_X1 U11190 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10055) );
  NOR2_X1 U11191 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10053) );
  NOR2_X1 U11192 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10051) );
  NOR2_X1 U11193 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10049) );
  NAND2_X1 U11194 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10047) );
  XOR2_X1 U11195 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10616) );
  NAND2_X1 U11196 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10045) );
  AOI21_X1 U11197 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10261) );
  INV_X1 U11198 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10374) );
  INV_X1 U11199 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10264) );
  NOR2_X1 U11200 ( .A1(n10374), .A2(n10264), .ZN(n10263) );
  AND2_X1 U11201 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n10263), .ZN(n10260) );
  NOR2_X1 U11202 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10260), .ZN(n10043) );
  NOR2_X1 U11203 ( .A1(n10261), .A2(n10043), .ZN(n10614) );
  XOR2_X1 U11204 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10613) );
  NAND2_X1 U11205 ( .A1(n10614), .A2(n10613), .ZN(n10044) );
  NAND2_X1 U11206 ( .A1(n10045), .A2(n10044), .ZN(n10615) );
  NAND2_X1 U11207 ( .A1(n10616), .A2(n10615), .ZN(n10046) );
  NAND2_X1 U11208 ( .A1(n10047), .A2(n10046), .ZN(n10618) );
  XNOR2_X1 U11209 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10617) );
  NOR2_X1 U11210 ( .A1(n10618), .A2(n10617), .ZN(n10048) );
  NOR2_X1 U11211 ( .A1(n10049), .A2(n10048), .ZN(n10606) );
  XNOR2_X1 U11212 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10605) );
  NOR2_X1 U11213 ( .A1(n10606), .A2(n10605), .ZN(n10050) );
  NOR2_X1 U11214 ( .A1(n10051), .A2(n10050), .ZN(n10604) );
  XNOR2_X1 U11215 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10603) );
  NOR2_X1 U11216 ( .A1(n10604), .A2(n10603), .ZN(n10052) );
  NOR2_X1 U11217 ( .A1(n10053), .A2(n10052), .ZN(n10610) );
  XNOR2_X1 U11218 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10609) );
  NOR2_X1 U11219 ( .A1(n10610), .A2(n10609), .ZN(n10054) );
  NOR2_X1 U11220 ( .A1(n10055), .A2(n10054), .ZN(n10612) );
  XNOR2_X1 U11221 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10611) );
  NOR2_X1 U11222 ( .A1(n10612), .A2(n10611), .ZN(n10056) );
  NOR2_X1 U11223 ( .A1(n10057), .A2(n10056), .ZN(n10608) );
  XNOR2_X1 U11224 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10607) );
  NOR2_X1 U11225 ( .A1(n10608), .A2(n10607), .ZN(n10058) );
  XNOR2_X1 U11226 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10282) );
  NOR2_X1 U11227 ( .A1(n10283), .A2(n10282), .ZN(n10060) );
  XNOR2_X1 U11228 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10280) );
  NOR2_X1 U11229 ( .A1(n10281), .A2(n10280), .ZN(n10062) );
  XNOR2_X1 U11230 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10278) );
  NOR2_X1 U11231 ( .A1(n10279), .A2(n10278), .ZN(n10064) );
  XNOR2_X1 U11232 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10276) );
  NOR2_X1 U11233 ( .A1(n10277), .A2(n10276), .ZN(n10066) );
  XNOR2_X1 U11234 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10274) );
  NOR2_X1 U11235 ( .A1(n10275), .A2(n10274), .ZN(n10068) );
  XNOR2_X1 U11236 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10272) );
  NOR2_X1 U11237 ( .A1(n10273), .A2(n10272), .ZN(n10070) );
  NOR2_X1 U11238 ( .A1(n10071), .A2(n10070), .ZN(n10271) );
  INV_X1 U11239 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n10072) );
  AOI22_X1 U11240 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n10567), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n10072), .ZN(n10270) );
  NOR2_X1 U11241 ( .A1(n10271), .A2(n10270), .ZN(n10073) );
  NOR2_X1 U11242 ( .A1(n10074), .A2(n10073), .ZN(n10269) );
  INV_X1 U11243 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10135) );
  INV_X1 U11244 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n10075) );
  AOI22_X1 U11245 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n10135), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n10075), .ZN(n10268) );
  NOR2_X1 U11246 ( .A1(n10269), .A2(n10268), .ZN(n10076) );
  NOR2_X1 U11247 ( .A1(n10077), .A2(n10076), .ZN(n10078) );
  NOR2_X1 U11248 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10078), .ZN(n10266) );
  AND2_X1 U11249 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10078), .ZN(n10265) );
  NOR2_X1 U11250 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10265), .ZN(n10079) );
  NOR2_X1 U11251 ( .A1(n10266), .A2(n10079), .ZN(n10081) );
  XNOR2_X1 U11252 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n10080) );
  XNOR2_X1 U11253 ( .A(n10081), .B(n10080), .ZN(ADD_1068_U4) );
  XNOR2_X1 U11254 ( .A(P1_WR_REG_SCAN_IN), .B(P2_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11255 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11256 ( .A(n10082), .ZN(n10084) );
  NAND2_X1 U11257 ( .A1(n4413), .A2(n10083), .ZN(n10085) );
  NAND2_X1 U11258 ( .A1(n10084), .A2(n10085), .ZN(n10086) );
  MUX2_X1 U11259 ( .A(n10086), .B(n10085), .S(n4764), .Z(n10088) );
  NAND2_X1 U11260 ( .A1(n10088), .A2(n10087), .ZN(n10091) );
  AOI22_X1 U11261 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n10089), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n4401), .ZN(n10090) );
  OAI21_X1 U11262 ( .B1(n10092), .B2(n10091), .A(n10090), .ZN(P1_U3243) );
  INV_X1 U11263 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10107) );
  AOI211_X1 U11264 ( .C1(n10095), .C2(n10094), .A(n10093), .B(n10137), .ZN(
        n10103) );
  AOI211_X1 U11265 ( .C1(n10098), .C2(n10097), .A(n10096), .B(n10141), .ZN(
        n10102) );
  NOR2_X1 U11266 ( .A1(n10100), .A2(n10099), .ZN(n10101) );
  NOR4_X1 U11267 ( .A1(n10104), .A2(n10103), .A3(n10102), .A4(n10101), .ZN(
        n10106) );
  OAI211_X1 U11268 ( .C1(n10107), .C2(n10148), .A(n10106), .B(n10105), .ZN(
        P1_U3247) );
  AOI211_X1 U11269 ( .C1(n10110), .C2(n10109), .A(n10108), .B(n10141), .ZN(
        n10111) );
  AOI21_X1 U11270 ( .B1(n10146), .B2(n10112), .A(n10111), .ZN(n10117) );
  OAI21_X1 U11271 ( .B1(n10114), .B2(n4522), .A(n10113), .ZN(n10115) );
  NAND2_X1 U11272 ( .A1(n10115), .A2(n10131), .ZN(n10116) );
  AND2_X1 U11273 ( .A1(n10117), .A2(n10116), .ZN(n10119) );
  OAI211_X1 U11274 ( .C1(n10148), .C2(n10567), .A(n10119), .B(n10118), .ZN(
        P1_U3259) );
  OAI21_X1 U11275 ( .B1(n10122), .B2(n10121), .A(n10120), .ZN(n10132) );
  OAI21_X1 U11276 ( .B1(n10125), .B2(n10124), .A(n10123), .ZN(n10126) );
  AOI22_X1 U11277 ( .A1(n10128), .A2(n10146), .B1(n10127), .B2(n10126), .ZN(
        n10129) );
  INV_X1 U11278 ( .A(n10129), .ZN(n10130) );
  AOI21_X1 U11279 ( .B1(n10132), .B2(n10131), .A(n10130), .ZN(n10134) );
  OAI211_X1 U11280 ( .C1(n10148), .C2(n10135), .A(n10134), .B(n10133), .ZN(
        P1_U3260) );
  INV_X1 U11281 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10542) );
  INV_X1 U11282 ( .A(n10136), .ZN(n10138) );
  AOI211_X1 U11283 ( .C1(n10140), .C2(n10139), .A(n10138), .B(n10137), .ZN(
        n10144) );
  AND2_X1 U11284 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10150), .ZN(P1_U3294) );
  INV_X1 U11285 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10407) );
  NOR2_X1 U11286 ( .A1(n10149), .A2(n10407), .ZN(P1_U3295) );
  INV_X1 U11287 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10383) );
  NOR2_X1 U11288 ( .A1(n10149), .A2(n10383), .ZN(P1_U3296) );
  AND2_X1 U11289 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10150), .ZN(P1_U3297) );
  AND2_X1 U11290 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10150), .ZN(P1_U3298) );
  AND2_X1 U11291 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10150), .ZN(P1_U3299) );
  AND2_X1 U11292 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10150), .ZN(P1_U3300) );
  AND2_X1 U11293 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10150), .ZN(P1_U3301) );
  AND2_X1 U11294 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10150), .ZN(P1_U3302) );
  INV_X1 U11295 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10559) );
  NOR2_X1 U11296 ( .A1(n10149), .A2(n10559), .ZN(P1_U3303) );
  INV_X1 U11297 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10464) );
  NOR2_X1 U11298 ( .A1(n10149), .A2(n10464), .ZN(P1_U3304) );
  AND2_X1 U11299 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10150), .ZN(P1_U3305) );
  AND2_X1 U11300 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10150), .ZN(P1_U3306) );
  AND2_X1 U11301 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10150), .ZN(P1_U3307) );
  INV_X1 U11302 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10485) );
  NOR2_X1 U11303 ( .A1(n10149), .A2(n10485), .ZN(P1_U3308) );
  AND2_X1 U11304 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10150), .ZN(P1_U3309) );
  INV_X1 U11305 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10430) );
  NOR2_X1 U11306 ( .A1(n10149), .A2(n10430), .ZN(P1_U3310) );
  AND2_X1 U11307 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10150), .ZN(P1_U3311) );
  AND2_X1 U11308 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10150), .ZN(P1_U3312) );
  AND2_X1 U11309 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10150), .ZN(P1_U3313) );
  AND2_X1 U11310 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10150), .ZN(P1_U3314) );
  AND2_X1 U11311 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10150), .ZN(P1_U3315) );
  AND2_X1 U11312 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10150), .ZN(P1_U3316) );
  AND2_X1 U11313 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10150), .ZN(P1_U3317) );
  AND2_X1 U11314 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10150), .ZN(P1_U3318) );
  AND2_X1 U11315 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10150), .ZN(P1_U3319) );
  AND2_X1 U11316 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10150), .ZN(P1_U3320) );
  AND2_X1 U11317 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10150), .ZN(P1_U3321) );
  AND2_X1 U11318 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10150), .ZN(P1_U3322) );
  AND2_X1 U11319 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10150), .ZN(P1_U3323) );
  INV_X1 U11320 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U11321 ( .A1(n10161), .A2(n10151), .B1(n10386), .B2(n10160), .ZN(
        P1_U3459) );
  AOI21_X1 U11322 ( .B1(n10154), .B2(n10153), .A(n10152), .ZN(n10155) );
  OAI211_X1 U11323 ( .C1(n10158), .C2(n10157), .A(n10156), .B(n10155), .ZN(
        n10159) );
  INV_X1 U11324 ( .A(n10159), .ZN(n10163) );
  AOI22_X1 U11325 ( .A1(n10161), .A2(n10163), .B1(n5539), .B2(n10160), .ZN(
        P1_U3465) );
  AOI22_X1 U11326 ( .A1(n10164), .A2(n10163), .B1(n7368), .B2(n10162), .ZN(
        P1_U3526) );
  XNOR2_X1 U11327 ( .A(n10165), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n10166) );
  AOI22_X1 U11328 ( .A1(n5231), .A2(n10166), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        P2_U3151), .ZN(n10181) );
  AOI21_X1 U11329 ( .B1(n10169), .B2(n10168), .A(n10167), .ZN(n10175) );
  NAND2_X1 U11330 ( .A1(n10170), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n10174) );
  OAI211_X1 U11331 ( .C1(n10289), .C2(n10172), .A(n10288), .B(n10171), .ZN(
        n10173) );
  OAI211_X1 U11332 ( .C1(n10176), .C2(n10175), .A(n10174), .B(n10173), .ZN(
        n10177) );
  AOI21_X1 U11333 ( .B1(n10179), .B2(n10178), .A(n10177), .ZN(n10180) );
  NAND2_X1 U11334 ( .A1(n10181), .A2(n10180), .ZN(P2_U3183) );
  INV_X1 U11335 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10203) );
  XOR2_X1 U11336 ( .A(n10183), .B(n10182), .Z(n10201) );
  NOR2_X1 U11337 ( .A1(n10298), .A2(n10184), .ZN(n10200) );
  AOI21_X1 U11338 ( .B1(n10187), .B2(n10186), .A(n10185), .ZN(n10198) );
  AND3_X1 U11339 ( .A1(n10190), .A2(n10189), .A3(n10188), .ZN(n10192) );
  OAI21_X1 U11340 ( .B1(n10193), .B2(n10192), .A(n10191), .ZN(n10196) );
  INV_X1 U11341 ( .A(n10194), .ZN(n10195) );
  OAI211_X1 U11342 ( .C1(n10198), .C2(n10197), .A(n10196), .B(n10195), .ZN(
        n10199) );
  AOI211_X1 U11343 ( .C1(n10201), .C2(n10288), .A(n10200), .B(n10199), .ZN(
        n10202) );
  OAI21_X1 U11344 ( .B1(n10294), .B2(n10203), .A(n10202), .ZN(P2_U3186) );
  OAI21_X1 U11345 ( .B1(n10205), .B2(n10210), .A(n10204), .ZN(n10227) );
  OAI22_X1 U11346 ( .A1(n10208), .A2(n10207), .B1(n10224), .B2(n10206), .ZN(
        n10219) );
  XNOR2_X1 U11347 ( .A(n10209), .B(n10210), .ZN(n10217) );
  OAI22_X1 U11348 ( .A1(n10213), .A2(n10212), .B1(n6633), .B2(n10211), .ZN(
        n10214) );
  AOI21_X1 U11349 ( .B1(n10227), .B2(n10215), .A(n10214), .ZN(n10216) );
  OAI21_X1 U11350 ( .B1(n10218), .B2(n10217), .A(n10216), .ZN(n10225) );
  AOI211_X1 U11351 ( .C1(n10220), .C2(n10227), .A(n10219), .B(n10225), .ZN(
        n10222) );
  AOI22_X1 U11352 ( .A1(n10223), .A2(n10441), .B1(n10222), .B2(n10221), .ZN(
        P2_U3231) );
  NOR2_X1 U11353 ( .A1(n10224), .A2(n10242), .ZN(n10226) );
  AOI211_X1 U11354 ( .C1(n10228), .C2(n10227), .A(n10226), .B(n10225), .ZN(
        n10251) );
  AOI22_X1 U11355 ( .A1(n10249), .A2(n6195), .B1(n10251), .B2(n10247), .ZN(
        P2_U3396) );
  INV_X1 U11356 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10234) );
  INV_X1 U11357 ( .A(n10229), .ZN(n10233) );
  OAI21_X1 U11358 ( .B1(n10231), .B2(n10242), .A(n10230), .ZN(n10232) );
  AOI21_X1 U11359 ( .B1(n10233), .B2(n10245), .A(n10232), .ZN(n10253) );
  AOI22_X1 U11360 ( .A1(n10249), .A2(n10234), .B1(n10253), .B2(n10247), .ZN(
        P2_U3399) );
  INV_X1 U11361 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10239) );
  NOR2_X1 U11362 ( .A1(n10235), .A2(n10242), .ZN(n10237) );
  AOI211_X1 U11363 ( .C1(n10238), .C2(n10245), .A(n10237), .B(n10236), .ZN(
        n10256) );
  AOI22_X1 U11364 ( .A1(n10249), .A2(n10239), .B1(n10256), .B2(n10247), .ZN(
        P2_U3402) );
  INV_X1 U11365 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10248) );
  INV_X1 U11366 ( .A(n10240), .ZN(n10246) );
  OAI21_X1 U11367 ( .B1(n10243), .B2(n10242), .A(n10241), .ZN(n10244) );
  AOI21_X1 U11368 ( .B1(n10246), .B2(n10245), .A(n10244), .ZN(n10258) );
  AOI22_X1 U11369 ( .A1(n10249), .A2(n10248), .B1(n10258), .B2(n10247), .ZN(
        P2_U3405) );
  AOI22_X1 U11370 ( .A1(n10254), .A2(n10251), .B1(n10250), .B2(n10257), .ZN(
        P2_U3461) );
  INV_X1 U11371 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10252) );
  AOI22_X1 U11372 ( .A1(n10254), .A2(n10253), .B1(n10252), .B2(n10257), .ZN(
        P2_U3462) );
  AOI22_X1 U11373 ( .A1(n10259), .A2(n10256), .B1(n10255), .B2(n10257), .ZN(
        P2_U3463) );
  AOI22_X1 U11374 ( .A1(n10259), .A2(n10258), .B1(n6827), .B2(n10257), .ZN(
        P2_U3464) );
  NOR2_X1 U11375 ( .A1(n10261), .A2(n10260), .ZN(n10262) );
  XOR2_X1 U11376 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10262), .Z(ADD_1068_U5) );
  AOI21_X1 U11377 ( .B1(n10374), .B2(n10264), .A(n10263), .ZN(ADD_1068_U46) );
  NOR2_X1 U11378 ( .A1(n10266), .A2(n10265), .ZN(n10267) );
  XOR2_X1 U11379 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n10267), .Z(ADD_1068_U55)
         );
  XNOR2_X1 U11380 ( .A(n10269), .B(n10268), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11381 ( .A(n10271), .B(n10270), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11382 ( .A(n10273), .B(n10272), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11383 ( .A(n10275), .B(n10274), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11384 ( .A(n10277), .B(n10276), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11385 ( .A(n10279), .B(n10278), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11386 ( .A(n10281), .B(n10280), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11387 ( .A(n10283), .B(n10282), .ZN(ADD_1068_U63) );
  INV_X1 U11388 ( .A(n10284), .ZN(n10285) );
  AND2_X1 U11389 ( .A1(n10286), .A2(n10285), .ZN(n10287) );
  OR2_X1 U11390 ( .A1(n10288), .A2(n10287), .ZN(n10293) );
  NOR2_X1 U11391 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7531), .ZN(n10291) );
  AOI21_X1 U11392 ( .B1(n10293), .B2(n10292), .A(n10291), .ZN(n10296) );
  OR2_X1 U11393 ( .A1(n10294), .A2(n10264), .ZN(n10295) );
  OAI211_X1 U11394 ( .C1(n10298), .C2(n10297), .A(n10296), .B(n10295), .ZN(
        n10299) );
  INV_X1 U11395 ( .A(n10299), .ZN(n10602) );
  NOR4_X1 U11396 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(P1_REG1_REG_26__SCAN_IN), 
        .A3(P1_REG0_REG_2__SCAN_IN), .A4(P1_ADDR_REG_10__SCAN_IN), .ZN(n10301)
         );
  NAND3_X1 U11397 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(n10301), .A3(n10300), .ZN(
        n10315) );
  NAND4_X1 U11398 ( .A1(n10303), .A2(n10302), .A3(SI_21_), .A4(
        P2_IR_REG_30__SCAN_IN), .ZN(n10304) );
  NOR3_X1 U11399 ( .A1(n10304), .A2(P1_REG0_REG_9__SCAN_IN), .A3(n10407), .ZN(
        n10313) );
  NAND4_X1 U11400 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(n10529), .A3(n10520), 
        .A4(n10526), .ZN(n10305) );
  NOR3_X1 U11401 ( .A1(n10306), .A2(P2_DATAO_REG_10__SCAN_IN), .A3(n10305), 
        .ZN(n10307) );
  INV_X1 U11402 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10510) );
  NAND3_X1 U11403 ( .A1(n10307), .A2(P1_REG0_REG_8__SCAN_IN), .A3(n10510), 
        .ZN(n10311) );
  NAND4_X1 U11404 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), 
        .A3(n10508), .A4(n10308), .ZN(n10310) );
  NAND4_X1 U11405 ( .A1(n10362), .A2(SI_23_), .A3(SI_2_), .A4(
        P2_REG0_REG_23__SCAN_IN), .ZN(n10309) );
  NOR3_X1 U11406 ( .A1(n10311), .A2(n10310), .A3(n10309), .ZN(n10312) );
  NAND4_X1 U11407 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(n10313), .A3(n10312), 
        .A4(n10394), .ZN(n10314) );
  NOR4_X1 U11408 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(SI_14_), .A3(n10315), 
        .A4(n10314), .ZN(n10361) );
  NAND4_X1 U11409 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), 
        .A3(P1_IR_REG_30__SCAN_IN), .A4(n10544), .ZN(n10325) );
  NAND4_X1 U11410 ( .A1(SI_1_), .A2(n10558), .A3(n5552), .A4(n10542), .ZN(
        n10324) );
  INV_X1 U11411 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10554) );
  NOR4_X1 U11412 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), 
        .A3(P1_WR_REG_SCAN_IN), .A4(n10554), .ZN(n10322) );
  NOR4_X1 U11413 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .A3(P1_ADDR_REG_3__SCAN_IN), .A4(n10452), .ZN(n10321) );
  INV_X1 U11414 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10545) );
  INV_X1 U11415 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10423) );
  NOR3_X1 U11416 ( .A1(n10545), .A2(n6395), .A3(n10423), .ZN(n10316) );
  NAND3_X1 U11417 ( .A1(n10317), .A2(P2_IR_REG_18__SCAN_IN), .A3(n10316), .ZN(
        n10319) );
  INV_X1 U11418 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n10318) );
  NOR4_X1 U11419 ( .A1(n10374), .A2(n10319), .A3(P2_IR_REG_7__SCAN_IN), .A4(
        n10318), .ZN(n10320) );
  NAND3_X1 U11420 ( .A1(n10322), .A2(n10321), .A3(n10320), .ZN(n10323) );
  NOR3_X1 U11421 ( .A1(n10325), .A2(n10324), .A3(n10323), .ZN(n10326) );
  NAND4_X1 U11422 ( .A1(n10328), .A2(P1_DATAO_REG_8__SCAN_IN), .A3(n10327), 
        .A4(n10326), .ZN(n10359) );
  INV_X1 U11423 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10484) );
  NOR4_X1 U11424 ( .A1(n6179), .A2(n10496), .A3(n5414), .A4(n10484), .ZN(
        n10335) );
  NAND4_X1 U11425 ( .A1(n10330), .A2(n10329), .A3(P1_DATAO_REG_18__SCAN_IN), 
        .A4(P2_REG3_REG_25__SCAN_IN), .ZN(n10333) );
  NOR4_X1 U11426 ( .A1(P2_REG1_REG_5__SCAN_IN), .A2(P1_REG1_REG_13__SCAN_IN), 
        .A3(n10482), .A4(n10523), .ZN(n10331) );
  NAND3_X1 U11427 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P1_REG1_REG_2__SCAN_IN), 
        .A3(n10331), .ZN(n10332) );
  NOR4_X1 U11428 ( .A1(n10333), .A2(n10332), .A3(n10498), .A4(
        P1_REG2_REG_10__SCAN_IN), .ZN(n10334) );
  NAND2_X1 U11429 ( .A1(n10335), .A2(n10334), .ZN(n10358) );
  NOR4_X1 U11430 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG1_REG_30__SCAN_IN), 
        .A3(n10572), .A4(n10567), .ZN(n10344) );
  NOR4_X1 U11431 ( .A1(n10581), .A2(n10539), .A3(n8831), .A4(n5136), .ZN(
        n10343) );
  NOR4_X1 U11432 ( .A1(P2_REG0_REG_17__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), 
        .A3(P2_ADDR_REG_18__SCAN_IN), .A4(n10336), .ZN(n10337) );
  NAND3_X1 U11433 ( .A1(n10339), .A2(n10338), .A3(n10337), .ZN(n10341) );
  NOR3_X1 U11434 ( .A1(n10341), .A2(P2_REG3_REG_13__SCAN_IN), .A3(n10340), 
        .ZN(n10342) );
  NAND3_X1 U11435 ( .A1(n10344), .A2(n10343), .A3(n10342), .ZN(n10357) );
  NAND4_X1 U11436 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_17__SCAN_IN), 
        .A3(P1_REG0_REG_18__SCAN_IN), .A4(n7736), .ZN(n10345) );
  NOR3_X1 U11437 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_REG2_REG_30__SCAN_IN), 
        .A3(n10345), .ZN(n10355) );
  NOR4_X1 U11438 ( .A1(n4952), .A2(n10346), .A3(P2_REG2_REG_13__SCAN_IN), .A4(
        SI_13_), .ZN(n10347) );
  NAND3_X1 U11439 ( .A1(n10347), .A2(P1_REG3_REG_3__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .ZN(n10353) );
  NOR4_X1 U11440 ( .A1(SI_17_), .A2(P2_DATAO_REG_6__SCAN_IN), .A3(
        P2_REG1_REG_8__SCAN_IN), .A4(P1_REG2_REG_23__SCAN_IN), .ZN(n10351) );
  NOR4_X1 U11441 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .A3(n5458), .A4(n10410), .ZN(n10350) );
  INV_X1 U11442 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n10456) );
  NOR4_X1 U11443 ( .A1(SI_12_), .A2(P2_REG1_REG_12__SCAN_IN), .A3(
        P2_REG2_REG_4__SCAN_IN), .A4(n10456), .ZN(n10349) );
  NOR4_X1 U11444 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(P2_REG1_REG_9__SCAN_IN), 
        .A3(P2_REG2_REG_2__SCAN_IN), .A4(P1_REG1_REG_27__SCAN_IN), .ZN(n10348)
         );
  NAND4_X1 U11445 ( .A1(n10351), .A2(n10350), .A3(n10349), .A4(n10348), .ZN(
        n10352) );
  NOR4_X1 U11446 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P1_DATAO_REG_16__SCAN_IN), 
        .A3(n10353), .A4(n10352), .ZN(n10354) );
  NAND4_X1 U11447 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_DATAO_REG_15__SCAN_IN), 
        .A3(n10355), .A4(n10354), .ZN(n10356) );
  NOR4_X1 U11448 ( .A1(n10359), .A2(n10358), .A3(n10357), .A4(n10356), .ZN(
        n10360) );
  AOI21_X1 U11449 ( .B1(n10361), .B2(n10360), .A(P2_IR_REG_11__SCAN_IN), .ZN(
        n10600) );
  XNOR2_X1 U11450 ( .A(n10362), .B(keyinput10), .ZN(n10367) );
  XNOR2_X1 U11451 ( .A(n10363), .B(keyinput45), .ZN(n10366) );
  XNOR2_X1 U11452 ( .A(n10364), .B(keyinput0), .ZN(n10365) );
  NOR3_X1 U11453 ( .A1(n10367), .A2(n10366), .A3(n10365), .ZN(n10370) );
  XNOR2_X1 U11454 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput47), .ZN(n10369)
         );
  XNOR2_X1 U11455 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput126), .ZN(n10368)
         );
  NAND3_X1 U11456 ( .A1(n10370), .A2(n10369), .A3(n10368), .ZN(n10377) );
  AOI22_X1 U11457 ( .A1(n10373), .A2(keyinput103), .B1(n10372), .B2(
        keyinput104), .ZN(n10371) );
  OAI221_X1 U11458 ( .B1(n10373), .B2(keyinput103), .C1(n10372), .C2(
        keyinput104), .A(n10371), .ZN(n10376) );
  XNOR2_X1 U11459 ( .A(n10374), .B(keyinput115), .ZN(n10375) );
  NOR3_X1 U11460 ( .A1(n10377), .A2(n10376), .A3(n10375), .ZN(n10421) );
  INV_X1 U11461 ( .A(SI_14_), .ZN(n10380) );
  INV_X1 U11462 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n10379) );
  AOI22_X1 U11463 ( .A1(n10380), .A2(keyinput111), .B1(n10379), .B2(keyinput72), .ZN(n10378) );
  OAI221_X1 U11464 ( .B1(n10380), .B2(keyinput111), .C1(n10379), .C2(
        keyinput72), .A(n10378), .ZN(n10392) );
  AOI22_X1 U11465 ( .A1(n10383), .A2(keyinput73), .B1(keyinput51), .B2(n10382), 
        .ZN(n10381) );
  OAI221_X1 U11466 ( .B1(n10383), .B2(keyinput73), .C1(n10382), .C2(keyinput51), .A(n10381), .ZN(n10391) );
  INV_X1 U11467 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n10385) );
  AOI22_X1 U11468 ( .A1(n10386), .A2(keyinput96), .B1(n10385), .B2(keyinput18), 
        .ZN(n10384) );
  OAI221_X1 U11469 ( .B1(n10386), .B2(keyinput96), .C1(n10385), .C2(keyinput18), .A(n10384), .ZN(n10390) );
  XNOR2_X1 U11470 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput16), .ZN(n10388) );
  XNOR2_X1 U11471 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput106), .ZN(n10387)
         );
  NAND2_X1 U11472 ( .A1(n10388), .A2(n10387), .ZN(n10389) );
  NOR4_X1 U11473 ( .A1(n10392), .A2(n10391), .A3(n10390), .A4(n10389), .ZN(
        n10420) );
  AOI22_X1 U11474 ( .A1(n10395), .A2(keyinput113), .B1(n10394), .B2(keyinput75), .ZN(n10393) );
  OAI221_X1 U11475 ( .B1(n10395), .B2(keyinput113), .C1(n10394), .C2(
        keyinput75), .A(n10393), .ZN(n10405) );
  AOI22_X1 U11476 ( .A1(n10303), .A2(keyinput116), .B1(keyinput17), .B2(n10397), .ZN(n10396) );
  OAI221_X1 U11477 ( .B1(n10303), .B2(keyinput116), .C1(n10397), .C2(
        keyinput17), .A(n10396), .ZN(n10404) );
  AOI22_X1 U11478 ( .A1(n4958), .A2(keyinput35), .B1(keyinput69), .B2(n10399), 
        .ZN(n10398) );
  OAI221_X1 U11479 ( .B1(n4958), .B2(keyinput35), .C1(n10399), .C2(keyinput69), 
        .A(n10398), .ZN(n10403) );
  XOR2_X1 U11480 ( .A(n8971), .B(keyinput92), .Z(n10401) );
  XNOR2_X1 U11481 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput109), .ZN(n10400) );
  NAND2_X1 U11482 ( .A1(n10401), .A2(n10400), .ZN(n10402) );
  NOR4_X1 U11483 ( .A1(n10405), .A2(n10404), .A3(n10403), .A4(n10402), .ZN(
        n10419) );
  AOI22_X1 U11484 ( .A1(n10407), .A2(keyinput114), .B1(n5458), .B2(keyinput3), 
        .ZN(n10406) );
  OAI221_X1 U11485 ( .B1(n10407), .B2(keyinput114), .C1(n5458), .C2(keyinput3), 
        .A(n10406), .ZN(n10417) );
  AOI22_X1 U11486 ( .A1(n10410), .A2(keyinput2), .B1(n10409), .B2(keyinput102), 
        .ZN(n10408) );
  OAI221_X1 U11487 ( .B1(n10410), .B2(keyinput2), .C1(n10409), .C2(keyinput102), .A(n10408), .ZN(n10416) );
  XOR2_X1 U11488 ( .A(n6266), .B(keyinput27), .Z(n10414) );
  XOR2_X1 U11489 ( .A(n9657), .B(keyinput28), .Z(n10413) );
  XNOR2_X1 U11490 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput81), .ZN(n10412) );
  XNOR2_X1 U11491 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput68), .ZN(n10411)
         );
  NAND4_X1 U11492 ( .A1(n10414), .A2(n10413), .A3(n10412), .A4(n10411), .ZN(
        n10415) );
  NOR3_X1 U11493 ( .A1(n10417), .A2(n10416), .A3(n10415), .ZN(n10418) );
  NAND4_X1 U11494 ( .A1(n10421), .A2(n10420), .A3(n10419), .A4(n10418), .ZN(
        n10598) );
  AOI22_X1 U11495 ( .A1(n10424), .A2(keyinput15), .B1(keyinput22), .B2(n10423), 
        .ZN(n10422) );
  OAI221_X1 U11496 ( .B1(n10424), .B2(keyinput15), .C1(n10423), .C2(keyinput22), .A(n10422), .ZN(n10434) );
  AOI22_X1 U11497 ( .A1(n10426), .A2(keyinput117), .B1(keyinput61), .B2(n9568), 
        .ZN(n10425) );
  OAI221_X1 U11498 ( .B1(n10426), .B2(keyinput117), .C1(n9568), .C2(keyinput61), .A(n10425), .ZN(n10433) );
  XNOR2_X1 U11499 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput1), .ZN(n10429) );
  XNOR2_X1 U11500 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput34), .ZN(n10428)
         );
  XNOR2_X1 U11501 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput93), .ZN(n10427) );
  NAND3_X1 U11502 ( .A1(n10429), .A2(n10428), .A3(n10427), .ZN(n10432) );
  XNOR2_X1 U11503 ( .A(n10430), .B(keyinput40), .ZN(n10431) );
  NOR4_X1 U11504 ( .A1(n10434), .A2(n10433), .A3(n10432), .A4(n10431), .ZN(
        n10479) );
  AOI22_X1 U11505 ( .A1(n10436), .A2(keyinput14), .B1(keyinput55), .B2(n7736), 
        .ZN(n10435) );
  OAI221_X1 U11506 ( .B1(n10436), .B2(keyinput14), .C1(n7736), .C2(keyinput55), 
        .A(n10435), .ZN(n10448) );
  AOI22_X1 U11507 ( .A1(n10439), .A2(keyinput71), .B1(n10438), .B2(keyinput23), 
        .ZN(n10437) );
  OAI221_X1 U11508 ( .B1(n10439), .B2(keyinput71), .C1(n10438), .C2(keyinput23), .A(n10437), .ZN(n10447) );
  INV_X1 U11509 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10442) );
  AOI22_X1 U11510 ( .A1(n10442), .A2(keyinput33), .B1(n10441), .B2(keyinput97), 
        .ZN(n10440) );
  OAI221_X1 U11511 ( .B1(n10442), .B2(keyinput33), .C1(n10441), .C2(keyinput97), .A(n10440), .ZN(n10446) );
  XNOR2_X1 U11512 ( .A(P2_REG1_REG_12__SCAN_IN), .B(keyinput82), .ZN(n10444)
         );
  XNOR2_X1 U11513 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput9), .ZN(n10443) );
  NAND2_X1 U11514 ( .A1(n10444), .A2(n10443), .ZN(n10445) );
  NOR4_X1 U11515 ( .A1(n10448), .A2(n10447), .A3(n10446), .A4(n10445), .ZN(
        n10478) );
  AOI22_X1 U11516 ( .A1(n10450), .A2(keyinput83), .B1(n6395), .B2(keyinput12), 
        .ZN(n10449) );
  OAI221_X1 U11517 ( .B1(n10450), .B2(keyinput83), .C1(n6395), .C2(keyinput12), 
        .A(n10449), .ZN(n10462) );
  AOI22_X1 U11518 ( .A1(n10453), .A2(keyinput101), .B1(keyinput52), .B2(n10452), .ZN(n10451) );
  OAI221_X1 U11519 ( .B1(n10453), .B2(keyinput101), .C1(n10452), .C2(
        keyinput52), .A(n10451), .ZN(n10461) );
  INV_X1 U11520 ( .A(SI_13_), .ZN(n10455) );
  AOI22_X1 U11521 ( .A1(n10456), .A2(keyinput70), .B1(n10455), .B2(keyinput25), 
        .ZN(n10454) );
  OAI221_X1 U11522 ( .B1(n10456), .B2(keyinput70), .C1(n10455), .C2(keyinput25), .A(n10454), .ZN(n10460) );
  XNOR2_X1 U11523 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(keyinput59), .ZN(n10458)
         );
  XNOR2_X1 U11524 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput37), .ZN(n10457) );
  NAND2_X1 U11525 ( .A1(n10458), .A2(n10457), .ZN(n10459) );
  NOR4_X1 U11526 ( .A1(n10462), .A2(n10461), .A3(n10460), .A4(n10459), .ZN(
        n10477) );
  AOI22_X1 U11527 ( .A1(n10465), .A2(keyinput74), .B1(keyinput78), .B2(n10464), 
        .ZN(n10463) );
  OAI221_X1 U11528 ( .B1(n10465), .B2(keyinput74), .C1(n10464), .C2(keyinput78), .A(n10463), .ZN(n10475) );
  AOI22_X1 U11529 ( .A1(n10468), .A2(keyinput79), .B1(n10467), .B2(keyinput31), 
        .ZN(n10466) );
  OAI221_X1 U11530 ( .B1(n10468), .B2(keyinput79), .C1(n10467), .C2(keyinput31), .A(n10466), .ZN(n10474) );
  XOR2_X1 U11531 ( .A(n7846), .B(keyinput100), .Z(n10472) );
  XNOR2_X1 U11532 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(keyinput8), .ZN(n10471) );
  XNOR2_X1 U11533 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput87), .ZN(n10470) );
  XNOR2_X1 U11534 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput124), .ZN(n10469) );
  NAND4_X1 U11535 ( .A1(n10472), .A2(n10471), .A3(n10470), .A4(n10469), .ZN(
        n10473) );
  NOR3_X1 U11536 ( .A1(n10475), .A2(n10474), .A3(n10473), .ZN(n10476) );
  NAND4_X1 U11537 ( .A1(n10479), .A2(n10478), .A3(n10477), .A4(n10476), .ZN(
        n10597) );
  AOI22_X1 U11538 ( .A1(n10482), .A2(keyinput46), .B1(keyinput30), .B2(n10481), 
        .ZN(n10480) );
  OAI221_X1 U11539 ( .B1(n10482), .B2(keyinput46), .C1(n10481), .C2(keyinput30), .A(n10480), .ZN(n10494) );
  AOI22_X1 U11540 ( .A1(n10485), .A2(keyinput121), .B1(keyinput120), .B2(
        n10484), .ZN(n10483) );
  OAI221_X1 U11541 ( .B1(n10485), .B2(keyinput121), .C1(n10484), .C2(
        keyinput120), .A(n10483), .ZN(n10493) );
  AOI22_X1 U11542 ( .A1(n10488), .A2(keyinput88), .B1(keyinput84), .B2(n10487), 
        .ZN(n10486) );
  OAI221_X1 U11543 ( .B1(n10488), .B2(keyinput88), .C1(n10487), .C2(keyinput84), .A(n10486), .ZN(n10492) );
  XNOR2_X1 U11544 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(keyinput5), .ZN(n10490)
         );
  XNOR2_X1 U11545 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(keyinput108), .ZN(n10489)
         );
  NAND2_X1 U11546 ( .A1(n10490), .A2(n10489), .ZN(n10491) );
  NOR4_X1 U11547 ( .A1(n10494), .A2(n10493), .A3(n10492), .A4(n10491), .ZN(
        n10537) );
  AOI22_X1 U11548 ( .A1(n10496), .A2(keyinput118), .B1(keyinput39), .B2(n5414), 
        .ZN(n10495) );
  OAI221_X1 U11549 ( .B1(n10496), .B2(keyinput118), .C1(n5414), .C2(keyinput39), .A(n10495), .ZN(n10505) );
  AOI22_X1 U11550 ( .A1(n10498), .A2(keyinput99), .B1(n5689), .B2(keyinput53), 
        .ZN(n10497) );
  OAI221_X1 U11551 ( .B1(n10498), .B2(keyinput99), .C1(n5689), .C2(keyinput53), 
        .A(n10497), .ZN(n10504) );
  XOR2_X1 U11552 ( .A(n6179), .B(keyinput41), .Z(n10502) );
  XNOR2_X1 U11553 ( .A(P1_REG1_REG_2__SCAN_IN), .B(keyinput94), .ZN(n10501) );
  XNOR2_X1 U11554 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput62), .ZN(n10500) );
  XNOR2_X1 U11555 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput107), .ZN(n10499)
         );
  NAND4_X1 U11556 ( .A1(n10502), .A2(n10501), .A3(n10500), .A4(n10499), .ZN(
        n10503) );
  NOR3_X1 U11557 ( .A1(n10505), .A2(n10504), .A3(n10503), .ZN(n10536) );
  AOI22_X1 U11558 ( .A1(n10508), .A2(keyinput44), .B1(keyinput98), .B2(n10507), 
        .ZN(n10506) );
  OAI221_X1 U11559 ( .B1(n10508), .B2(keyinput44), .C1(n10507), .C2(keyinput98), .A(n10506), .ZN(n10518) );
  AOI22_X1 U11560 ( .A1(n10511), .A2(keyinput57), .B1(n10510), .B2(keyinput85), 
        .ZN(n10509) );
  OAI221_X1 U11561 ( .B1(n10511), .B2(keyinput57), .C1(n10510), .C2(keyinput85), .A(n10509), .ZN(n10517) );
  XNOR2_X1 U11562 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput127), .ZN(n10515)
         );
  XNOR2_X1 U11563 ( .A(P2_REG0_REG_23__SCAN_IN), .B(keyinput54), .ZN(n10514)
         );
  XNOR2_X1 U11564 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput67), .ZN(n10513) );
  XNOR2_X1 U11565 ( .A(keyinput60), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n10512) );
  NAND4_X1 U11566 ( .A1(n10515), .A2(n10514), .A3(n10513), .A4(n10512), .ZN(
        n10516) );
  NOR3_X1 U11567 ( .A1(n10518), .A2(n10517), .A3(n10516), .ZN(n10535) );
  AOI22_X1 U11568 ( .A1(n10521), .A2(keyinput19), .B1(n10520), .B2(keyinput26), 
        .ZN(n10519) );
  OAI221_X1 U11569 ( .B1(n10521), .B2(keyinput19), .C1(n10520), .C2(keyinput26), .A(n10519), .ZN(n10533) );
  AOI22_X1 U11570 ( .A1(n10523), .A2(keyinput48), .B1(n6827), .B2(keyinput122), 
        .ZN(n10522) );
  OAI221_X1 U11571 ( .B1(n10523), .B2(keyinput48), .C1(n6827), .C2(keyinput122), .A(n10522), .ZN(n10532) );
  AOI22_X1 U11572 ( .A1(n10526), .A2(keyinput24), .B1(keyinput21), .B2(n10525), 
        .ZN(n10524) );
  OAI221_X1 U11573 ( .B1(n10526), .B2(keyinput24), .C1(n10525), .C2(keyinput21), .A(n10524), .ZN(n10531) );
  AOI22_X1 U11574 ( .A1(n10529), .A2(keyinput20), .B1(n10528), .B2(keyinput119), .ZN(n10527) );
  OAI221_X1 U11575 ( .B1(n10529), .B2(keyinput20), .C1(n10528), .C2(
        keyinput119), .A(n10527), .ZN(n10530) );
  NOR4_X1 U11576 ( .A1(n10533), .A2(n10532), .A3(n10531), .A4(n10530), .ZN(
        n10534) );
  NAND4_X1 U11577 ( .A1(n10537), .A2(n10536), .A3(n10535), .A4(n10534), .ZN(
        n10596) );
  AOI22_X1 U11578 ( .A1(n8831), .A2(keyinput58), .B1(n10539), .B2(keyinput36), 
        .ZN(n10538) );
  OAI221_X1 U11579 ( .B1(n8831), .B2(keyinput58), .C1(n10539), .C2(keyinput36), 
        .A(n10538), .ZN(n10551) );
  AOI22_X1 U11580 ( .A1(n10542), .A2(keyinput65), .B1(n10541), .B2(keyinput42), 
        .ZN(n10540) );
  OAI221_X1 U11581 ( .B1(n10542), .B2(keyinput65), .C1(n10541), .C2(keyinput42), .A(n10540), .ZN(n10550) );
  AOI22_X1 U11582 ( .A1(n10545), .A2(keyinput29), .B1(n10544), .B2(keyinput11), 
        .ZN(n10543) );
  OAI221_X1 U11583 ( .B1(n10545), .B2(keyinput29), .C1(n10544), .C2(keyinput11), .A(n10543), .ZN(n10549) );
  XOR2_X1 U11584 ( .A(n5400), .B(keyinput63), .Z(n10547) );
  XNOR2_X1 U11585 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(keyinput80), .ZN(n10546)
         );
  NAND2_X1 U11586 ( .A1(n10547), .A2(n10546), .ZN(n10548) );
  NOR4_X1 U11587 ( .A1(n10551), .A2(n10550), .A3(n10549), .A4(n10548), .ZN(
        n10594) );
  INV_X1 U11588 ( .A(P1_WR_REG_SCAN_IN), .ZN(n10553) );
  AOI22_X1 U11589 ( .A1(n10554), .A2(keyinput64), .B1(keyinput66), .B2(n10553), 
        .ZN(n10552) );
  OAI221_X1 U11590 ( .B1(n10554), .B2(keyinput64), .C1(n10553), .C2(keyinput66), .A(n10552), .ZN(n10565) );
  AOI22_X1 U11591 ( .A1(keyinput86), .A2(n10556), .B1(keyinput7), .B2(n6353), 
        .ZN(n10555) );
  OAI21_X1 U11592 ( .B1(n10556), .B2(keyinput86), .A(n10555), .ZN(n10564) );
  AOI22_X1 U11593 ( .A1(n10559), .A2(keyinput89), .B1(n10558), .B2(keyinput77), 
        .ZN(n10557) );
  OAI221_X1 U11594 ( .B1(n10559), .B2(keyinput89), .C1(n10558), .C2(keyinput77), .A(n10557), .ZN(n10563) );
  XOR2_X1 U11595 ( .A(n5552), .B(keyinput56), .Z(n10561) );
  XNOR2_X1 U11596 ( .A(SI_1_), .B(keyinput43), .ZN(n10560) );
  NAND2_X1 U11597 ( .A1(n10561), .A2(n10560), .ZN(n10562) );
  NOR4_X1 U11598 ( .A1(n10565), .A2(n10564), .A3(n10563), .A4(n10562), .ZN(
        n10593) );
  AOI22_X1 U11599 ( .A1(n10567), .A2(keyinput49), .B1(n6217), .B2(keyinput90), 
        .ZN(n10566) );
  OAI221_X1 U11600 ( .B1(n10567), .B2(keyinput49), .C1(n6217), .C2(keyinput90), 
        .A(n10566), .ZN(n10579) );
  INV_X1 U11601 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10569) );
  AOI22_X1 U11602 ( .A1(n10570), .A2(keyinput105), .B1(keyinput50), .B2(n10569), .ZN(n10568) );
  OAI221_X1 U11603 ( .B1(n10570), .B2(keyinput105), .C1(n10569), .C2(
        keyinput50), .A(n10568), .ZN(n10578) );
  AOI22_X1 U11604 ( .A1(n10573), .A2(keyinput6), .B1(keyinput38), .B2(n10572), 
        .ZN(n10571) );
  OAI221_X1 U11605 ( .B1(n10573), .B2(keyinput6), .C1(n10572), .C2(keyinput38), 
        .A(n10571), .ZN(n10577) );
  XNOR2_X1 U11606 ( .A(P1_REG0_REG_26__SCAN_IN), .B(keyinput13), .ZN(n10575)
         );
  XNOR2_X1 U11607 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput4), .ZN(n10574) );
  NAND2_X1 U11608 ( .A1(n10575), .A2(n10574), .ZN(n10576) );
  NOR4_X1 U11609 ( .A1(n10579), .A2(n10578), .A3(n10577), .A4(n10576), .ZN(
        n10592) );
  AOI22_X1 U11610 ( .A1(n10581), .A2(keyinput95), .B1(keyinput123), .B2(n5136), 
        .ZN(n10580) );
  OAI221_X1 U11611 ( .B1(n10581), .B2(keyinput95), .C1(n5136), .C2(keyinput123), .A(n10580), .ZN(n10590) );
  AOI22_X1 U11612 ( .A1(n10583), .A2(keyinput76), .B1(keyinput110), .B2(n10339), .ZN(n10582) );
  OAI221_X1 U11613 ( .B1(n10583), .B2(keyinput76), .C1(n10339), .C2(
        keyinput110), .A(n10582), .ZN(n10589) );
  XOR2_X1 U11614 ( .A(n6578), .B(keyinput112), .Z(n10587) );
  XNOR2_X1 U11615 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(keyinput32), .ZN(n10586)
         );
  XNOR2_X1 U11616 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput91), .ZN(n10585) );
  XNOR2_X1 U11617 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput125), .ZN(n10584) );
  NAND4_X1 U11618 ( .A1(n10587), .A2(n10586), .A3(n10585), .A4(n10584), .ZN(
        n10588) );
  NOR3_X1 U11619 ( .A1(n10590), .A2(n10589), .A3(n10588), .ZN(n10591) );
  NAND4_X1 U11620 ( .A1(n10594), .A2(n10593), .A3(n10592), .A4(n10591), .ZN(
        n10595) );
  NOR4_X1 U11621 ( .A1(n10598), .A2(n10597), .A3(n10596), .A4(n10595), .ZN(
        n10599) );
  OAI21_X1 U11622 ( .B1(keyinput7), .B2(n10600), .A(n10599), .ZN(n10601) );
  XOR2_X1 U11623 ( .A(n10602), .B(n10601), .Z(P2_U3182) );
  XNOR2_X1 U11624 ( .A(n10604), .B(n10603), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11625 ( .A(n10606), .B(n10605), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11626 ( .A(n10608), .B(n10607), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11627 ( .A(n10610), .B(n10609), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11628 ( .A(n10612), .B(n10611), .ZN(ADD_1068_U48) );
  XOR2_X1 U11629 ( .A(n10614), .B(n10613), .Z(ADD_1068_U54) );
  XOR2_X1 U11630 ( .A(n10616), .B(n10615), .Z(ADD_1068_U53) );
  XNOR2_X1 U11631 ( .A(n10618), .B(n10617), .ZN(ADD_1068_U52) );
  NAND2_X1 U4916 ( .A1(n4577), .A2(n6176), .ZN(n6238) );
endmodule

