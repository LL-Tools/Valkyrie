

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16036;

  NAND2_X1 U7285 ( .A1(n13208), .A2(n13207), .ZN(n14926) );
  INV_X1 U7286 ( .A(n14503), .ZN(n14540) );
  NOR2_X1 U7287 ( .A1(n7999), .A2(n7007), .ZN(n7006) );
  NAND2_X1 U7288 ( .A1(n9729), .A2(n9728), .ZN(n14732) );
  NAND2_X2 U7289 ( .A1(n10871), .A2(n10790), .ZN(n11908) );
  INV_X1 U7291 ( .A(n14107), .ZN(n15924) );
  NAND2_X2 U7292 ( .A1(n10871), .A2(n10957), .ZN(n13195) );
  CLKBUF_X1 U7293 ( .A(n8174), .Z(n6549) );
  CLKBUF_X2 U7294 ( .A(n8863), .Z(n9308) );
  NOR2_X2 U7295 ( .A1(n8160), .A2(n8159), .ZN(n10860) );
  NAND4_X1 U7296 ( .A1(n9436), .A2(n9435), .A3(n9434), .A4(n9882), .ZN(n9878)
         );
  NAND3_X1 U7297 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n8937) );
  AOI21_X1 U7298 ( .B1(n6957), .B2(n6956), .A(n13652), .ZN(n13128) );
  NOR2_X1 U7299 ( .A1(n6807), .A2(n9878), .ZN(n6806) );
  INV_X2 U7300 ( .A(n9020), .ZN(n9131) );
  INV_X1 U7302 ( .A(n8136), .ZN(n7166) );
  INV_X2 U7303 ( .A(n13101), .ZN(n13124) );
  INV_X1 U7304 ( .A(n13223), .ZN(n13235) );
  INV_X4 U7305 ( .A(n13224), .ZN(n13189) );
  AND4_X1 U7306 ( .A1(n8685), .A2(n8683), .A3(n8684), .A4(n9016), .ZN(n8690)
         );
  INV_X2 U7307 ( .A(n12261), .ZN(n6545) );
  AND2_X1 U7308 ( .A1(n13638), .A2(n13833), .ZN(n13642) );
  CLKBUF_X3 U7309 ( .A(n7166), .Z(n6538) );
  AND2_X1 U7310 ( .A1(n6797), .A2(n7285), .ZN(n14367) );
  INV_X1 U7311 ( .A(n14214), .ZN(n12104) );
  NOR2_X1 U7312 ( .A1(n7165), .A2(n15941), .ZN(n7106) );
  INV_X1 U7313 ( .A(n14620), .ZN(n14759) );
  NAND2_X1 U7314 ( .A1(n8855), .A2(n15674), .ZN(n8843) );
  INV_X1 U7315 ( .A(n15591), .ZN(n8753) );
  NAND2_X1 U7316 ( .A1(n15165), .A2(n15169), .ZN(n15204) );
  INV_X1 U7317 ( .A(n12001), .ZN(n15821) );
  NAND2_X2 U7319 ( .A1(n9468), .A2(n9467), .ZN(n14705) );
  NAND2_X2 U7320 ( .A1(n9265), .A2(n9264), .ZN(n15488) );
  INV_X1 U7321 ( .A(n15392), .ZN(n15748) );
  XNOR2_X1 U7322 ( .A(n9066), .B(n9065), .ZN(n10783) );
  NAND2_X1 U7323 ( .A1(n8178), .A2(n7169), .ZN(n13462) );
  NAND2_X1 U7324 ( .A1(n8126), .A2(n14001), .ZN(n14008) );
  AND2_X1 U7325 ( .A1(n9655), .A2(n9654), .ZN(n14816) );
  INV_X1 U7326 ( .A(n9461), .ZN(n14828) );
  INV_X1 U7327 ( .A(n11860), .ZN(n14332) );
  INV_X1 U7328 ( .A(n12426), .ZN(n15828) );
  NAND2_X1 U7329 ( .A1(n9013), .A2(n8990), .ZN(n10657) );
  OR2_X2 U7331 ( .A1(n7816), .A2(n11519), .ZN(n7424) );
  XNOR2_X2 U7334 ( .A(n8700), .B(n8698), .ZN(n15591) );
  NAND2_X1 U7335 ( .A1(n11504), .A2(n9384), .ZN(n15750) );
  AOI21_X2 U7336 ( .B1(n15647), .B2(n15646), .A(n15645), .ZN(n15655) );
  NOR2_X2 U7337 ( .A1(n10729), .A2(n10730), .ZN(n10728) );
  OAI222_X1 U7338 ( .A1(n15597), .A2(n13277), .B1(P1_U3086), .B2(n13276), .C1(
        n15595), .C2(n13278), .ZN(P1_U3325) );
  OR2_X1 U7339 ( .A1(n13276), .A2(n8753), .ZN(n9273) );
  AOI22_X2 U7340 ( .A1(n11845), .A2(n11844), .B1(n8264), .B2(n13456), .ZN(
        n12193) );
  NAND2_X2 U7341 ( .A1(n8253), .A2(n7709), .ZN(n11280) );
  NAND2_X2 U7342 ( .A1(n8066), .A2(n8064), .ZN(n8068) );
  INV_X2 U7343 ( .A(n7924), .ZN(n8066) );
  NAND2_X1 U7344 ( .A1(n8128), .A2(n14008), .ZN(n8175) );
  INV_X1 U7345 ( .A(n8546), .ZN(n11630) );
  CLKBUF_X1 U7346 ( .A(n7166), .Z(n6537) );
  XNOR2_X1 U7348 ( .A(n8713), .B(n8712), .ZN(n15392) );
  AND2_X1 U7349 ( .A1(n10808), .A2(n10807), .ZN(n6540) );
  AND2_X2 U7350 ( .A1(n10375), .A2(n9853), .ZN(n11861) );
  OAI22_X2 U7354 ( .A1(n9231), .A2(n8662), .B1(n9229), .B2(SI_23_), .ZN(n8663)
         );
  XNOR2_X1 U7355 ( .A(n8548), .B(P3_IR_REG_22__SCAN_IN), .ZN(n13146) );
  OAI211_X1 U7356 ( .C1(n6943), .C2(n14918), .A(n14916), .B(n6940), .ZN(n14967) );
  NAND2_X1 U7357 ( .A1(n9806), .A2(n9805), .ZN(n14369) );
  NAND2_X1 U7358 ( .A1(n12707), .A2(n9394), .ZN(n15235) );
  NAND2_X1 U7359 ( .A1(n9282), .A2(n9281), .ZN(n15482) );
  NAND2_X1 U7361 ( .A1(n9747), .A2(n9746), .ZN(n14515) );
  NAND2_X1 U7362 ( .A1(n8997), .A2(n8996), .ZN(n12426) );
  NAND2_X1 U7363 ( .A1(n9615), .A2(n9614), .ZN(n12242) );
  NAND2_X1 U7364 ( .A1(n8836), .A2(n8835), .ZN(n15812) );
  NAND2_X1 U7365 ( .A1(n10900), .A2(n15991), .ZN(n7938) );
  INV_X2 U7366 ( .A(n15764), .ZN(n6544) );
  INV_X2 U7367 ( .A(n15439), .ZN(n15780) );
  NOR2_X1 U7368 ( .A1(n10450), .A2(n13274), .ZN(n10417) );
  INV_X1 U7369 ( .A(n15745), .ZN(n10985) );
  NAND2_X2 U7370 ( .A1(n11434), .A2(n10876), .ZN(n13223) );
  INV_X4 U7371 ( .A(n13195), .ZN(n10876) );
  BUF_X1 U7372 ( .A(n8175), .Z(n6547) );
  INV_X4 U7373 ( .A(n6793), .ZN(n10321) );
  INV_X2 U7374 ( .A(n9517), .ZN(n7527) );
  NAND2_X2 U7375 ( .A1(n9484), .A2(n9478), .ZN(n9507) );
  NAND2_X2 U7376 ( .A1(n8136), .A2(n7219), .ZN(n12950) );
  CLKBUF_X2 U7377 ( .A(n8906), .Z(n9296) );
  NAND2_X1 U7378 ( .A1(n7182), .A2(n7179), .ZN(n15674) );
  NAND2_X1 U7379 ( .A1(n8614), .A2(SI_6_), .ZN(n8829) );
  AND2_X1 U7381 ( .A1(n9421), .A2(n9420), .ZN(n9625) );
  INV_X4 U7382 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  OR2_X1 U7383 ( .A1(n10401), .A2(n10372), .ZN(n10403) );
  AND2_X1 U7384 ( .A1(n7874), .A2(n7877), .ZN(n7873) );
  OAI21_X1 U7385 ( .B1(n13637), .B2(n13636), .A(n13635), .ZN(n13643) );
  NOR2_X1 U7386 ( .A1(n14336), .A2(n14658), .ZN(n14676) );
  NAND2_X1 U7387 ( .A1(n12735), .A2(n12734), .ZN(n12737) );
  NAND2_X1 U7388 ( .A1(n14941), .A2(n13201), .ZN(n14860) );
  NOR2_X1 U7389 ( .A1(n7565), .A2(n7240), .ZN(n7457) );
  OR3_X1 U7390 ( .A1(n14719), .A2(n14718), .A3(n14717), .ZN(n14795) );
  NAND2_X1 U7391 ( .A1(n14072), .A2(n7536), .ZN(n14096) );
  OR2_X1 U7392 ( .A1(n10306), .A2(n7566), .ZN(n7565) );
  NAND2_X1 U7393 ( .A1(n6792), .A2(n7282), .ZN(n7882) );
  NAND2_X1 U7394 ( .A1(n13317), .A2(n8460), .ZN(n10153) );
  NAND2_X1 U7395 ( .A1(n12897), .A2(n12896), .ZN(n13717) );
  AOI211_X1 U7396 ( .C1(n13417), .C2(n6577), .A(n6639), .B(n6553), .ZN(n7381)
         );
  NAND2_X1 U7397 ( .A1(n14157), .A2(n12777), .ZN(n14032) );
  OAI21_X1 U7398 ( .B1(n6569), .B2(n6664), .A(n7947), .ZN(n7946) );
  OAI21_X1 U7399 ( .B1(n14423), .B2(n6560), .A(n7281), .ZN(n7280) );
  AND2_X1 U7400 ( .A1(n7082), .A2(n13492), .ZN(n13471) );
  XNOR2_X1 U7401 ( .A(n8759), .B(n8758), .ZN(n14825) );
  NAND2_X1 U7402 ( .A1(n12690), .A2(n12689), .ZN(n15402) );
  XNOR2_X1 U7403 ( .A(n14705), .B(n14077), .ZN(n14428) );
  NAND2_X1 U7404 ( .A1(n13796), .A2(n13079), .ZN(n13785) );
  NAND2_X1 U7405 ( .A1(n7155), .A2(n8673), .ZN(n8759) );
  NAND2_X1 U7406 ( .A1(n13470), .A2(n13486), .ZN(n13492) );
  OAI21_X1 U7407 ( .B1(n9831), .B2(n7886), .A(n6696), .ZN(n6795) );
  NAND2_X1 U7408 ( .A1(n9311), .A2(n9310), .ZN(n15213) );
  AND2_X1 U7409 ( .A1(n9288), .A2(n10335), .ZN(n7564) );
  XNOR2_X1 U7410 ( .A(n14700), .B(n14169), .ZN(n14417) );
  NAND2_X1 U7411 ( .A1(n12602), .A2(n12608), .ZN(n12690) );
  NAND2_X1 U7412 ( .A1(n9302), .A2(n9301), .ZN(n14998) );
  OR2_X1 U7413 ( .A1(n9332), .A2(n9331), .ZN(n7155) );
  XNOR2_X1 U7414 ( .A(n9332), .B(n9331), .ZN(n13258) );
  NAND2_X1 U7415 ( .A1(n6914), .A2(n6915), .ZN(n13798) );
  NAND2_X1 U7416 ( .A1(n12220), .A2(n10335), .ZN(n9468) );
  OR2_X2 U7417 ( .A1(n14581), .A2(n14566), .ZN(n14564) );
  AND2_X1 U7418 ( .A1(n9263), .A2(n9262), .ZN(n12220) );
  NAND2_X1 U7419 ( .A1(n11625), .A2(n11624), .ZN(n11825) );
  NAND2_X1 U7420 ( .A1(n13386), .A2(n8340), .ZN(n7905) );
  NAND2_X1 U7421 ( .A1(n7159), .A2(n12530), .ZN(n12885) );
  XNOR2_X1 U7422 ( .A(n9280), .B(n9279), .ZN(n12477) );
  NAND2_X1 U7423 ( .A1(n7906), .A2(n13329), .ZN(n13386) );
  NAND2_X1 U7424 ( .A1(n15369), .A2(n12716), .ZN(n15405) );
  NAND2_X1 U7425 ( .A1(n7164), .A2(SI_24_), .ZN(n7572) );
  NAND2_X1 U7426 ( .A1(n7571), .A2(n9259), .ZN(n7570) );
  NAND2_X1 U7427 ( .A1(n9234), .A2(n9233), .ZN(n15265) );
  INV_X1 U7428 ( .A(n14754), .ZN(n14605) );
  OR2_X1 U7429 ( .A1(n15543), .A2(n15412), .ZN(n15370) );
  NAND2_X1 U7430 ( .A1(n6794), .A2(n9821), .ZN(n7292) );
  AND2_X1 U7431 ( .A1(n9823), .A2(n7898), .ZN(n6794) );
  NAND2_X1 U7432 ( .A1(n7734), .A2(n9679), .ZN(n14754) );
  AND2_X1 U7433 ( .A1(n9054), .A2(n9053), .ZN(n15419) );
  NOR2_X1 U7434 ( .A1(n14632), .A2(n7902), .ZN(n7901) );
  NAND2_X1 U7435 ( .A1(n12057), .A2(n7548), .ZN(n12346) );
  XNOR2_X1 U7436 ( .A(n9211), .B(n9210), .ZN(n11550) );
  AND2_X1 U7437 ( .A1(n12275), .A2(n12236), .ZN(n9823) );
  NAND2_X1 U7438 ( .A1(n7016), .A2(n12049), .ZN(n12057) );
  AOI21_X1 U7439 ( .B1(n7384), .B2(n7389), .A(n8327), .ZN(n7383) );
  AND2_X1 U7440 ( .A1(n9064), .A2(n9048), .ZN(n10776) );
  NAND2_X1 U7441 ( .A1(n9019), .A2(n9018), .ZN(n15559) );
  XNOR2_X1 U7442 ( .A(n7404), .B(n9153), .ZN(n11346) );
  NAND2_X1 U7443 ( .A1(n9207), .A2(n9191), .ZN(n12824) );
  NAND2_X1 U7444 ( .A1(n7406), .A2(n7405), .ZN(n7404) );
  NAND2_X1 U7445 ( .A1(n9710), .A2(n9709), .ZN(n14566) );
  OR2_X1 U7446 ( .A1(n9190), .A2(n9189), .ZN(n9207) );
  NAND2_X1 U7447 ( .A1(n9105), .A2(n9104), .ZN(n15531) );
  NAND3_X1 U7448 ( .A1(n10991), .A2(n10990), .A3(n10995), .ZN(n11351) );
  NOR2_X1 U7449 ( .A1(n11760), .A2(n15812), .ZN(n11950) );
  OR2_X1 U7450 ( .A1(n9150), .A2(SI_18_), .ZN(n7405) );
  NOR2_X1 U7451 ( .A1(n9606), .A2(n10388), .ZN(n9607) );
  XNOR2_X1 U7452 ( .A(n8774), .B(n6786), .ZN(n10646) );
  AOI21_X1 U7453 ( .B1(n9099), .B2(n8646), .A(n6558), .ZN(n9149) );
  INV_X1 U7454 ( .A(n12366), .ZN(n12468) );
  NAND2_X2 U7455 ( .A1(n11859), .A2(n14642), .ZN(n14645) );
  NAND2_X1 U7456 ( .A1(n11234), .A2(n11327), .ZN(n11337) );
  NAND2_X1 U7457 ( .A1(n7135), .A2(n7133), .ZN(n9099) );
  AND2_X1 U7458 ( .A1(n9596), .A2(n9595), .ZN(n12366) );
  NAND2_X1 U7459 ( .A1(n7745), .A2(n8624), .ZN(n8987) );
  AND2_X1 U7460 ( .A1(n8914), .A2(n11507), .ZN(n11539) );
  NAND2_X1 U7461 ( .A1(n8949), .A2(n8948), .ZN(n11742) );
  XNOR2_X1 U7462 ( .A(n8978), .B(n8979), .ZN(n10621) );
  INV_X1 U7463 ( .A(n11521), .ZN(n11525) );
  INV_X1 U7464 ( .A(n12407), .ZN(n6802) );
  AND2_X1 U7465 ( .A1(n13028), .A2(n13027), .ZN(n13025) );
  XNOR2_X1 U7466 ( .A(n14216), .B(n12099), .ZN(n12091) );
  AND2_X1 U7467 ( .A1(n7748), .A2(n6601), .ZN(n8979) );
  AND2_X1 U7468 ( .A1(n8928), .A2(n8927), .ZN(n11521) );
  NAND2_X1 U7469 ( .A1(n8806), .A2(n8621), .ZN(n7748) );
  INV_X1 U7470 ( .A(n13462), .ZN(n15991) );
  AND2_X1 U7471 ( .A1(n6803), .A2(n9516), .ZN(n12407) );
  NOR2_X1 U7472 ( .A1(n13464), .A2(n11399), .ZN(n15980) );
  NAND2_X1 U7473 ( .A1(n7122), .A2(n8611), .ZN(n8790) );
  AND2_X1 U7474 ( .A1(n7134), .A2(n8641), .ZN(n7133) );
  NAND3_X1 U7475 ( .A1(n8158), .A2(n8157), .A3(n8156), .ZN(n8160) );
  INV_X1 U7476 ( .A(n12085), .ZN(n14215) );
  AND4_X1 U7477 ( .A1(n9506), .A2(n9505), .A3(n9504), .A4(n9503), .ZN(n12085)
         );
  NAND4_X1 U7478 ( .A1(n9533), .A2(n9532), .A3(n9531), .A4(n9530), .ZN(n14213)
         );
  NAND4_X1 U7479 ( .A1(n9493), .A2(n9492), .A3(n9491), .A4(n9490), .ZN(n10168)
         );
  AND4_X1 U7480 ( .A1(n9500), .A2(n9499), .A3(n9498), .A4(n9497), .ZN(n13274)
         );
  NAND4_X1 U7481 ( .A1(n9522), .A2(n9521), .A3(n9520), .A4(n9519), .ZN(n14214)
         );
  OAI211_X1 U7482 ( .C1(n8136), .C2(n11125), .A(n7064), .B(n7062), .ZN(n15972)
         );
  NAND3_X1 U7483 ( .A1(n9499), .A2(n7528), .A3(n9500), .ZN(n14216) );
  NAND4_X1 U7484 ( .A1(n8891), .A2(n8890), .A3(n8889), .A4(n8888), .ZN(n15745)
         );
  INV_X2 U7485 ( .A(n8579), .ZN(n13101) );
  INV_X2 U7486 ( .A(n9793), .ZN(n10335) );
  AND3_X1 U7487 ( .A1(n8188), .A2(n8187), .A3(n8186), .ZN(n10929) );
  NAND4_X1 U7488 ( .A1(n8932), .A2(n8931), .A3(n8930), .A4(n8929), .ZN(n15018)
         );
  NAND2_X1 U7489 ( .A1(n7021), .A2(n14332), .ZN(n7019) );
  AOI21_X1 U7490 ( .B1(n7559), .B2(n7557), .A(n7556), .ZN(n7555) );
  INV_X2 U7491 ( .A(n6547), .ZN(n12939) );
  AND2_X1 U7492 ( .A1(n12938), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8159) );
  CLKBUF_X1 U7493 ( .A(n8175), .Z(n6548) );
  AND2_X2 U7494 ( .A1(n13255), .A2(n8127), .ZN(n12938) );
  CLKBUF_X2 U7495 ( .A(n12951), .Z(n7252) );
  INV_X2 U7496 ( .A(n12950), .ZN(n12935) );
  INV_X2 U7497 ( .A(n10325), .ZN(n10328) );
  NAND2_X2 U7498 ( .A1(n10957), .A2(n6953), .ZN(n13224) );
  CLKBUF_X1 U7499 ( .A(n8886), .Z(n9323) );
  NAND2_X1 U7500 ( .A1(n8886), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n8867) );
  INV_X2 U7501 ( .A(n8897), .ZN(n9333) );
  AOI21_X1 U7502 ( .B1(n8640), .B2(n9118), .A(n8639), .ZN(n8641) );
  XNOR2_X1 U7503 ( .A(n9430), .B(n9429), .ZN(n9433) );
  NAND2_X1 U7504 ( .A1(n8843), .A2(n7219), .ZN(n8897) );
  INV_X2 U7505 ( .A(n8843), .ZN(n9154) );
  NAND2_X4 U7506 ( .A1(n14828), .A2(n13279), .ZN(n6793) );
  AOI22_X1 U7507 ( .A1(n8650), .A2(n8649), .B1(n10967), .B2(n9152), .ZN(n8651)
         );
  CLKBUF_X1 U7508 ( .A(n9273), .Z(n7213) );
  NAND2_X1 U7509 ( .A1(n14828), .A2(n7108), .ZN(n10325) );
  INV_X1 U7510 ( .A(n9035), .ZN(n8634) );
  NAND2_X1 U7511 ( .A1(n8078), .A2(n8547), .ZN(n11492) );
  OAI21_X1 U7512 ( .B1(n8614), .B2(SI_6_), .A(n8829), .ZN(n8787) );
  NAND2_X1 U7513 ( .A1(n8204), .A2(n8220), .ZN(n11302) );
  NAND2_X1 U7514 ( .A1(n9871), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9430) );
  OAI21_X1 U7515 ( .B1(n8633), .B2(SI_13_), .A(n8635), .ZN(n9035) );
  INV_X1 U7516 ( .A(n7109), .ZN(n13279) );
  NAND2_X4 U7517 ( .A1(n12879), .A2(n13576), .ZN(n8136) );
  NAND2_X1 U7518 ( .A1(n8075), .A2(n8074), .ZN(n8547) );
  XNOR2_X1 U7519 ( .A(n8642), .B(SI_16_), .ZN(n9120) );
  XNOR2_X1 U7520 ( .A(n9432), .B(P2_IR_REG_19__SCAN_IN), .ZN(n11860) );
  OR2_X1 U7521 ( .A1(n9425), .A2(n9693), .ZN(n9427) );
  MUX2_X1 U7522 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8124), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n8126) );
  OAI21_X1 U7523 ( .B1(n8622), .B2(SI_9_), .A(n8624), .ZN(n8978) );
  NAND2_X1 U7524 ( .A1(n8633), .A2(SI_13_), .ZN(n8635) );
  XNOR2_X1 U7525 ( .A(n9424), .B(P2_IR_REG_21__SCAN_IN), .ZN(n10375) );
  NAND2_X1 U7526 ( .A1(n7769), .A2(n7768), .ZN(n9871) );
  XNOR2_X1 U7527 ( .A(n9460), .B(P2_IR_REG_29__SCAN_IN), .ZN(n9461) );
  NAND2_X1 U7528 ( .A1(n8068), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8065) );
  NAND2_X1 U7529 ( .A1(n9431), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9432) );
  AND2_X1 U7530 ( .A1(n8085), .A2(n8088), .ZN(n8094) );
  INV_X2 U7531 ( .A(n13999), .ZN(n13257) );
  XNOR2_X1 U7532 ( .A(n9372), .B(n9371), .ZN(n12222) );
  NAND2_X1 U7533 ( .A1(n9370), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9372) );
  NAND2_X2 U7534 ( .A1(n7176), .A2(P3_U3151), .ZN(n14006) );
  NOR2_X1 U7535 ( .A1(n8597), .A2(n8844), .ZN(n8850) );
  OR2_X1 U7536 ( .A1(n8125), .A2(n8121), .ZN(n8122) );
  NAND2_X2 U7537 ( .A1(n6542), .A2(P1_U3086), .ZN(n15597) );
  NAND2_X1 U7538 ( .A1(n15586), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7823) );
  NAND2_X1 U7539 ( .A1(n8695), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8693) );
  BUF_X4 U7540 ( .A(n6541), .Z(n7176) );
  OAI21_X1 U7541 ( .B1(n8556), .B2(n8081), .A(n8080), .ZN(n8085) );
  NAND2_X2 U7542 ( .A1(n8069), .A2(P1_U3086), .ZN(n15595) );
  OR2_X1 U7543 ( .A1(n9366), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n9370) );
  OR2_X1 U7544 ( .A1(n6987), .A2(n6986), .ZN(n9122) );
  INV_X1 U7545 ( .A(n9422), .ZN(n7894) );
  AND2_X2 U7546 ( .A1(n7126), .A2(n7124), .ZN(n8615) );
  AND3_X1 U7547 ( .A1(n8690), .A2(n8689), .A3(n8925), .ZN(n9067) );
  AND2_X1 U7548 ( .A1(n8072), .A2(n7998), .ZN(n7923) );
  NAND2_X1 U7549 ( .A1(n8063), .A2(n7998), .ZN(n8315) );
  AND3_X1 U7550 ( .A1(n8079), .A2(n8082), .A3(n8058), .ZN(n7922) );
  AND4_X1 U7551 ( .A1(n8062), .A2(n8059), .A3(n8061), .A4(n8060), .ZN(n8063)
         );
  AND3_X1 U7552 ( .A1(n8054), .A2(n8053), .A3(n8052), .ZN(n8072) );
  AND2_X1 U7553 ( .A1(n8688), .A2(n8781), .ZN(n8689) );
  AND2_X1 U7554 ( .A1(n7834), .A2(n8251), .ZN(n7998) );
  AND2_X1 U7555 ( .A1(n8057), .A2(n8056), .ZN(n8079) );
  AND3_X1 U7556 ( .A1(n7523), .A2(n7522), .A3(n9416), .ZN(n9419) );
  AND2_X1 U7557 ( .A1(n7167), .A2(n8055), .ZN(n8082) );
  AND2_X2 U7558 ( .A1(n8686), .A2(n8687), .ZN(n8925) );
  AND3_X1 U7559 ( .A1(n9651), .A2(n6819), .A3(n6818), .ZN(n7983) );
  NOR2_X1 U7560 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n8781) );
  INV_X1 U7561 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9016) );
  INV_X1 U7562 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n9438) );
  INV_X1 U7563 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8712) );
  INV_X4 U7564 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U7565 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7522) );
  NOR2_X1 U7566 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n7523) );
  NOR2_X1 U7567 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n8686) );
  NOR2_X1 U7568 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n8687) );
  INV_X1 U7569 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9371) );
  NOR2_X1 U7570 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .ZN(
        n8052) );
  NOR2_X1 U7571 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), .ZN(
        n8053) );
  NOR2_X1 U7572 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_14__SCAN_IN), .ZN(
        n8054) );
  NOR2_X1 U7573 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n8056) );
  NOR2_X1 U7574 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_22__SCAN_IN), .ZN(
        n8057) );
  NOR2_X1 U7575 ( .A1(P3_IR_REG_23__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), .ZN(
        n7167) );
  NOR2_X1 U7576 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n8251) );
  NOR2_X1 U7577 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n7834) );
  NOR2_X1 U7578 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n8060) );
  NOR2_X1 U7579 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n8061) );
  NOR2_X1 U7580 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8059) );
  NOR2_X1 U7581 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n8062) );
  INV_X1 U7582 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8120) );
  XNOR2_X2 U7583 ( .A(n8076), .B(P3_IR_REG_21__SCAN_IN), .ZN(n8546) );
  NOR2_X2 U7584 ( .A1(n7924), .A2(n7953), .ZN(n8125) );
  AND2_X4 U7585 ( .A1(n11864), .A2(n9853), .ZN(n10450) );
  NAND3_X1 U7586 ( .A1(n7020), .A2(n10412), .A3(n7019), .ZN(n6546) );
  AND2_X2 U7587 ( .A1(n7938), .A2(n13014), .ZN(n15965) );
  OAI211_X2 U7588 ( .C1(n13787), .C2(n7077), .A(n7075), .B(n12856), .ZN(n12858) );
  OAI22_X4 U7589 ( .A1(n13800), .A2(n13797), .B1(n13361), .B2(n13812), .ZN(
        n13787) );
  AOI21_X2 U7590 ( .B1(n7207), .B2(n15963), .A(n10906), .ZN(n11406) );
  AND2_X1 U7591 ( .A1(n8128), .A2(n8127), .ZN(n8174) );
  NAND2_X1 U7592 ( .A1(n12850), .A2(n13829), .ZN(n7970) );
  NAND4_X1 U7593 ( .A1(n8681), .A2(n8710), .A3(n8712), .A4(n9918), .ZN(n8715)
         );
  NOR2_X1 U7594 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n8681) );
  XNOR2_X1 U7595 ( .A(n13958), .B(n13760), .ZN(n7852) );
  OR2_X1 U7596 ( .A1(n13344), .A2(n13388), .ZN(n13061) );
  NOR2_X1 U7597 ( .A1(n8012), .A2(n7672), .ZN(n7671) );
  AND2_X1 U7598 ( .A1(n10527), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8012) );
  INV_X1 U7599 ( .A(n8011), .ZN(n7672) );
  NAND2_X1 U7600 ( .A1(n14422), .A2(n7279), .ZN(n7277) );
  NAND2_X1 U7601 ( .A1(n14690), .A2(n7884), .ZN(n7883) );
  AND2_X1 U7602 ( .A1(n7983), .A2(n7797), .ZN(n7796) );
  AND2_X1 U7603 ( .A1(n9438), .A2(n9439), .ZN(n7797) );
  NAND2_X1 U7604 ( .A1(n15482), .A2(n15212), .ZN(n12707) );
  INV_X1 U7605 ( .A(n9331), .ZN(n7156) );
  NAND2_X1 U7606 ( .A1(n8670), .A2(n8669), .ZN(n9332) );
  NAND2_X1 U7607 ( .A1(n9314), .A2(n8668), .ZN(n8670) );
  AOI21_X1 U7608 ( .B1(n7139), .B2(n7570), .A(n7140), .ZN(n9314) );
  NOR2_X1 U7609 ( .A1(n7143), .A2(n7141), .ZN(n7140) );
  AND2_X1 U7610 ( .A1(n7572), .A2(n6761), .ZN(n7139) );
  INV_X1 U7611 ( .A(n8666), .ZN(n7141) );
  OAI21_X1 U7612 ( .B1(n8546), .B2(n13599), .A(n11492), .ZN(n7392) );
  NAND3_X1 U7613 ( .A1(n11630), .A2(n8096), .A3(n6604), .ZN(n7390) );
  INV_X1 U7614 ( .A(n12938), .ZN(n12264) );
  OR2_X1 U7615 ( .A1(n8572), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n13625) );
  OR2_X1 U7616 ( .A1(n12857), .A2(n13760), .ZN(n7994) );
  AND2_X1 U7617 ( .A1(n7961), .A2(n7960), .ZN(n7959) );
  OR2_X1 U7618 ( .A1(n13996), .A2(n13811), .ZN(n7960) );
  INV_X1 U7619 ( .A(n7967), .ZN(n7962) );
  XNOR2_X1 U7620 ( .A(n13921), .B(n13448), .ZN(n13635) );
  NAND2_X1 U7621 ( .A1(n7688), .A2(n7689), .ZN(n12947) );
  AOI21_X1 U7622 ( .B1(n7691), .B2(n12869), .A(n7690), .ZN(n7689) );
  INV_X1 U7623 ( .A(n12928), .ZN(n7690) );
  NOR2_X1 U7624 ( .A1(n14681), .A2(n10380), .ZN(n7617) );
  NOR2_X1 U7625 ( .A1(n14383), .A2(n14369), .ZN(n14359) );
  NAND2_X1 U7626 ( .A1(n14695), .A2(n14196), .ZN(n9804) );
  NOR2_X2 U7627 ( .A1(n9878), .A2(n6809), .ZN(n9441) );
  OR2_X1 U7628 ( .A1(n13221), .A2(n13220), .ZN(n13222) );
  NAND2_X1 U7629 ( .A1(n7732), .A2(n6586), .ZN(n6944) );
  OAI21_X1 U7630 ( .B1(n10345), .B2(n12412), .A(n10201), .ZN(n7476) );
  INV_X1 U7631 ( .A(n10210), .ZN(n7787) );
  NAND2_X1 U7632 ( .A1(n9090), .A2(n9134), .ZN(n7200) );
  NAND2_X1 U7633 ( .A1(n12528), .A2(n13101), .ZN(n7265) );
  INV_X1 U7634 ( .A(n7784), .ZN(n7782) );
  OAI21_X1 U7635 ( .B1(n10217), .B2(n10216), .A(n10215), .ZN(n10218) );
  NAND2_X1 U7636 ( .A1(n6675), .A2(n7784), .ZN(n7779) );
  OAI21_X1 U7637 ( .B1(n7564), .B2(n7563), .A(n7561), .ZN(n10246) );
  AND2_X1 U7638 ( .A1(n13116), .A2(n13683), .ZN(n7267) );
  CLKBUF_X1 U7639 ( .A(n10194), .Z(n10345) );
  INV_X1 U7640 ( .A(n9266), .ZN(n7614) );
  NAND2_X1 U7641 ( .A1(n13125), .A2(n13124), .ZN(n6956) );
  NAND2_X1 U7642 ( .A1(n6958), .A2(n13126), .ZN(n6957) );
  OR2_X1 U7643 ( .A1(n12959), .A2(n13624), .ZN(n13134) );
  NOR2_X1 U7644 ( .A1(n6896), .A2(n7708), .ZN(n6895) );
  AND2_X1 U7645 ( .A1(n13782), .A2(n13759), .ZN(n12889) );
  AND2_X1 U7646 ( .A1(n13974), .A2(n13773), .ZN(n13751) );
  OR2_X1 U7647 ( .A1(n13817), .A2(n13831), .ZN(n13074) );
  NOR2_X1 U7648 ( .A1(n10353), .A2(n7218), .ZN(n10399) );
  AND2_X1 U7649 ( .A1(n10367), .A2(n14193), .ZN(n7218) );
  NAND2_X1 U7650 ( .A1(n9248), .A2(n9247), .ZN(n9267) );
  OR2_X1 U7651 ( .A1(n9244), .A2(n9243), .ZN(n9248) );
  AND2_X1 U7652 ( .A1(n12011), .A2(n12006), .ZN(n12007) );
  OR2_X1 U7653 ( .A1(n15821), .A2(n14840), .ZN(n12006) );
  NOR2_X1 U7654 ( .A1(n8661), .A2(n11615), .ZN(n8662) );
  NAND2_X1 U7655 ( .A1(n7554), .A2(n7552), .ZN(n8657) );
  AND2_X1 U7656 ( .A1(n7553), .A2(n8656), .ZN(n7552) );
  AND2_X1 U7657 ( .A1(n8655), .A2(n9208), .ZN(n8656) );
  NAND2_X1 U7658 ( .A1(n8988), .A2(n10578), .ZN(n8769) );
  NAND2_X1 U7659 ( .A1(n8790), .A2(n7120), .ZN(n8806) );
  NOR2_X1 U7660 ( .A1(n8787), .A2(n7121), .ZN(n7120) );
  INV_X1 U7661 ( .A(n8617), .ZN(n7121) );
  INV_X1 U7662 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10536) );
  XNOR2_X1 U7663 ( .A(n13874), .B(n12911), .ZN(n8458) );
  NAND2_X1 U7664 ( .A1(n7376), .A2(n8487), .ZN(n7375) );
  NAND2_X1 U7665 ( .A1(n12970), .A2(n6581), .ZN(n7183) );
  NAND2_X1 U7666 ( .A1(n11255), .A2(n11233), .ZN(n11234) );
  INV_X1 U7667 ( .A(n6893), .ZN(n6890) );
  INV_X1 U7668 ( .A(n13491), .ZN(n13489) );
  NAND2_X1 U7669 ( .A1(n8115), .A2(n8114), .ZN(n8507) );
  INV_X1 U7670 ( .A(n8491), .ZN(n8115) );
  AND2_X1 U7671 ( .A1(n6743), .A2(n7326), .ZN(n7325) );
  INV_X1 U7672 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n7326) );
  NOR2_X1 U7673 ( .A1(n13635), .A2(n13636), .ZN(n12868) );
  NOR2_X1 U7674 ( .A1(n13751), .A2(n12889), .ZN(n7168) );
  INV_X1 U7675 ( .A(n13785), .ZN(n6919) );
  OR2_X1 U7676 ( .A1(n13964), .A2(n13772), .ZN(n13092) );
  INV_X1 U7677 ( .A(n13831), .ZN(n7969) );
  AND2_X1 U7678 ( .A1(n9469), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n9784) );
  NAND2_X1 U7679 ( .A1(n7131), .A2(n7129), .ZN(n10368) );
  AND2_X1 U7680 ( .A1(n7130), .A2(n10320), .ZN(n7129) );
  INV_X1 U7681 ( .A(n14193), .ZN(n7130) );
  INV_X1 U7682 ( .A(n11041), .ZN(n7305) );
  OR3_X1 U7683 ( .A1(n9808), .A2(n12820), .A3(n9807), .ZN(n9858) );
  AOI21_X1 U7684 ( .B1(n7279), .B2(n6560), .A(n6706), .ZN(n7278) );
  NAND2_X1 U7685 ( .A1(n14540), .A2(n7414), .ZN(n7413) );
  INV_X1 U7686 ( .A(n8003), .ZN(n7414) );
  OR2_X1 U7687 ( .A1(n14737), .A2(n14563), .ZN(n14505) );
  NOR2_X1 U7688 ( .A1(n14592), .A2(n7888), .ZN(n7887) );
  INV_X1 U7689 ( .A(n9830), .ZN(n7888) );
  OR2_X1 U7690 ( .A1(n12232), .A2(n7532), .ZN(n14622) );
  NAND2_X1 U7691 ( .A1(n7534), .A2(n7533), .ZN(n7532) );
  INV_X1 U7692 ( .A(n9648), .ZN(n7534) );
  NOR2_X2 U7693 ( .A1(n12277), .A2(n12468), .ZN(n12241) );
  NAND2_X1 U7694 ( .A1(n9821), .A2(n7898), .ZN(n12324) );
  NAND2_X1 U7695 ( .A1(n11973), .A2(n9818), .ZN(n12126) );
  NAND2_X1 U7696 ( .A1(n9484), .A2(n6642), .ZN(n9512) );
  NAND4_X1 U7697 ( .A1(n7893), .A2(n7894), .A3(n9441), .A4(n7535), .ZN(n9459)
         );
  NOR2_X1 U7698 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n7535) );
  NOR2_X1 U7699 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n9421) );
  NOR2_X1 U7700 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n9420) );
  AND2_X1 U7701 ( .A1(n11892), .A2(n6633), .ZN(n6937) );
  INV_X1 U7702 ( .A(n7725), .ZN(n6949) );
  NAND2_X1 U7703 ( .A1(n6789), .A2(n6787), .ZN(n7641) );
  AOI21_X1 U7704 ( .B1(n7981), .B2(n7005), .A(n6698), .ZN(n6789) );
  NAND2_X1 U7705 ( .A1(n7981), .A2(n6788), .ZN(n6787) );
  INV_X1 U7706 ( .A(n12711), .ZN(n7007) );
  NAND2_X1 U7707 ( .A1(n15543), .A2(n15412), .ZN(n12717) );
  INV_X1 U7708 ( .A(n12697), .ZN(n7804) );
  NAND2_X1 U7709 ( .A1(n12010), .A2(n7656), .ZN(n7658) );
  NOR2_X1 U7710 ( .A1(n12011), .A2(n7657), .ZN(n7656) );
  INV_X1 U7711 ( .A(n12009), .ZN(n7657) );
  NAND2_X1 U7712 ( .A1(n15231), .A2(n7826), .ZN(n15196) );
  NOR2_X1 U7713 ( .A1(n15462), .A2(n7828), .ZN(n7826) );
  XNOR2_X1 U7714 ( .A(n8671), .B(SI_28_), .ZN(n9331) );
  NAND2_X1 U7715 ( .A1(n7142), .A2(n7570), .ZN(n7144) );
  NOR2_X2 U7716 ( .A1(n8715), .A2(n8682), .ZN(n8717) );
  NOR2_X1 U7717 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n8683) );
  NOR2_X1 U7718 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n8684) );
  NAND2_X1 U7719 ( .A1(n8622), .A2(SI_9_), .ZN(n8624) );
  NAND2_X1 U7720 ( .A1(n10559), .A2(n10558), .ZN(n10561) );
  AND2_X1 U7721 ( .A1(n13464), .A2(n12677), .ZN(n10904) );
  NAND2_X1 U7722 ( .A1(n12226), .A2(n6551), .ZN(n12945) );
  INV_X1 U7723 ( .A(n13625), .ZN(n12226) );
  NAND2_X1 U7724 ( .A1(n7701), .A2(n7700), .ZN(n11326) );
  AOI21_X1 U7725 ( .B1(n7707), .B2(n7705), .A(n6693), .ZN(n7700) );
  NAND2_X1 U7726 ( .A1(n11218), .A2(n7704), .ZN(n7701) );
  NAND2_X1 U7727 ( .A1(n7350), .A2(n7349), .ZN(n13514) );
  NOR2_X1 U7728 ( .A1(n13500), .A2(n13501), .ZN(n7349) );
  OAI21_X1 U7729 ( .B1(n13471), .B2(n7081), .A(n7080), .ZN(n13526) );
  AOI21_X1 U7730 ( .B1(n13492), .B2(n7581), .A(n13499), .ZN(n7080) );
  AND2_X1 U7731 ( .A1(n13526), .A2(n13525), .ZN(n13527) );
  NAND2_X1 U7732 ( .A1(n6708), .A2(n6573), .ZN(n7072) );
  NOR2_X1 U7733 ( .A1(n7864), .A2(n13118), .ZN(n7863) );
  INV_X1 U7734 ( .A(n7866), .ZN(n7864) );
  OR2_X1 U7735 ( .A1(n8435), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8451) );
  INV_X1 U7736 ( .A(n13452), .ZN(n13811) );
  INV_X1 U7737 ( .A(n7842), .ZN(n7841) );
  AND2_X1 U7738 ( .A1(n12970), .A2(n12954), .ZN(n12926) );
  XNOR2_X1 U7739 ( .A(n13927), .B(n13666), .ZN(n13649) );
  NOR2_X1 U7740 ( .A1(n6684), .A2(n7951), .ZN(n7950) );
  INV_X1 U7741 ( .A(n7994), .ZN(n7951) );
  NAND2_X1 U7742 ( .A1(n12853), .A2(n7076), .ZN(n7075) );
  NAND2_X1 U7743 ( .A1(n12853), .A2(n7079), .ZN(n7077) );
  NOR2_X1 U7744 ( .A1(n12888), .A2(n7861), .ZN(n7860) );
  INV_X1 U7745 ( .A(n12886), .ZN(n7861) );
  OR2_X1 U7746 ( .A1(n13996), .A2(n13452), .ZN(n7862) );
  NAND2_X1 U7747 ( .A1(n7966), .A2(n7970), .ZN(n7965) );
  INV_X1 U7748 ( .A(n7968), .ZN(n7966) );
  AOI21_X1 U7749 ( .B1(n12983), .B2(n6552), .A(n6671), .ZN(n7968) );
  XNOR2_X1 U7750 ( .A(n13996), .B(n13811), .ZN(n13826) );
  OR2_X1 U7751 ( .A1(n13124), .A2(n10909), .ZN(n15990) );
  OR2_X1 U7752 ( .A1(n13124), .A2(n8569), .ZN(n15992) );
  NAND2_X1 U7753 ( .A1(n6764), .A2(n11389), .ZN(n13833) );
  NAND2_X1 U7754 ( .A1(n12947), .A2(n12946), .ZN(n12949) );
  NAND2_X1 U7755 ( .A1(n12829), .A2(n12828), .ZN(n12870) );
  OR2_X1 U7756 ( .A1(n12827), .A2(n12826), .ZN(n12829) );
  OAI21_X1 U7757 ( .B1(n8502), .B2(n7696), .A(n7694), .ZN(n12827) );
  INV_X1 U7758 ( .A(n7697), .ZN(n7696) );
  AOI21_X1 U7759 ( .B1(n7697), .B2(n7695), .A(n6773), .ZN(n7694) );
  AOI21_X1 U7760 ( .B1(n8501), .B2(n8050), .A(n6772), .ZN(n7697) );
  OAI21_X1 U7761 ( .B1(n8035), .B2(n7001), .A(n6998), .ZN(n8477) );
  INV_X1 U7762 ( .A(n7002), .ZN(n7001) );
  AND2_X1 U7763 ( .A1(n7684), .A2(n6999), .ZN(n6998) );
  NAND2_X1 U7764 ( .A1(n7002), .A2(n7000), .ZN(n6999) );
  NAND2_X1 U7765 ( .A1(n8041), .A2(n6740), .ZN(n8464) );
  NAND2_X1 U7766 ( .A1(n8547), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8076) );
  NAND2_X1 U7767 ( .A1(n6966), .A2(n6968), .ZN(n6964) );
  NAND2_X1 U7768 ( .A1(n8014), .A2(n8013), .ZN(n8249) );
  NAND2_X1 U7769 ( .A1(n7667), .A2(n7665), .ZN(n8014) );
  AOI21_X1 U7770 ( .B1(n7668), .B2(n7670), .A(n7666), .ZN(n7665) );
  XNOR2_X1 U7771 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n8233) );
  XNOR2_X1 U7772 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8200) );
  AOI21_X1 U7773 ( .B1(n12815), .B2(n12814), .A(n14049), .ZN(n12816) );
  NAND2_X1 U7774 ( .A1(n7018), .A2(n11861), .ZN(n7020) );
  AND2_X1 U7775 ( .A1(n7538), .A2(n7031), .ZN(n7030) );
  AOI21_X1 U7776 ( .B1(n6599), .B2(n7541), .A(n7539), .ZN(n7538) );
  NAND2_X1 U7777 ( .A1(n6599), .A2(n7032), .ZN(n7031) );
  INV_X1 U7778 ( .A(n14055), .ZN(n7539) );
  INV_X1 U7779 ( .A(n6599), .ZN(n7033) );
  OR3_X1 U7780 ( .A1(n12225), .A2(n12484), .A3(n12478), .ZN(n11021) );
  NAND2_X1 U7781 ( .A1(n7882), .A2(n7883), .ZN(n9857) );
  AOI21_X1 U7782 ( .B1(n14391), .B2(n14392), .A(n7284), .ZN(n14377) );
  OR2_X1 U7783 ( .A1(n14457), .A2(n14199), .ZN(n7988) );
  NAND2_X1 U7784 ( .A1(n9867), .A2(n7626), .ZN(n14581) );
  AND3_X1 U7785 ( .A1(n14605), .A2(n7627), .A3(n7628), .ZN(n7626) );
  NAND2_X1 U7786 ( .A1(n6707), .A2(n6796), .ZN(n9831) );
  NAND2_X1 U7787 ( .A1(n12502), .A2(n7287), .ZN(n6796) );
  XNOR2_X1 U7788 ( .A(n14759), .B(n14637), .ZN(n14625) );
  INV_X1 U7789 ( .A(n7288), .ZN(n7287) );
  OAI21_X1 U7790 ( .B1(n7289), .B2(n9825), .A(n7899), .ZN(n7288) );
  AOI21_X1 U7791 ( .B1(n7901), .B2(n9826), .A(n7900), .ZN(n7899) );
  INV_X1 U7792 ( .A(n9828), .ZN(n7900) );
  NAND2_X1 U7793 ( .A1(n6843), .A2(n7292), .ZN(n12501) );
  NOR2_X1 U7794 ( .A1(n7982), .A2(n6844), .ZN(n6843) );
  NAND2_X1 U7795 ( .A1(n7290), .A2(n9824), .ZN(n6844) );
  XNOR2_X1 U7796 ( .A(n12104), .B(n12407), .ZN(n6842) );
  NAND2_X1 U7797 ( .A1(n14369), .A2(n14355), .ZN(n14344) );
  NAND2_X1 U7798 ( .A1(n7101), .A2(n7407), .ZN(n9815) );
  AOI21_X1 U7799 ( .B1(n7408), .B2(n7410), .A(n6705), .ZN(n7407) );
  NAND2_X1 U7800 ( .A1(n14404), .A2(n7408), .ZN(n7101) );
  AND2_X1 U7801 ( .A1(n10398), .A2(n7883), .ZN(n7881) );
  OR2_X1 U7802 ( .A1(n9815), .A2(n9856), .ZN(n7412) );
  OR2_X1 U7803 ( .A1(n10482), .A2(n10485), .ZN(n15931) );
  AND2_X1 U7804 ( .A1(n9484), .A2(n11007), .ZN(n9487) );
  XNOR2_X1 U7805 ( .A(n9458), .B(P2_IR_REG_30__SCAN_IN), .ZN(n7109) );
  NAND2_X1 U7806 ( .A1(n9459), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9460) );
  AND2_X1 U7807 ( .A1(n13187), .A2(n13188), .ZN(n7727) );
  XNOR2_X1 U7808 ( .A(n13218), .B(n11908), .ZN(n13221) );
  NAND2_X1 U7809 ( .A1(n6944), .A2(n6680), .ZN(n6942) );
  NOR2_X1 U7810 ( .A1(n7730), .A2(n6946), .ZN(n6945) );
  INV_X1 U7811 ( .A(n12634), .ZN(n6946) );
  NAND2_X1 U7812 ( .A1(n7732), .A2(n7731), .ZN(n7730) );
  NAND2_X1 U7813 ( .A1(n9082), .A2(n9081), .ZN(n14965) );
  INV_X2 U7814 ( .A(n8863), .ZN(n9324) );
  INV_X1 U7815 ( .A(n13276), .ZN(n7008) );
  OR2_X1 U7816 ( .A1(n7490), .A2(n7489), .ZN(n15080) );
  INV_X1 U7817 ( .A(n15068), .ZN(n7489) );
  NAND2_X1 U7818 ( .A1(n15080), .A2(n7488), .ZN(n15082) );
  OR2_X1 U7819 ( .A1(n15081), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7488) );
  NOR2_X1 U7820 ( .A1(n15196), .A2(n15175), .ZN(n15174) );
  NAND2_X1 U7821 ( .A1(n15242), .A2(n12732), .ZN(n15236) );
  OR2_X1 U7822 ( .A1(n15482), .A2(n15212), .ZN(n9394) );
  AOI21_X1 U7823 ( .B1(n7807), .B2(n7811), .A(n6691), .ZN(n7805) );
  INV_X1 U7824 ( .A(n12705), .ZN(n7811) );
  NAND2_X1 U7825 ( .A1(n7443), .A2(n12701), .ZN(n7442) );
  NAND2_X1 U7826 ( .A1(n15329), .A2(n7444), .ZN(n7443) );
  NOR2_X1 U7827 ( .A1(n15330), .A2(n15329), .ZN(n7448) );
  INV_X2 U7828 ( .A(n8898), .ZN(n9155) );
  NAND2_X1 U7829 ( .A1(n15473), .A2(n6654), .ZN(n15201) );
  XNOR2_X1 U7830 ( .A(n8727), .B(n8726), .ZN(n13275) );
  NAND2_X1 U7831 ( .A1(n7149), .A2(n7152), .ZN(n8727) );
  NAND2_X1 U7832 ( .A1(n7157), .A2(n7150), .ZN(n7149) );
  XNOR2_X1 U7833 ( .A(n9314), .B(n9313), .ZN(n12908) );
  NAND2_X1 U7834 ( .A1(n10830), .A2(n10829), .ZN(n10841) );
  OR2_X1 U7835 ( .A1(n11323), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7767) );
  NAND2_X1 U7836 ( .A1(n7041), .A2(n7498), .ZN(n7766) );
  NOR2_X1 U7837 ( .A1(n7501), .A2(n6579), .ZN(n7498) );
  NAND2_X1 U7838 ( .A1(n7762), .A2(n15623), .ZN(n15632) );
  NAND2_X1 U7839 ( .A1(n7509), .A2(n10129), .ZN(n7508) );
  NAND2_X1 U7840 ( .A1(n8578), .A2(n8577), .ZN(n13448) );
  NAND2_X1 U7841 ( .A1(n6683), .A2(n7618), .ZN(n14343) );
  OR2_X1 U7842 ( .A1(n11858), .A2(n11857), .ZN(n11859) );
  NAND2_X1 U7843 ( .A1(n15620), .A2(n15621), .ZN(n7762) );
  NAND2_X1 U7844 ( .A1(n15632), .A2(n15631), .ZN(n7512) );
  NAND2_X1 U7845 ( .A1(n8933), .A2(n8868), .ZN(n7242) );
  NAND2_X1 U7846 ( .A1(n15980), .A2(n11630), .ZN(n7210) );
  NAND2_X1 U7847 ( .A1(n6802), .A2(n10232), .ZN(n10192) );
  AOI21_X1 U7848 ( .B1(n10194), .B2(n6802), .A(n6798), .ZN(n10195) );
  NOR2_X1 U7849 ( .A1(n12104), .A2(n10194), .ZN(n6798) );
  NAND2_X1 U7850 ( .A1(n10179), .A2(n10180), .ZN(n10188) );
  MUX2_X1 U7851 ( .A(n11955), .B(n11761), .S(n9076), .Z(n8963) );
  INV_X1 U7852 ( .A(n9005), .ZN(n7605) );
  MUX2_X1 U7853 ( .A(n15828), .B(n12170), .S(n9344), .Z(n9005) );
  OAI21_X1 U7854 ( .B1(n7476), .B2(n7475), .A(n6695), .ZN(n7474) );
  NAND2_X1 U7855 ( .A1(n7476), .A2(n7475), .ZN(n7471) );
  NAND2_X1 U7856 ( .A1(n7772), .A2(n7771), .ZN(n7770) );
  OR2_X1 U7857 ( .A1(n7605), .A2(n7601), .ZN(n7600) );
  NAND2_X1 U7858 ( .A1(n7478), .A2(n7477), .ZN(n10213) );
  AOI21_X1 U7859 ( .B1(n7479), .B2(n7481), .A(n6689), .ZN(n7477) );
  AND2_X1 U7860 ( .A1(n10207), .A2(n10209), .ZN(n7481) );
  INV_X1 U7861 ( .A(n7595), .ZN(n7594) );
  OAI21_X1 U7862 ( .B1(n9142), .B2(n9141), .A(n9139), .ZN(n7595) );
  INV_X1 U7863 ( .A(n7200), .ZN(n9139) );
  OAI211_X1 U7864 ( .C1(n7200), .C2(n9137), .A(n9136), .B(n9135), .ZN(n9138)
         );
  NAND2_X1 U7865 ( .A1(n10224), .A2(n10223), .ZN(n6833) );
  INV_X1 U7866 ( .A(n7783), .ZN(n7778) );
  NOR2_X1 U7867 ( .A1(n7783), .A2(n10223), .ZN(n7780) );
  NAND2_X1 U7868 ( .A1(n6997), .A2(n9214), .ZN(n6996) );
  NAND2_X1 U7869 ( .A1(n10288), .A2(n10289), .ZN(n10293) );
  NAND2_X1 U7870 ( .A1(n10237), .A2(n7468), .ZN(n7463) );
  INV_X1 U7871 ( .A(n7463), .ZN(n7459) );
  AND2_X1 U7872 ( .A1(n10307), .A2(n10308), .ZN(n7566) );
  AND2_X1 U7873 ( .A1(n7465), .A2(n7462), .ZN(n7461) );
  NAND2_X1 U7874 ( .A1(n7467), .A2(n7466), .ZN(n7465) );
  NAND2_X1 U7875 ( .A1(n7464), .A2(n7463), .ZN(n7462) );
  NOR2_X1 U7876 ( .A1(n10237), .A2(n7468), .ZN(n7464) );
  NAND2_X1 U7877 ( .A1(n6824), .A2(n6822), .ZN(n10235) );
  NAND2_X1 U7878 ( .A1(n6823), .A2(n10230), .ZN(n6822) );
  OR2_X1 U7879 ( .A1(n7470), .A2(n6589), .ZN(n6824) );
  INV_X1 U7880 ( .A(n10231), .ZN(n6823) );
  AND2_X1 U7881 ( .A1(n15749), .A2(n8869), .ZN(n8868) );
  NOR2_X1 U7882 ( .A1(n6558), .A2(n8647), .ZN(n7559) );
  INV_X1 U7883 ( .A(n13517), .ZN(n6896) );
  INV_X1 U7884 ( .A(n8029), .ZN(n7664) );
  OR2_X1 U7885 ( .A1(n7614), .A2(n9268), .ZN(n7613) );
  INV_X1 U7886 ( .A(n12712), .ZN(n6788) );
  NAND2_X1 U7887 ( .A1(n6620), .A2(n11712), .ZN(n7632) );
  INV_X1 U7888 ( .A(n7137), .ZN(n7136) );
  OAI21_X1 U7889 ( .B1(n8634), .B2(n7138), .A(n6687), .ZN(n7137) );
  OAI21_X1 U7890 ( .B1(n6542), .B2(n7199), .A(n7198), .ZN(n8630) );
  NAND2_X1 U7891 ( .A1(n7195), .A2(n6644), .ZN(n8628) );
  INV_X1 U7892 ( .A(n9014), .ZN(n7195) );
  NOR2_X1 U7893 ( .A1(n8458), .A2(n13744), .ZN(n8459) );
  NOR2_X1 U7894 ( .A1(n13377), .A2(n7916), .ZN(n7915) );
  INV_X1 U7895 ( .A(n8432), .ZN(n7916) );
  AOI21_X1 U7896 ( .B1(n8298), .B2(n7388), .A(n6646), .ZN(n7387) );
  INV_X1 U7897 ( .A(n12194), .ZN(n7388) );
  INV_X1 U7898 ( .A(n8373), .ZN(n7928) );
  OR2_X1 U7899 ( .A1(n13927), .A2(n13639), .ZN(n7268) );
  NOR2_X1 U7900 ( .A1(n13135), .A2(n13136), .ZN(n6994) );
  INV_X1 U7901 ( .A(n11492), .ZN(n10908) );
  AND2_X1 U7902 ( .A1(n12926), .A2(n7846), .ZN(n7845) );
  OR2_X1 U7903 ( .A1(n13635), .A2(n7847), .ZN(n7846) );
  NAND2_X1 U7904 ( .A1(n7845), .A2(n7847), .ZN(n7843) );
  NAND2_X1 U7905 ( .A1(n7059), .A2(n7058), .ZN(n7336) );
  NOR2_X1 U7906 ( .A1(n6676), .A2(n7060), .ZN(n7059) );
  NOR2_X1 U7907 ( .A1(n7332), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7331) );
  NAND2_X1 U7908 ( .A1(n11262), .A2(n11145), .ZN(n11186) );
  INV_X1 U7909 ( .A(n7372), .ZN(n7369) );
  AND2_X1 U7910 ( .A1(n11205), .A2(n7371), .ZN(n7370) );
  NAND2_X1 U7911 ( .A1(n11295), .A2(n11199), .ZN(n7371) );
  INV_X1 U7912 ( .A(n11229), .ZN(n7358) );
  INV_X1 U7913 ( .A(n6739), .ZN(n7343) );
  NAND2_X1 U7914 ( .A1(n7347), .A2(n7345), .ZN(n7344) );
  INV_X1 U7915 ( .A(n13564), .ZN(n7345) );
  NAND2_X1 U7916 ( .A1(n7074), .A2(n7072), .ZN(n7070) );
  INV_X1 U7917 ( .A(n7072), .ZN(n7071) );
  AND2_X1 U7918 ( .A1(n8110), .A2(n7322), .ZN(n7321) );
  INV_X1 U7919 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n7322) );
  INV_X1 U7920 ( .A(n8394), .ZN(n8111) );
  AND2_X1 U7921 ( .A1(n8108), .A2(n7319), .ZN(n7318) );
  INV_X1 U7922 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n7319) );
  INV_X1 U7923 ( .A(n13826), .ZN(n7964) );
  INV_X1 U7924 ( .A(n8333), .ZN(n8109) );
  INV_X1 U7925 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n7327) );
  INV_X1 U7926 ( .A(n8273), .ZN(n8106) );
  OR2_X1 U7927 ( .A1(n7959), .A2(n12984), .ZN(n7956) );
  INV_X1 U7928 ( .A(n7862), .ZN(n7859) );
  INV_X1 U7929 ( .A(n13074), .ZN(n7855) );
  NAND2_X1 U7930 ( .A1(n7857), .A2(n12884), .ZN(n6916) );
  NAND2_X1 U7931 ( .A1(n6934), .A2(n7944), .ZN(n6933) );
  INV_X1 U7932 ( .A(n6935), .ZN(n6934) );
  INV_X1 U7933 ( .A(n8461), .ZN(n7687) );
  INV_X1 U7934 ( .A(n8200), .ZN(n6975) );
  AOI21_X1 U7935 ( .B1(n6974), .B2(n8200), .A(n6701), .ZN(n6973) );
  INV_X1 U7936 ( .A(n8007), .ZN(n6974) );
  INV_X1 U7937 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n8009) );
  INV_X1 U7938 ( .A(n10465), .ZN(n7039) );
  NOR2_X1 U7939 ( .A1(n9774), .A2(n14098), .ZN(n9469) );
  NAND2_X1 U7940 ( .A1(n7037), .A2(n7039), .ZN(n7036) );
  INV_X1 U7941 ( .A(n7038), .ZN(n7037) );
  OAI21_X1 U7942 ( .B1(n6610), .B2(n7039), .A(n14142), .ZN(n7038) );
  INV_X1 U7943 ( .A(n12759), .ZN(n7544) );
  INV_X1 U7944 ( .A(n7546), .ZN(n7545) );
  OAI21_X1 U7945 ( .B1(n14141), .B2(n7547), .A(n14063), .ZN(n7546) );
  INV_X1 U7946 ( .A(n14062), .ZN(n7547) );
  INV_X1 U7947 ( .A(n9721), .ZN(n9451) );
  INV_X1 U7948 ( .A(n14625), .ZN(n6810) );
  NOR2_X1 U7949 ( .A1(n6817), .A2(n10399), .ZN(n6816) );
  NAND2_X1 U7950 ( .A1(n10398), .A2(n10396), .ZN(n6817) );
  NAND2_X1 U7951 ( .A1(n10341), .A2(n10362), .ZN(n7255) );
  OR2_X1 U7952 ( .A1(n10399), .A2(n10361), .ZN(n7253) );
  NOR2_X1 U7953 ( .A1(n7624), .A2(n14491), .ZN(n7623) );
  INV_X1 U7954 ( .A(n7625), .ZN(n7624) );
  INV_X1 U7955 ( .A(n7629), .ZN(n7628) );
  NAND2_X1 U7956 ( .A1(n14620), .A2(n14816), .ZN(n7629) );
  NOR2_X1 U7957 ( .A1(n9433), .A2(n11861), .ZN(n7021) );
  NAND2_X1 U7958 ( .A1(n15583), .A2(n10335), .ZN(n7131) );
  NAND2_X1 U7959 ( .A1(n14436), .A2(n7621), .ZN(n14383) );
  AND2_X1 U7960 ( .A1(n6572), .A2(n7622), .ZN(n7621) );
  NAND4_X1 U7961 ( .A1(n9439), .A2(n9440), .A3(n9438), .A4(n9437), .ZN(n6809)
         );
  NAND2_X1 U7962 ( .A1(n9444), .A2(n9459), .ZN(n9478) );
  NAND2_X1 U7963 ( .A1(n6805), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9443) );
  INV_X1 U7964 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9882) );
  OAI21_X1 U7965 ( .B1(n9871), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9883) );
  NOR2_X1 U7966 ( .A1(n7550), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n7549) );
  NAND2_X1 U7967 ( .A1(n9426), .A2(n7551), .ZN(n7550) );
  INV_X1 U7968 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n7551) );
  INV_X1 U7969 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6819) );
  OR2_X1 U7970 ( .A1(n12572), .A2(n7980), .ZN(n12441) );
  OAI22_X1 U7971 ( .A1(n11541), .A2(n13195), .B1(n11498), .B2(n13224), .ZN(
        n10992) );
  INV_X1 U7972 ( .A(n14937), .ZN(n7724) );
  NAND2_X1 U7973 ( .A1(n14966), .A2(n6649), .ZN(n6948) );
  INV_X1 U7974 ( .A(n6952), .ZN(n6951) );
  INV_X1 U7975 ( .A(n9336), .ZN(n7598) );
  INV_X1 U7976 ( .A(n15222), .ZN(n13225) );
  AND2_X1 U7977 ( .A1(n7805), .A2(n7435), .ZN(n7434) );
  INV_X1 U7978 ( .A(n15235), .ZN(n7435) );
  NAND2_X1 U7979 ( .A1(n12705), .A2(n7810), .ZN(n7809) );
  INV_X1 U7980 ( .A(n12704), .ZN(n7810) );
  AOI21_X1 U7981 ( .B1(n7647), .B2(n6571), .A(n15245), .ZN(n7646) );
  INV_X1 U7982 ( .A(n7647), .ZN(n7644) );
  AND2_X1 U7983 ( .A1(n7648), .A2(n7650), .ZN(n7647) );
  INV_X1 U7984 ( .A(n15259), .ZN(n7648) );
  OR2_X1 U7985 ( .A1(n15289), .A2(n7444), .ZN(n7440) );
  NAND2_X1 U7986 ( .A1(n15337), .A2(n15336), .ZN(n12721) );
  NOR2_X1 U7987 ( .A1(n6908), .A2(n12001), .ZN(n6907) );
  NAND2_X1 U7988 ( .A1(n12007), .A2(n6663), .ZN(n7423) );
  NAND2_X1 U7989 ( .A1(n11525), .A2(n15018), .ZN(n11520) );
  INV_X1 U7990 ( .A(n15425), .ZN(n11498) );
  AND3_X1 U7991 ( .A1(n8861), .A2(n8860), .A3(n8859), .ZN(n11501) );
  OAI21_X1 U7992 ( .B1(n10676), .B2(n15150), .A(n8856), .ZN(n8860) );
  NAND2_X1 U7993 ( .A1(n10642), .A2(n8854), .ZN(n8861) );
  AOI21_X1 U7994 ( .B1(n12737), .B2(n12738), .A(n12739), .ZN(n7636) );
  AND2_X1 U7995 ( .A1(n8722), .A2(n10788), .ZN(n10807) );
  INV_X1 U7996 ( .A(n7570), .ZN(n7569) );
  INV_X1 U7997 ( .A(n8663), .ZN(n7164) );
  NAND2_X1 U7998 ( .A1(n7231), .A2(n7230), .ZN(n7132) );
  INV_X1 U7999 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8705) );
  NAND2_X1 U8000 ( .A1(n8690), .A2(n8925), .ZN(n6987) );
  NAND2_X1 U8001 ( .A1(n9038), .A2(n8635), .ZN(n9115) );
  AOI21_X1 U8002 ( .B1(n8628), .B2(n8772), .A(n8627), .ZN(n8629) );
  AOI21_X1 U8003 ( .B1(n8806), .B2(n7119), .A(n6617), .ZN(n7416) );
  XNOR2_X1 U8004 ( .A(n8630), .B(SI_12_), .ZN(n8627) );
  INV_X1 U8005 ( .A(n8628), .ZN(n8770) );
  NAND2_X1 U8006 ( .A1(n7748), .A2(n7746), .ZN(n7745) );
  INV_X1 U8007 ( .A(n7747), .ZN(n7746) );
  INV_X1 U8008 ( .A(n8609), .ZN(n7735) );
  AND2_X1 U8009 ( .A1(n8925), .A2(n8775), .ZN(n8926) );
  NAND2_X1 U8010 ( .A1(n7219), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7997) );
  XNOR2_X1 U8011 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n7040) );
  AND2_X1 U8012 ( .A1(n7503), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n10555) );
  INV_X1 U8013 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7503) );
  AND2_X1 U8014 ( .A1(n10539), .A2(n10538), .ZN(n10558) );
  XNOR2_X1 U8015 ( .A(n10814), .B(n11194), .ZN(n10545) );
  INV_X1 U8016 ( .A(n7915), .ZN(n7914) );
  AOI21_X1 U8017 ( .B1(n7915), .B2(n7913), .A(n6748), .ZN(n7912) );
  INV_X1 U8018 ( .A(n13310), .ZN(n7913) );
  AND2_X1 U8019 ( .A1(n10925), .A2(n10926), .ZN(n8196) );
  NAND2_X1 U8020 ( .A1(n7403), .A2(n8199), .ZN(n7909) );
  INV_X1 U8021 ( .A(n11104), .ZN(n7403) );
  NAND2_X1 U8022 ( .A1(n10154), .A2(n13731), .ZN(n7918) );
  AND2_X1 U8023 ( .A1(n7398), .A2(n7925), .ZN(n7397) );
  NAND2_X1 U8024 ( .A1(n7926), .A2(n7399), .ZN(n7398) );
  AOI21_X1 U8025 ( .B1(n7926), .B2(n7928), .A(n6694), .ZN(n7925) );
  INV_X1 U8026 ( .A(n7400), .ZN(n7399) );
  INV_X1 U8027 ( .A(n13366), .ZN(n7395) );
  AND4_X1 U8028 ( .A1(n8324), .A2(n8323), .A3(n8322), .A4(n8321), .ZN(n13388)
         );
  AND4_X2 U8029 ( .A1(n8214), .A2(n8213), .A3(n8212), .A4(n8211), .ZN(n11408)
         );
  OR2_X1 U8030 ( .A1(n6545), .A2(n8210), .ZN(n8211) );
  NAND2_X1 U8031 ( .A1(n8151), .A2(n6583), .ZN(n7574) );
  NAND2_X1 U8032 ( .A1(n7574), .A2(n7573), .ZN(n11177) );
  AND2_X1 U8033 ( .A1(n11151), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7573) );
  NAND2_X1 U8034 ( .A1(n11281), .A2(n6660), .ZN(n11216) );
  NAND2_X1 U8035 ( .A1(n7092), .A2(n11201), .ZN(n11192) );
  INV_X1 U8036 ( .A(n11191), .ZN(n7092) );
  NAND2_X1 U8037 ( .A1(n7364), .A2(n7374), .ZN(n7363) );
  INV_X1 U8038 ( .A(n7367), .ZN(n7364) );
  AOI21_X1 U8039 ( .B1(n7370), .B2(n7369), .A(n7368), .ZN(n7367) );
  INV_X1 U8040 ( .A(n11247), .ZN(n7368) );
  INV_X1 U8041 ( .A(n11245), .ZN(n7705) );
  AOI21_X1 U8042 ( .B1(n11337), .B2(n7586), .A(n6779), .ZN(n7584) );
  NAND2_X1 U8043 ( .A1(n6899), .A2(n6897), .ZN(n11557) );
  NAND2_X1 U8044 ( .A1(n11328), .A2(n6648), .ZN(n6899) );
  OAI21_X1 U8045 ( .B1(n6901), .B2(n11465), .A(n6744), .ZN(n6898) );
  AND2_X1 U8046 ( .A1(n11873), .A2(n12141), .ZN(n11874) );
  NAND2_X1 U8047 ( .A1(n11872), .A2(n12145), .ZN(n12141) );
  AOI21_X1 U8048 ( .B1(n11887), .B2(n11886), .A(n6741), .ZN(n12135) );
  NOR2_X1 U8049 ( .A1(n13477), .A2(n13478), .ZN(n7351) );
  XNOR2_X1 U8050 ( .A(n13527), .B(n13534), .ZN(n13528) );
  OAI21_X1 U8051 ( .B1(n13527), .B2(n7095), .A(n7093), .ZN(n13568) );
  AOI21_X1 U8052 ( .B1(n6557), .B2(n7708), .A(n6597), .ZN(n7095) );
  NAND2_X1 U8053 ( .A1(n13528), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n13548) );
  OAI211_X1 U8054 ( .C1(n13489), .C2(n6891), .A(P3_REG1_REG_15__SCAN_IN), .B(
        n6888), .ZN(n13535) );
  NAND2_X1 U8055 ( .A1(n6893), .A2(n6894), .ZN(n6891) );
  NOR2_X1 U8056 ( .A1(n6890), .A2(n6892), .ZN(n6889) );
  INV_X1 U8057 ( .A(n7344), .ZN(n7341) );
  AOI21_X1 U8058 ( .B1(n6565), .B2(n7348), .A(n6765), .ZN(n7347) );
  AOI21_X1 U8059 ( .B1(n13582), .B2(P3_REG1_REG_17__SCAN_IN), .A(n7260), .ZN(
        n13609) );
  AND2_X1 U8060 ( .A1(n13580), .A2(n13581), .ZN(n7260) );
  NAND2_X1 U8061 ( .A1(n8118), .A2(n8117), .ZN(n8572) );
  NAND2_X1 U8062 ( .A1(n8523), .A2(n8522), .ZN(n13672) );
  NAND2_X1 U8063 ( .A1(n13123), .A2(n13120), .ZN(n13663) );
  INV_X1 U8064 ( .A(n13663), .ZN(n13667) );
  AOI21_X1 U8065 ( .B1(n13683), .B2(n6924), .A(n6923), .ZN(n6922) );
  INV_X1 U8066 ( .A(n13113), .ZN(n6924) );
  INV_X1 U8067 ( .A(n13121), .ZN(n6923) );
  NAND2_X1 U8068 ( .A1(n16036), .A2(n7073), .ZN(n7069) );
  NAND2_X1 U8069 ( .A1(n7066), .A2(n6562), .ZN(n13677) );
  OR2_X1 U8070 ( .A1(n16036), .A2(n7071), .ZN(n7066) );
  NAND2_X1 U8071 ( .A1(n8111), .A2(n7321), .ZN(n8423) );
  NAND2_X1 U8072 ( .A1(n7964), .A2(n7965), .ZN(n7963) );
  OAI21_X1 U8073 ( .B1(n7841), .B2(n6564), .A(n13041), .ZN(n7840) );
  NAND2_X1 U8074 ( .A1(n13038), .A2(n6608), .ZN(n7842) );
  NAND3_X1 U8075 ( .A1(n8104), .A2(n6609), .A3(n8105), .ZN(n8257) );
  INV_X1 U8076 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n8105) );
  NAND2_X1 U8077 ( .A1(n8189), .A2(n7316), .ZN(n8209) );
  INV_X1 U8078 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n7316) );
  AND4_X1 U8079 ( .A1(n8149), .A2(n8148), .A3(n8147), .A4(n8146), .ZN(n11664)
         );
  NAND2_X1 U8080 ( .A1(n7063), .A2(n6785), .ZN(n7062) );
  NAND2_X1 U8081 ( .A1(n7065), .A2(n10506), .ZN(n7064) );
  INV_X1 U8082 ( .A(n12950), .ZN(n7063) );
  OAI21_X1 U8083 ( .B1(n10905), .B2(n10904), .A(n10903), .ZN(n15963) );
  INV_X1 U8084 ( .A(n10866), .ZN(n15982) );
  NAND2_X1 U8085 ( .A1(n12285), .A2(n12935), .ZN(n6962) );
  NAND2_X1 U8086 ( .A1(n8506), .A2(n8505), .ZN(n13119) );
  NAND2_X1 U8087 ( .A1(n8490), .A2(n8489), .ZN(n12898) );
  AOI21_X1 U8088 ( .B1(n7851), .B2(n13086), .A(n7850), .ZN(n7849) );
  INV_X1 U8089 ( .A(n13096), .ZN(n7850) );
  AND2_X1 U8090 ( .A1(n7851), .A2(n7168), .ZN(n6918) );
  INV_X1 U8091 ( .A(n7852), .ZN(n12895) );
  NAND2_X1 U8092 ( .A1(n6919), .A2(n7168), .ZN(n12894) );
  AND2_X1 U8093 ( .A1(n8441), .A2(n8440), .ZN(n13760) );
  AND2_X1 U8094 ( .A1(n7970), .A2(n6552), .ZN(n7967) );
  INV_X1 U8095 ( .A(n12885), .ZN(n6917) );
  INV_X1 U8096 ( .A(n7943), .ZN(n7942) );
  OAI21_X1 U8097 ( .B1(n11805), .B2(n7944), .A(n12069), .ZN(n7943) );
  INV_X1 U8098 ( .A(n15990), .ZN(n13828) );
  NAND2_X1 U8099 ( .A1(n13048), .A2(n6936), .ZN(n6935) );
  INV_X1 U8100 ( .A(n13047), .ZN(n6936) );
  AOI21_X1 U8101 ( .B1(n7839), .B2(n7841), .A(n7836), .ZN(n7835) );
  INV_X1 U8102 ( .A(n13042), .ZN(n7836) );
  AND2_X1 U8103 ( .A1(n6931), .A2(n6933), .ZN(n12527) );
  INV_X1 U8104 ( .A(n15992), .ZN(n13830) );
  INV_X1 U8105 ( .A(n12872), .ZN(n7692) );
  OR2_X1 U8106 ( .A1(n8046), .A2(n12223), .ZN(n8047) );
  NAND2_X1 U8107 ( .A1(n8444), .A2(n8037), .ZN(n8041) );
  NAND2_X1 U8108 ( .A1(n8035), .A2(n8034), .ZN(n8444) );
  INV_X1 U8109 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8074) );
  INV_X1 U8110 ( .A(n8102), .ZN(n8075) );
  XNOR2_X1 U8111 ( .A(n8444), .B(n11311), .ZN(n8443) );
  NAND2_X1 U8112 ( .A1(n8032), .A2(n8031), .ZN(n8420) );
  NAND2_X1 U8113 ( .A1(n7674), .A2(n8025), .ZN(n8360) );
  NAND2_X1 U8114 ( .A1(n8342), .A2(n7675), .ZN(n7674) );
  NAND2_X1 U8115 ( .A1(n8020), .A2(n8019), .ZN(n8314) );
  NAND2_X1 U8116 ( .A1(n7678), .A2(n7679), .ZN(n8281) );
  AOI21_X1 U8117 ( .B1(n7681), .B2(n7683), .A(n6700), .ZN(n7679) );
  XNOR2_X1 U8118 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n8280) );
  XNOR2_X1 U8119 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n8265) );
  AOI21_X1 U8120 ( .B1(n7671), .B2(n7669), .A(n6699), .ZN(n7668) );
  INV_X1 U8121 ( .A(n8134), .ZN(n7669) );
  INV_X1 U8122 ( .A(n7671), .ZN(n7670) );
  XNOR2_X1 U8123 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n8134) );
  OAI21_X1 U8124 ( .B1(n8008), .B2(n6975), .A(n6973), .ZN(n8135) );
  NAND2_X1 U8125 ( .A1(n8006), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8007) );
  INV_X1 U8126 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8006) );
  NAND2_X1 U8127 ( .A1(n6954), .A2(n8005), .ZN(n8183) );
  NAND2_X1 U8128 ( .A1(n8593), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8005) );
  XNOR2_X1 U8129 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8182) );
  NAND2_X1 U8130 ( .A1(n7575), .A2(n9960), .ZN(n8253) );
  NAND2_X1 U8131 ( .A1(n7085), .A2(n7084), .ZN(n11150) );
  INV_X1 U8132 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7085) );
  INV_X1 U8133 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7084) );
  XNOR2_X1 U8134 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8152) );
  NAND2_X1 U8135 ( .A1(n9494), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8168) );
  NAND3_X1 U8136 ( .A1(n6866), .A2(n9447), .A3(P2_REG3_REG_5__SCAN_IN), .ZN(
        n9584) );
  AND2_X1 U8137 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n9447) );
  OAI21_X1 U8138 ( .B1(n12476), .B2(n7039), .A(n7037), .ZN(n10470) );
  XNOR2_X1 U8139 ( .A(n6546), .B(n12688), .ZN(n10419) );
  NAND2_X1 U8140 ( .A1(n6866), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9571) );
  AND3_X1 U8141 ( .A1(n10478), .A2(n15914), .A3(n10487), .ZN(n10486) );
  AOI21_X1 U8142 ( .B1(n6561), .B2(n12802), .A(n14076), .ZN(n7027) );
  AND2_X1 U8143 ( .A1(n6623), .A2(n6561), .ZN(n7026) );
  NAND2_X1 U8144 ( .A1(n12792), .A2(n6752), .ZN(n14073) );
  AND4_X1 U8145 ( .A1(n9661), .A2(n9660), .A3(n9659), .A4(n9658), .ZN(n14205)
         );
  AND4_X1 U8146 ( .A1(n9604), .A2(n9603), .A3(n9602), .A4(n9601), .ZN(n12329)
         );
  NAND2_X1 U8147 ( .A1(n10321), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n9499) );
  NAND2_X1 U8148 ( .A1(n7527), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9500) );
  NOR2_X1 U8149 ( .A1(n7108), .A2(n9477), .ZN(n7531) );
  AND2_X1 U8150 ( .A1(n7108), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7529) );
  NAND2_X1 U8151 ( .A1(n7301), .A2(n7299), .ZN(n11086) );
  NOR2_X1 U8152 ( .A1(n7300), .A2(n11044), .ZN(n7299) );
  INV_X1 U8153 ( .A(n7303), .ZN(n7300) );
  INV_X1 U8154 ( .A(n15887), .ZN(n7308) );
  NOR2_X1 U8155 ( .A1(n11090), .A2(n7310), .ZN(n7309) );
  INV_X1 U8156 ( .A(n11088), .ZN(n7310) );
  OR2_X1 U8157 ( .A1(n14301), .A2(n14312), .ZN(n7298) );
  NAND2_X1 U8158 ( .A1(n7297), .A2(n7296), .ZN(n14321) );
  INV_X1 U8159 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n7296) );
  INV_X1 U8160 ( .A(n14304), .ZN(n7297) );
  NOR2_X1 U8161 ( .A1(n14381), .A2(n7283), .ZN(n7282) );
  NAND2_X1 U8162 ( .A1(n7277), .A2(n7276), .ZN(n6792) );
  NOR2_X1 U8163 ( .A1(n14392), .A2(n7284), .ZN(n7283) );
  AND2_X1 U8164 ( .A1(n9809), .A2(n9858), .ZN(n14366) );
  NOR2_X1 U8165 ( .A1(n10396), .A2(n7409), .ZN(n7408) );
  NOR2_X1 U8166 ( .A1(n14403), .A2(n7410), .ZN(n7409) );
  INV_X1 U8167 ( .A(n9804), .ZN(n7410) );
  XNOR2_X1 U8168 ( .A(n14695), .B(n12818), .ZN(n14403) );
  NAND2_X1 U8169 ( .A1(n14416), .A2(n9792), .ZN(n14404) );
  NAND2_X1 U8170 ( .A1(n14404), .A2(n14403), .ZN(n14402) );
  NAND2_X1 U8171 ( .A1(n14436), .A2(n6572), .ZN(n14396) );
  INV_X1 U8172 ( .A(n14403), .ZN(n14392) );
  NAND2_X1 U8173 ( .A1(n7277), .A2(n7278), .ZN(n14391) );
  NAND2_X1 U8174 ( .A1(n14427), .A2(n7239), .ZN(n14418) );
  NAND2_X1 U8175 ( .A1(n14705), .A2(n14198), .ZN(n7239) );
  NAND2_X1 U8176 ( .A1(n14418), .A2(n14417), .ZN(n14416) );
  NAND2_X1 U8177 ( .A1(n9764), .A2(n9763), .ZN(n12751) );
  AND2_X1 U8178 ( .A1(n7754), .A2(n9758), .ZN(n7753) );
  NAND2_X1 U8179 ( .A1(n7526), .A2(n8003), .ZN(n7525) );
  NOR2_X1 U8180 ( .A1(n14544), .A2(n14506), .ZN(n14523) );
  NAND2_X1 U8181 ( .A1(n14523), .A2(n14522), .ZN(n14521) );
  NAND2_X1 U8182 ( .A1(n14607), .A2(n9690), .ZN(n9692) );
  AND2_X1 U8183 ( .A1(n7749), .A2(n7117), .ZN(n7116) );
  NAND2_X1 U8184 ( .A1(n7118), .A2(n9706), .ZN(n7117) );
  INV_X1 U8185 ( .A(n7750), .ZN(n7749) );
  INV_X1 U8186 ( .A(n9691), .ZN(n7118) );
  NAND2_X1 U8187 ( .A1(n6795), .A2(n9834), .ZN(n14502) );
  NOR2_X1 U8188 ( .A1(n14502), .A2(n14561), .ZN(n14560) );
  NAND2_X1 U8189 ( .A1(n9692), .A2(n9691), .ZN(n14587) );
  XNOR2_X1 U8190 ( .A(n14754), .B(n14576), .ZN(n14609) );
  NAND2_X1 U8191 ( .A1(n9831), .A2(n7887), .ZN(n14596) );
  INV_X1 U8192 ( .A(n9827), .ZN(n7902) );
  OR2_X1 U8193 ( .A1(n14651), .A2(n9826), .ZN(n7903) );
  NOR2_X1 U8194 ( .A1(n14639), .A2(n14641), .ZN(n14640) );
  AND2_X1 U8195 ( .A1(n14823), .A2(n7619), .ZN(n7620) );
  NAND2_X1 U8196 ( .A1(n12502), .A2(n9825), .ZN(n14651) );
  OR2_X1 U8197 ( .A1(n9630), .A2(n14145), .ZN(n9641) );
  INV_X1 U8198 ( .A(n9822), .ZN(n7293) );
  NAND2_X1 U8199 ( .A1(n12241), .A2(n9865), .ZN(n9866) );
  NAND2_X1 U8200 ( .A1(n12126), .A2(n9819), .ZN(n9821) );
  NOR2_X1 U8201 ( .A1(n6847), .A2(n11971), .ZN(n6845) );
  NOR2_X1 U8202 ( .A1(n10386), .A2(n6848), .ZN(n6847) );
  XNOR2_X1 U8203 ( .A(n14211), .B(n15932), .ZN(n11971) );
  NAND2_X1 U8204 ( .A1(n11967), .A2(n11971), .ZN(n11966) );
  NAND2_X1 U8205 ( .A1(n12104), .A2(n6802), .ZN(n11991) );
  NAND2_X1 U8206 ( .A1(n12091), .A2(n12084), .ZN(n12107) );
  OR2_X1 U8207 ( .A1(n11022), .A2(n7295), .ZN(n14638) );
  AND2_X1 U8208 ( .A1(n10414), .A2(n12688), .ZN(n12113) );
  NAND2_X1 U8209 ( .A1(n9496), .A2(n12089), .ZN(n12093) );
  INV_X1 U8210 ( .A(n14638), .ZN(n14654) );
  INV_X1 U8211 ( .A(n10482), .ZN(n11864) );
  OR2_X1 U8212 ( .A1(n12254), .A2(n6842), .ZN(n12255) );
  AND2_X1 U8213 ( .A1(n11026), .A2(n9485), .ZN(n9486) );
  NAND2_X1 U8214 ( .A1(n9883), .A2(n9882), .ZN(n9885) );
  AND2_X1 U8215 ( .A1(n9423), .A2(n9440), .ZN(n6820) );
  INV_X1 U8216 ( .A(n9707), .ZN(n6821) );
  INV_X1 U8217 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9551) );
  NAND2_X1 U8218 ( .A1(n6938), .A2(n6937), .ZN(n11905) );
  AOI21_X1 U8219 ( .B1(n7716), .B2(n7715), .A(n6611), .ZN(n7714) );
  INV_X1 U8220 ( .A(n7718), .ZN(n7715) );
  NAND2_X1 U8221 ( .A1(n11303), .A2(n11304), .ZN(n10991) );
  INV_X1 U8222 ( .A(n10988), .ZN(n10989) );
  OR2_X1 U8223 ( .A1(n13181), .A2(n13182), .ZN(n6952) );
  INV_X1 U8224 ( .A(n7727), .ZN(n7726) );
  AND2_X1 U8225 ( .A1(n10874), .A2(n8000), .ZN(n10879) );
  OR2_X1 U8226 ( .A1(n13223), .A2(n15749), .ZN(n10874) );
  INV_X1 U8227 ( .A(n6948), .ZN(n14867) );
  INV_X1 U8228 ( .A(n9216), .ZN(n8749) );
  NAND2_X1 U8229 ( .A1(n6942), .A2(n6947), .ZN(n6940) );
  AND2_X1 U8230 ( .A1(n11787), .A2(n11786), .ZN(n11897) );
  NAND2_X1 U8231 ( .A1(n8751), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n9321) );
  OAI22_X1 U8232 ( .A1(n13225), .A2(n13224), .B1(n14852), .B2(n13223), .ZN(
        n13229) );
  NAND2_X1 U8233 ( .A1(n7609), .A2(n9303), .ZN(n7608) );
  OR2_X1 U8234 ( .A1(n7609), .A2(n9303), .ZN(n7607) );
  NOR2_X1 U8235 ( .A1(n9364), .A2(n9360), .ZN(n9352) );
  AND2_X1 U8236 ( .A1(n10958), .A2(n10955), .ZN(n11438) );
  AND4_X1 U8237 ( .A1(n8977), .A2(n8976), .A3(n8975), .A4(n8974), .ZN(n12432)
         );
  NAND2_X1 U8238 ( .A1(n10711), .A2(n6878), .ZN(n6877) );
  INV_X1 U8239 ( .A(n7486), .ZN(n6878) );
  OR2_X1 U8240 ( .A1(n15065), .A2(n7491), .ZN(n7490) );
  AND2_X1 U8241 ( .A1(n15066), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7491) );
  NAND2_X1 U8242 ( .A1(n6835), .A2(n6834), .ZN(n15105) );
  INV_X1 U8243 ( .A(n15094), .ZN(n6834) );
  INV_X1 U8244 ( .A(n15095), .ZN(n6835) );
  NOR2_X1 U8245 ( .A1(n15083), .A2(n15721), .ZN(n6872) );
  NOR2_X1 U8246 ( .A1(n6872), .A2(n15085), .ZN(n6869) );
  XNOR2_X1 U8247 ( .A(n15135), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n15145) );
  NOR2_X1 U8248 ( .A1(n15134), .A2(n15133), .ZN(n15135) );
  NAND2_X1 U8249 ( .A1(n8697), .A2(n8696), .ZN(n15152) );
  NAND2_X1 U8250 ( .A1(n8761), .A2(n8760), .ZN(n15175) );
  XNOR2_X1 U8251 ( .A(n15175), .B(n14997), .ZN(n15168) );
  NAND2_X1 U8252 ( .A1(n7633), .A2(n6672), .ZN(n15191) );
  INV_X1 U8253 ( .A(n7434), .ZN(n7433) );
  AOI21_X1 U8254 ( .B1(n7434), .B2(n7808), .A(n7432), .ZN(n7431) );
  INV_X1 U8255 ( .A(n12707), .ZN(n7432) );
  NAND2_X1 U8256 ( .A1(n15236), .A2(n15235), .ZN(n15209) );
  NAND2_X1 U8257 ( .A1(n7652), .A2(n7654), .ZN(n7650) );
  NAND2_X1 U8258 ( .A1(n7653), .A2(n12729), .ZN(n7652) );
  INV_X1 U8259 ( .A(n12728), .ZN(n7653) );
  OR2_X1 U8260 ( .A1(n7651), .A2(n6571), .ZN(n7649) );
  INV_X1 U8261 ( .A(n15290), .ZN(n7651) );
  AND2_X1 U8262 ( .A1(n7649), .A2(n7647), .ZN(n15243) );
  NOR2_X1 U8264 ( .A1(n12727), .A2(n15507), .ZN(n12728) );
  NAND2_X1 U8265 ( .A1(n15298), .A2(n12726), .ZN(n15290) );
  NAND2_X1 U8266 ( .A1(n15512), .A2(n15003), .ZN(n12726) );
  INV_X1 U8267 ( .A(n7446), .ZN(n7444) );
  NAND2_X1 U8268 ( .A1(n7641), .A2(n7640), .ZN(n15298) );
  AND2_X1 U8269 ( .A1(n12725), .A2(n15299), .ZN(n7640) );
  NAND2_X1 U8270 ( .A1(n12700), .A2(n7447), .ZN(n7446) );
  NAND2_X1 U8271 ( .A1(n7800), .A2(n7799), .ZN(n12699) );
  AOI21_X1 U8272 ( .B1(n7801), .B2(n7803), .A(n6677), .ZN(n7799) );
  NAND2_X1 U8273 ( .A1(n7004), .A2(n7981), .ZN(n12724) );
  NAND2_X1 U8274 ( .A1(n12712), .A2(n7006), .ZN(n7004) );
  OR2_X1 U8275 ( .A1(n9108), .A2(n8746), .ZN(n9093) );
  AND2_X1 U8276 ( .A1(n9165), .A2(n9164), .ZN(n15341) );
  NAND2_X1 U8277 ( .A1(n12713), .A2(n12717), .ZN(n12715) );
  AND2_X1 U8278 ( .A1(n15363), .A2(n15345), .ZN(n15343) );
  INV_X1 U8279 ( .A(n14965), .ZN(n15345) );
  AOI21_X1 U8280 ( .B1(n6567), .B2(n7802), .A(n6678), .ZN(n7801) );
  INV_X1 U8281 ( .A(n15376), .ZN(n7802) );
  INV_X1 U8282 ( .A(n6567), .ZN(n7803) );
  OR2_X1 U8283 ( .A1(n12697), .A2(n6678), .ZN(n15357) );
  NAND2_X1 U8284 ( .A1(n15402), .A2(n7419), .ZN(n7418) );
  NAND2_X1 U8285 ( .A1(n15375), .A2(n15376), .ZN(n15374) );
  NAND2_X1 U8286 ( .A1(n9055), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9108) );
  NAND2_X1 U8287 ( .A1(n12165), .A2(n6554), .ZN(n12617) );
  NAND2_X1 U8288 ( .A1(n12165), .A2(n14964), .ZN(n12387) );
  NAND2_X1 U8289 ( .A1(n11958), .A2(n11957), .ZN(n12010) );
  NAND2_X1 U8290 ( .A1(n8740), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n8824) );
  INV_X1 U8291 ( .A(n8822), .ZN(n8740) );
  NAND2_X1 U8292 ( .A1(n6681), .A2(n6905), .ZN(n11760) );
  XNOR2_X1 U8293 ( .A(n11742), .B(n15017), .ZN(n11709) );
  NOR2_X1 U8294 ( .A1(n6902), .A2(n15435), .ZN(n11532) );
  NAND2_X1 U8295 ( .A1(n6903), .A2(n11534), .ZN(n6902) );
  NAND2_X1 U8296 ( .A1(n8869), .A2(n15753), .ZN(n15738) );
  INV_X1 U8297 ( .A(n15159), .ZN(n15447) );
  NAND2_X1 U8298 ( .A1(n9157), .A2(n9156), .ZN(n15519) );
  NAND2_X1 U8299 ( .A1(n9332), .A2(n6556), .ZN(n7147) );
  AOI21_X1 U8300 ( .B1(n6556), .B2(n7151), .A(n6774), .ZN(n7148) );
  AND2_X1 U8301 ( .A1(n8717), .A2(n6716), .ZN(n7822) );
  NAND2_X1 U8302 ( .A1(n6886), .A2(n7821), .ZN(n8695) );
  AND2_X1 U8303 ( .A1(n8717), .A2(n7427), .ZN(n6886) );
  NOR2_X1 U8304 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n7427) );
  INV_X1 U8305 ( .A(n8695), .ZN(n7181) );
  NOR2_X1 U8306 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n7180) );
  INV_X1 U8307 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7426) );
  NAND2_X1 U8308 ( .A1(n7821), .A2(n8717), .ZN(n9373) );
  INV_X1 U8309 ( .A(n9124), .ZN(n8714) );
  INV_X1 U8310 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8710) );
  OR2_X1 U8311 ( .A1(n6987), .A2(n6983), .ZN(n9124) );
  NAND2_X1 U8312 ( .A1(n8689), .A2(n6612), .ZN(n6983) );
  NAND2_X1 U8313 ( .A1(n9064), .A2(n9063), .ZN(n9066) );
  AND2_X1 U8314 ( .A1(n8810), .A2(n8809), .ZN(n10617) );
  OR2_X1 U8315 ( .A1(n8808), .A2(n8807), .ZN(n8809) );
  NAND2_X1 U8316 ( .A1(n7123), .A2(n8605), .ZN(n8918) );
  NAND2_X1 U8317 ( .A1(n8858), .A2(n8857), .ZN(n8880) );
  INV_X1 U8318 ( .A(n7056), .ZN(n7055) );
  INV_X1 U8319 ( .A(n10547), .ZN(n7057) );
  NAND2_X1 U8320 ( .A1(n10545), .A2(n10544), .ZN(n10816) );
  NAND2_X1 U8321 ( .A1(n7497), .A2(n10820), .ZN(n10828) );
  OAI21_X1 U8322 ( .B1(n11319), .B2(n11318), .A(n11321), .ZN(n11620) );
  OAI21_X1 U8323 ( .B1(n10842), .B2(n7502), .A(n11317), .ZN(n7501) );
  NAND2_X1 U8324 ( .A1(n8479), .A2(n8478), .ZN(n13710) );
  NAND2_X1 U8325 ( .A1(n13415), .A2(n8418), .ZN(n13311) );
  INV_X1 U8326 ( .A(n7930), .ZN(n7929) );
  NAND2_X1 U8327 ( .A1(n7933), .A2(n7932), .ZN(n7931) );
  OAI21_X1 U8328 ( .B1(n12063), .B2(n7993), .A(n7935), .ZN(n7930) );
  AND2_X1 U8329 ( .A1(n8497), .A2(n8496), .ZN(n13704) );
  NAND2_X1 U8330 ( .A1(n10853), .A2(n8196), .ZN(n10924) );
  NOR2_X1 U8331 ( .A1(n7907), .A2(n7909), .ZN(n11103) );
  INV_X1 U8332 ( .A(n10924), .ZN(n7907) );
  NAND2_X1 U8333 ( .A1(n8331), .A2(n8330), .ZN(n13389) );
  AND2_X1 U8334 ( .A1(n8457), .A2(n8456), .ZN(n13398) );
  AND2_X1 U8335 ( .A1(n8429), .A2(n8428), .ZN(n13772) );
  AND3_X1 U8336 ( .A1(n8378), .A2(n8377), .A3(n8376), .ZN(n13812) );
  AND2_X1 U8337 ( .A1(n8565), .A2(n11374), .ZN(n13437) );
  NAND2_X1 U8338 ( .A1(n8513), .A2(n8512), .ZN(n13665) );
  INV_X1 U8339 ( .A(n13398), .ZN(n13744) );
  OAI211_X1 U8340 ( .C1(n12264), .C2(n13898), .A(n8371), .B(n8370), .ZN(n13831) );
  OAI211_X1 U8341 ( .C1(n12264), .C2(n13901), .A(n8356), .B(n8355), .ZN(n13452) );
  NAND4_X1 U8342 ( .A1(n8338), .A2(n8337), .A3(n8336), .A4(n8335), .ZN(n13829)
         );
  XNOR2_X1 U8343 ( .A(n11326), .B(n11225), .ZN(n11328) );
  NAND2_X1 U8344 ( .A1(n11328), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n6900) );
  XNOR2_X1 U8345 ( .A(n11557), .B(n11483), .ZN(n11561) );
  NAND2_X1 U8346 ( .A1(n13538), .A2(n13537), .ZN(n13557) );
  AND2_X1 U8347 ( .A1(n13621), .A2(n7089), .ZN(n7088) );
  OAI22_X1 U8348 ( .A1(n13609), .A2(n13608), .B1(n13607), .B2(n13887), .ZN(
        n13611) );
  NAND2_X1 U8349 ( .A1(n8450), .A2(n8449), .ZN(n13874) );
  AND3_X1 U8350 ( .A1(n8207), .A2(n8206), .A3(n8205), .ZN(n16006) );
  OR2_X1 U8351 ( .A1(n15981), .A2(n8567), .ZN(n15985) );
  AND2_X1 U8352 ( .A1(n13911), .A2(n16011), .ZN(n13893) );
  NAND2_X1 U8353 ( .A1(n12953), .A2(n12952), .ZN(n13915) );
  OR2_X1 U8354 ( .A1(n13256), .A2(n12950), .ZN(n12953) );
  NAND2_X1 U8355 ( .A1(n7977), .A2(n7976), .ZN(n7975) );
  XNOR2_X1 U8356 ( .A(n12927), .B(n12926), .ZN(n13845) );
  AOI21_X1 U8357 ( .B1(n6928), .B2(n6930), .A(n7847), .ZN(n6925) );
  NAND2_X1 U8358 ( .A1(n12878), .A2(n12877), .ZN(n13844) );
  OR2_X1 U8359 ( .A1(n14009), .A2(n12950), .ZN(n12878) );
  NAND2_X1 U8360 ( .A1(n12867), .A2(n12866), .ZN(n13921) );
  XNOR2_X1 U8361 ( .A(n13634), .B(n13635), .ZN(n13922) );
  NAND2_X1 U8362 ( .A1(n8466), .A2(n8465), .ZN(n13948) );
  AND2_X1 U8363 ( .A1(n8393), .A2(n8392), .ZN(n13974) );
  NAND2_X1 U8364 ( .A1(n8350), .A2(n8349), .ZN(n13996) );
  AND2_X1 U8365 ( .A1(n8239), .A2(n8238), .ZN(n15950) );
  OR2_X1 U8366 ( .A1(n16018), .A2(n15981), .ZN(n13997) );
  NAND2_X1 U8367 ( .A1(n8101), .A2(n8102), .ZN(n13599) );
  NAND2_X1 U8368 ( .A1(n12908), .A2(n10335), .ZN(n9446) );
  INV_X1 U8369 ( .A(n12816), .ZN(n7225) );
  NAND2_X1 U8370 ( .A1(n14023), .A2(n14022), .ZN(n14072) );
  XNOR2_X1 U8371 ( .A(n14073), .B(n14071), .ZN(n14023) );
  NAND2_X1 U8372 ( .A1(n9772), .A2(n9771), .ZN(n14710) );
  AND2_X1 U8373 ( .A1(n14189), .A2(n6802), .ZN(n6799) );
  NAND2_X1 U8374 ( .A1(n7228), .A2(n7227), .ZN(n14109) );
  INV_X1 U8375 ( .A(n11675), .ZN(n7227) );
  NAND2_X1 U8376 ( .A1(n11346), .A2(n10335), .ZN(n9729) );
  AND2_X1 U8377 ( .A1(n12813), .A2(n12812), .ZN(n14049) );
  AND2_X1 U8378 ( .A1(n14042), .A2(n14180), .ZN(n14050) );
  NAND2_X1 U8379 ( .A1(n10416), .A2(n13269), .ZN(n11681) );
  NAND2_X1 U8380 ( .A1(n12767), .A2(n12766), .ZN(n12849) );
  OR2_X1 U8381 ( .A1(n12824), .A2(n9793), .ZN(n9747) );
  AND4_X1 U8382 ( .A1(n9672), .A2(n9671), .A3(n9670), .A4(n9669), .ZN(n14637)
         );
  AND2_X1 U8383 ( .A1(n10493), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14168) );
  INV_X1 U8384 ( .A(n14168), .ZN(n14186) );
  INV_X1 U8385 ( .A(n14154), .ZN(n14180) );
  OR2_X1 U8386 ( .A1(n14167), .A2(n9517), .ZN(n9803) );
  NAND2_X1 U8387 ( .A1(n6857), .A2(n9745), .ZN(n14200) );
  NAND2_X1 U8388 ( .A1(n6858), .A2(n7527), .ZN(n6857) );
  INV_X1 U8389 ( .A(n12548), .ZN(n14210) );
  NAND2_X1 U8390 ( .A1(n14235), .A2(n11032), .ZN(n15862) );
  NAND2_X1 U8391 ( .A1(n7752), .A2(n9705), .ZN(n14748) );
  INV_X1 U8392 ( .A(n14587), .ZN(n7752) );
  AND2_X1 U8393 ( .A1(n14672), .A2(n12303), .ZN(n6801) );
  NAND2_X1 U8394 ( .A1(n15914), .A2(n10483), .ZN(n14642) );
  INV_X1 U8395 ( .A(n14664), .ZN(n14433) );
  AND2_X1 U8396 ( .A1(n9853), .A2(n11860), .ZN(n11866) );
  OAI21_X1 U8397 ( .B1(n14348), .B2(n7742), .A(n7741), .ZN(n7740) );
  NOR2_X1 U8398 ( .A1(n9856), .A2(n7743), .ZN(n7742) );
  NAND2_X1 U8399 ( .A1(n14348), .A2(n14344), .ZN(n7741) );
  NAND2_X1 U8400 ( .A1(n9815), .A2(n6632), .ZN(n7736) );
  NAND2_X1 U8401 ( .A1(n7739), .A2(n6650), .ZN(n7738) );
  INV_X1 U8402 ( .A(n9815), .ZN(n7739) );
  AND2_X1 U8403 ( .A1(n7878), .A2(n14356), .ZN(n7876) );
  INV_X1 U8404 ( .A(n14687), .ZN(n7878) );
  NAND2_X1 U8405 ( .A1(n14350), .A2(n14657), .ZN(n14357) );
  AOI21_X1 U8406 ( .B1(n7881), .B2(n14381), .A(n6682), .ZN(n7880) );
  NOR2_X1 U8407 ( .A1(n7106), .A2(n6753), .ZN(n7104) );
  AND2_X1 U8408 ( .A1(n14345), .A2(n6594), .ZN(n7102) );
  NAND2_X1 U8409 ( .A1(n15944), .A2(n14770), .ZN(n14781) );
  NAND2_X1 U8410 ( .A1(n13275), .A2(n10335), .ZN(n10327) );
  OR2_X1 U8411 ( .A1(n7876), .A2(n15938), .ZN(n7874) );
  NAND2_X1 U8412 ( .A1(n15938), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7877) );
  INV_X1 U8413 ( .A(n14357), .ZN(n7871) );
  NOR2_X1 U8414 ( .A1(n6634), .A2(n6804), .ZN(n6803) );
  NAND2_X1 U8415 ( .A1(n9903), .A2(n9902), .ZN(n15910) );
  NAND2_X1 U8416 ( .A1(n9876), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9442) );
  AND2_X1 U8417 ( .A1(n9088), .A2(n9087), .ZN(n15321) );
  NAND2_X1 U8418 ( .A1(n7189), .A2(n7720), .ZN(n7188) );
  NAND2_X1 U8419 ( .A1(n14926), .A2(n14927), .ZN(n7189) );
  NAND2_X1 U8420 ( .A1(n12477), .A2(n9333), .ZN(n9282) );
  NAND2_X1 U8421 ( .A1(n12220), .A2(n9333), .ZN(n9265) );
  OR2_X1 U8422 ( .A1(n12824), .A2(n8897), .ZN(n9193) );
  NAND3_X1 U8423 ( .A1(n8885), .A2(n8884), .A3(n8883), .ZN(n15439) );
  NAND2_X1 U8424 ( .A1(n7713), .A2(n7716), .ZN(n14977) );
  NAND2_X1 U8425 ( .A1(n6977), .A2(n6976), .ZN(n9357) );
  AOI21_X1 U8426 ( .B1(n6978), .B2(n6981), .A(n6588), .ZN(n6976) );
  NAND2_X1 U8427 ( .A1(n9318), .A2(n6978), .ZN(n6977) );
  AND2_X1 U8428 ( .A1(n9319), .A2(n6982), .ZN(n6981) );
  INV_X1 U8429 ( .A(n15274), .ZN(n15000) );
  INV_X1 U8430 ( .A(n14839), .ZN(n15016) );
  NAND2_X1 U8431 ( .A1(n8887), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n8864) );
  NAND2_X1 U8432 ( .A1(n7187), .A2(n7186), .ZN(n15026) );
  NAND2_X1 U8433 ( .A1(n10678), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7186) );
  OR2_X1 U8434 ( .A1(n10678), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7187) );
  NOR2_X1 U8435 ( .A1(n11768), .A2(n11769), .ZN(n15065) );
  XNOR2_X1 U8436 ( .A(n15082), .B(n7487), .ZN(n15719) );
  INV_X1 U8437 ( .A(n15721), .ZN(n7487) );
  NAND2_X1 U8438 ( .A1(n15718), .A2(n15717), .ZN(n15716) );
  NAND2_X1 U8439 ( .A1(n13258), .A2(n9333), .ZN(n9335) );
  AND2_X1 U8440 ( .A1(n6710), .A2(n12741), .ZN(n7451) );
  AND2_X1 U8441 ( .A1(n12740), .A2(n15471), .ZN(n6913) );
  INV_X1 U8442 ( .A(n7451), .ZN(n7450) );
  NOR2_X1 U8443 ( .A1(n15792), .A2(n7453), .ZN(n7452) );
  NAND2_X1 U8444 ( .A1(n15473), .A2(n12708), .ZN(n12709) );
  NAND2_X1 U8445 ( .A1(n10562), .A2(n10563), .ZN(n15668) );
  AND2_X1 U8446 ( .A1(n7504), .A2(n16026), .ZN(n15603) );
  NAND2_X1 U8447 ( .A1(n16025), .A2(n16027), .ZN(n7504) );
  XNOR2_X1 U8448 ( .A(n10841), .B(n10839), .ZN(n15609) );
  AND2_X1 U8449 ( .A1(n7765), .A2(n7767), .ZN(n7764) );
  INV_X1 U8450 ( .A(n11624), .ZN(n7765) );
  NAND2_X1 U8451 ( .A1(n11832), .A2(n11831), .ZN(n12290) );
  AND2_X1 U8452 ( .A1(n7046), .A2(n7044), .ZN(n12582) );
  AND2_X1 U8453 ( .A1(n12296), .A2(n11831), .ZN(n7045) );
  OR2_X1 U8454 ( .A1(n12591), .A2(n12590), .ZN(n7521) );
  NAND3_X1 U8455 ( .A1(n7521), .A2(n15610), .A3(n7755), .ZN(n15611) );
  INV_X1 U8456 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7755) );
  INV_X1 U8457 ( .A(n15631), .ZN(n7510) );
  INV_X1 U8458 ( .A(n7508), .ZN(n7507) );
  OAI21_X1 U8459 ( .B1(n9131), .B2(n7243), .A(n7242), .ZN(n8873) );
  NOR2_X1 U8460 ( .A1(n7208), .A2(n7207), .ZN(n7206) );
  INV_X1 U8461 ( .A(n13009), .ZN(n7208) );
  NAND2_X1 U8462 ( .A1(n10194), .A2(n12114), .ZN(n10178) );
  AND2_X1 U8463 ( .A1(n13037), .A2(n13036), .ZN(n7261) );
  NAND2_X1 U8464 ( .A1(n6613), .A2(n7484), .ZN(n7482) );
  AND2_X1 U8465 ( .A1(n8958), .A2(n8957), .ZN(n8959) );
  INV_X1 U8466 ( .A(n7776), .ZN(n7772) );
  NAND2_X1 U8467 ( .A1(n7795), .A2(n6606), .ZN(n7794) );
  INV_X1 U8468 ( .A(n7474), .ZN(n7473) );
  AND2_X1 U8469 ( .A1(n7480), .A2(n6643), .ZN(n7479) );
  OR2_X1 U8470 ( .A1(n10207), .A2(n10209), .ZN(n7480) );
  AND2_X1 U8471 ( .A1(n9023), .A2(n6970), .ZN(n6969) );
  INV_X1 U8472 ( .A(n9021), .ZN(n6970) );
  AND3_X1 U8473 ( .A1(n7602), .A2(n7604), .A3(n7600), .ZN(n9022) );
  AND2_X1 U8474 ( .A1(n13069), .A2(n13826), .ZN(n7263) );
  NAND2_X1 U8475 ( .A1(n10212), .A2(n6830), .ZN(n6829) );
  NAND2_X1 U8476 ( .A1(n10220), .A2(n7785), .ZN(n7784) );
  NAND2_X1 U8477 ( .A1(n9166), .A2(n9382), .ZN(n7592) );
  NAND2_X1 U8478 ( .A1(n9176), .A2(n9175), .ZN(n7591) );
  AND2_X1 U8479 ( .A1(n9143), .A2(n12720), .ZN(n7596) );
  NOR2_X1 U8480 ( .A1(n7785), .A2(n10220), .ZN(n7783) );
  INV_X1 U8481 ( .A(n9794), .ZN(n7563) );
  OAI22_X1 U8482 ( .A1(n6614), .A2(n6832), .B1(n10226), .B2(n7485), .ZN(n6831)
         );
  INV_X1 U8483 ( .A(n10225), .ZN(n7485) );
  NAND2_X1 U8484 ( .A1(n6833), .A2(n6636), .ZN(n6832) );
  NAND2_X1 U8485 ( .A1(n10229), .A2(n7792), .ZN(n7791) );
  NAND2_X1 U8486 ( .A1(n7788), .A2(n7789), .ZN(n7470) );
  NAND2_X1 U8487 ( .A1(n10228), .A2(n7790), .ZN(n7789) );
  NAND2_X1 U8488 ( .A1(n6831), .A2(n7791), .ZN(n7788) );
  INV_X1 U8489 ( .A(n10229), .ZN(n7790) );
  NAND2_X1 U8490 ( .A1(n7205), .A2(n13101), .ZN(n7204) );
  NAND2_X1 U8491 ( .A1(n7266), .A2(n13667), .ZN(n6959) );
  INV_X1 U8492 ( .A(n13120), .ZN(n7205) );
  AND2_X1 U8493 ( .A1(n6842), .A2(n10382), .ZN(n6841) );
  AND2_X1 U8494 ( .A1(n12236), .A2(n12275), .ZN(n6811) );
  INV_X1 U8495 ( .A(n14632), .ZN(n6812) );
  NAND2_X1 U8496 ( .A1(n10293), .A2(n10250), .ZN(n10297) );
  INV_X1 U8497 ( .A(n7565), .ZN(n10305) );
  NAND2_X1 U8498 ( .A1(n7241), .A2(n7458), .ZN(n7240) );
  INV_X1 U8499 ( .A(n10271), .ZN(n7241) );
  NAND2_X1 U8500 ( .A1(n7461), .A2(n7459), .ZN(n7458) );
  OR2_X1 U8501 ( .A1(n12650), .A2(n12569), .ZN(n12437) );
  INV_X1 U8502 ( .A(n9226), .ZN(n7588) );
  INV_X1 U8503 ( .A(n8635), .ZN(n7138) );
  NAND2_X1 U8504 ( .A1(n8831), .A2(n8618), .ZN(n8617) );
  NAND2_X1 U8505 ( .A1(n10153), .A2(n6635), .ZN(n7376) );
  OAI22_X1 U8506 ( .A1(n13914), .A2(n13447), .B1(n12958), .B2(n13915), .ZN(
        n12969) );
  INV_X1 U8507 ( .A(n8068), .ZN(n7332) );
  NOR2_X1 U8508 ( .A1(n12859), .A2(n13731), .ZN(n12860) );
  INV_X1 U8509 ( .A(n16006), .ZN(n11407) );
  INV_X1 U8510 ( .A(n13777), .ZN(n13739) );
  INV_X1 U8511 ( .A(n8043), .ZN(n7686) );
  NAND2_X1 U8512 ( .A1(n10358), .A2(n10359), .ZN(n7254) );
  NAND2_X1 U8513 ( .A1(n7457), .A2(n7460), .ZN(n7455) );
  INV_X1 U8514 ( .A(n7461), .ZN(n7460) );
  INV_X1 U8515 ( .A(n7280), .ZN(n7279) );
  INV_X1 U8516 ( .A(n14417), .ZN(n7281) );
  NOR2_X1 U8517 ( .A1(n6856), .A2(n6855), .ZN(n6854) );
  AND2_X1 U8518 ( .A1(n14491), .A2(n14200), .ZN(n6856) );
  INV_X1 U8519 ( .A(n9736), .ZN(n6855) );
  NOR2_X1 U8520 ( .A1(n9666), .A2(n11694), .ZN(n6861) );
  NAND2_X1 U8521 ( .A1(n6808), .A2(n9455), .ZN(n6807) );
  INV_X1 U8522 ( .A(n6809), .ZN(n6808) );
  INV_X1 U8523 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n9439) );
  NAND2_X1 U8524 ( .A1(n8733), .A2(n8732), .ZN(n8933) );
  NAND2_X1 U8525 ( .A1(n8736), .A2(n10793), .ZN(n8733) );
  NAND2_X1 U8526 ( .A1(n8731), .A2(n10808), .ZN(n8736) );
  INV_X1 U8527 ( .A(n7006), .ZN(n7005) );
  NAND2_X1 U8528 ( .A1(n15780), .A2(n15745), .ZN(n9383) );
  INV_X1 U8529 ( .A(n9279), .ZN(n7145) );
  NOR2_X1 U8530 ( .A1(n8654), .A2(SI_21_), .ZN(n8653) );
  INV_X1 U8531 ( .A(n8646), .ZN(n7557) );
  INV_X1 U8532 ( .A(n8651), .ZN(n7556) );
  INV_X1 U8533 ( .A(n7559), .ZN(n7558) );
  INV_X1 U8534 ( .A(n9120), .ZN(n8639) );
  NAND2_X1 U8535 ( .A1(n7136), .A2(n7138), .ZN(n7134) );
  OAI21_X1 U8536 ( .B1(n6542), .B2(n7257), .A(n7256), .ZN(n8626) );
  NAND2_X1 U8537 ( .A1(n6542), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7256) );
  AND2_X1 U8538 ( .A1(n8805), .A2(n7411), .ZN(n8621) );
  NAND2_X1 U8539 ( .A1(n8619), .A2(SI_8_), .ZN(n7411) );
  NAND2_X1 U8540 ( .A1(n7567), .A2(n8617), .ZN(n8805) );
  NAND2_X1 U8541 ( .A1(n8829), .A2(n8618), .ZN(n7567) );
  NAND2_X1 U8542 ( .A1(n7912), .A2(n7914), .ZN(n7911) );
  INV_X1 U8543 ( .A(n8418), .ZN(n7380) );
  NOR2_X1 U8544 ( .A1(n8357), .A2(n8339), .ZN(n7400) );
  INV_X1 U8545 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8559) );
  NOR2_X1 U8546 ( .A1(n7373), .A2(n11206), .ZN(n7372) );
  NOR2_X1 U8547 ( .A1(n11245), .A2(n11200), .ZN(n7704) );
  OR2_X1 U8548 ( .A1(n11234), .A2(n11327), .ZN(n11235) );
  INV_X1 U8549 ( .A(n13547), .ZN(n7096) );
  NOR2_X1 U8550 ( .A1(n13498), .A2(n13534), .ZN(n6892) );
  AOI21_X1 U8551 ( .B1(n13498), .B2(n6895), .A(n6755), .ZN(n6893) );
  INV_X1 U8552 ( .A(n6895), .ZN(n6894) );
  NAND2_X1 U8553 ( .A1(n13557), .A2(n13558), .ZN(n13580) );
  NAND2_X1 U8554 ( .A1(n8116), .A2(n9957), .ZN(n8521) );
  INV_X1 U8555 ( .A(n8507), .ZN(n8116) );
  NOR2_X1 U8556 ( .A1(n7949), .A2(n12860), .ZN(n7948) );
  INV_X1 U8557 ( .A(n7950), .ZN(n7949) );
  INV_X1 U8558 ( .A(n12860), .ZN(n7947) );
  OR2_X1 U8559 ( .A1(n13710), .A2(n13693), .ZN(n13112) );
  NAND2_X1 U8560 ( .A1(n12971), .A2(n13106), .ZN(n7870) );
  NAND2_X1 U8561 ( .A1(n8113), .A2(n6771), .ZN(n8491) );
  INV_X1 U8562 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n7328) );
  XNOR2_X1 U8563 ( .A(n13710), .B(n13720), .ZN(n13702) );
  OR2_X1 U8564 ( .A1(n13948), .A2(n13731), .ZN(n13106) );
  AND2_X1 U8565 ( .A1(n8112), .A2(n7330), .ZN(n7329) );
  INV_X1 U8566 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n7330) );
  INV_X1 U8567 ( .A(n8451), .ZN(n8113) );
  INV_X1 U8568 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n11480) );
  INV_X1 U8569 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n7323) );
  INV_X1 U8570 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8103) );
  INV_X1 U8571 ( .A(n8209), .ZN(n8104) );
  INV_X1 U8572 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n8189) );
  NAND2_X1 U8573 ( .A1(n13422), .A2(n13654), .ZN(n13120) );
  NAND2_X1 U8574 ( .A1(n6922), .A2(n13678), .ZN(n6921) );
  NAND2_X1 U8575 ( .A1(n6961), .A2(n6960), .ZN(n13123) );
  AND2_X1 U8576 ( .A1(n13739), .A2(n13741), .ZN(n12853) );
  NOR2_X1 U8577 ( .A1(n13750), .A2(n7078), .ZN(n7076) );
  INV_X1 U8578 ( .A(n12889), .ZN(n13083) );
  AND2_X1 U8579 ( .A1(n13371), .A2(n13801), .ZN(n12890) );
  AND2_X1 U8580 ( .A1(n12526), .A2(n13060), .ZN(n7160) );
  NOR2_X1 U8581 ( .A1(n13041), .A2(n7940), .ZN(n7939) );
  INV_X1 U8582 ( .A(n11633), .ZN(n7940) );
  NAND2_X1 U8583 ( .A1(n11634), .A2(n11633), .ZN(n11635) );
  INV_X1 U8584 ( .A(n8050), .ZN(n7695) );
  NAND2_X1 U8585 ( .A1(n8477), .A2(n8045), .ZN(n8046) );
  NOR2_X1 U8586 ( .A1(n7003), .A2(n7686), .ZN(n7002) );
  INV_X1 U8587 ( .A(n8037), .ZN(n7003) );
  INV_X1 U8588 ( .A(n8034), .ZN(n7000) );
  AND2_X1 U8589 ( .A1(n7685), .A2(n8474), .ZN(n7684) );
  OR2_X1 U8590 ( .A1(n6740), .A2(n7686), .ZN(n7685) );
  INV_X1 U8591 ( .A(n8027), .ZN(n6968) );
  NOR2_X1 U8592 ( .A1(n7663), .A2(n6967), .ZN(n6966) );
  NOR2_X1 U8593 ( .A1(n8359), .A2(n6968), .ZN(n6967) );
  AOI21_X1 U8594 ( .B1(n7662), .B2(n7664), .A(n6754), .ZN(n7660) );
  INV_X1 U8595 ( .A(n7676), .ZN(n7675) );
  OAI21_X1 U8596 ( .B1(P1_DATAO_REG_13__SCAN_IN), .B2(n10651), .A(n8023), .ZN(
        n7676) );
  INV_X1 U8597 ( .A(n7682), .ZN(n7681) );
  OAI21_X1 U8598 ( .B1(n8015), .B2(n7683), .A(n8265), .ZN(n7682) );
  INV_X1 U8599 ( .A(n8016), .ZN(n7683) );
  INV_X1 U8600 ( .A(n8233), .ZN(n7666) );
  NAND2_X1 U8601 ( .A1(n6972), .A2(n6640), .ZN(n7667) );
  NAND2_X1 U8602 ( .A1(n6973), .A2(n6975), .ZN(n6971) );
  INV_X1 U8603 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n8593) );
  AND2_X1 U8604 ( .A1(n14332), .A2(n9433), .ZN(n7018) );
  INV_X1 U8605 ( .A(n14031), .ZN(n7032) );
  XNOR2_X1 U8606 ( .A(n10413), .B(n6802), .ZN(n10427) );
  INV_X1 U8607 ( .A(n9539), .ZN(n6866) );
  AOI21_X1 U8608 ( .B1(n7030), .B2(n7033), .A(n6704), .ZN(n7029) );
  NOR2_X1 U8609 ( .A1(n14130), .A2(n14132), .ZN(n12790) );
  NAND2_X1 U8610 ( .A1(n9784), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n9808) );
  OR2_X1 U8611 ( .A1(n9773), .A2(n9452), .ZN(n9774) );
  NAND2_X1 U8612 ( .A1(n6575), .A2(n14522), .ZN(n7754) );
  NAND2_X1 U8613 ( .A1(n9451), .A2(n6859), .ZN(n9749) );
  NOR2_X1 U8614 ( .A1(n6751), .A2(n6860), .ZN(n6859) );
  NOR2_X1 U8615 ( .A1(n14732), .A2(n14515), .ZN(n7625) );
  AOI21_X1 U8616 ( .B1(n7116), .B2(n7751), .A(n6627), .ZN(n7115) );
  OAI21_X1 U8617 ( .B1(n9705), .B2(n7751), .A(n14561), .ZN(n7750) );
  INV_X1 U8618 ( .A(n9832), .ZN(n7886) );
  OR2_X1 U8619 ( .A1(n7887), .A2(n7886), .ZN(n7885) );
  NAND2_X1 U8620 ( .A1(n6861), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9699) );
  NAND2_X1 U8621 ( .A1(n7287), .A2(n7289), .ZN(n7286) );
  INV_X1 U8622 ( .A(n6861), .ZN(n9681) );
  OR2_X1 U8623 ( .A1(n14823), .A2(n14653), .ZN(n9825) );
  AND2_X1 U8624 ( .A1(n12319), .A2(n9820), .ZN(n7898) );
  NAND2_X1 U8625 ( .A1(n9448), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n9599) );
  INV_X1 U8626 ( .A(n9584), .ZN(n9448) );
  NAND2_X1 U8627 ( .A1(n6853), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n9617) );
  INV_X1 U8628 ( .A(n9599), .ZN(n6853) );
  NAND2_X1 U8629 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n9539) );
  AOI22_X1 U8630 ( .A1(n14215), .A2(n12114), .B1(n6802), .B2(n14214), .ZN(
        n9523) );
  AND2_X1 U8631 ( .A1(n11861), .A2(n9433), .ZN(n10371) );
  INV_X1 U8632 ( .A(n10490), .ZN(n10478) );
  AND2_X1 U8633 ( .A1(n14548), .A2(n7623), .ZN(n14490) );
  INV_X1 U8634 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n9651) );
  INV_X1 U8635 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n9416) );
  INV_X1 U8636 ( .A(n12637), .ZN(n7731) );
  OAI21_X1 U8637 ( .B1(n9267), .B2(n6568), .A(n6692), .ZN(n7246) );
  MUX2_X1 U8638 ( .A(n9346), .B(n9345), .S(n9344), .Z(n9405) );
  NOR2_X1 U8639 ( .A1(n15122), .A2(n7494), .ZN(n15132) );
  AND2_X1 U8640 ( .A1(n15123), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7494) );
  OR2_X1 U8641 ( .A1(n15462), .A2(n15181), .ZN(n15165) );
  NOR2_X1 U8642 ( .A1(n12739), .A2(n7635), .ZN(n7634) );
  NAND2_X1 U8643 ( .A1(n12736), .A2(n7638), .ZN(n7637) );
  INV_X1 U8644 ( .A(n12738), .ZN(n7638) );
  NAND2_X1 U8645 ( .A1(n15209), .A2(n15210), .ZN(n12735) );
  NAND2_X1 U8646 ( .A1(n15493), .A2(n7833), .ZN(n7832) );
  NOR2_X1 U8647 ( .A1(n15500), .A2(n15507), .ZN(n7833) );
  NOR2_X1 U8648 ( .A1(n15318), .A2(n15305), .ZN(n6911) );
  AND2_X1 U8649 ( .A1(n12694), .A2(n12691), .ZN(n7419) );
  AND2_X1 U8650 ( .A1(n8745), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9055) );
  INV_X1 U8651 ( .A(n9057), .ZN(n8745) );
  INV_X1 U8652 ( .A(n12713), .ZN(n15369) );
  NOR2_X1 U8653 ( .A1(n7632), .A2(n7015), .ZN(n7014) );
  INV_X1 U8654 ( .A(n11526), .ZN(n7015) );
  NAND2_X1 U8655 ( .A1(n6702), .A2(n11520), .ZN(n7815) );
  INV_X1 U8656 ( .A(n6904), .ZN(n6903) );
  NAND2_X1 U8657 ( .A1(n11541), .A2(n11521), .ZN(n6904) );
  NAND2_X1 U8658 ( .A1(n15231), .A2(n7827), .ZN(n15195) );
  INV_X1 U8659 ( .A(n15405), .ZN(n15408) );
  OR2_X1 U8660 ( .A1(n12605), .A2(n12604), .ZN(n12606) );
  NAND2_X1 U8661 ( .A1(n12611), .A2(n12610), .ZN(n12712) );
  NAND2_X1 U8662 ( .A1(n11950), .A2(n6907), .ZN(n12031) );
  AND2_X2 U8663 ( .A1(n11506), .A2(n9383), .ZN(n15429) );
  AND2_X1 U8664 ( .A1(n11502), .A2(n11501), .ZN(n15739) );
  INV_X1 U8665 ( .A(n9332), .ZN(n7157) );
  INV_X1 U8666 ( .A(n7153), .ZN(n7152) );
  OAI21_X1 U8667 ( .B1(n8673), .B2(n7154), .A(n8675), .ZN(n7153) );
  INV_X1 U8668 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9342) );
  AND2_X1 U8669 ( .A1(n7146), .A2(n6742), .ZN(n7143) );
  XNOR2_X1 U8670 ( .A(n8664), .B(SI_25_), .ZN(n9279) );
  NAND2_X1 U8671 ( .A1(n6984), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8716) );
  INV_X1 U8672 ( .A(n8715), .ZN(n6985) );
  INV_X1 U8673 ( .A(n9366), .ZN(n7236) );
  OAI21_X1 U8674 ( .B1(n9099), .B2(n7558), .A(n7555), .ZN(n9186) );
  NAND2_X1 U8675 ( .A1(n9148), .A2(n9078), .ZN(n7406) );
  NOR2_X1 U8676 ( .A1(n9065), .A2(n8638), .ZN(n9116) );
  NAND2_X1 U8677 ( .A1(n8636), .A2(n10661), .ZN(n9118) );
  OAI21_X1 U8678 ( .B1(n6542), .B2(n10571), .A(n7568), .ZN(n8614) );
  NAND2_X1 U8679 ( .A1(n6541), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7568) );
  INV_X1 U8680 ( .A(n8926), .ZN(n8946) );
  NAND4_X1 U8681 ( .A1(n15661), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(n7125), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n7124) );
  NAND4_X1 U8682 ( .A1(n15147), .A2(n7128), .A3(P3_ADDR_REG_19__SCAN_IN), .A4(
        n7127), .ZN(n7126) );
  INV_X1 U8683 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7128) );
  NAND2_X1 U8684 ( .A1(n10561), .A2(n6653), .ZN(n7760) );
  INV_X1 U8685 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7759) );
  NAND2_X1 U8686 ( .A1(n7760), .A2(n15035), .ZN(n7056) );
  NAND2_X1 U8687 ( .A1(n10550), .A2(n10543), .ZN(n10814) );
  NAND2_X1 U8688 ( .A1(n10835), .A2(n10834), .ZN(n10845) );
  OR2_X1 U8689 ( .A1(n10832), .A2(n10831), .ZN(n10835) );
  OR2_X1 U8690 ( .A1(n11620), .A2(n11619), .ZN(n11622) );
  INV_X1 U8691 ( .A(n7934), .ZN(n7933) );
  INV_X1 U8692 ( .A(n12063), .ZN(n7932) );
  NAND2_X1 U8693 ( .A1(n13347), .A2(n13348), .ZN(n8515) );
  OR2_X1 U8694 ( .A1(n6548), .A2(n15962), .ZN(n8227) );
  NAND2_X1 U8695 ( .A1(n12193), .A2(n12194), .ZN(n13297) );
  NOR2_X1 U8696 ( .A1(n7995), .A2(n7385), .ZN(n7384) );
  INV_X1 U8697 ( .A(n7387), .ZN(n7385) );
  INV_X1 U8698 ( .A(n8298), .ZN(n7389) );
  NAND2_X1 U8699 ( .A1(n7386), .A2(n7387), .ZN(n13331) );
  OR2_X1 U8700 ( .A1(n12193), .A2(n7389), .ZN(n7386) );
  NAND2_X1 U8701 ( .A1(n7937), .A2(n11661), .ZN(n7934) );
  NAND2_X1 U8702 ( .A1(n8109), .A2(n7318), .ZN(n8368) );
  INV_X1 U8703 ( .A(n6994), .ZN(n6993) );
  NAND3_X1 U8704 ( .A1(n6989), .A2(n6991), .A3(n6992), .ZN(n6988) );
  NOR2_X1 U8705 ( .A1(n6994), .A2(n7183), .ZN(n6989) );
  NAND2_X1 U8706 ( .A1(n13130), .A2(n6629), .ZN(n6991) );
  AND2_X1 U8707 ( .A1(n12993), .A2(n7996), .ZN(n12963) );
  NOR2_X1 U8708 ( .A1(n12966), .A2(n6764), .ZN(n12967) );
  NOR2_X1 U8709 ( .A1(n12965), .A2(n13616), .ZN(n12966) );
  AND2_X1 U8710 ( .A1(n12945), .A2(n12944), .ZN(n13624) );
  NAND2_X1 U8711 ( .A1(n8151), .A2(n6659), .ZN(n6909) );
  INV_X1 U8712 ( .A(n7333), .ZN(n11171) );
  OAI21_X1 U8713 ( .B1(n7336), .B2(n7335), .A(n7334), .ZN(n7333) );
  XNOR2_X1 U8714 ( .A(n11186), .B(n7100), .ZN(n11184) );
  NAND2_X1 U8715 ( .A1(n11154), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n11289) );
  NAND2_X1 U8716 ( .A1(n11153), .A2(n11185), .ZN(n11287) );
  NAND2_X1 U8717 ( .A1(n7582), .A2(n7090), .ZN(n11255) );
  NAND2_X1 U8718 ( .A1(n11252), .A2(n7091), .ZN(n7090) );
  INV_X1 U8719 ( .A(n11192), .ZN(n7091) );
  NAND2_X1 U8720 ( .A1(n7366), .A2(n7370), .ZN(n11248) );
  NAND2_X1 U8721 ( .A1(n11297), .A2(n7372), .ZN(n7366) );
  NAND2_X1 U8722 ( .A1(n6767), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n11338) );
  NAND2_X1 U8723 ( .A1(n7357), .A2(n7356), .ZN(n11334) );
  AOI21_X1 U8724 ( .B1(n7362), .B2(n7365), .A(n7358), .ZN(n7357) );
  AND2_X1 U8725 ( .A1(n7363), .A2(n11224), .ZN(n7362) );
  NAND2_X1 U8726 ( .A1(n7099), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7098) );
  NAND2_X1 U8727 ( .A1(n11874), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n12142) );
  NAND2_X1 U8728 ( .A1(n7355), .A2(n7354), .ZN(n7353) );
  INV_X1 U8729 ( .A(n12148), .ZN(n7355) );
  INV_X1 U8730 ( .A(n12147), .ZN(n7354) );
  NAND2_X1 U8731 ( .A1(n13465), .A2(n6766), .ZN(n7699) );
  NAND2_X1 U8732 ( .A1(n13471), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n13493) );
  OAI211_X1 U8733 ( .C1(n13489), .C2(n6894), .A(n6893), .B(n6887), .ZN(n13519)
         );
  NAND2_X1 U8734 ( .A1(n13489), .A2(n6892), .ZN(n6887) );
  NAND2_X1 U8735 ( .A1(n13514), .A2(n13513), .ZN(n13539) );
  NOR2_X1 U8736 ( .A1(n13568), .A2(n7251), .ZN(n13571) );
  NOR2_X1 U8737 ( .A1(n13556), .A2(n13803), .ZN(n7251) );
  NOR2_X1 U8738 ( .A1(n13571), .A2(n13570), .ZN(n13590) );
  XNOR2_X1 U8739 ( .A(n13580), .B(n13570), .ZN(n13582) );
  NAND2_X1 U8740 ( .A1(n7344), .A2(n6739), .ZN(n7340) );
  NOR2_X1 U8741 ( .A1(n7343), .A2(n13561), .ZN(n7342) );
  OR2_X1 U8742 ( .A1(n8521), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8523) );
  NAND2_X1 U8743 ( .A1(n7068), .A2(n7067), .ZN(n13664) );
  AOI21_X1 U8744 ( .B1(n6562), .B2(n7071), .A(n6679), .ZN(n7067) );
  AOI21_X1 U8745 ( .B1(n7869), .B2(n7868), .A(n7867), .ZN(n7866) );
  INV_X1 U8746 ( .A(n13106), .ZN(n7868) );
  INV_X1 U8747 ( .A(n13112), .ZN(n7867) );
  NAND2_X1 U8748 ( .A1(n8113), .A2(n7329), .ZN(n8480) );
  NAND2_X1 U8749 ( .A1(n8111), .A2(n6596), .ZN(n8435) );
  INV_X1 U8750 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n7320) );
  AND2_X1 U8751 ( .A1(n13752), .A2(n13083), .ZN(n13777) );
  AOI21_X1 U8752 ( .B1(n13792), .B2(n6551), .A(n8398), .ZN(n13773) );
  NAND2_X1 U8753 ( .A1(n8111), .A2(n8110), .ZN(n8409) );
  NAND2_X1 U8754 ( .A1(n8109), .A2(n6595), .ZN(n8374) );
  INV_X1 U8755 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n7317) );
  OR2_X1 U8756 ( .A1(n8374), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8394) );
  NAND2_X1 U8757 ( .A1(n8109), .A2(n8108), .ZN(n8351) );
  NAND2_X1 U8758 ( .A1(n8106), .A2(n7324), .ZN(n8333) );
  AND2_X1 U8759 ( .A1(n7325), .A2(n8107), .ZN(n7324) );
  NAND2_X1 U8760 ( .A1(n8106), .A2(n6743), .ZN(n8307) );
  NAND2_X1 U8761 ( .A1(n8106), .A2(n11480), .ZN(n8289) );
  OR2_X1 U8762 ( .A1(n8257), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8273) );
  AND2_X1 U8763 ( .A1(n13039), .A2(n13038), .ZN(n13037) );
  INV_X1 U8764 ( .A(n13037), .ZN(n11429) );
  NAND2_X1 U8765 ( .A1(n11584), .A2(n12973), .ZN(n11631) );
  NAND2_X1 U8766 ( .A1(n8104), .A2(n6609), .ZN(n8240) );
  NAND2_X1 U8767 ( .A1(n8104), .A2(n8103), .ZN(n8224) );
  NAND2_X1 U8768 ( .A1(n11452), .A2(n13022), .ZN(n11421) );
  NAND2_X1 U8769 ( .A1(n12937), .A2(n12936), .ZN(n12959) );
  NOR2_X1 U8770 ( .A1(n13624), .A2(n13623), .ZN(n13912) );
  AOI21_X1 U8771 ( .B1(n12868), .B2(n13649), .A(n6686), .ZN(n7977) );
  INV_X1 U8772 ( .A(n12926), .ZN(n7976) );
  AND2_X1 U8773 ( .A1(n13635), .A2(n6929), .ZN(n6928) );
  OR2_X1 U8774 ( .A1(n13649), .A2(n6930), .ZN(n6929) );
  AND2_X1 U8775 ( .A1(n8415), .A2(n8414), .ZN(n13759) );
  AND2_X1 U8776 ( .A1(n13092), .A2(n13091), .ZN(n13755) );
  OR2_X1 U8777 ( .A1(n7963), .A2(n12984), .ZN(n7957) );
  AND2_X1 U8778 ( .A1(n7854), .A2(n6916), .ZN(n6915) );
  NAND2_X1 U8779 ( .A1(n12885), .A2(n7857), .ZN(n6914) );
  AOI21_X1 U8780 ( .B1(n7857), .B2(n7859), .A(n7855), .ZN(n7854) );
  AND2_X1 U8781 ( .A1(n13078), .A2(n13079), .ZN(n13797) );
  NAND2_X1 U8782 ( .A1(n11803), .A2(n12979), .ZN(n11837) );
  INV_X1 U8783 ( .A(n11835), .ZN(n11803) );
  INV_X1 U8784 ( .A(n7941), .ZN(n12070) );
  AOI21_X1 U8785 ( .B1(n11837), .B2(n11805), .A(n7944), .ZN(n7941) );
  OR2_X1 U8786 ( .A1(n8550), .A2(n8549), .ZN(n10933) );
  XNOR2_X1 U8787 ( .A(n8094), .B(n8086), .ZN(n8092) );
  NAND2_X1 U8788 ( .A1(n8096), .A2(n8095), .ZN(n11372) );
  AND2_X1 U8789 ( .A1(n8120), .A2(n8064), .ZN(n7952) );
  NAND2_X2 U8790 ( .A1(n7163), .A2(n7162), .ZN(n7061) );
  NAND2_X1 U8791 ( .A1(n8064), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7162) );
  XNOR2_X1 U8792 ( .A(n8046), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n8488) );
  NAND2_X1 U8793 ( .A1(n8098), .A2(n8073), .ZN(n8102) );
  AND2_X1 U8794 ( .A1(n8328), .A2(n8072), .ZN(n8098) );
  NAND2_X1 U8795 ( .A1(n7677), .A2(n8022), .ZN(n8342) );
  XNOR2_X1 U8796 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8300) );
  OR2_X1 U8797 ( .A1(n8220), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n8235) );
  NAND2_X1 U8798 ( .A1(n7250), .A2(n8184), .ZN(n8202) );
  NAND2_X1 U8799 ( .A1(n6955), .A2(n8004), .ZN(n8181) );
  NAND2_X1 U8800 ( .A1(n10525), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8004) );
  INV_X1 U8801 ( .A(n8168), .ZN(n7659) );
  XNOR2_X1 U8802 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8180) );
  OR2_X1 U8803 ( .A1(n14030), .A2(n7541), .ZN(n7540) );
  INV_X1 U8804 ( .A(n14118), .ZN(n7541) );
  AND2_X1 U8805 ( .A1(n6732), .A2(n7036), .ZN(n7035) );
  INV_X1 U8806 ( .A(n14209), .ZN(n12471) );
  NAND2_X1 U8807 ( .A1(n14032), .A2(n14031), .ZN(n12782) );
  NAND2_X1 U8808 ( .A1(n9449), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9656) );
  INV_X1 U8809 ( .A(n9641), .ZN(n9449) );
  OR2_X1 U8810 ( .A1(n9656), .A2(n11607), .ZN(n9666) );
  OAI21_X1 U8811 ( .B1(n10470), .B2(n7547), .A(n7545), .ZN(n12760) );
  NAND2_X1 U8812 ( .A1(n9739), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n9773) );
  INV_X1 U8813 ( .A(n9749), .ZN(n9739) );
  NAND2_X1 U8814 ( .A1(n9451), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9748) );
  AND2_X1 U8815 ( .A1(n10443), .A2(n10438), .ZN(n7548) );
  AND2_X1 U8816 ( .A1(n6813), .A2(n11551), .ZN(n7171) );
  XNOR2_X1 U8817 ( .A(n6814), .B(n11860), .ZN(n6813) );
  NAND2_X1 U8818 ( .A1(n7184), .A2(n10370), .ZN(n10401) );
  INV_X1 U8819 ( .A(n9861), .ZN(n10329) );
  AND4_X1 U8820 ( .A1(n9687), .A2(n9686), .A3(n9685), .A4(n9684), .ZN(n14089)
         );
  NAND2_X1 U8821 ( .A1(n14236), .A2(n14237), .ZN(n14235) );
  NOR2_X1 U8822 ( .A1(n7304), .A2(n6667), .ZN(n7303) );
  NOR2_X1 U8823 ( .A1(n11056), .A2(n7305), .ZN(n7304) );
  OR2_X1 U8824 ( .A1(n14277), .A2(n7305), .ZN(n7301) );
  OR2_X1 U8825 ( .A1(n11112), .A2(n11113), .ZN(n11110) );
  OR2_X1 U8826 ( .A1(n11119), .A2(n11118), .ZN(n11116) );
  NAND2_X1 U8827 ( .A1(n11116), .A2(n7309), .ZN(n15889) );
  OR2_X1 U8828 ( .A1(n11606), .A2(n11605), .ZN(n11693) );
  OR2_X1 U8829 ( .A1(n11599), .A2(n11600), .ZN(n11700) );
  NAND2_X1 U8830 ( .A1(n14321), .A2(n7298), .ZN(n14323) );
  AND2_X1 U8831 ( .A1(n14436), .A2(n14415), .ZN(n14395) );
  OR2_X1 U8832 ( .A1(n14457), .A2(n12795), .ZN(n7990) );
  NAND2_X1 U8833 ( .A1(n14548), .A2(n6655), .ZN(n14451) );
  OR2_X2 U8834 ( .A1(n14451), .A2(n14710), .ZN(n14452) );
  OR2_X1 U8835 ( .A1(n14481), .A2(n14469), .ZN(n14482) );
  AND2_X1 U8836 ( .A1(n14531), .A2(n9736), .ZN(n14499) );
  OR2_X1 U8837 ( .A1(n14499), .A2(n14498), .ZN(n14501) );
  NAND2_X1 U8838 ( .A1(n14548), .A2(n7625), .ZN(n14513) );
  AOI21_X1 U8839 ( .B1(n9726), .B2(n14503), .A(n8003), .ZN(n14533) );
  NOR3_X1 U8840 ( .A1(n14560), .A2(n14504), .A3(n14503), .ZN(n14544) );
  NAND2_X1 U8841 ( .A1(n9450), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9712) );
  INV_X1 U8842 ( .A(n9699), .ZN(n9450) );
  OR2_X1 U8843 ( .A1(n9712), .A2(n9711), .ZN(n9721) );
  NAND2_X1 U8844 ( .A1(n14596), .A2(n9832), .ZN(n14573) );
  OR2_X1 U8845 ( .A1(n9689), .A2(n14625), .ZN(n14606) );
  NAND2_X1 U8846 ( .A1(n9867), .A2(n6749), .ZN(n14599) );
  NAND2_X1 U8847 ( .A1(n6852), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9630) );
  INV_X1 U8848 ( .A(n9617), .ZN(n6852) );
  AOI21_X1 U8849 ( .B1(n9608), .B2(n7113), .A(n9607), .ZN(n7110) );
  NAND2_X1 U8850 ( .A1(n11966), .A2(n9565), .ZN(n12123) );
  NAND2_X1 U8851 ( .A1(n7615), .A2(n15932), .ZN(n12130) );
  NAND2_X1 U8852 ( .A1(n7891), .A2(n7889), .ZN(n6849) );
  NAND2_X1 U8853 ( .A1(n12178), .A2(n12181), .ZN(n12177) );
  AOI21_X1 U8854 ( .B1(n11990), .B2(n11991), .A(n11992), .ZN(n7892) );
  OR2_X1 U8855 ( .A1(n10482), .A2(n10400), .ZN(n10488) );
  OAI21_X1 U8856 ( .B1(n10371), .B2(n7021), .A(n14332), .ZN(n11968) );
  INV_X1 U8857 ( .A(n14344), .ZN(n7743) );
  NAND2_X1 U8858 ( .A1(n7131), .A2(n10320), .ZN(n10367) );
  NAND2_X1 U8859 ( .A1(n13258), .A2(n10335), .ZN(n9806) );
  AND2_X1 U8860 ( .A1(n14384), .A2(n14383), .ZN(n14689) );
  NOR2_X1 U8861 ( .A1(n9793), .A2(n10630), .ZN(n6804) );
  NAND2_X1 U8862 ( .A1(n12251), .A2(n6802), .ZN(n12252) );
  AND2_X1 U8863 ( .A1(n11021), .A2(n11020), .ZN(n10492) );
  INV_X1 U8864 ( .A(n9759), .ZN(n7229) );
  INV_X1 U8865 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7768) );
  INV_X1 U8866 ( .A(n9428), .ZN(n7769) );
  CLKBUF_X1 U8867 ( .A(n9509), .Z(n9510) );
  INV_X1 U8868 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9494) );
  OR2_X1 U8869 ( .A1(n12636), .A2(n12637), .ZN(n7733) );
  INV_X1 U8870 ( .A(n12568), .ZN(n12570) );
  NAND2_X1 U8871 ( .A1(n14836), .A2(n14837), .ZN(n11915) );
  NAND2_X1 U8872 ( .A1(n6697), .A2(n11351), .ZN(n6938) );
  INV_X1 U8873 ( .A(n11350), .ZN(n6939) );
  NAND2_X1 U8874 ( .A1(n8743), .A2(n8742), .ZN(n9029) );
  INV_X1 U8875 ( .A(n9007), .ZN(n8743) );
  NAND2_X1 U8876 ( .A1(n8744), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9057) );
  INV_X1 U8877 ( .A(n9029), .ZN(n8744) );
  INV_X1 U8878 ( .A(n7723), .ZN(n7722) );
  NAND2_X1 U8879 ( .A1(n6948), .A2(n6584), .ZN(n7721) );
  OAI21_X1 U8880 ( .B1(n7725), .B2(n7724), .A(n13193), .ZN(n7723) );
  NAND2_X1 U8881 ( .A1(n14942), .A2(n14943), .ZN(n14941) );
  XNOR2_X1 U8882 ( .A(n7212), .B(n13233), .ZN(n10981) );
  AND2_X1 U8883 ( .A1(n11651), .A2(n11650), .ZN(n11894) );
  INV_X1 U8884 ( .A(n9270), .ZN(n8750) );
  NOR2_X1 U8885 ( .A1(n14898), .A2(n7719), .ZN(n7718) );
  INV_X1 U8886 ( .A(n14927), .ZN(n7719) );
  INV_X1 U8887 ( .A(n9317), .ZN(n6982) );
  AND2_X1 U8888 ( .A1(n7597), .A2(n6979), .ZN(n6978) );
  NAND2_X1 U8889 ( .A1(n6980), .A2(n9317), .ZN(n6979) );
  NAND2_X1 U8890 ( .A1(n9337), .A2(n7598), .ZN(n7597) );
  AND2_X1 U8891 ( .A1(n9222), .A2(n9221), .ZN(n13194) );
  AND4_X1 U8892 ( .A1(n8802), .A2(n8801), .A3(n8800), .A4(n8799), .ZN(n14839)
         );
  NAND2_X1 U8893 ( .A1(n10687), .A2(n10686), .ZN(n15689) );
  AOI21_X1 U8894 ( .B1(n15689), .B2(n10736), .A(n10735), .ZN(n10734) );
  NOR2_X1 U8895 ( .A1(n10688), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7486) );
  OR2_X1 U8896 ( .A1(n8946), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n8792) );
  OAI21_X1 U8897 ( .B1(n10734), .B2(n10704), .A(n10703), .ZN(n10716) );
  NAND2_X1 U8898 ( .A1(n8780), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8993) );
  OR2_X1 U8899 ( .A1(n8811), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n8780) );
  NOR2_X1 U8900 ( .A1(n11072), .A2(n6883), .ZN(n6882) );
  INV_X1 U8901 ( .A(n6607), .ZN(n6883) );
  OR2_X1 U8902 ( .A1(n15719), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6873) );
  NAND2_X1 U8903 ( .A1(n15105), .A2(n6770), .ZN(n15109) );
  NOR2_X1 U8904 ( .A1(n15124), .A2(n15125), .ZN(n15134) );
  XNOR2_X1 U8905 ( .A(n15132), .B(n15131), .ZN(n15124) );
  NAND2_X1 U8906 ( .A1(n15462), .A2(n15181), .ZN(n15169) );
  AND2_X1 U8907 ( .A1(n9322), .A2(n15176), .ZN(n15192) );
  AND2_X1 U8908 ( .A1(n15231), .A2(n13225), .ZN(n15216) );
  NAND2_X1 U8909 ( .A1(n9291), .A2(n9290), .ZN(n15222) );
  OR2_X1 U8910 ( .A1(n12486), .A2(n8897), .ZN(n9291) );
  NAND2_X1 U8911 ( .A1(n6911), .A2(n6910), .ZN(n15250) );
  NOR2_X1 U8912 ( .A1(n15488), .A2(n7832), .ZN(n6910) );
  NAND2_X1 U8913 ( .A1(n15290), .A2(n7646), .ZN(n7645) );
  AND2_X1 U8914 ( .A1(n7643), .A2(n15244), .ZN(n7642) );
  NAND2_X1 U8915 ( .A1(n7646), .A2(n7644), .ZN(n7643) );
  OR2_X1 U8916 ( .A1(n7442), .A2(n15289), .ZN(n7441) );
  INV_X1 U8917 ( .A(n7439), .ZN(n7438) );
  OAI21_X1 U8918 ( .B1(n7442), .B2(n7440), .A(n12702), .ZN(n7439) );
  NOR2_X1 U8919 ( .A1(n15302), .A2(n7831), .ZN(n15270) );
  INV_X1 U8920 ( .A(n7833), .ZN(n7831) );
  NOR2_X1 U8921 ( .A1(n15302), .A2(n15507), .ZN(n15286) );
  INV_X1 U8922 ( .A(n6911), .ZN(n15302) );
  NAND2_X1 U8923 ( .A1(n8747), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9159) );
  AND3_X1 U8924 ( .A1(n9097), .A2(n9096), .A3(n9095), .ZN(n15340) );
  NAND2_X1 U8925 ( .A1(n12712), .A2(n12711), .ZN(n15409) );
  AND2_X1 U8926 ( .A1(n15414), .A2(n6592), .ZN(n15363) );
  NAND2_X1 U8927 ( .A1(n15414), .A2(n6566), .ZN(n15377) );
  NAND2_X1 U8928 ( .A1(n15414), .A2(n12742), .ZN(n15385) );
  AND3_X1 U8929 ( .A1(n9075), .A2(n9074), .A3(n9073), .ZN(n15412) );
  OR2_X1 U8930 ( .A1(n8999), .A2(n8998), .ZN(n9007) );
  AND2_X1 U8931 ( .A1(n11950), .A2(n6720), .ZN(n12165) );
  NAND2_X1 U8932 ( .A1(n7658), .A2(n6576), .ZN(n12158) );
  NOR2_X1 U8933 ( .A1(n7421), .A2(n6656), .ZN(n7420) );
  INV_X1 U8934 ( .A(n7423), .ZN(n7421) );
  NAND2_X1 U8935 ( .A1(n8741), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8972) );
  INV_X1 U8936 ( .A(n8824), .ZN(n8741) );
  OR2_X1 U8937 ( .A1(n8972), .A2(n8971), .ZN(n8999) );
  NAND2_X1 U8938 ( .A1(n12010), .A2(n12009), .ZN(n12012) );
  AND2_X1 U8939 ( .A1(n7422), .A2(n7423), .ZN(n12023) );
  XNOR2_X1 U8940 ( .A(n12001), .B(n15014), .ZN(n11959) );
  NAND2_X1 U8941 ( .A1(n11950), .A2(n15821), .ZN(n12029) );
  INV_X1 U8942 ( .A(n7815), .ZN(n7817) );
  NAND2_X1 U8943 ( .A1(n8739), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8822) );
  INV_X1 U8944 ( .A(n8937), .ZN(n8739) );
  AND2_X1 U8945 ( .A1(n10789), .A2(n10676), .ZN(n15426) );
  NAND2_X1 U8946 ( .A1(n7818), .A2(n11520), .ZN(n11748) );
  NAND2_X1 U8947 ( .A1(n7820), .A2(n7819), .ZN(n7818) );
  INV_X1 U8948 ( .A(n11519), .ZN(n7820) );
  OR2_X1 U8949 ( .A1(n6904), .A2(n15435), .ZN(n11533) );
  AND2_X1 U8950 ( .A1(n10789), .A2(n8855), .ZN(n15746) );
  NAND2_X1 U8951 ( .A1(n6540), .A2(n6539), .ZN(n11434) );
  INV_X1 U8952 ( .A(n15746), .ZN(n15411) );
  NAND2_X1 U8953 ( .A1(n7009), .A2(n15754), .ZN(n12741) );
  NAND2_X1 U8954 ( .A1(n7011), .A2(n7010), .ZN(n7009) );
  NAND2_X1 U8955 ( .A1(n12737), .A2(n6652), .ZN(n7010) );
  INV_X1 U8956 ( .A(n7636), .ZN(n7011) );
  INV_X1 U8957 ( .A(n15265), .ZN(n15493) );
  AND2_X1 U8958 ( .A1(n10943), .A2(n10942), .ZN(n15813) );
  NAND2_X1 U8959 ( .A1(n7144), .A2(n7143), .ZN(n9289) );
  NAND2_X1 U8960 ( .A1(n7144), .A2(n6742), .ZN(n9287) );
  INV_X1 U8961 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9367) );
  NAND2_X1 U8962 ( .A1(n7572), .A2(n7569), .ZN(n9263) );
  NAND2_X1 U8963 ( .A1(n7237), .A2(n7234), .ZN(n10788) );
  NOR2_X1 U8964 ( .A1(n7236), .A2(n7235), .ZN(n7234) );
  OR2_X1 U8965 ( .A1(n8716), .A2(n7238), .ZN(n7237) );
  NOR2_X1 U8966 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n7235) );
  NAND2_X1 U8967 ( .A1(n7728), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8706) );
  NAND2_X1 U8968 ( .A1(n8689), .A2(n8705), .ZN(n6986) );
  NAND2_X1 U8969 ( .A1(n8714), .A2(n8710), .ZN(n9079) );
  NAND2_X1 U8970 ( .A1(n7201), .A2(n9063), .ZN(n9047) );
  OAI211_X1 U8971 ( .C1(n7416), .C2(n7417), .A(n8632), .B(n7415), .ZN(n9036)
         );
  NAND2_X1 U8972 ( .A1(n6791), .A2(n8634), .ZN(n9038) );
  INV_X1 U8973 ( .A(n8627), .ZN(n6786) );
  OAI21_X1 U8974 ( .B1(n6542), .B2(P2_DATAO_REG_10__SCAN_IN), .A(n7196), .ZN(
        n8988) );
  NAND2_X1 U8975 ( .A1(n6542), .A2(n10658), .ZN(n7196) );
  OAI21_X1 U8976 ( .B1(SI_10_), .B2(n8987), .A(n9012), .ZN(n8989) );
  NAND2_X1 U8977 ( .A1(n8790), .A2(n8789), .ZN(n8830) );
  INV_X1 U8978 ( .A(n8787), .ZN(n8789) );
  NOR2_X1 U8979 ( .A1(n8926), .A2(n7495), .ZN(n15684) );
  OAI22_X1 U8980 ( .A1(n8925), .A2(n7496), .B1(P1_IR_REG_4__SCAN_IN), .B2(
        P1_IR_REG_31__SCAN_IN), .ZN(n7495) );
  NAND2_X1 U8981 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n7496) );
  NAND3_X1 U8982 ( .A1(n8603), .A2(n8876), .A3(n8602), .ZN(n7123) );
  NAND2_X1 U8983 ( .A1(n8598), .A2(SI_1_), .ZN(n8874) );
  NAND2_X1 U8984 ( .A1(n7519), .A2(n10557), .ZN(n10562) );
  NAND2_X1 U8985 ( .A1(n16029), .A2(n16030), .ZN(n7519) );
  AND2_X1 U8986 ( .A1(n12296), .A2(n15901), .ZN(n7047) );
  NAND2_X1 U8987 ( .A1(n7508), .A2(n7512), .ZN(n15644) );
  NAND2_X1 U8988 ( .A1(n13297), .A2(n8298), .ZN(n13298) );
  NAND2_X1 U8989 ( .A1(n13311), .A2(n13310), .ZN(n13309) );
  AND4_X1 U8990 ( .A1(n8246), .A2(n8245), .A3(n8244), .A4(n8243), .ZN(n11851)
         );
  NAND2_X1 U8991 ( .A1(n6537), .A2(n7335), .ZN(n8154) );
  NAND2_X1 U8992 ( .A1(n7910), .A2(n7912), .ZN(n13318) );
  OR2_X1 U8993 ( .A1(n13311), .A2(n7914), .ZN(n7910) );
  NAND2_X1 U8994 ( .A1(n7402), .A2(n7908), .ZN(n11365) );
  NAND2_X1 U8995 ( .A1(n7909), .A2(n8216), .ZN(n7402) );
  OR2_X1 U8996 ( .A1(n7905), .A2(n7927), .ZN(n7393) );
  NAND2_X1 U8997 ( .A1(n6621), .A2(n13347), .ZN(n7919) );
  NAND2_X1 U8998 ( .A1(n13347), .A2(n13693), .ZN(n7920) );
  INV_X1 U8999 ( .A(n13456), .ZN(n12198) );
  INV_X1 U9000 ( .A(n7918), .ZN(n7917) );
  NAND2_X1 U9001 ( .A1(n10154), .A2(n10155), .ZN(n13395) );
  NAND2_X1 U9002 ( .A1(n7396), .A2(n7394), .ZN(n8401) );
  AOI21_X1 U9003 ( .B1(n7397), .B2(n7927), .A(n7395), .ZN(n7394) );
  NAND2_X1 U9004 ( .A1(n13417), .A2(n13416), .ZN(n13415) );
  OR2_X1 U9005 ( .A1(n11363), .A2(n7934), .ZN(n11660) );
  AND2_X1 U9006 ( .A1(n8568), .A2(n15985), .ZN(n13446) );
  NAND2_X1 U9007 ( .A1(n7401), .A2(n6582), .ZN(n13436) );
  AND2_X1 U9008 ( .A1(n12945), .A2(n12230), .ZN(n13640) );
  NAND2_X1 U9009 ( .A1(n8133), .A2(n8132), .ZN(n13666) );
  INV_X1 U9010 ( .A(n13704), .ZN(n13449) );
  INV_X1 U9011 ( .A(n13772), .ZN(n13743) );
  INV_X1 U9012 ( .A(n13759), .ZN(n13789) );
  INV_X1 U9013 ( .A(n11851), .ZN(n13457) );
  INV_X1 U9014 ( .A(P3_U3897), .ZN(n13463) );
  INV_X1 U9015 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n11165) );
  AND2_X1 U9016 ( .A1(n6615), .A2(n6909), .ZN(n11176) );
  AND2_X1 U9017 ( .A1(n7574), .A2(n11151), .ZN(n11178) );
  NAND2_X1 U9018 ( .A1(n6775), .A2(n11192), .ZN(n11253) );
  NAND2_X1 U9019 ( .A1(n7359), .A2(n7363), .ZN(n11250) );
  NAND2_X1 U9020 ( .A1(n7360), .A2(n7361), .ZN(n7359) );
  AND2_X1 U9021 ( .A1(n7703), .A2(n7702), .ZN(n11244) );
  INV_X1 U9022 ( .A(n7707), .ZN(n7703) );
  NAND2_X1 U9023 ( .A1(n11218), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7702) );
  OAI211_X1 U9024 ( .C1(n7707), .C2(n11218), .A(n7706), .B(n7705), .ZN(n11242)
         );
  OR2_X1 U9025 ( .A1(n7707), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7706) );
  OR2_X1 U9026 ( .A1(n7098), .A2(n7097), .ZN(n11576) );
  OAI22_X1 U9027 ( .A1(n11561), .A2(n11560), .B1(n11559), .B2(n11558), .ZN(
        n11887) );
  INV_X1 U9028 ( .A(n12141), .ZN(n7578) );
  AOI21_X1 U9029 ( .B1(n12141), .B2(n7577), .A(n6780), .ZN(n7576) );
  INV_X1 U9030 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n7577) );
  XNOR2_X1 U9031 ( .A(n7699), .B(n13496), .ZN(n13487) );
  AOI21_X1 U9032 ( .B1(n13487), .B2(P3_REG1_REG_13__SCAN_IN), .A(n7698), .ZN(
        n13491) );
  AND2_X1 U9033 ( .A1(n7699), .A2(n13486), .ZN(n7698) );
  NAND2_X1 U9034 ( .A1(n7094), .A2(n13534), .ZN(n13546) );
  INV_X1 U9035 ( .A(n13527), .ZN(n7094) );
  NOR2_X1 U9036 ( .A1(n13540), .A2(n6565), .ZN(n13562) );
  NAND2_X1 U9037 ( .A1(n13535), .A2(n13536), .ZN(n13538) );
  NAND2_X1 U9038 ( .A1(n13518), .A2(n13517), .ZN(n13533) );
  NAND2_X1 U9039 ( .A1(n7346), .A2(n7347), .ZN(n13563) );
  NAND2_X1 U9040 ( .A1(n13540), .A2(n7348), .ZN(n7346) );
  XNOR2_X1 U9041 ( .A(n13668), .B(n13667), .ZN(n13855) );
  NAND2_X1 U9042 ( .A1(n7069), .A2(n7072), .ZN(n13679) );
  NAND2_X1 U9043 ( .A1(n13684), .A2(n13683), .ZN(n13682) );
  NAND2_X1 U9044 ( .A1(n13694), .A2(n13113), .ZN(n13684) );
  NAND2_X1 U9045 ( .A1(n12858), .A2(n7994), .ZN(n13729) );
  NAND2_X1 U9046 ( .A1(n8408), .A2(n8407), .ZN(n13782) );
  OAI21_X1 U9047 ( .B1(n12523), .B2(n7963), .A(n7959), .ZN(n13809) );
  NAND2_X1 U9048 ( .A1(n7837), .A2(n7835), .ZN(n11834) );
  NAND2_X1 U9049 ( .A1(n7842), .A2(n7838), .ZN(n11632) );
  NAND2_X1 U9050 ( .A1(n11584), .A2(n6564), .ZN(n7838) );
  AND3_X1 U9051 ( .A1(n8143), .A2(n8142), .A3(n8141), .ZN(n16012) );
  INV_X1 U9052 ( .A(n15985), .ZN(n15977) );
  AND2_X1 U9053 ( .A1(n8256), .A2(n8255), .ZN(n11800) );
  INV_X1 U9054 ( .A(n13893), .ZN(n13905) );
  INV_X1 U9055 ( .A(n12959), .ZN(n13914) );
  NAND2_X1 U9056 ( .A1(n8071), .A2(n8070), .ZN(n13927) );
  NAND2_X1 U9057 ( .A1(n12394), .A2(n12935), .ZN(n8071) );
  AOI21_X1 U9058 ( .B1(n13657), .B2(n13833), .A(n13656), .ZN(n13925) );
  OAI21_X1 U9059 ( .B1(n13653), .B2(n13652), .A(n13651), .ZN(n13657) );
  XNOR2_X1 U9060 ( .A(n13648), .B(n13649), .ZN(n13928) );
  AOI21_X1 U9061 ( .B1(n12858), .B2(n7950), .A(n6569), .ZN(n13719) );
  NAND2_X1 U9062 ( .A1(n7848), .A2(n7849), .ZN(n13727) );
  NAND2_X1 U9063 ( .A1(n8434), .A2(n8433), .ZN(n13958) );
  NAND2_X1 U9064 ( .A1(n7853), .A2(n7851), .ZN(n13737) );
  AND2_X1 U9065 ( .A1(n7853), .A2(n13091), .ZN(n13738) );
  NAND2_X1 U9066 ( .A1(n12894), .A2(n13085), .ZN(n7853) );
  NAND2_X1 U9067 ( .A1(n8422), .A2(n8421), .ZN(n13964) );
  NAND2_X1 U9068 ( .A1(n8383), .A2(n8382), .ZN(n13980) );
  NAND2_X1 U9069 ( .A1(n12887), .A2(n7860), .ZN(n7856) );
  NAND2_X1 U9070 ( .A1(n7958), .A2(n7965), .ZN(n13827) );
  NAND2_X1 U9071 ( .A1(n12523), .A2(n7967), .ZN(n7958) );
  NAND2_X1 U9072 ( .A1(n12887), .A2(n12886), .ZN(n13822) );
  OAI21_X1 U9073 ( .B1(n12523), .B2(n12983), .A(n6552), .ZN(n12851) );
  NAND2_X1 U9074 ( .A1(n8318), .A2(n8317), .ZN(n13344) );
  NAND2_X1 U9075 ( .A1(n8288), .A2(n8287), .ZN(n13308) );
  NAND2_X1 U9076 ( .A1(n6932), .A2(n6935), .ZN(n7979) );
  INV_X1 U9077 ( .A(n11800), .ZN(n11853) );
  INV_X1 U9078 ( .A(n11372), .ZN(n8097) );
  INV_X1 U9079 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7954) );
  OR2_X1 U9080 ( .A1(n12947), .A2(n12946), .ZN(n12948) );
  NAND2_X1 U9081 ( .A1(n7693), .A2(n7691), .ZN(n12929) );
  NAND2_X1 U9082 ( .A1(n7693), .A2(n12872), .ZN(n12875) );
  XNOR2_X1 U9083 ( .A(n8519), .B(n8518), .ZN(n12285) );
  NAND2_X1 U9084 ( .A1(n8504), .A2(n8050), .ZN(n8519) );
  NAND2_X1 U9085 ( .A1(n8464), .A2(n8043), .ZN(n8475) );
  NAND2_X1 U9086 ( .A1(n8041), .A2(n8040), .ZN(n8462) );
  NAND2_X1 U9087 ( .A1(n7661), .A2(n8029), .ZN(n8387) );
  NAND2_X1 U9088 ( .A1(n8380), .A2(n8028), .ZN(n7661) );
  NAND2_X1 U9089 ( .A1(n7680), .A2(n8016), .ZN(n8266) );
  NAND2_X1 U9090 ( .A1(n8249), .A2(n8015), .ZN(n7680) );
  OAI21_X1 U9091 ( .B1(n8135), .B2(n7670), .A(n7668), .ZN(n8234) );
  NAND2_X1 U9092 ( .A1(n7673), .A2(n8011), .ZN(n8219) );
  NAND2_X1 U9093 ( .A1(n8135), .A2(n8134), .ZN(n7673) );
  NAND2_X1 U9094 ( .A1(n8008), .A2(n8007), .ZN(n8201) );
  AOI21_X1 U9095 ( .B1(n11150), .B2(n6662), .A(n7710), .ZN(n7709) );
  NOR2_X1 U9096 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n7710) );
  NOR2_X1 U9097 ( .A1(n10481), .A2(n10480), .ZN(n14012) );
  NAND2_X1 U9098 ( .A1(n12476), .A2(n6610), .ZN(n12659) );
  NAND2_X1 U9099 ( .A1(n12476), .A2(n10460), .ZN(n12658) );
  OAI21_X1 U9100 ( .B1(n14032), .B2(n7033), .A(n7030), .ZN(n14129) );
  AND4_X1 U9101 ( .A1(n9635), .A2(n9634), .A3(n9633), .A4(n9632), .ZN(n14066)
         );
  NAND2_X1 U9102 ( .A1(n10470), .A2(n14141), .ZN(n14064) );
  NAND2_X1 U9103 ( .A1(n7022), .A2(n7027), .ZN(n14163) );
  NAND2_X1 U9104 ( .A1(n14073), .A2(n6561), .ZN(n7022) );
  AND2_X1 U9105 ( .A1(n9796), .A2(n9786), .ZN(n14413) );
  INV_X1 U9106 ( .A(n14213), .ZN(n12179) );
  INV_X1 U9107 ( .A(n14211), .ZN(n12336) );
  NAND2_X1 U9108 ( .A1(n7537), .A2(n14071), .ZN(n7536) );
  INV_X1 U9109 ( .A(n14073), .ZN(n7537) );
  OR2_X1 U9110 ( .A1(n10450), .A2(n12086), .ZN(n10415) );
  NAND2_X1 U9111 ( .A1(n12782), .A2(n14030), .ZN(n14120) );
  NAND2_X1 U9112 ( .A1(n12659), .A2(n10465), .ZN(n14143) );
  NAND2_X1 U9113 ( .A1(n12849), .A2(n12771), .ZN(n14156) );
  NAND2_X1 U9114 ( .A1(n12057), .A2(n10438), .ZN(n12348) );
  AND4_X1 U9115 ( .A1(n9545), .A2(n9544), .A3(n9543), .A4(n9542), .ZN(n14104)
         );
  AND4_X1 U9116 ( .A1(n9576), .A2(n9575), .A3(n9574), .A4(n9573), .ZN(n12548)
         );
  OR2_X1 U9117 ( .A1(n14147), .A2(n14636), .ZN(n14185) );
  NAND2_X1 U9118 ( .A1(n7025), .A2(n7023), .ZN(n14175) );
  NAND2_X1 U9119 ( .A1(n7024), .A2(n6623), .ZN(n7023) );
  INV_X1 U9120 ( .A(n7027), .ZN(n7024) );
  NAND2_X1 U9121 ( .A1(n10783), .A2(n10335), .ZN(n7734) );
  NOR2_X1 U9122 ( .A1(n15911), .A2(n7271), .ZN(n10406) );
  NAND2_X1 U9123 ( .A1(n14652), .A2(n7272), .ZN(n7271) );
  NAND2_X1 U9124 ( .A1(n9814), .A2(n9813), .ZN(n14355) );
  INV_X1 U9125 ( .A(n14104), .ZN(n14212) );
  AND2_X1 U9126 ( .A1(n9497), .A2(n9498), .ZN(n7528) );
  NAND2_X1 U9127 ( .A1(n7302), .A2(n11041), .ZN(n11058) );
  NAND2_X1 U9128 ( .A1(n14277), .A2(n11056), .ZN(n7302) );
  OR2_X1 U9129 ( .A1(n11018), .A2(n11019), .ZN(n11096) );
  NAND2_X1 U9130 ( .A1(n11116), .A2(n11088), .ZN(n11091) );
  AOI21_X1 U9131 ( .B1(n7309), .B2(n11118), .A(n7308), .ZN(n7307) );
  INV_X1 U9132 ( .A(n15873), .ZN(n15896) );
  NAND2_X1 U9133 ( .A1(n7298), .A2(n14302), .ZN(n14304) );
  AOI21_X1 U9134 ( .B1(n15851), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n14334), .ZN(
        n7313) );
  OAI22_X1 U9135 ( .A1(n14331), .A2(n14330), .B1(n14329), .B2(n15873), .ZN(
        n7314) );
  INV_X1 U9136 ( .A(n14045), .ZN(n7285) );
  NAND2_X1 U9137 ( .A1(n7882), .A2(n7881), .ZN(n14347) );
  NAND2_X1 U9138 ( .A1(n14402), .A2(n9804), .ZN(n14382) );
  AOI21_X1 U9139 ( .B1(n14379), .B2(n14657), .A(n14378), .ZN(n14692) );
  AOI21_X1 U9140 ( .B1(n14394), .B2(n14657), .A(n14393), .ZN(n14697) );
  AOI21_X1 U9141 ( .B1(n14422), .B2(n14423), .A(n6560), .ZN(n14408) );
  INV_X1 U9142 ( .A(n12751), .ZN(n14716) );
  NAND2_X1 U9143 ( .A1(n7524), .A2(n6574), .ZN(n14465) );
  AOI21_X1 U9144 ( .B1(n14521), .B2(n6851), .A(n6850), .ZN(n14510) );
  AND2_X1 U9145 ( .A1(n14508), .A2(n14507), .ZN(n6851) );
  INV_X1 U9146 ( .A(n14509), .ZN(n6850) );
  OAI21_X1 U9147 ( .B1(n9692), .B2(n7751), .A(n7116), .ZN(n14558) );
  NAND2_X1 U9148 ( .A1(n14748), .A2(n9706), .ZN(n14559) );
  NOR2_X1 U9149 ( .A1(n14560), .A2(n6670), .ZN(n14562) );
  NAND2_X1 U9150 ( .A1(n9831), .A2(n9830), .ZN(n14593) );
  OAI21_X1 U9151 ( .B1(n12502), .B2(n7289), .A(n7287), .ZN(n14613) );
  NAND2_X1 U9152 ( .A1(n7903), .A2(n9827), .ZN(n14631) );
  INV_X1 U9153 ( .A(n9866), .ZN(n12506) );
  NAND2_X1 U9154 ( .A1(n11966), .A2(n7112), .ZN(n12274) );
  NAND2_X1 U9155 ( .A1(n9821), .A2(n9820), .ZN(n12326) );
  NAND2_X1 U9156 ( .A1(n9582), .A2(n9581), .ZN(n12331) );
  OR2_X1 U9157 ( .A1(n14752), .A2(n14751), .ZN(n14810) );
  INV_X1 U9158 ( .A(n12331), .ZN(n12554) );
  NAND2_X1 U9159 ( .A1(n7295), .A2(n9485), .ZN(n7294) );
  AND2_X1 U9160 ( .A1(n10492), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15914) );
  NOR2_X1 U9161 ( .A1(n7896), .A2(n9422), .ZN(n7895) );
  NAND2_X1 U9162 ( .A1(n9457), .A2(n7897), .ZN(n7896) );
  AND2_X1 U9163 ( .A1(n9456), .A2(n9455), .ZN(n9457) );
  NAND2_X1 U9164 ( .A1(n9885), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9873) );
  INV_X1 U9165 ( .A(n10375), .ZN(n11551) );
  NOR2_X1 U9166 ( .A1(n9431), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n9425) );
  AND2_X1 U9167 ( .A1(n9613), .A2(n9623), .ZN(n11114) );
  INV_X1 U9168 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10527) );
  AND2_X1 U9169 ( .A1(n9553), .A2(n9566), .ZN(n15869) );
  NOR2_X1 U9170 ( .A1(n9511), .A2(n9418), .ZN(n14231) );
  NOR2_X1 U9171 ( .A1(n9481), .A2(n9693), .ZN(n9508) );
  INV_X1 U9172 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10525) );
  INV_X1 U9173 ( .A(n9481), .ZN(n9482) );
  NAND2_X1 U9174 ( .A1(n9316), .A2(n9315), .ZN(n15469) );
  NAND2_X1 U9175 ( .A1(n12908), .A2(n9333), .ZN(n9316) );
  AOI21_X1 U9176 ( .B1(n7714), .B2(n7717), .A(n6690), .ZN(n7711) );
  NAND2_X1 U9177 ( .A1(n12635), .A2(n12634), .ZN(n12636) );
  NAND2_X1 U9178 ( .A1(n10991), .A2(n10990), .ZN(n10993) );
  NAND2_X1 U9179 ( .A1(n14966), .A2(n6952), .ZN(n14868) );
  AND4_X1 U9180 ( .A1(n8828), .A2(n8827), .A3(n8826), .A4(n8825), .ZN(n11955)
         );
  NOR2_X1 U9181 ( .A1(n14936), .A2(n7727), .ZN(n14876) );
  OR2_X1 U9182 ( .A1(n14936), .A2(n7725), .ZN(n14875) );
  AND2_X1 U9183 ( .A1(n7191), .A2(n7190), .ZN(n12447) );
  NAND2_X1 U9184 ( .A1(n6943), .A2(n6944), .ZN(n14910) );
  INV_X1 U9185 ( .A(n6942), .ZN(n6941) );
  NAND2_X1 U9186 ( .A1(n11351), .A2(n11350), .ZN(n11644) );
  NAND2_X1 U9187 ( .A1(n10642), .A2(n15600), .ZN(n8847) );
  NOR2_X1 U9188 ( .A1(n6559), .A2(n14937), .ZN(n14936) );
  AND2_X1 U9189 ( .A1(n9355), .A2(n9354), .ZN(n7233) );
  NAND4_X1 U9190 ( .A1(n8910), .A2(n8909), .A3(n8908), .A4(n8907), .ZN(n15425)
         );
  OR2_X1 U9191 ( .A1(n9273), .A2(n7249), .ZN(n8908) );
  INV_X1 U9192 ( .A(P1_U4016), .ZN(n15019) );
  OR2_X1 U9193 ( .A1(n10728), .A2(n6877), .ZN(n10710) );
  NAND2_X1 U9194 ( .A1(n6876), .A2(n6874), .ZN(n10721) );
  AOI21_X1 U9195 ( .B1(n6877), .B2(n6600), .A(n6875), .ZN(n6874) );
  INV_X1 U9196 ( .A(n10722), .ZN(n6875) );
  NAND2_X1 U9197 ( .A1(n10710), .A2(n6600), .ZN(n10723) );
  NOR2_X1 U9198 ( .A1(n10672), .A2(n10673), .ZN(n10745) );
  AOI21_X1 U9199 ( .B1(n10716), .B2(n10715), .A(n10714), .ZN(n10727) );
  AOI21_X1 U9200 ( .B1(n10747), .B2(n10746), .A(n10745), .ZN(n10748) );
  NOR2_X1 U9201 ( .A1(n10748), .A2(n10749), .ZN(n11067) );
  AOI21_X1 U9202 ( .B1(n11068), .B2(n11075), .A(n11067), .ZN(n15050) );
  NAND2_X1 U9203 ( .A1(n15050), .A2(n15049), .ZN(n15048) );
  INV_X1 U9204 ( .A(n7493), .ZN(n11765) );
  NAND2_X1 U9205 ( .A1(n15048), .A2(n6607), .ZN(n11071) );
  NOR2_X1 U9206 ( .A1(n11770), .A2(n6628), .ZN(n15706) );
  AND2_X1 U9207 ( .A1(n7493), .A2(n7492), .ZN(n15709) );
  NAND2_X1 U9208 ( .A1(n11767), .A2(n11766), .ZN(n7492) );
  NAND2_X1 U9209 ( .A1(n15706), .A2(n15707), .ZN(n15705) );
  OAI22_X1 U9210 ( .A1(n15709), .A2(n15708), .B1(n15710), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n11768) );
  NOR2_X1 U9211 ( .A1(n11774), .A2(n11773), .ZN(n15075) );
  NAND2_X1 U9212 ( .A1(n15705), .A2(n6836), .ZN(n11774) );
  OR2_X1 U9213 ( .A1(n15710), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6836) );
  INV_X1 U9214 ( .A(n7490), .ZN(n15067) );
  NAND2_X1 U9215 ( .A1(n15716), .A2(n15091), .ZN(n15095) );
  NAND2_X1 U9216 ( .A1(n6873), .A2(n6871), .ZN(n15084) );
  INV_X1 U9217 ( .A(n6872), .ZN(n6871) );
  OAI21_X1 U9218 ( .B1(n6869), .B2(n6870), .A(n6867), .ZN(n15104) );
  OR2_X1 U9219 ( .A1(n15719), .A2(n6868), .ZN(n6867) );
  OR2_X1 U9220 ( .A1(n6870), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6868) );
  INV_X1 U9221 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n15147) );
  OAI21_X1 U9222 ( .B1(n15144), .B2(n15142), .A(n6839), .ZN(n6838) );
  AOI21_X1 U9223 ( .B1(n15143), .B2(n15723), .A(n15720), .ZN(n6839) );
  NAND2_X1 U9224 ( .A1(n6881), .A2(n6880), .ZN(n6879) );
  NAND2_X1 U9225 ( .A1(n15145), .A2(n15723), .ZN(n6881) );
  NAND2_X1 U9226 ( .A1(n15144), .A2(n15724), .ZN(n6880) );
  NAND2_X1 U9227 ( .A1(n15149), .A2(n10870), .ZN(n15444) );
  NAND2_X1 U9228 ( .A1(n8729), .A2(n8728), .ZN(n15159) );
  NAND2_X1 U9229 ( .A1(n7428), .A2(n7431), .ZN(n15225) );
  OR2_X1 U9230 ( .A1(n15258), .A2(n7433), .ZN(n7428) );
  NAND2_X1 U9231 ( .A1(n7436), .A2(n7805), .ZN(n15228) );
  NAND2_X1 U9232 ( .A1(n15258), .A2(n7807), .ZN(n7436) );
  AND2_X1 U9233 ( .A1(n9270), .A2(n9251), .ZN(n15252) );
  NAND2_X1 U9234 ( .A1(n7806), .A2(n12705), .ZN(n15241) );
  NAND2_X1 U9235 ( .A1(n15258), .A2(n12704), .ZN(n7806) );
  NAND2_X1 U9236 ( .A1(n7649), .A2(n7650), .ZN(n15260) );
  AOI21_X1 U9237 ( .B1(n15290), .B2(n15289), .A(n12728), .ZN(n15269) );
  INV_X1 U9238 ( .A(n7437), .ZN(n15285) );
  AOI21_X1 U9239 ( .B1(n15330), .B2(n7444), .A(n7442), .ZN(n7437) );
  AND2_X1 U9240 ( .A1(n7639), .A2(n12725), .ZN(n15300) );
  INV_X1 U9241 ( .A(n12700), .ZN(n7445) );
  INV_X1 U9242 ( .A(n15519), .ZN(n15327) );
  NAND2_X1 U9243 ( .A1(n12724), .A2(n12723), .ZN(n15316) );
  OAI21_X1 U9244 ( .B1(n15375), .B2(n7803), .A(n7801), .ZN(n15335) );
  NAND2_X1 U9245 ( .A1(n15374), .A2(n12696), .ZN(n15352) );
  NAND2_X1 U9246 ( .A1(n10783), .A2(n9333), .ZN(n6790) );
  AND2_X1 U9247 ( .A1(n7655), .A2(n6709), .ZN(n12027) );
  OR2_X1 U9248 ( .A1(n11440), .A2(n11439), .ZN(n15393) );
  INV_X1 U9249 ( .A(n11532), .ZN(n11717) );
  NAND2_X1 U9250 ( .A1(n7630), .A2(n11712), .ZN(n11754) );
  NAND2_X1 U9251 ( .A1(n6544), .A2(n15743), .ZN(n15418) );
  AND2_X1 U9252 ( .A1(n6544), .A2(n11446), .ZN(n15383) );
  INV_X1 U9253 ( .A(n15418), .ZN(n15730) );
  OR2_X1 U9254 ( .A1(n10969), .A2(n11436), .ZN(n15848) );
  NOR2_X1 U9255 ( .A1(n15453), .A2(n15452), .ZN(n15456) );
  AND2_X1 U9256 ( .A1(n15464), .A2(n15463), .ZN(n15465) );
  INV_X1 U9257 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n7454) );
  NAND3_X1 U9258 ( .A1(n7822), .A2(n7821), .A3(n8698), .ZN(n15586) );
  XNOR2_X1 U9259 ( .A(n8680), .B(n8679), .ZN(n15583) );
  NAND2_X1 U9260 ( .A1(n7147), .A2(n7148), .ZN(n8680) );
  NAND2_X1 U9261 ( .A1(n8699), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8700) );
  OR2_X1 U9262 ( .A1(n8694), .A2(n8691), .ZN(n7182) );
  NOR2_X1 U9263 ( .A1(n7181), .A2(n7180), .ZN(n7179) );
  NAND2_X1 U9264 ( .A1(n9373), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9374) );
  NAND2_X1 U9265 ( .A1(n9289), .A2(n9288), .ZN(n12486) );
  INV_X1 U9266 ( .A(n10788), .ZN(n15598) );
  XNOR2_X1 U9267 ( .A(n9223), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15599) );
  NAND2_X1 U9268 ( .A1(n8707), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8708) );
  INV_X1 U9269 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10622) );
  INV_X1 U9270 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10618) );
  INV_X1 U9271 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10583) );
  NAND2_X1 U9272 ( .A1(n8924), .A2(n8943), .ZN(n10626) );
  AND2_X1 U9273 ( .A1(n8902), .A2(n8901), .ZN(n15040) );
  NAND2_X1 U9274 ( .A1(n8899), .A2(n6884), .ZN(n10683) );
  AOI21_X1 U9275 ( .B1(n8880), .B2(n6661), .A(n6885), .ZN(n6884) );
  NOR2_X1 U9276 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n6885) );
  OAI211_X1 U9277 ( .C1(P1_IR_REG_31__SCAN_IN), .C2(P1_IR_REG_1__SCAN_IN), .A(
        n8880), .B(n6840), .ZN(n10678) );
  XNOR2_X1 U9278 ( .A(n10556), .B(n7520), .ZN(n16029) );
  INV_X1 U9279 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7520) );
  INV_X1 U9280 ( .A(n10567), .ZN(n7505) );
  NAND2_X1 U9281 ( .A1(n10566), .A2(n15669), .ZN(n7506) );
  NAND2_X1 U9282 ( .A1(n7517), .A2(n7756), .ZN(n7758) );
  NAND2_X1 U9283 ( .A1(n10546), .A2(n10816), .ZN(n7756) );
  NAND2_X1 U9284 ( .A1(n7757), .A2(n6624), .ZN(n7517) );
  AND2_X1 U9285 ( .A1(n6624), .A2(n10816), .ZN(n7518) );
  XNOR2_X1 U9286 ( .A(n10818), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(n15605) );
  XNOR2_X1 U9287 ( .A(n10828), .B(n10821), .ZN(n15607) );
  XNOR2_X1 U9288 ( .A(n11620), .B(n11322), .ZN(n11323) );
  INV_X1 U9289 ( .A(n7501), .ZN(n7500) );
  INV_X1 U9290 ( .A(n11831), .ZN(n7763) );
  XNOR2_X1 U9291 ( .A(n15644), .B(n15642), .ZN(n15647) );
  INV_X1 U9292 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n15661) );
  NAND2_X1 U9293 ( .A1(n10924), .A2(n8199), .ZN(n11105) );
  AND2_X1 U9294 ( .A1(n6901), .A2(n6900), .ZN(n11466) );
  OAI211_X1 U9295 ( .C1(n13613), .C2(n13612), .A(n7158), .B(n6912), .ZN(
        P3_U3201) );
  NAND2_X1 U9296 ( .A1(n6637), .A2(n13503), .ZN(n7158) );
  AND2_X1 U9297 ( .A1(n7086), .A2(n6758), .ZN(n6912) );
  MUX2_X1 U9298 ( .A(n10125), .B(n13842), .S(n15995), .Z(n13633) );
  AOI21_X1 U9299 ( .B1(n13922), .B2(n13837), .A(n7214), .ZN(n7220) );
  INV_X1 U9300 ( .A(n13646), .ZN(n7214) );
  AOI22_X1 U9301 ( .A1(n13845), .A2(n13902), .B1(n13893), .B2(n13844), .ZN(
        n13846) );
  AND2_X1 U9302 ( .A1(n13921), .A2(n13893), .ZN(n7172) );
  NAND2_X1 U9303 ( .A1(n13844), .A2(n13981), .ZN(n7174) );
  AND2_X1 U9304 ( .A1(n13921), .A2(n13981), .ZN(n7173) );
  AND2_X1 U9305 ( .A1(n12823), .A2(n7222), .ZN(n7221) );
  NAND2_X1 U9306 ( .A1(n14690), .A2(n14189), .ZN(n7222) );
  NOR2_X1 U9307 ( .A1(n11674), .A2(n6799), .ZN(n11679) );
  NAND2_X1 U9308 ( .A1(n14052), .A2(n6747), .ZN(n7217) );
  NAND2_X1 U9309 ( .A1(n7315), .A2(n7311), .ZN(P2_U3233) );
  AOI21_X1 U9310 ( .B1(n7314), .B2(n14332), .A(n7312), .ZN(n7311) );
  NAND2_X1 U9311 ( .A1(n14333), .A2(n11860), .ZN(n7315) );
  INV_X1 U9312 ( .A(n7313), .ZN(n7312) );
  AOI21_X1 U9313 ( .B1(n14433), .B2(n6802), .A(n6801), .ZN(n12260) );
  AOI21_X1 U9314 ( .B1(n14682), .B2(n14681), .A(n14680), .ZN(n14683) );
  AND2_X1 U9315 ( .A1(n7740), .A2(n15929), .ZN(n7737) );
  INV_X1 U9316 ( .A(n10149), .ZN(n7107) );
  NAND2_X1 U9317 ( .A1(n7105), .A2(n7104), .ZN(n7103) );
  AOI21_X1 U9318 ( .B1(n14682), .B2(n6802), .A(n6800), .ZN(n12306) );
  NOR2_X1 U9319 ( .A1(n15944), .A2(n9518), .ZN(n6800) );
  AOI21_X1 U9320 ( .B1(n12906), .B2(n14681), .A(n12905), .ZN(n12907) );
  NAND2_X1 U9321 ( .A1(n14818), .A2(n15929), .ZN(n7875) );
  NAND2_X1 U9322 ( .A1(n7871), .A2(n14818), .ZN(n7872) );
  NAND2_X1 U9323 ( .A1(n6863), .A2(n6862), .ZN(P2_U3495) );
  NAND2_X1 U9324 ( .A1(n15938), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6862) );
  NAND2_X1 U9325 ( .A1(n6864), .A2(n14818), .ZN(n6863) );
  NAND2_X1 U9326 ( .A1(n6865), .A2(n7165), .ZN(n6864) );
  OAI21_X1 U9327 ( .B1(n15594), .B2(n12909), .A(n7273), .ZN(P2_U3300) );
  NOR2_X1 U9328 ( .A1(n7275), .A2(n7274), .ZN(n7273) );
  NOR2_X1 U9329 ( .A1(n14826), .A2(n12910), .ZN(n7275) );
  XNOR2_X1 U9330 ( .A(n7188), .B(n14898), .ZN(n14904) );
  OAI21_X1 U9331 ( .B1(n7245), .B2(n14994), .A(n14984), .ZN(P1_U3240) );
  XNOR2_X1 U9332 ( .A(n14977), .B(n6611), .ZN(n7245) );
  NAND2_X1 U9333 ( .A1(n7177), .A2(n6837), .ZN(P1_U3262) );
  AOI21_X1 U9334 ( .B1(n6879), .B2(n6539), .A(n7178), .ZN(n7177) );
  NAND2_X1 U9335 ( .A1(n6838), .A2(n15748), .ZN(n6837) );
  OAI21_X1 U9336 ( .B1(n15728), .B2(n15147), .A(n15146), .ZN(n7178) );
  AOI21_X1 U9337 ( .B1(n7450), .B2(n15838), .A(n6598), .ZN(n7449) );
  NAND2_X1 U9338 ( .A1(n10843), .A2(n10842), .ZN(n11314) );
  NAND2_X1 U9339 ( .A1(n12582), .A2(n7042), .ZN(n12297) );
  NAND2_X1 U9340 ( .A1(n7521), .A2(n15610), .ZN(n12592) );
  AND2_X1 U9341 ( .A1(n15623), .A2(n15620), .ZN(n15622) );
  NAND2_X1 U9342 ( .A1(n7761), .A2(n15623), .ZN(n15624) );
  INV_X1 U9343 ( .A(n7762), .ZN(n7761) );
  NAND2_X1 U9344 ( .A1(n7507), .A2(n7512), .ZN(n15635) );
  NAND2_X1 U9345 ( .A1(n7509), .A2(n7512), .ZN(n15633) );
  NAND2_X1 U9346 ( .A1(n7052), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n7051) );
  INV_X2 U9347 ( .A(n10340), .ZN(n10339) );
  OAI21_X1 U9348 ( .B1(n6582), .B2(n7928), .A(n13359), .ZN(n7927) );
  OR2_X1 U9349 ( .A1(n12522), .A2(n13388), .ZN(n6552) );
  NAND2_X1 U9350 ( .A1(n7911), .A2(n13319), .ZN(n6553) );
  AND2_X1 U9351 ( .A1(n14964), .A2(n7830), .ZN(n6554) );
  AND4_X1 U9352 ( .A1(n10391), .A2(n6722), .A3(n6590), .A4(n14586), .ZN(n6555)
         );
  AND2_X1 U9353 ( .A1(n7152), .A2(n8726), .ZN(n6556) );
  AND2_X1 U9354 ( .A1(n7096), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n6557) );
  INV_X1 U9355 ( .A(n10194), .ZN(n10340) );
  CLKBUF_X3 U9356 ( .A(n9678), .Z(n10336) );
  INV_X1 U9358 ( .A(n10413), .ZN(n12750) );
  NOR2_X1 U9359 ( .A1(n8645), .A2(n9100), .ZN(n6558) );
  NOR2_X1 U9360 ( .A1(n14867), .A2(n7987), .ZN(n6559) );
  AND2_X1 U9361 ( .A1(n14705), .A2(n14077), .ZN(n6560) );
  INV_X1 U9362 ( .A(n8332), .ZN(n12911) );
  AND2_X1 U9363 ( .A1(n12800), .A2(n12801), .ZN(n6561) );
  AND2_X1 U9364 ( .A1(n13678), .A2(n7070), .ZN(n6562) );
  NAND2_X1 U9365 ( .A1(n14695), .A2(n12818), .ZN(n6563) );
  AND2_X1 U9366 ( .A1(n13038), .A2(n12973), .ZN(n6564) );
  AND2_X1 U9367 ( .A1(n13541), .A2(n7708), .ZN(n6565) );
  AND2_X1 U9368 ( .A1(n12742), .A2(n7825), .ZN(n6566) );
  AND2_X1 U9369 ( .A1(n7804), .A2(n12696), .ZN(n6567) );
  AND2_X1 U9370 ( .A1(n9268), .A2(n7614), .ZN(n6568) );
  AND2_X1 U9371 ( .A1(n13061), .A2(n13067), .ZN(n12983) );
  NOR2_X1 U9372 ( .A1(n13874), .A2(n13744), .ZN(n6569) );
  INV_X1 U9373 ( .A(n10203), .ZN(n7475) );
  AND2_X1 U9374 ( .A1(n9564), .A2(n9563), .ZN(n15932) );
  INV_X1 U9375 ( .A(n7927), .ZN(n7926) );
  AND2_X1 U9376 ( .A1(n13710), .A2(n13720), .ZN(n6570) );
  NAND2_X1 U9377 ( .A1(n7654), .A2(n15289), .ZN(n6571) );
  AND2_X1 U9378 ( .A1(n14401), .A2(n14415), .ZN(n6572) );
  OR2_X1 U9379 ( .A1(n12898), .A2(n13449), .ZN(n6573) );
  AND2_X1 U9380 ( .A1(n7753), .A2(n7525), .ZN(n6574) );
  XNOR2_X1 U9381 ( .A(n10380), .B(n10379), .ZN(n14348) );
  INV_X1 U9382 ( .A(n14348), .ZN(n6815) );
  AND2_X1 U9383 ( .A1(n6750), .A2(n6854), .ZN(n6575) );
  NAND2_X1 U9384 ( .A1(n15599), .A2(n10642), .ZN(n15277) );
  AND2_X1 U9385 ( .A1(n12026), .A2(n6709), .ZN(n6576) );
  INV_X1 U9386 ( .A(n13133), .ZN(n7847) );
  XNOR2_X1 U9387 ( .A(n8706), .B(P1_IR_REG_21__SCAN_IN), .ZN(n8720) );
  AND2_X1 U9388 ( .A1(n7912), .A2(n13416), .ZN(n6577) );
  INV_X1 U9389 ( .A(n14198), .ZN(n14077) );
  OR2_X1 U9390 ( .A1(n15302), .A2(n7832), .ZN(n6578) );
  AND2_X1 U9391 ( .A1(n11323), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n6579) );
  INV_X1 U9392 ( .A(n7717), .ZN(n7716) );
  OAI21_X1 U9393 ( .B1(n14898), .B2(n7720), .A(n13222), .ZN(n7717) );
  INV_X1 U9394 ( .A(n12242), .ZN(n9865) );
  AND2_X1 U9395 ( .A1(n8804), .A2(n8803), .ZN(n6580) );
  OR2_X1 U9396 ( .A1(n13921), .A2(n13655), .ZN(n6581) );
  NOR2_X1 U9397 ( .A1(n13434), .A2(n13433), .ZN(n6582) );
  NAND2_X1 U9398 ( .A1(n9335), .A2(n9334), .ZN(n15462) );
  AND2_X1 U9399 ( .A1(n6619), .A2(n11150), .ZN(n6583) );
  AND2_X1 U9400 ( .A1(n6949), .A2(n6950), .ZN(n6584) );
  AND3_X1 U9401 ( .A1(n8712), .A2(n8710), .A3(n9918), .ZN(n6585) );
  NAND2_X1 U9402 ( .A1(n13172), .A2(n13164), .ZN(n6586) );
  NAND2_X2 U9403 ( .A1(n8136), .A2(n6542), .ZN(n12951) );
  NAND2_X1 U9404 ( .A1(n9044), .A2(n9043), .ZN(n15553) );
  INV_X1 U9405 ( .A(n15553), .ZN(n7829) );
  NOR2_X1 U9406 ( .A1(n7448), .A2(n7445), .ZN(n6587) );
  AND2_X1 U9407 ( .A1(n7599), .A2(n9336), .ZN(n6588) );
  AND2_X1 U9408 ( .A1(n7469), .A2(n10231), .ZN(n6589) );
  AND3_X1 U9409 ( .A1(n6812), .A2(n6811), .A3(n14668), .ZN(n6590) );
  AND2_X1 U9410 ( .A1(n10262), .A2(n10261), .ZN(n6591) );
  AND2_X1 U9411 ( .A1(n6566), .A2(n7824), .ZN(n6592) );
  AND2_X1 U9412 ( .A1(n11926), .A2(n11914), .ZN(n6593) );
  AOI21_X1 U9413 ( .B1(n13672), .B2(n6551), .A(n8526), .ZN(n13654) );
  INV_X1 U9414 ( .A(n13654), .ZN(n6960) );
  INV_X1 U9415 ( .A(n10269), .ZN(n7466) );
  AND2_X1 U9416 ( .A1(n15944), .A2(n15929), .ZN(n6594) );
  NAND2_X1 U9417 ( .A1(n11915), .A2(n11914), .ZN(n11925) );
  INV_X1 U9418 ( .A(n7151), .ZN(n7150) );
  NAND2_X1 U9419 ( .A1(n7156), .A2(n8758), .ZN(n7151) );
  AND2_X1 U9420 ( .A1(n7318), .A2(n7317), .ZN(n6595) );
  AND2_X1 U9421 ( .A1(n7321), .A2(n7320), .ZN(n6596) );
  NOR2_X1 U9422 ( .A1(n13547), .A2(n7708), .ZN(n6597) );
  NOR2_X1 U9423 ( .A1(n15838), .A2(n7454), .ZN(n6598) );
  XNOR2_X1 U9424 ( .A(n11216), .B(n11201), .ZN(n11218) );
  AND2_X1 U9425 ( .A1(n7540), .A2(n14119), .ZN(n6599) );
  OR2_X1 U9426 ( .A1(n10670), .A2(n11723), .ZN(n6600) );
  NAND2_X1 U9427 ( .A1(n6927), .A2(n13127), .ZN(n13634) );
  XNOR2_X1 U9428 ( .A(n13119), .B(n13665), .ZN(n13683) );
  NAND2_X1 U9429 ( .A1(n14548), .A2(n14530), .ZN(n14512) );
  AOI21_X1 U9430 ( .B1(n13787), .B2(n13750), .A(n7078), .ZN(n13768) );
  AOI21_X1 U9431 ( .B1(n14502), .B2(n9841), .A(n9840), .ZN(n14441) );
  NAND2_X1 U9432 ( .A1(n7411), .A2(n8620), .ZN(n6601) );
  NAND2_X1 U9433 ( .A1(n7733), .A2(n13164), .ZN(n6602) );
  NAND2_X1 U9434 ( .A1(n7821), .A2(n7425), .ZN(n6603) );
  XNOR2_X1 U9435 ( .A(n12242), .B(n14207), .ZN(n12236) );
  INV_X1 U9436 ( .A(n12236), .ZN(n7533) );
  XNOR2_X1 U9437 ( .A(n15469), .B(n15213), .ZN(n12736) );
  AND2_X1 U9438 ( .A1(n10908), .A2(n8095), .ZN(n6604) );
  NAND2_X1 U9439 ( .A1(n8106), .A2(n7325), .ZN(n6605) );
  AND2_X1 U9440 ( .A1(n10205), .A2(n10204), .ZN(n6606) );
  INV_X1 U9441 ( .A(n9706), .ZN(n7751) );
  OR2_X1 U9442 ( .A1(n11069), .A2(n11070), .ZN(n6607) );
  NAND2_X1 U9443 ( .A1(n13034), .A2(n13039), .ZN(n6608) );
  INV_X1 U9444 ( .A(n14196), .ZN(n12818) );
  NAND2_X1 U9445 ( .A1(n9803), .A2(n9802), .ZN(n14196) );
  XNOR2_X1 U9446 ( .A(n8708), .B(n7729), .ZN(n8722) );
  NAND2_X1 U9447 ( .A1(n8367), .A2(n8366), .ZN(n13817) );
  AND2_X1 U9448 ( .A1(n8103), .A2(n7323), .ZN(n6609) );
  INV_X1 U9449 ( .A(n10219), .ZN(n7785) );
  AND2_X1 U9450 ( .A1(n10462), .A2(n10460), .ZN(n6610) );
  XNOR2_X1 U9451 ( .A(n13229), .B(n13230), .ZN(n6611) );
  INV_X1 U9452 ( .A(n9509), .ZN(n9418) );
  AND2_X1 U9453 ( .A1(n8705), .A2(n8709), .ZN(n6612) );
  AND2_X1 U9454 ( .A1(n10193), .A2(n10192), .ZN(n6613) );
  AND2_X1 U9455 ( .A1(n7777), .A2(n10222), .ZN(n6614) );
  OR3_X1 U9456 ( .A1(n11123), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n6615) );
  NOR2_X1 U9457 ( .A1(n9675), .A2(n14632), .ZN(n6616) );
  NAND2_X1 U9458 ( .A1(n8772), .A2(n8769), .ZN(n6617) );
  NOR2_X1 U9459 ( .A1(n9591), .A2(n12317), .ZN(n6618) );
  OR2_X1 U9460 ( .A1(n11149), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n6619) );
  NAND2_X1 U9461 ( .A1(n15731), .A2(n14839), .ZN(n6620) );
  NAND2_X1 U9462 ( .A1(n10159), .A2(n10158), .ZN(n6621) );
  NAND2_X1 U9463 ( .A1(n6965), .A2(n8027), .ZN(n8380) );
  NAND2_X1 U9464 ( .A1(n7336), .A2(n7335), .ZN(n7334) );
  XNOR2_X1 U9465 ( .A(n15222), .B(n14998), .ZN(n12734) );
  INV_X1 U9466 ( .A(n12734), .ZN(n7635) );
  AND4_X1 U9467 ( .A1(n10387), .A2(n10386), .A3(n12319), .A4(n12125), .ZN(
        n6622) );
  NAND2_X1 U9468 ( .A1(n7393), .A2(n7397), .ZN(n13368) );
  AND2_X1 U9469 ( .A1(n14177), .A2(n12807), .ZN(n6623) );
  NAND2_X1 U9470 ( .A1(n10568), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n6624) );
  NOR2_X1 U9471 ( .A1(n8653), .A2(n8652), .ZN(n6625) );
  INV_X1 U9472 ( .A(n10211), .ZN(n7786) );
  NAND2_X1 U9473 ( .A1(n10276), .A2(n10275), .ZN(n6626) );
  AND2_X1 U9474 ( .A1(n14566), .A2(n14575), .ZN(n6627) );
  NAND2_X1 U9475 ( .A1(n13436), .A2(n8373), .ZN(n13358) );
  NAND2_X1 U9476 ( .A1(n13309), .A2(n8432), .ZN(n13376) );
  NOR2_X1 U9477 ( .A1(n8315), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n8328) );
  AND2_X1 U9478 ( .A1(n11771), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6628) );
  AND2_X1 U9479 ( .A1(n13133), .A2(n8579), .ZN(n6629) );
  AND2_X1 U9480 ( .A1(n10383), .A2(n6842), .ZN(n6630) );
  AND2_X1 U9481 ( .A1(n11645), .A2(n11646), .ZN(n6631) );
  INV_X1 U9482 ( .A(SI_12_), .ZN(n10639) );
  INV_X1 U9483 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n13260) );
  AND2_X1 U9484 ( .A1(n14348), .A2(n9856), .ZN(n6632) );
  XNOR2_X1 U9485 ( .A(n15507), .B(n15002), .ZN(n15289) );
  INV_X1 U9486 ( .A(n9864), .ZN(n15917) );
  OR2_X1 U9487 ( .A1(n11645), .A2(n11646), .ZN(n6633) );
  AND2_X1 U9488 ( .A1(n9727), .A2(n15855), .ZN(n6634) );
  OR2_X1 U9489 ( .A1(n10152), .A2(n13731), .ZN(n6635) );
  NAND2_X1 U9490 ( .A1(n7375), .A2(n8500), .ZN(n13347) );
  INV_X1 U9491 ( .A(n13347), .ZN(n7921) );
  OR2_X1 U9492 ( .A1(n10227), .A2(n10225), .ZN(n6636) );
  XNOR2_X1 U9493 ( .A(n13604), .B(n13603), .ZN(n6637) );
  XNOR2_X1 U9494 ( .A(n14351), .B(n14681), .ZN(n6638) );
  NAND2_X1 U9495 ( .A1(n9466), .A2(n9465), .ZN(n14195) );
  INV_X1 U9496 ( .A(n14195), .ZN(n7884) );
  AND2_X1 U9497 ( .A1(n12710), .A2(n15201), .ZN(n15472) );
  NAND2_X1 U9498 ( .A1(n14533), .A2(n14532), .ZN(n14531) );
  AND2_X1 U9499 ( .A1(n7912), .A2(n7380), .ZN(n6639) );
  NAND2_X1 U9500 ( .A1(n8795), .A2(n8794), .ZN(n15731) );
  AND2_X1 U9501 ( .A1(n7668), .A2(n6971), .ZN(n6640) );
  NAND4_X1 U9502 ( .A1(n8295), .A2(n8294), .A3(n8293), .A4(n8292), .ZN(n13455)
         );
  NAND2_X1 U9503 ( .A1(n9791), .A2(n9790), .ZN(n14197) );
  OR2_X1 U9504 ( .A1(n10157), .A2(n10156), .ZN(n6641) );
  INV_X1 U9505 ( .A(n12984), .ZN(n13814) );
  AND2_X1 U9506 ( .A1(n13074), .A2(n13075), .ZN(n12984) );
  INV_X1 U9507 ( .A(n12315), .ZN(n12412) );
  NAND2_X1 U9508 ( .A1(n9555), .A2(n9554), .ZN(n12315) );
  NAND2_X1 U9509 ( .A1(n8720), .A2(n8722), .ZN(n10871) );
  INV_X1 U9510 ( .A(n10871), .ZN(n6953) );
  AND2_X1 U9511 ( .A1(n9478), .A2(n14231), .ZN(n6642) );
  INV_X1 U9512 ( .A(n10396), .ZN(n14381) );
  XNOR2_X1 U9513 ( .A(n14690), .B(n14195), .ZN(n10396) );
  NAND2_X1 U9514 ( .A1(n7787), .A2(n7786), .ZN(n6643) );
  OR2_X1 U9515 ( .A1(n8988), .A2(n10578), .ZN(n6644) );
  NAND2_X1 U9516 ( .A1(n8151), .A2(n11150), .ZN(n11183) );
  INV_X1 U9517 ( .A(n11183), .ZN(n7335) );
  INV_X1 U9518 ( .A(n14732), .ZN(n14530) );
  INV_X1 U9519 ( .A(n14816), .ZN(n14641) );
  OR2_X1 U9520 ( .A1(n15812), .A2(n11955), .ZN(n6645) );
  INV_X1 U9521 ( .A(n10214), .ZN(n6830) );
  AND2_X1 U9522 ( .A1(n8299), .A2(n13455), .ZN(n6646) );
  NAND2_X1 U9523 ( .A1(n8814), .A2(n8813), .ZN(n12001) );
  AND2_X1 U9524 ( .A1(n7865), .A2(n7866), .ZN(n6647) );
  NOR2_X1 U9525 ( .A1(n11465), .A2(n11642), .ZN(n6648) );
  NOR2_X1 U9526 ( .A1(n14869), .A2(n6951), .ZN(n6649) );
  NOR2_X1 U9527 ( .A1(n14348), .A2(n7743), .ZN(n6650) );
  AND2_X1 U9528 ( .A1(n12983), .A2(n7160), .ZN(n6651) );
  AND2_X1 U9529 ( .A1(n12739), .A2(n12738), .ZN(n6652) );
  AND2_X1 U9530 ( .A1(n10539), .A2(n7759), .ZN(n6653) );
  AND2_X1 U9531 ( .A1(n12739), .A2(n12708), .ZN(n6654) );
  INV_X1 U9532 ( .A(n12884), .ZN(n7258) );
  AND2_X1 U9533 ( .A1(n7623), .A2(n14716), .ZN(n6655) );
  NOR2_X1 U9534 ( .A1(n12655), .A2(n15013), .ZN(n6656) );
  INV_X1 U9535 ( .A(n9285), .ZN(n7612) );
  AND2_X1 U9536 ( .A1(n7053), .A2(n15656), .ZN(n6657) );
  AND2_X1 U9537 ( .A1(n12898), .A2(n13449), .ZN(n6658) );
  NAND2_X1 U9538 ( .A1(n9418), .A2(n9419), .ZN(n9577) );
  INV_X1 U9539 ( .A(n7808), .ZN(n7807) );
  NAND2_X1 U9540 ( .A1(n12706), .A2(n7809), .ZN(n7808) );
  AND2_X1 U9541 ( .A1(n11150), .A2(n11144), .ZN(n6659) );
  AND2_X1 U9542 ( .A1(n13043), .A2(n13042), .ZN(n13041) );
  AND4_X1 U9543 ( .A1(n8194), .A2(n8193), .A3(n8192), .A4(n8191), .ZN(n15967)
         );
  OR2_X1 U9544 ( .A1(n11195), .A2(n16021), .ZN(n6660) );
  AND2_X1 U9545 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n6661) );
  AND2_X1 U9546 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n6662) );
  INV_X1 U9547 ( .A(n9215), .ZN(n6997) );
  NAND2_X1 U9548 ( .A1(n12004), .A2(n12003), .ZN(n6663) );
  INV_X1 U9549 ( .A(n7113), .ZN(n7112) );
  NAND2_X1 U9550 ( .A1(n6618), .A2(n9565), .ZN(n7113) );
  INV_X1 U9551 ( .A(n7365), .ZN(n7361) );
  NAND2_X1 U9552 ( .A1(n7370), .A2(n7374), .ZN(n7365) );
  NOR2_X1 U9553 ( .A1(n13948), .A2(n13450), .ZN(n6664) );
  AND2_X1 U9554 ( .A1(n12490), .A2(n13454), .ZN(n6665) );
  AND2_X1 U9555 ( .A1(n7903), .A2(n7901), .ZN(n6666) );
  INV_X1 U9556 ( .A(n7663), .ZN(n7662) );
  OAI21_X1 U9557 ( .B1(n8028), .B2(n7664), .A(n8386), .ZN(n7663) );
  AND2_X1 U9558 ( .A1(n11042), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6667) );
  INV_X1 U9559 ( .A(n8339), .ZN(n7904) );
  OR2_X1 U9560 ( .A1(n9027), .A2(n9028), .ZN(n6668) );
  INV_X1 U9561 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9693) );
  AND2_X1 U9562 ( .A1(n7341), .A2(n7346), .ZN(n6669) );
  AND2_X1 U9563 ( .A1(n14502), .A2(n14561), .ZN(n6670) );
  AND2_X1 U9564 ( .A1(n13389), .A2(n13284), .ZN(n6671) );
  AND2_X1 U9565 ( .A1(n7986), .A2(n7637), .ZN(n6672) );
  AND2_X1 U9566 ( .A1(n7917), .A2(n10155), .ZN(n6673) );
  INV_X1 U9567 ( .A(n11804), .ZN(n7944) );
  NAND2_X1 U9568 ( .A1(n8616), .A2(SI_7_), .ZN(n8618) );
  INV_X1 U9569 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n7729) );
  INV_X1 U9570 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8709) );
  INV_X1 U9571 ( .A(n7079), .ZN(n7078) );
  NAND2_X1 U9572 ( .A1(n13974), .A2(n13801), .ZN(n7079) );
  INV_X1 U9573 ( .A(n7982), .ZN(n7291) );
  NOR2_X1 U9574 ( .A1(n7533), .A2(n12234), .ZN(n7982) );
  NAND2_X1 U9575 ( .A1(n8969), .A2(n8968), .ZN(n6674) );
  AND2_X1 U9576 ( .A1(n10217), .A2(n10216), .ZN(n6675) );
  INV_X1 U9577 ( .A(n7858), .ZN(n7857) );
  OAI21_X1 U9578 ( .B1(n7860), .B2(n7859), .A(n12984), .ZN(n7858) );
  NOR2_X1 U9579 ( .A1(n8068), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n6676) );
  NOR2_X1 U9580 ( .A1(n14965), .A2(n15359), .ZN(n6677) );
  NAND2_X1 U9581 ( .A1(n8198), .A2(n10901), .ZN(n8199) );
  AND2_X1 U9582 ( .A1(n10338), .A2(n10337), .ZN(n14686) );
  INV_X1 U9583 ( .A(n14686), .ZN(n10380) );
  AND2_X1 U9584 ( .A1(n15531), .A2(n15005), .ZN(n6678) );
  NAND2_X1 U9585 ( .A1(n9193), .A2(n9192), .ZN(n15305) );
  INV_X1 U9586 ( .A(n15305), .ZN(n15512) );
  INV_X1 U9587 ( .A(n15965), .ZN(n7207) );
  INV_X1 U9588 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9598) );
  INV_X1 U9589 ( .A(n11246), .ZN(n7374) );
  AND2_X1 U9590 ( .A1(n13119), .A2(n13665), .ZN(n6679) );
  INV_X1 U9591 ( .A(n14918), .ZN(n6947) );
  NAND2_X1 U9592 ( .A1(n13174), .A2(n13173), .ZN(n6680) );
  AND3_X1 U9593 ( .A1(n6903), .A2(n11534), .A3(n11797), .ZN(n6681) );
  AND2_X1 U9594 ( .A1(n14346), .A2(n14355), .ZN(n6682) );
  AND2_X1 U9595 ( .A1(n12901), .A2(n10450), .ZN(n6683) );
  INV_X1 U9596 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n9455) );
  AND2_X1 U9597 ( .A1(n13874), .A2(n13744), .ZN(n6684) );
  NAND2_X1 U9598 ( .A1(n10240), .A2(n10168), .ZN(n6685) );
  AND2_X1 U9599 ( .A1(n13921), .A2(n13448), .ZN(n6686) );
  AND2_X1 U9600 ( .A1(n9118), .A2(n9114), .ZN(n6687) );
  OR2_X1 U9601 ( .A1(n14052), .A2(n14053), .ZN(n6688) );
  NOR2_X1 U9602 ( .A1(n7786), .A2(n7787), .ZN(n6689) );
  NOR2_X1 U9603 ( .A1(n13230), .A2(n13229), .ZN(n6690) );
  NOR2_X1 U9604 ( .A1(n15488), .A2(n14999), .ZN(n6691) );
  AND2_X1 U9605 ( .A1(n7613), .A2(n7612), .ZN(n6692) );
  INV_X1 U9606 ( .A(n7828), .ZN(n7827) );
  NAND2_X1 U9607 ( .A1(n15161), .A2(n13225), .ZN(n7828) );
  NOR2_X1 U9608 ( .A1(n11258), .A2(n11219), .ZN(n6693) );
  AND2_X1 U9609 ( .A1(n8385), .A2(n13788), .ZN(n6694) );
  OR2_X1 U9610 ( .A1(n7795), .A2(n6606), .ZN(n6695) );
  INV_X1 U9611 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n9423) );
  INV_X1 U9612 ( .A(n11541), .ZN(n15786) );
  AND3_X1 U9613 ( .A1(n8905), .A2(n8904), .A3(n8903), .ZN(n11541) );
  AND2_X1 U9614 ( .A1(n7885), .A2(n9833), .ZN(n6696) );
  INV_X1 U9615 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10571) );
  NOR2_X1 U9616 ( .A1(n6631), .A2(n6939), .ZN(n6697) );
  INV_X1 U9617 ( .A(n11150), .ZN(n7575) );
  OR2_X1 U9618 ( .A1(n15317), .A2(n12722), .ZN(n6698) );
  AND2_X1 U9619 ( .A1(n10571), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6699) );
  AND2_X1 U9620 ( .A1(n10622), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n6700) );
  AND2_X1 U9621 ( .A1(n8009), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6701) );
  INV_X1 U9622 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10655) );
  AND2_X1 U9623 ( .A1(n11745), .A2(n11743), .ZN(n6702) );
  NAND2_X1 U9624 ( .A1(n11804), .A2(n12979), .ZN(n6703) );
  OR2_X1 U9625 ( .A1(n12791), .A2(n12790), .ZN(n6704) );
  NOR2_X1 U9626 ( .A1(n7622), .A2(n7884), .ZN(n6705) );
  AND2_X1 U9627 ( .A1(n14700), .A2(n14169), .ZN(n6706) );
  NAND2_X1 U9628 ( .A1(n7905), .A2(n7400), .ZN(n7401) );
  AND2_X1 U9629 ( .A1(n7286), .A2(n9829), .ZN(n6707) );
  MUX2_X1 U9630 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8150), .S(
        P3_IR_REG_1__SCAN_IN), .Z(n8151) );
  INV_X1 U9631 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8064) );
  OR2_X1 U9632 ( .A1(n13844), .A2(n13640), .ZN(n12970) );
  INV_X1 U9633 ( .A(n7074), .ZN(n7073) );
  NAND2_X1 U9634 ( .A1(n6573), .A2(n12989), .ZN(n7074) );
  OR2_X1 U9635 ( .A1(n6570), .A2(n6658), .ZN(n6708) );
  INV_X1 U9636 ( .A(n13171), .ZN(n7732) );
  INV_X1 U9637 ( .A(n7937), .ZN(n7936) );
  NAND2_X1 U9638 ( .A1(n8217), .A2(n11664), .ZN(n7937) );
  INV_X1 U9639 ( .A(n9337), .ZN(n7599) );
  NAND2_X1 U9640 ( .A1(n14877), .A2(n7726), .ZN(n7725) );
  NAND2_X1 U9641 ( .A1(n12655), .A2(n12432), .ZN(n6709) );
  INV_X1 U9642 ( .A(n9006), .ZN(n7601) );
  NAND2_X1 U9643 ( .A1(n8608), .A2(SI_5_), .ZN(n8611) );
  AND2_X1 U9644 ( .A1(n15470), .A2(n6913), .ZN(n6710) );
  AND2_X1 U9645 ( .A1(n7944), .A2(n13048), .ZN(n6711) );
  AND3_X1 U9646 ( .A1(n12436), .A2(n14952), .A3(n12435), .ZN(n6712) );
  AND2_X1 U9647 ( .A1(n7555), .A2(n6625), .ZN(n6713) );
  OR2_X1 U9648 ( .A1(n13874), .A2(n13398), .ZN(n6714) );
  AND2_X1 U9649 ( .A1(n7849), .A2(n6714), .ZN(n6715) );
  INV_X1 U9650 ( .A(n12398), .ZN(n12342) );
  AND2_X1 U9651 ( .A1(n9569), .A2(n9568), .ZN(n12398) );
  NOR3_X1 U9652 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .A3(
        P1_IR_REG_27__SCAN_IN), .ZN(n6716) );
  INV_X1 U9653 ( .A(n10398), .ZN(n9856) );
  OAI21_X1 U9654 ( .B1(n14369), .B2(n14355), .A(n14344), .ZN(n10398) );
  NAND2_X1 U9655 ( .A1(n9446), .A2(n9445), .ZN(n14690) );
  INV_X1 U9656 ( .A(n14690), .ZN(n7622) );
  AND2_X1 U9657 ( .A1(n12758), .A2(n7543), .ZN(n6717) );
  AND2_X1 U9658 ( .A1(n12741), .A2(n12740), .ZN(n6718) );
  AND4_X1 U9659 ( .A1(n8230), .A2(n8229), .A3(n8228), .A4(n8227), .ZN(n12059)
         );
  AND2_X1 U9660 ( .A1(n10364), .A2(n10363), .ZN(n6719) );
  AND2_X1 U9661 ( .A1(n6907), .A2(n15828), .ZN(n6720) );
  AND2_X1 U9662 ( .A1(n12892), .A2(n13092), .ZN(n13085) );
  NOR2_X1 U9663 ( .A1(n7852), .A2(n12893), .ZN(n7851) );
  AND2_X1 U9664 ( .A1(n13019), .A2(n13018), .ZN(n6721) );
  AND2_X1 U9665 ( .A1(n6622), .A2(n10392), .ZN(n6722) );
  OR2_X1 U9666 ( .A1(n7448), .A2(n7446), .ZN(n6723) );
  OAI21_X1 U9667 ( .B1(n11992), .B2(n11991), .A(n12180), .ZN(n7890) );
  AND2_X1 U9668 ( .A1(n6964), .A2(n7660), .ZN(n6724) );
  AND2_X1 U9669 ( .A1(n12963), .A2(n7843), .ZN(n6725) );
  NAND2_X1 U9670 ( .A1(n10313), .A2(n10312), .ZN(n6726) );
  AND2_X1 U9671 ( .A1(n12772), .A2(n12771), .ZN(n6727) );
  INV_X1 U9672 ( .A(n11970), .ZN(n6848) );
  AND2_X1 U9673 ( .A1(n13040), .A2(n13041), .ZN(n6728) );
  OR2_X1 U9674 ( .A1(n6997), .A2(n9214), .ZN(n6729) );
  INV_X1 U9675 ( .A(n9319), .ZN(n6980) );
  AND2_X1 U9676 ( .A1(n6933), .A2(n6651), .ZN(n6730) );
  AND2_X1 U9677 ( .A1(n6626), .A2(n10257), .ZN(n6731) );
  AND2_X1 U9678 ( .A1(n7544), .A2(n7545), .ZN(n6732) );
  INV_X1 U9679 ( .A(n6563), .ZN(n7284) );
  AND2_X1 U9680 ( .A1(n6921), .A2(n13123), .ZN(n6733) );
  AND2_X1 U9681 ( .A1(n6585), .A2(n7729), .ZN(n6734) );
  INV_X1 U9682 ( .A(n11313), .ZN(n7502) );
  INV_X1 U9683 ( .A(n7987), .ZN(n6950) );
  INV_X1 U9684 ( .A(n9304), .ZN(n7609) );
  AND2_X1 U9685 ( .A1(n10250), .A2(n6626), .ZN(n6735) );
  AND2_X1 U9686 ( .A1(n6554), .A2(n7829), .ZN(n6736) );
  AND2_X1 U9687 ( .A1(n6612), .A2(n6985), .ZN(n6737) );
  AND2_X1 U9688 ( .A1(n13134), .A2(n12956), .ZN(n12993) );
  OR2_X1 U9689 ( .A1(n13817), .A2(n7969), .ZN(n6738) );
  INV_X1 U9690 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9918) );
  INV_X1 U9691 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n7238) );
  INV_X1 U9692 ( .A(n11518), .ZN(n7819) );
  AND2_X1 U9693 ( .A1(n13702), .A2(n7870), .ZN(n7869) );
  NAND2_X1 U9694 ( .A1(n6962), .A2(n8520), .ZN(n13422) );
  INV_X1 U9695 ( .A(n13422), .ZN(n6961) );
  AND2_X1 U9696 ( .A1(n6938), .A2(n6633), .ZN(n11893) );
  AND2_X1 U9697 ( .A1(n10808), .A2(n10807), .ZN(n10870) );
  NAND2_X1 U9698 ( .A1(n12635), .A2(n6945), .ZN(n6943) );
  INV_X1 U9699 ( .A(n14580), .ZN(n7627) );
  NAND2_X1 U9700 ( .A1(n10327), .A2(n10326), .ZN(n14681) );
  INV_X1 U9701 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7249) );
  INV_X1 U9702 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n7586) );
  INV_X1 U9703 ( .A(n10230), .ZN(n7469) );
  NAND2_X1 U9704 ( .A1(n12321), .A2(n12554), .ZN(n12277) );
  NAND2_X1 U9705 ( .A1(n6746), .A2(n9441), .ZN(n9874) );
  NAND2_X1 U9706 ( .A1(n6849), .A2(n10386), .ZN(n11969) );
  NAND2_X1 U9707 ( .A1(n12324), .A2(n9822), .ZN(n12233) );
  INV_X1 U9708 ( .A(n14994), .ZN(n14969) );
  NOR2_X1 U9709 ( .A1(n9707), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n9716) );
  INV_X1 U9710 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n7583) );
  INV_X1 U9711 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n7257) );
  NAND2_X1 U9712 ( .A1(n6917), .A2(n7258), .ZN(n12887) );
  NAND2_X1 U9713 ( .A1(n13581), .A2(n13577), .ZN(n6739) );
  INV_X1 U9714 ( .A(n10270), .ZN(n7467) );
  INV_X1 U9715 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n7338) );
  AND2_X1 U9716 ( .A1(n8040), .A2(n7687), .ZN(n6740) );
  AND2_X1 U9717 ( .A1(n11885), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n6741) );
  OR2_X1 U9718 ( .A1(n8664), .A2(SI_25_), .ZN(n6742) );
  XNOR2_X1 U9719 ( .A(n15305), .B(n15003), .ZN(n15299) );
  INV_X1 U9720 ( .A(n15299), .ZN(n7447) );
  AND2_X1 U9721 ( .A1(n11480), .A2(n7327), .ZN(n6743) );
  NAND2_X1 U9722 ( .A1(n7012), .A2(n7013), .ZN(n11954) );
  NAND2_X1 U9723 ( .A1(n7856), .A2(n7862), .ZN(n13813) );
  NAND2_X1 U9724 ( .A1(n11527), .A2(n11526), .ZN(n11710) );
  OR2_X1 U9725 ( .A1(n11464), .A2(n11740), .ZN(n6744) );
  AND2_X1 U9726 ( .A1(n6943), .A2(n6941), .ZN(n6745) );
  NOR2_X1 U9727 ( .A1(n9577), .A2(n9422), .ZN(n6746) );
  INV_X1 U9728 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7199) );
  INV_X1 U9729 ( .A(n13127), .ZN(n6930) );
  AND3_X1 U9730 ( .A1(n14044), .A2(n14043), .A3(n14180), .ZN(n6747) );
  NOR2_X1 U9731 ( .A1(n14639), .A2(n7629), .ZN(n14598) );
  AND2_X1 U9732 ( .A1(n7111), .A2(n7110), .ZN(n12232) );
  AND2_X1 U9733 ( .A1(n8442), .A2(n13760), .ZN(n6748) );
  INV_X1 U9734 ( .A(n8758), .ZN(n7154) );
  XNOR2_X1 U9735 ( .A(n8674), .B(SI_29_), .ZN(n8758) );
  INV_X1 U9736 ( .A(n10228), .ZN(n7792) );
  AND2_X1 U9737 ( .A1(n14605), .A2(n7628), .ZN(n6749) );
  NAND2_X1 U9738 ( .A1(n14515), .A2(n14484), .ZN(n6750) );
  NAND2_X1 U9739 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n6751) );
  INV_X1 U9740 ( .A(n7350), .ZN(n13502) );
  NAND2_X1 U9741 ( .A1(n7352), .A2(n7351), .ZN(n7350) );
  OR2_X1 U9742 ( .A1(n12793), .A2(n12794), .ZN(n6752) );
  NOR2_X1 U9743 ( .A1(n15944), .A2(n9904), .ZN(n6753) );
  AND2_X1 U9744 ( .A1(n10775), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n6754) );
  AND2_X1 U9745 ( .A1(n6896), .A2(n7708), .ZN(n6755) );
  INV_X1 U9746 ( .A(n7352), .ZN(n13479) );
  OR2_X1 U9747 ( .A1(n12149), .A2(n7353), .ZN(n7352) );
  AND2_X1 U9748 ( .A1(n13615), .A2(n13616), .ZN(n6756) );
  AND2_X1 U9749 ( .A1(n11660), .A2(n7993), .ZN(n6757) );
  NOR2_X1 U9750 ( .A1(n13614), .A2(n6756), .ZN(n6758) );
  AND2_X1 U9751 ( .A1(n6869), .A2(n6873), .ZN(n6759) );
  NAND2_X1 U9752 ( .A1(n6821), .A2(n6820), .ZN(n9431) );
  AND2_X1 U9753 ( .A1(n7905), .A2(n7904), .ZN(n6760) );
  AND2_X1 U9754 ( .A1(n7145), .A2(n8666), .ZN(n6761) );
  OR2_X1 U9755 ( .A1(n15836), .A2(n7452), .ZN(n6762) );
  AND2_X1 U9756 ( .A1(n6557), .A2(n13534), .ZN(n6763) );
  INV_X1 U9757 ( .A(n7892), .ZN(n11989) );
  NAND2_X1 U9758 ( .A1(n8546), .A2(n10908), .ZN(n6764) );
  NAND2_X1 U9759 ( .A1(n11866), .A2(n9433), .ZN(n10166) );
  NAND2_X1 U9760 ( .A1(n9127), .A2(n9126), .ZN(n15537) );
  INV_X1 U9761 ( .A(n15537), .ZN(n7825) );
  NAND2_X1 U9762 ( .A1(n8786), .A2(n8785), .ZN(n12605) );
  INV_X1 U9763 ( .A(n12605), .ZN(n7830) );
  NOR2_X1 U9764 ( .A1(n12251), .A2(n6802), .ZN(n11996) );
  INV_X1 U9765 ( .A(n15531), .ZN(n7824) );
  INV_X1 U9766 ( .A(n13731), .ZN(n13450) );
  AND2_X1 U9767 ( .A1(n8473), .A2(n8472), .ZN(n13731) );
  AND2_X1 U9768 ( .A1(n13556), .A2(n13542), .ZN(n6765) );
  AND2_X1 U9769 ( .A1(n11968), .A2(n10166), .ZN(n14774) );
  NAND2_X1 U9770 ( .A1(n9638), .A2(n9637), .ZN(n14769) );
  INV_X1 U9771 ( .A(n14769), .ZN(n7619) );
  NAND2_X1 U9772 ( .A1(n8486), .A2(n8485), .ZN(n13720) );
  OR2_X1 U9773 ( .A1(n13475), .A2(n13466), .ZN(n6766) );
  AND2_X1 U9774 ( .A1(n11235), .A2(n11337), .ZN(n6767) );
  NAND2_X1 U9775 ( .A1(n11470), .A2(n11483), .ZN(n7580) );
  INV_X1 U9776 ( .A(n7580), .ZN(n7097) );
  AND2_X1 U9777 ( .A1(n10484), .A2(n14642), .ZN(n14173) );
  INV_X1 U9778 ( .A(n9478), .ZN(n7295) );
  INV_X1 U9779 ( .A(n13534), .ZN(n7708) );
  INV_X1 U9780 ( .A(n13561), .ZN(n7348) );
  AND2_X1 U9781 ( .A1(n7099), .A2(n7580), .ZN(n6768) );
  INV_X1 U9782 ( .A(n14492), .ZN(n6858) );
  AND2_X1 U9783 ( .A1(n7301), .A2(n7303), .ZN(n6769) );
  INV_X1 U9784 ( .A(n15435), .ZN(n6905) );
  INV_X1 U9785 ( .A(n6906), .ZN(n11540) );
  OR2_X1 U9786 ( .A1(n15435), .A2(n15786), .ZN(n6906) );
  INV_X1 U9787 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6860) );
  OR2_X1 U9788 ( .A1(n15106), .A2(n15092), .ZN(n6770) );
  AND2_X1 U9789 ( .A1(n7329), .A2(n7328), .ZN(n6771) );
  OR2_X1 U9790 ( .A1(n12187), .A2(n12315), .ZN(n12186) );
  INV_X1 U9791 ( .A(n12186), .ZN(n7615) );
  AND2_X1 U9792 ( .A1(n12485), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6772) );
  AND2_X1 U9793 ( .A1(n12483), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6773) );
  AND2_X1 U9794 ( .A1(n8677), .A2(SI_30_), .ZN(n6774) );
  AND2_X1 U9795 ( .A1(n11252), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n6775) );
  AND2_X1 U9796 ( .A1(n14829), .A2(n9484), .ZN(n6776) );
  OR2_X1 U9797 ( .A1(n13618), .A2(n13620), .ZN(n6777) );
  NOR2_X1 U9798 ( .A1(n12874), .A2(n7692), .ZN(n7691) );
  AND2_X1 U9799 ( .A1(n11192), .A2(n11252), .ZN(n6778) );
  INV_X1 U9800 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7530) );
  INV_X1 U9801 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7897) );
  NAND3_X1 U9802 ( .A1(n7518), .A2(n10546), .A3(n7757), .ZN(n10812) );
  XOR2_X1 U9803 ( .A(n11464), .B(P3_REG2_REG_8__SCAN_IN), .Z(n6779) );
  XOR2_X1 U9804 ( .A(n13475), .B(P3_REG2_REG_12__SCAN_IN), .Z(n6780) );
  INV_X1 U9805 ( .A(n15815), .ZN(n7453) );
  XOR2_X1 U9806 ( .A(n11258), .B(P3_REG2_REG_6__SCAN_IN), .Z(n6781) );
  NOR2_X1 U9807 ( .A1(n11020), .A2(P2_U3088), .ZN(n6782) );
  AND2_X1 U9808 ( .A1(n7758), .A2(n10812), .ZN(n6783) );
  NOR2_X1 U9809 ( .A1(n10728), .A2(n7486), .ZN(n6784) );
  INV_X1 U9810 ( .A(n7391), .ZN(n13139) );
  NAND2_X1 U9811 ( .A1(n11492), .A2(n13599), .ZN(n7391) );
  INV_X1 U9812 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6818) );
  XOR2_X1 U9813 ( .A(n8181), .B(n8180), .Z(n6785) );
  NAND2_X1 U9814 ( .A1(n7575), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n11151) );
  INV_X1 U9815 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n7337) );
  INV_X1 U9816 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n7581) );
  INV_X2 U9817 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NAND2_X2 U9818 ( .A1(n8586), .A2(n8585), .ZN(n13443) );
  NAND2_X2 U9819 ( .A1(n6790), .A2(n9069), .ZN(n15543) );
  NAND2_X1 U9820 ( .A1(n6791), .A2(n7136), .ZN(n7135) );
  INV_X1 U9821 ( .A(n9036), .ZN(n6791) );
  NAND3_X1 U9822 ( .A1(n7201), .A2(n9063), .A3(n9045), .ZN(n9064) );
  NAND2_X1 U9823 ( .A1(n9852), .A2(n7988), .ZN(n14422) );
  AND2_X2 U9824 ( .A1(n14367), .A2(n9870), .ZN(n7165) );
  NAND2_X1 U9825 ( .A1(n9863), .A2(n14347), .ZN(n6797) );
  NAND3_X1 U9826 ( .A1(n7894), .A2(n7893), .A3(n6806), .ZN(n6805) );
  AND3_X2 U9827 ( .A1(n9418), .A2(n9419), .A3(n7897), .ZN(n7893) );
  NAND3_X1 U9828 ( .A1(n6555), .A2(n6810), .A3(n14609), .ZN(n10393) );
  NAND4_X1 U9829 ( .A1(n10397), .A2(n6816), .A3(n6815), .A4(n6638), .ZN(n6814)
         );
  INV_X2 U9830 ( .A(n10240), .ZN(n10194) );
  OR2_X2 U9831 ( .A1(n10166), .A2(n11551), .ZN(n10240) );
  OAI21_X1 U9832 ( .B1(n10235), .B2(n10234), .A(n10233), .ZN(n6825) );
  NAND2_X1 U9833 ( .A1(n6825), .A2(n10236), .ZN(n10239) );
  NAND2_X1 U9834 ( .A1(n6828), .A2(n6826), .ZN(n10217) );
  NAND2_X1 U9835 ( .A1(n10214), .A2(n6827), .ZN(n6826) );
  INV_X1 U9836 ( .A(n10212), .ZN(n6827) );
  NAND2_X1 U9837 ( .A1(n10213), .A2(n6829), .ZN(n6828) );
  MUX2_X1 U9838 ( .A(n10679), .B(P1_REG2_REG_1__SCAN_IN), .S(n10678), .Z(
        n15029) );
  NAND3_X1 U9839 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n6840) );
  NAND3_X1 U9840 ( .A1(n12102), .A2(n14784), .A3(n6841), .ZN(n10385) );
  NAND2_X1 U9841 ( .A1(n12254), .A2(n6842), .ZN(n11990) );
  XNOR2_X1 U9842 ( .A(n12250), .B(n6842), .ZN(n12299) );
  OR2_X2 U9843 ( .A1(n12501), .A2(n12504), .ZN(n12502) );
  NAND2_X1 U9844 ( .A1(n7891), .A2(n11970), .ZN(n6846) );
  OAI21_X1 U9845 ( .B1(n7890), .B2(n6846), .A(n6845), .ZN(n11973) );
  NAND3_X1 U9846 ( .A1(n7412), .A2(n15929), .A3(n14345), .ZN(n6865) );
  AND2_X1 U9847 ( .A1(n15101), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6870) );
  NAND2_X1 U9848 ( .A1(n10728), .A2(n6600), .ZN(n6876) );
  NAND2_X1 U9849 ( .A1(n15048), .A2(n6882), .ZN(n7493) );
  AND4_X2 U9850 ( .A1(n8690), .A2(n8689), .A3(n8925), .A4(n7992), .ZN(n7821)
         );
  NAND2_X1 U9851 ( .A1(n13489), .A2(n6889), .ZN(n6888) );
  NAND2_X1 U9852 ( .A1(n13489), .A2(n13488), .ZN(n13518) );
  INV_X1 U9853 ( .A(n6898), .ZN(n6897) );
  NAND2_X1 U9854 ( .A1(n11326), .A2(n11327), .ZN(n6901) );
  INV_X1 U9855 ( .A(n12019), .ZN(n6908) );
  NAND3_X1 U9856 ( .A1(n6615), .A2(n6909), .A3(P3_REG1_REG_1__SCAN_IN), .ZN(
        n11175) );
  NOR2_X2 U9857 ( .A1(n15250), .A2(n15482), .ZN(n15231) );
  NAND2_X1 U9858 ( .A1(n6919), .A2(n6918), .ZN(n7848) );
  OAI21_X1 U9859 ( .B1(n13694), .B2(n13678), .A(n6922), .ZN(n13668) );
  NAND2_X1 U9860 ( .A1(n6920), .A2(n6733), .ZN(n12899) );
  NAND2_X1 U9861 ( .A1(n13694), .A2(n6922), .ZN(n6920) );
  NAND2_X1 U9862 ( .A1(n6926), .A2(n6925), .ZN(n12927) );
  NAND2_X1 U9863 ( .A1(n13648), .A2(n6928), .ZN(n6926) );
  NAND2_X1 U9864 ( .A1(n13648), .A2(n13649), .ZN(n6927) );
  NAND2_X1 U9865 ( .A1(n6931), .A2(n6730), .ZN(n7159) );
  NAND3_X1 U9866 ( .A1(n7837), .A2(n7835), .A3(n6711), .ZN(n6931) );
  NAND3_X1 U9867 ( .A1(n7835), .A2(n7837), .A3(n13048), .ZN(n6932) );
  INV_X1 U9868 ( .A(n10957), .ZN(n10875) );
  NAND2_X2 U9869 ( .A1(n9376), .A2(n9377), .ZN(n10957) );
  NAND2_X1 U9870 ( .A1(n8181), .A2(n8180), .ZN(n6954) );
  NAND2_X1 U9871 ( .A1(n7659), .A2(n8152), .ZN(n6955) );
  NAND2_X1 U9872 ( .A1(n6959), .A2(n7204), .ZN(n6958) );
  NAND2_X1 U9873 ( .A1(n8360), .A2(n6966), .ZN(n6963) );
  NAND2_X1 U9874 ( .A1(n6963), .A2(n6724), .ZN(n8403) );
  NAND2_X1 U9875 ( .A1(n8360), .A2(n8359), .ZN(n6965) );
  OAI22_X2 U9876 ( .A1(n9022), .A2(n6969), .B1(n9023), .B2(n6970), .ZN(n9027)
         );
  NAND2_X1 U9877 ( .A1(n8008), .A2(n6973), .ZN(n6972) );
  NAND4_X1 U9878 ( .A1(n8690), .A2(n6737), .A3(n8925), .A4(n8689), .ZN(n6984)
         );
  AND2_X1 U9879 ( .A1(n6988), .A2(n6990), .ZN(n13138) );
  NAND3_X1 U9880 ( .A1(n6990), .A2(n6988), .A3(n15983), .ZN(n7270) );
  NAND2_X1 U9881 ( .A1(n13137), .A2(n6993), .ZN(n6990) );
  NAND3_X1 U9882 ( .A1(n13131), .A2(n13133), .A3(n13101), .ZN(n6992) );
  NAND3_X1 U9883 ( .A1(n9198), .A2(n9197), .A3(n6729), .ZN(n6995) );
  NAND2_X1 U9884 ( .A1(n6995), .A2(n6996), .ZN(n9227) );
  NAND2_X4 U9885 ( .A1(n7008), .A2(n8753), .ZN(n9295) );
  INV_X1 U9886 ( .A(n7631), .ZN(n7013) );
  NAND2_X1 U9887 ( .A1(n11527), .A2(n7014), .ZN(n7012) );
  NAND3_X1 U9888 ( .A1(n7012), .A2(n7013), .A3(n6645), .ZN(n11958) );
  NAND2_X1 U9889 ( .A1(n7822), .A2(n7821), .ZN(n8699) );
  NAND2_X1 U9890 ( .A1(n14108), .A2(n10434), .ZN(n7016) );
  NAND2_X1 U9891 ( .A1(n14109), .A2(n7017), .ZN(n14108) );
  AND2_X1 U9892 ( .A1(n14111), .A2(n10431), .ZN(n7017) );
  NAND3_X4 U9893 ( .A1(n7020), .A2(n10412), .A3(n7019), .ZN(n10413) );
  INV_X1 U9894 ( .A(n12688), .ZN(n12099) );
  AND3_X2 U9895 ( .A1(n9489), .A2(n9488), .A3(n7294), .ZN(n12688) );
  NAND2_X1 U9896 ( .A1(n14073), .A2(n7026), .ZN(n7025) );
  INV_X1 U9897 ( .A(n14163), .ZN(n12808) );
  NAND2_X1 U9898 ( .A1(n14032), .A2(n7030), .ZN(n7028) );
  NAND2_X1 U9899 ( .A1(n7028), .A2(n7029), .ZN(n12792) );
  NAND2_X1 U9900 ( .A1(n12476), .A2(n7037), .ZN(n7034) );
  NAND2_X1 U9901 ( .A1(n7034), .A2(n7035), .ZN(n7542) );
  OAI21_X1 U9902 ( .B1(n10555), .B2(n7040), .A(n10554), .ZN(n10556) );
  NAND2_X1 U9903 ( .A1(n10555), .A2(n7040), .ZN(n10554) );
  NAND2_X1 U9904 ( .A1(n7041), .A2(n7500), .ZN(n11324) );
  NAND2_X1 U9905 ( .A1(n7499), .A2(n11313), .ZN(n7041) );
  NAND3_X1 U9906 ( .A1(n12582), .A2(n7042), .A3(n7048), .ZN(n12583) );
  NAND3_X1 U9907 ( .A1(n7043), .A2(n7049), .A3(n12290), .ZN(n7042) );
  NAND2_X1 U9908 ( .A1(n12289), .A2(n15901), .ZN(n7043) );
  NAND2_X1 U9909 ( .A1(n11832), .A2(n7045), .ZN(n7044) );
  NAND2_X1 U9910 ( .A1(n12289), .A2(n7047), .ZN(n7046) );
  INV_X1 U9911 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7048) );
  INV_X1 U9912 ( .A(n12296), .ZN(n7049) );
  NAND2_X1 U9913 ( .A1(n7051), .A2(n7050), .ZN(SUB_1596_U62) );
  NAND2_X1 U9914 ( .A1(n7054), .A2(n6657), .ZN(n7050) );
  NAND2_X1 U9915 ( .A1(n7054), .A2(n7053), .ZN(n7052) );
  NAND2_X1 U9916 ( .A1(n15655), .A2(n15654), .ZN(n7053) );
  NAND2_X1 U9917 ( .A1(n7513), .A2(n15653), .ZN(n7054) );
  NAND2_X1 U9918 ( .A1(n7056), .A2(n10541), .ZN(n10548) );
  NAND2_X1 U9919 ( .A1(n7055), .A2(n10541), .ZN(n10552) );
  AND2_X1 U9920 ( .A1(n10541), .A2(n7760), .ZN(n10553) );
  NAND3_X1 U9921 ( .A1(n7056), .A2(n10541), .A3(n7057), .ZN(n10549) );
  NAND2_X1 U9922 ( .A1(n15611), .A2(n15610), .ZN(n15619) );
  NAND3_X1 U9923 ( .A1(n15610), .A2(n15611), .A3(n15617), .ZN(n15620) );
  NAND2_X4 U9924 ( .A1(n7061), .A2(n8068), .ZN(n13576) );
  NAND2_X1 U9925 ( .A1(n7331), .A2(n7061), .ZN(n7058) );
  NOR2_X1 U9926 ( .A1(n7061), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7060) );
  INV_X1 U9927 ( .A(n15972), .ZN(n10900) );
  INV_X2 U9928 ( .A(n12951), .ZN(n7065) );
  NAND2_X1 U9929 ( .A1(n16036), .A2(n6562), .ZN(n7068) );
  AOI21_X1 U9930 ( .B1(n16036), .B2(n12989), .A(n6570), .ZN(n13690) );
  AOI21_X2 U9931 ( .B1(n12492), .B2(n12491), .A(n6665), .ZN(n12523) );
  OAI21_X2 U9932 ( .B1(n11835), .B2(n6703), .A(n7942), .ZN(n12492) );
  INV_X1 U9933 ( .A(n13492), .ZN(n7081) );
  NAND2_X1 U9934 ( .A1(n7083), .A2(n13496), .ZN(n7082) );
  INV_X1 U9935 ( .A(n13470), .ZN(n7083) );
  OAI211_X1 U9936 ( .C1(n13619), .C2(n6777), .A(n7087), .B(n7088), .ZN(n7086)
         );
  NAND2_X1 U9937 ( .A1(n13619), .A2(n13620), .ZN(n7087) );
  NAND2_X1 U9938 ( .A1(n13618), .A2(n13620), .ZN(n7089) );
  NAND2_X1 U9939 ( .A1(n13527), .A2(n6763), .ZN(n7093) );
  NAND2_X1 U9940 ( .A1(n7579), .A2(n11559), .ZN(n7099) );
  NAND2_X1 U9941 ( .A1(n7098), .A2(n7580), .ZN(n11578) );
  INV_X1 U9942 ( .A(n11185), .ZN(n7100) );
  XNOR2_X1 U9943 ( .A(n11153), .B(n7100), .ZN(n11154) );
  NAND2_X1 U9944 ( .A1(n11289), .A2(n11287), .ZN(n11189) );
  NAND2_X1 U9945 ( .A1(n7412), .A2(n7102), .ZN(n7105) );
  XNOR2_X1 U9946 ( .A(n7103), .B(n7107), .ZN(P2_U3527) );
  NAND2_X1 U9947 ( .A1(n7412), .A2(n14345), .ZN(n14373) );
  CLKBUF_X1 U9948 ( .A(n7109), .Z(n7108) );
  NAND2_X2 U9949 ( .A1(n9461), .A2(n7109), .ZN(n9517) );
  NAND3_X1 U9950 ( .A1(n11967), .A2(n9608), .A3(n11971), .ZN(n7111) );
  NAND2_X1 U9951 ( .A1(n9692), .A2(n7116), .ZN(n7114) );
  NAND2_X1 U9952 ( .A1(n7114), .A2(n7115), .ZN(n14537) );
  AND2_X1 U9953 ( .A1(n8621), .A2(n8624), .ZN(n7119) );
  NAND2_X1 U9954 ( .A1(n8612), .A2(n8613), .ZN(n7122) );
  INV_X1 U9955 ( .A(n7123), .ZN(n8895) );
  INV_X1 U9956 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7125) );
  INV_X1 U9957 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7127) );
  INV_X1 U9958 ( .A(n10368), .ZN(n10353) );
  NAND3_X1 U9959 ( .A1(n7132), .A2(n7229), .A3(n8659), .ZN(n9762) );
  NAND2_X1 U9960 ( .A1(n8657), .A2(SI_22_), .ZN(n8659) );
  NAND2_X1 U9961 ( .A1(n7132), .A2(n8659), .ZN(n9760) );
  AND2_X1 U9962 ( .A1(n7572), .A2(n7145), .ZN(n7142) );
  NAND2_X1 U9963 ( .A1(n7570), .A2(n7572), .ZN(n9280) );
  INV_X1 U9964 ( .A(n9286), .ZN(n7146) );
  NAND2_X1 U9965 ( .A1(n8235), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8221) );
  INV_X1 U9966 ( .A(n8253), .ZN(n7250) );
  OAI21_X1 U9967 ( .B1(n7585), .B2(n11235), .A(n7584), .ZN(n11469) );
  NAND2_X1 U9968 ( .A1(n7997), .A2(n8595), .ZN(n8598) );
  OAI21_X2 U9969 ( .B1(n9196), .B2(n9195), .A(n9194), .ZN(n9198) );
  NAND2_X1 U9970 ( .A1(n9228), .A2(n7587), .ZN(n9244) );
  NAND2_X1 U9971 ( .A1(n6668), .A2(n9026), .ZN(n9140) );
  NAND2_X1 U9972 ( .A1(n7865), .A2(n7863), .ZN(n13694) );
  NAND2_X1 U9973 ( .A1(n10902), .A2(n10907), .ZN(n11402) );
  NAND2_X1 U9974 ( .A1(n8067), .A2(P3_IR_REG_27__SCAN_IN), .ZN(n7163) );
  NAND3_X1 U9975 ( .A1(n7161), .A2(n7607), .A3(n7246), .ZN(n7606) );
  NAND2_X1 U9976 ( .A1(n9284), .A2(n9283), .ZN(n7161) );
  NAND2_X1 U9977 ( .A1(n8596), .A2(n10517), .ZN(n8848) );
  INV_X1 U9978 ( .A(SI_22_), .ZN(n7230) );
  INV_X1 U9979 ( .A(n8661), .ZN(n9229) );
  NAND2_X1 U9980 ( .A1(n8623), .A2(n6601), .ZN(n7747) );
  NAND2_X1 U9981 ( .A1(n12863), .A2(n12862), .ZN(n13650) );
  NAND2_X1 U9983 ( .A1(n11428), .A2(n7215), .ZN(n11430) );
  NAND2_X1 U9984 ( .A1(n14889), .A2(n12452), .ZN(n12630) );
  NAND2_X1 U9985 ( .A1(n11987), .A2(n9537), .ZN(n12178) );
  NOR2_X2 U9986 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n9435) );
  NAND2_X1 U9987 ( .A1(n14429), .A2(n14428), .ZN(n14427) );
  NAND2_X1 U9988 ( .A1(n7712), .A2(n7711), .ZN(n14850) );
  NAND2_X1 U9989 ( .A1(n14828), .A2(n7529), .ZN(n9497) );
  OAI22_X1 U9990 ( .A1(n10950), .A2(n13224), .B1(n11501), .B2(n13195), .ZN(
        n7212) );
  NAND2_X1 U9991 ( .A1(n12417), .A2(n12416), .ZN(n12568) );
  NAND2_X1 U9992 ( .A1(n12568), .A2(n6712), .ZN(n7248) );
  AND3_X1 U9993 ( .A1(n8177), .A2(n8176), .A3(n8179), .ZN(n7169) );
  XNOR2_X2 U9994 ( .A(n8122), .B(n14002), .ZN(n13255) );
  NAND2_X1 U9995 ( .A1(n11402), .A2(n13016), .ZN(n11453) );
  NAND3_X1 U9996 ( .A1(n8154), .A2(n8153), .A3(n8155), .ZN(n10866) );
  NAND3_X1 U9997 ( .A1(n10403), .A2(n10402), .A3(n7170), .ZN(n10404) );
  OAI21_X1 U9998 ( .B1(n10401), .B2(n10400), .A(n7171), .ZN(n7170) );
  AOI21_X1 U9999 ( .B1(n13922), .B2(n13902), .A(n7172), .ZN(n13849) );
  AOI21_X1 U10000 ( .B1(n13922), .B2(n13992), .A(n7173), .ZN(n13923) );
  NAND2_X1 U10001 ( .A1(n13846), .A2(n13847), .ZN(P3_U3488) );
  NAND3_X1 U10002 ( .A1(n7175), .A2(n12900), .A3(n7174), .ZN(P3_U3456) );
  NAND2_X1 U10003 ( .A1(n13845), .A2(n13992), .ZN(n7175) );
  OAI21_X1 U10004 ( .B1(n7269), .B2(n13141), .A(n13140), .ZN(n13148) );
  NAND2_X1 U10005 ( .A1(n15982), .A2(n8170), .ZN(n13008) );
  NAND2_X1 U10006 ( .A1(n11802), .A2(n11801), .ZN(n11835) );
  NAND2_X1 U10007 ( .A1(n15038), .A2(n15039), .ZN(n15691) );
  AND2_X2 U10008 ( .A1(n13035), .A2(n13034), .ZN(n12973) );
  NAND2_X1 U10009 ( .A1(n11667), .A2(n13458), .ZN(n13035) );
  AOI21_X1 U10010 ( .B1(n11427), .B2(n13025), .A(n7216), .ZN(n7215) );
  NAND2_X1 U10011 ( .A1(n7247), .A2(n9177), .ZN(n9196) );
  NAND2_X1 U10012 ( .A1(n6542), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7198) );
  AOI21_X1 U10013 ( .B1(n8958), .B2(n6580), .A(n6674), .ZN(n7194) );
  NAND2_X1 U10014 ( .A1(n8048), .A2(n8047), .ZN(n8502) );
  NAND2_X1 U10015 ( .A1(n10365), .A2(n10366), .ZN(n7184) );
  OAI21_X1 U10016 ( .B1(n8615), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n7185), .ZN(
        n8597) );
  NAND2_X1 U10017 ( .A1(n8615), .A2(n9494), .ZN(n7185) );
  NAND2_X1 U10018 ( .A1(n8183), .A2(n8182), .ZN(n8008) );
  NAND2_X1 U10019 ( .A1(n8314), .A2(n8021), .ZN(n7677) );
  NAND2_X1 U10020 ( .A1(n8420), .A2(n8033), .ZN(n8035) );
  NAND2_X1 U10021 ( .A1(n8018), .A2(n8017), .ZN(n8301) );
  NAND3_X1 U10022 ( .A1(n7758), .A2(n15880), .A3(n10812), .ZN(n10813) );
  NAND2_X1 U10023 ( .A1(n12442), .A2(n14887), .ZN(n7190) );
  OAI21_X1 U10024 ( .B1(n12442), .B2(n14887), .A(n14888), .ZN(n7191) );
  NAND2_X1 U10025 ( .A1(n12448), .A2(n7248), .ZN(n14889) );
  NAND2_X1 U10026 ( .A1(n7192), .A2(n8872), .ZN(n8893) );
  NAND3_X1 U10027 ( .A1(n7193), .A2(n11504), .A3(n8871), .ZN(n7192) );
  INV_X1 U10028 ( .A(n9227), .ZN(n7589) );
  INV_X1 U10029 ( .A(n11505), .ZN(n7243) );
  NAND2_X1 U10030 ( .A1(n8970), .A2(n7194), .ZN(n8983) );
  INV_X1 U10031 ( .A(n8873), .ZN(n7193) );
  NAND2_X1 U10032 ( .A1(n7197), .A2(n7590), .ZN(n7247) );
  NAND3_X1 U10033 ( .A1(n9144), .A2(n7596), .A3(n7593), .ZN(n7197) );
  AOI22_X1 U10034 ( .A1(n7255), .A2(n7254), .B1(n10368), .B2(n10342), .ZN(
        n10343) );
  NAND2_X1 U10035 ( .A1(n7202), .A2(n10663), .ZN(n7201) );
  INV_X1 U10036 ( .A(n9115), .ZN(n7202) );
  NAND2_X1 U10037 ( .A1(n7203), .A2(n6728), .ZN(n13046) );
  NAND2_X1 U10038 ( .A1(n7262), .A2(n7261), .ZN(n7203) );
  NAND2_X1 U10039 ( .A1(n7264), .A2(n7263), .ZN(n13073) );
  NAND2_X1 U10040 ( .A1(n7209), .A2(n7206), .ZN(n13013) );
  NAND2_X1 U10041 ( .A1(n13005), .A2(n7210), .ZN(n7209) );
  NAND2_X1 U10042 ( .A1(n7211), .A2(n10982), .ZN(n11303) );
  NAND2_X1 U10043 ( .A1(n10977), .A2(n10978), .ZN(n7211) );
  NAND2_X2 U10044 ( .A1(n10456), .A2(n12469), .ZN(n12476) );
  NAND2_X1 U10045 ( .A1(n10449), .A2(n12333), .ZN(n12546) );
  NAND2_X1 U10046 ( .A1(n9716), .A2(n7549), .ZN(n9428) );
  NAND2_X1 U10047 ( .A1(n10421), .A2(n10420), .ZN(n11688) );
  NAND2_X1 U10048 ( .A1(n10426), .A2(n10425), .ZN(n11676) );
  NAND2_X1 U10049 ( .A1(n11422), .A2(n13028), .ZN(n11584) );
  INV_X1 U10050 ( .A(n15959), .ZN(n11667) );
  AND2_X1 U10051 ( .A1(n13458), .A2(n15959), .ZN(n7216) );
  NAND2_X1 U10052 ( .A1(n12546), .A2(n10452), .ZN(n12555) );
  NAND3_X1 U10053 ( .A1(n6688), .A2(n7217), .A3(n14051), .ZN(P2_U3192) );
  NAND2_X1 U10054 ( .A1(n12346), .A2(n10444), .ZN(n10449) );
  INV_X1 U10055 ( .A(n11676), .ZN(n7228) );
  NOR2_X1 U10056 ( .A1(n14175), .A2(n7989), .ZN(n12817) );
  NAND3_X1 U10057 ( .A1(n8848), .A2(n8877), .A3(n8850), .ZN(n8603) );
  NAND2_X1 U10058 ( .A1(n9762), .A2(n8659), .ZN(n9231) );
  INV_X2 U10059 ( .A(n8615), .ZN(n7219) );
  NOR2_X2 U10060 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n9434) );
  NAND2_X1 U10061 ( .A1(n13647), .A2(n7220), .ZN(P3_U3205) );
  NAND2_X1 U10062 ( .A1(n7223), .A2(n7221), .ZN(P2_U3186) );
  NAND3_X1 U10063 ( .A1(n7224), .A2(n14052), .A3(n14180), .ZN(n7223) );
  NAND2_X1 U10064 ( .A1(n7226), .A2(n7225), .ZN(n7224) );
  INV_X1 U10065 ( .A(n12817), .ZN(n7226) );
  NAND2_X1 U10066 ( .A1(n11681), .A2(n11680), .ZN(n10421) );
  NAND2_X1 U10067 ( .A1(n7645), .A2(n7642), .ZN(n15242) );
  OAI21_X1 U10068 ( .B1(n15472), .B2(n7452), .A(n7451), .ZN(n15567) );
  AOI21_X1 U10069 ( .B1(n10360), .B2(n7253), .A(n6719), .ZN(n10365) );
  INV_X1 U10070 ( .A(n8657), .ZN(n7231) );
  OAI211_X1 U10071 ( .C1(n9357), .C2(n9358), .A(n7232), .B(n9356), .ZN(n9415)
         );
  NAND2_X1 U10072 ( .A1(n9357), .A2(n7233), .ZN(n7232) );
  NAND2_X1 U10073 ( .A1(n7511), .A2(n7510), .ZN(n7509) );
  NAND2_X1 U10074 ( .A1(n15966), .A2(n15965), .ZN(n15964) );
  NOR2_X1 U10075 ( .A1(n12973), .A2(n11585), .ZN(n11427) );
  INV_X1 U10076 ( .A(n7840), .ZN(n7839) );
  NAND2_X1 U10077 ( .A1(n7259), .A2(n7869), .ZN(n7865) );
  NAND3_X1 U10078 ( .A1(n11826), .A2(n11825), .A3(n7763), .ZN(n12289) );
  INV_X1 U10079 ( .A(n15632), .ZN(n7511) );
  AOI21_X2 U10080 ( .B1(n14622), .B2(n9676), .A(n6616), .ZN(n14607) );
  NAND2_X1 U10081 ( .A1(n9726), .A2(n7526), .ZN(n7524) );
  NAND2_X1 U10082 ( .A1(n11634), .A2(n7939), .ZN(n11802) );
  MUX2_X1 U10083 ( .A(n13644), .B(n13919), .S(n15995), .Z(n13647) );
  NAND2_X1 U10084 ( .A1(n11430), .A2(n11429), .ZN(n11634) );
  NAND2_X1 U10085 ( .A1(n6591), .A2(n6726), .ZN(n10306) );
  NAND2_X1 U10086 ( .A1(n7572), .A2(n7571), .ZN(n9261) );
  NAND3_X1 U10087 ( .A1(n6731), .A2(n10250), .A3(n10293), .ZN(n10300) );
  NAND3_X1 U10088 ( .A1(n7244), .A2(n7603), .A3(n8982), .ZN(n7602) );
  NAND2_X1 U10089 ( .A1(n8983), .A2(n8984), .ZN(n7244) );
  INV_X2 U10090 ( .A(n8933), .ZN(n9020) );
  OAI21_X2 U10091 ( .B1(n9122), .B2(n8711), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8713) );
  INV_X2 U10092 ( .A(n9273), .ZN(n9252) );
  NAND2_X1 U10093 ( .A1(n11871), .A2(n11870), .ZN(n11872) );
  AOI21_X1 U10094 ( .B1(n13594), .B2(n13593), .A(n13592), .ZN(n13619) );
  INV_X1 U10095 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8055) );
  OAI211_X1 U10096 ( .C1(n12523), .C2(n7957), .A(n6738), .B(n7956), .ZN(n7955)
         );
  INV_X1 U10097 ( .A(n7955), .ZN(n13800) );
  OR2_X2 U10098 ( .A1(n13650), .A2(n13649), .ZN(n13651) );
  NAND2_X1 U10099 ( .A1(n7589), .A2(n7588), .ZN(n7587) );
  NOR2_X1 U10100 ( .A1(n8944), .A2(n8610), .ZN(n8612) );
  OAI21_X1 U10101 ( .B1(n8615), .B2(n8607), .A(n8606), .ZN(n8608) );
  INV_X1 U10102 ( .A(n13717), .ZN(n7259) );
  NAND2_X1 U10103 ( .A1(n7924), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8067) );
  NAND3_X2 U10104 ( .A1(n7923), .A2(n7922), .A3(n8063), .ZN(n7924) );
  NAND2_X1 U10105 ( .A1(n7848), .A2(n6715), .ZN(n12897) );
  XNOR2_X1 U10106 ( .A(n12135), .B(n12145), .ZN(n11888) );
  NAND2_X1 U10107 ( .A1(n12139), .A2(n12140), .ZN(n13465) );
  XNOR2_X2 U10108 ( .A(n8185), .B(n8184), .ZN(n11185) );
  NAND2_X1 U10109 ( .A1(n13033), .A2(n13032), .ZN(n7262) );
  NAND3_X1 U10110 ( .A1(n13099), .A2(n13098), .A3(n13728), .ZN(n13105) );
  NAND3_X1 U10111 ( .A1(n13066), .A2(n13065), .A3(n7265), .ZN(n7264) );
  OAI21_X1 U10112 ( .B1(n13021), .B2(n13020), .A(n6721), .ZN(n13026) );
  OR2_X1 U10113 ( .A1(n12950), .A2(n10516), .ZN(n8153) );
  OAI21_X1 U10114 ( .B1(n13117), .B2(n13118), .A(n7267), .ZN(n7266) );
  NAND2_X1 U10115 ( .A1(n13129), .A2(n7268), .ZN(n13130) );
  OAI21_X1 U10116 ( .B1(n13138), .B2(n7391), .A(n7270), .ZN(n7269) );
  NOR2_X1 U10117 ( .A1(n9484), .A2(n12902), .ZN(n14352) );
  NOR2_X1 U10118 ( .A1(n10405), .A2(n9484), .ZN(n7272) );
  NOR2_X1 U10119 ( .A1(n9484), .A2(P2_U3088), .ZN(n7274) );
  AND2_X1 U10120 ( .A1(n7278), .A2(n6563), .ZN(n7276) );
  INV_X1 U10121 ( .A(n7901), .ZN(n7289) );
  AND3_X1 U10122 ( .A1(n7292), .A2(n7290), .A3(n7291), .ZN(n12235) );
  NAND2_X1 U10123 ( .A1(n9823), .A2(n7293), .ZN(n7290) );
  NAND3_X1 U10124 ( .A1(n7893), .A2(n7894), .A3(n9441), .ZN(n9876) );
  MUX2_X1 U10125 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n11028), .S(n14231), .Z(
        n14237) );
  NAND2_X1 U10126 ( .A1(n7306), .A2(n7307), .ZN(n11602) );
  NAND2_X1 U10127 ( .A1(n11119), .A2(n7309), .ZN(n7306) );
  NAND2_X1 U10128 ( .A1(n8113), .A2(n8112), .ZN(n8467) );
  NAND2_X1 U10129 ( .A1(n7340), .A2(n7339), .ZN(n13602) );
  NAND2_X1 U10130 ( .A1(n13540), .A2(n7342), .ZN(n7339) );
  INV_X1 U10131 ( .A(n11297), .ZN(n7360) );
  NAND2_X1 U10132 ( .A1(n7362), .A2(n11297), .ZN(n7356) );
  AOI21_X1 U10133 ( .B1(n11297), .B2(n11296), .A(n11295), .ZN(n11299) );
  INV_X1 U10134 ( .A(n11296), .ZN(n7373) );
  NAND2_X1 U10135 ( .A1(n7377), .A2(n8592), .ZN(P3_U3154) );
  NAND2_X1 U10136 ( .A1(n7378), .A2(n13437), .ZN(n7377) );
  NAND2_X1 U10137 ( .A1(n12924), .A2(n7379), .ZN(n7378) );
  OR2_X1 U10138 ( .A1(n8530), .A2(n8531), .ZN(n7379) );
  NAND2_X1 U10139 ( .A1(n8530), .A2(n8531), .ZN(n12924) );
  INV_X1 U10140 ( .A(n7381), .ZN(n13317) );
  NAND2_X1 U10141 ( .A1(n7382), .A2(n7383), .ZN(n7906) );
  NAND2_X1 U10142 ( .A1(n12193), .A2(n7384), .ZN(n7382) );
  NAND2_X1 U10143 ( .A1(n11630), .A2(n10908), .ZN(n12995) );
  NAND2_X4 U10144 ( .A1(n7390), .A2(n7392), .ZN(n8332) );
  NAND2_X1 U10145 ( .A1(n7905), .A2(n7397), .ZN(n7396) );
  INV_X1 U10146 ( .A(n7401), .ZN(n13435) );
  NOR2_X2 U10147 ( .A1(n11365), .A2(n11364), .ZN(n11363) );
  OAI21_X1 U10148 ( .B1(n14404), .B2(n7410), .A(n7408), .ZN(n14380) );
  OAI21_X1 U10149 ( .B1(n8619), .B2(SI_8_), .A(n7411), .ZN(n8620) );
  NAND3_X1 U10150 ( .A1(n7747), .A2(n8629), .A3(n8624), .ZN(n7415) );
  INV_X1 U10151 ( .A(n8629), .ZN(n7417) );
  NAND3_X1 U10152 ( .A1(n6574), .A2(n7524), .A3(n14470), .ZN(n14467) );
  NAND2_X2 U10153 ( .A1(n7418), .A2(n12695), .ZN(n15375) );
  NAND2_X1 U10154 ( .A1(n7422), .A2(n7420), .ZN(n12025) );
  NAND4_X1 U10155 ( .A1(n7814), .A2(n7424), .A3(n11755), .A4(n12007), .ZN(
        n7422) );
  NAND3_X1 U10156 ( .A1(n7814), .A2(n7424), .A3(n11755), .ZN(n12005) );
  AND2_X1 U10157 ( .A1(n8717), .A2(n7426), .ZN(n7425) );
  NAND2_X1 U10158 ( .A1(n15258), .A2(n7431), .ZN(n7430) );
  NAND2_X2 U10159 ( .A1(n7430), .A2(n7429), .ZN(n15473) );
  AOI21_X2 U10160 ( .B1(n7431), .B2(n7433), .A(n12734), .ZN(n7429) );
  OAI21_X2 U10161 ( .B1(n15330), .B2(n7441), .A(n7438), .ZN(n15281) );
  OAI21_X1 U10162 ( .B1(n15472), .B2(n6762), .A(n7449), .ZN(P1_U3523) );
  OAI21_X1 U10163 ( .B1(n15472), .B2(n15433), .A(n6718), .ZN(n15468) );
  NAND2_X1 U10164 ( .A1(n10239), .A2(n7457), .ZN(n7456) );
  NAND3_X1 U10165 ( .A1(n7456), .A2(n8001), .A3(n7455), .ZN(n10352) );
  INV_X1 U10166 ( .A(n10238), .ZN(n7468) );
  NAND3_X1 U10167 ( .A1(n7770), .A2(n7773), .A3(n7471), .ZN(n7472) );
  NAND2_X1 U10168 ( .A1(n7472), .A2(n7473), .ZN(n7793) );
  NAND2_X1 U10169 ( .A1(n10208), .A2(n7479), .ZN(n7478) );
  NAND3_X1 U10170 ( .A1(n10179), .A2(n10180), .A3(n10187), .ZN(n10185) );
  INV_X2 U10171 ( .A(n9507), .ZN(n9727) );
  XNOR2_X2 U10172 ( .A(n9442), .B(n9455), .ZN(n9484) );
  OAI21_X1 U10173 ( .B1(n10196), .B2(n7483), .A(n7482), .ZN(n7776) );
  NOR2_X1 U10174 ( .A1(n6613), .A2(n7484), .ZN(n7483) );
  INV_X1 U10175 ( .A(n10195), .ZN(n7484) );
  NAND2_X1 U10176 ( .A1(n15607), .A2(n15608), .ZN(n10830) );
  NAND2_X1 U10177 ( .A1(n15605), .A2(n15606), .ZN(n7497) );
  INV_X1 U10178 ( .A(n10843), .ZN(n7499) );
  NAND3_X1 U10179 ( .A1(n10566), .A2(n15669), .A3(n10567), .ZN(n16025) );
  NAND2_X1 U10180 ( .A1(n7506), .A2(n7505), .ZN(n16026) );
  INV_X1 U10181 ( .A(n15655), .ZN(n7513) );
  OAI21_X1 U10182 ( .B1(n15655), .B2(n7515), .A(n7514), .ZN(n7516) );
  OR2_X1 U10183 ( .A1(n15654), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n7514) );
  NOR2_X1 U10184 ( .A1(n15653), .A2(n15656), .ZN(n7515) );
  XNOR2_X1 U10185 ( .A(n7516), .B(n15665), .ZN(SUB_1596_U4) );
  NAND2_X1 U10186 ( .A1(n12591), .A2(n12590), .ZN(n15610) );
  NAND2_X2 U10187 ( .A1(n9461), .A2(n13279), .ZN(n9861) );
  NAND2_X1 U10188 ( .A1(n9461), .A2(n7531), .ZN(n9498) );
  OAI21_X1 U10189 ( .B1(n12782), .B2(n7541), .A(n6599), .ZN(n14054) );
  NAND2_X1 U10190 ( .A1(n7542), .A2(n6717), .ZN(n12767) );
  NAND3_X1 U10191 ( .A1(n7544), .A2(n7545), .A3(n7547), .ZN(n7543) );
  NAND2_X1 U10192 ( .A1(n12849), .A2(n6727), .ZN(n14157) );
  NAND2_X1 U10193 ( .A1(n9099), .A2(n6713), .ZN(n7554) );
  NAND3_X1 U10194 ( .A1(n7555), .A2(n7558), .A3(n6625), .ZN(n7553) );
  AND2_X1 U10195 ( .A1(n10293), .A2(n6735), .ZN(n10283) );
  NAND2_X1 U10196 ( .A1(n7564), .A2(n9289), .ZN(n7560) );
  NAND2_X2 U10197 ( .A1(n7560), .A2(n9794), .ZN(n14695) );
  INV_X1 U10198 ( .A(n7562), .ZN(n7561) );
  OAI21_X1 U10199 ( .B1(n9289), .B2(n7563), .A(n10339), .ZN(n7562) );
  NAND2_X1 U10200 ( .A1(n8663), .A2(n11812), .ZN(n7571) );
  OAI21_X2 U10201 ( .B1(n11874), .B2(n7578), .A(n7576), .ZN(n13469) );
  INV_X1 U10202 ( .A(n11470), .ZN(n7579) );
  AOI21_X1 U10203 ( .B1(n11252), .B2(n7583), .A(n6781), .ZN(n7582) );
  INV_X1 U10204 ( .A(n11337), .ZN(n7585) );
  INV_X1 U10205 ( .A(n8790), .ZN(n8788) );
  NAND2_X1 U10206 ( .A1(n8830), .A2(n8829), .ZN(n8832) );
  NOR2_X1 U10207 ( .A1(n7592), .A2(n7591), .ZN(n7590) );
  NAND2_X1 U10208 ( .A1(n9140), .A2(n7594), .ZN(n7593) );
  NAND2_X1 U10209 ( .A1(n7605), .A2(n7601), .ZN(n7603) );
  NAND3_X1 U10210 ( .A1(n8986), .A2(n8985), .A3(n7603), .ZN(n7604) );
  NAND2_X1 U10211 ( .A1(n7606), .A2(n7608), .ZN(n9318) );
  NAND2_X1 U10212 ( .A1(n9267), .A2(n7613), .ZN(n7610) );
  NAND2_X1 U10213 ( .A1(n7610), .A2(n7611), .ZN(n9284) );
  AOI21_X1 U10214 ( .B1(n6568), .B2(n7613), .A(n7612), .ZN(n7611) );
  NAND2_X1 U10215 ( .A1(n15932), .A2(n12398), .ZN(n7616) );
  NOR2_X2 U10216 ( .A1(n12186), .A2(n7616), .ZN(n12321) );
  NAND2_X1 U10217 ( .A1(n14359), .A2(n7617), .ZN(n7618) );
  NAND2_X1 U10218 ( .A1(n14359), .A2(n14686), .ZN(n14358) );
  INV_X1 U10219 ( .A(n7618), .ZN(n14335) );
  NAND2_X1 U10220 ( .A1(n14343), .A2(n14337), .ZN(n14679) );
  NAND3_X1 U10221 ( .A1(n9865), .A2(n12241), .A3(n14823), .ZN(n14659) );
  AND3_X2 U10222 ( .A1(n7620), .A2(n9865), .A3(n12241), .ZN(n9867) );
  INV_X2 U10223 ( .A(n8933), .ZN(n9076) );
  NAND2_X1 U10224 ( .A1(n9481), .A2(n9417), .ZN(n9509) );
  INV_X1 U10225 ( .A(n15429), .ZN(n11495) );
  NAND2_X1 U10226 ( .A1(n15428), .A2(n15429), .ZN(n15427) );
  NAND2_X1 U10227 ( .A1(n10985), .A2(n15439), .ZN(n11506) );
  NAND2_X1 U10228 ( .A1(n11710), .A2(n11709), .ZN(n7630) );
  OAI21_X1 U10229 ( .B1(n11709), .B2(n7632), .A(n11753), .ZN(n7631) );
  NAND2_X1 U10230 ( .A1(n12735), .A2(n7634), .ZN(n7633) );
  CLKBUF_X1 U10231 ( .A(n7641), .Z(n7639) );
  INV_X1 U10232 ( .A(n7639), .ZN(n15315) );
  NAND2_X1 U10233 ( .A1(n15500), .A2(n13194), .ZN(n7654) );
  CLKBUF_X1 U10234 ( .A(n7658), .Z(n7655) );
  NAND2_X1 U10235 ( .A1(n8249), .A2(n7681), .ZN(n7678) );
  NAND2_X1 U10236 ( .A1(n12870), .A2(n7691), .ZN(n7688) );
  OR2_X1 U10237 ( .A1(n12870), .A2(n12869), .ZN(n7693) );
  OR2_X1 U10238 ( .A1(n8502), .A2(n8501), .ZN(n8504) );
  AND2_X1 U10239 ( .A1(n11216), .A2(n11217), .ZN(n7707) );
  NAND2_X1 U10240 ( .A1(n14926), .A2(n7714), .ZN(n7712) );
  NAND2_X1 U10241 ( .A1(n14926), .A2(n7718), .ZN(n7713) );
  NAND2_X1 U10242 ( .A1(n13213), .A2(n13214), .ZN(n7720) );
  NAND2_X1 U10243 ( .A1(n11915), .A2(n6593), .ZN(n12417) );
  NAND2_X1 U10244 ( .A1(n7721), .A2(n7722), .ZN(n14942) );
  NAND2_X1 U10245 ( .A1(n8714), .A2(n6585), .ZN(n8707) );
  NAND2_X1 U10246 ( .A1(n8714), .A2(n6734), .ZN(n7728) );
  INV_X1 U10247 ( .A(n7733), .ZN(n13165) );
  NAND2_X1 U10248 ( .A1(n7735), .A2(n10501), .ZN(n8919) );
  MUX2_X1 U10249 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n8069), .Z(n8609) );
  NAND2_X1 U10250 ( .A1(n9815), .A2(n9856), .ZN(n14345) );
  NAND3_X1 U10251 ( .A1(n7744), .A2(n14357), .A3(n7876), .ZN(n14789) );
  NAND3_X1 U10252 ( .A1(n7738), .A2(n7740), .A3(n7736), .ZN(n14684) );
  NAND3_X1 U10253 ( .A1(n7738), .A2(n7737), .A3(n7736), .ZN(n7744) );
  NAND2_X1 U10254 ( .A1(n15604), .A2(n15603), .ZN(n7757) );
  NAND2_X1 U10255 ( .A1(n10561), .A2(n10539), .ZN(n10540) );
  NAND2_X1 U10256 ( .A1(n11826), .A2(n11825), .ZN(n11832) );
  NAND2_X1 U10257 ( .A1(n7766), .A2(n7767), .ZN(n11625) );
  NAND2_X1 U10258 ( .A1(n7766), .A2(n7764), .ZN(n11824) );
  NAND2_X1 U10259 ( .A1(n11324), .A2(n11323), .ZN(n11617) );
  OR2_X1 U10260 ( .A1(n11324), .A2(n11323), .ZN(n11618) );
  INV_X1 U10261 ( .A(n10200), .ZN(n7771) );
  NAND2_X1 U10262 ( .A1(n7775), .A2(n7774), .ZN(n7773) );
  INV_X1 U10263 ( .A(n10199), .ZN(n7774) );
  NAND2_X1 U10264 ( .A1(n7776), .A2(n10200), .ZN(n7775) );
  OR2_X1 U10265 ( .A1(n10218), .A2(n7782), .ZN(n7781) );
  NAND3_X1 U10266 ( .A1(n7781), .A2(n7780), .A3(n7779), .ZN(n7777) );
  NAND3_X1 U10267 ( .A1(n7781), .A2(n7779), .A3(n7778), .ZN(n10224) );
  NAND2_X1 U10268 ( .A1(n7793), .A2(n7794), .ZN(n10208) );
  INV_X1 U10269 ( .A(n10206), .ZN(n7795) );
  INV_X2 U10270 ( .A(n10194), .ZN(n10232) );
  NAND4_X1 U10271 ( .A1(n7796), .A2(n9419), .A3(n9418), .A4(n9625), .ZN(n9707)
         );
  NAND2_X1 U10272 ( .A1(n9625), .A2(n7983), .ZN(n9422) );
  NOR2_X1 U10273 ( .A1(n9577), .A2(n7798), .ZN(n9694) );
  NAND3_X1 U10274 ( .A1(n9625), .A2(n9438), .A3(n7983), .ZN(n7798) );
  NAND2_X1 U10275 ( .A1(n15375), .A2(n7801), .ZN(n7800) );
  NAND3_X1 U10276 ( .A1(n7813), .A2(n11747), .A3(n7812), .ZN(n11749) );
  NAND2_X1 U10277 ( .A1(n7817), .A2(n11518), .ZN(n7812) );
  NAND2_X1 U10278 ( .A1(n11519), .A2(n7817), .ZN(n7813) );
  NAND2_X1 U10279 ( .A1(n7815), .A2(n11747), .ZN(n7814) );
  NAND2_X1 U10280 ( .A1(n7819), .A2(n11747), .ZN(n7816) );
  NAND2_X1 U10281 ( .A1(n8753), .A2(n13276), .ZN(n8863) );
  XNOR2_X2 U10282 ( .A(n7823), .B(n10123), .ZN(n13276) );
  NAND2_X1 U10283 ( .A1(n6736), .A2(n12165), .ZN(n15415) );
  NAND3_X1 U10284 ( .A1(n8251), .A2(n7834), .A3(n8250), .ZN(n8252) );
  NAND2_X1 U10285 ( .A1(n11584), .A2(n7839), .ZN(n7837) );
  OAI21_X1 U10286 ( .B1(n11584), .B2(n7841), .A(n7839), .ZN(n11798) );
  OAI21_X1 U10287 ( .B1(n13634), .B2(n7847), .A(n7845), .ZN(n12964) );
  NAND2_X1 U10288 ( .A1(n7844), .A2(n6725), .ZN(n12968) );
  NAND2_X1 U10289 ( .A1(n13634), .A2(n7845), .ZN(n7844) );
  OAI21_X1 U10290 ( .B1(n13717), .B2(n12971), .A(n13106), .ZN(n13701) );
  OAI211_X1 U10291 ( .C1(n7875), .C2(n14684), .A(n7873), .B(n7872), .ZN(
        P2_U3496) );
  NAND2_X1 U10292 ( .A1(n14357), .A2(n14356), .ZN(n14688) );
  NAND2_X1 U10293 ( .A1(n7879), .A2(n7880), .ZN(n14349) );
  NAND2_X1 U10294 ( .A1(n14377), .A2(n7881), .ZN(n7879) );
  INV_X1 U10295 ( .A(n7890), .ZN(n7889) );
  NAND2_X1 U10296 ( .A1(n12254), .A2(n6630), .ZN(n7891) );
  NAND3_X1 U10297 ( .A1(n9441), .A2(n7895), .A3(n9626), .ZN(n13265) );
  NAND3_X1 U10298 ( .A1(n8216), .A2(n10853), .A3(n8196), .ZN(n7908) );
  NAND2_X1 U10299 ( .A1(n7918), .A2(n10155), .ZN(n10157) );
  OAI211_X1 U10300 ( .C1(n13288), .C2(n7920), .A(n7919), .B(n13437), .ZN(
        n10165) );
  OR2_X1 U10301 ( .A1(n13288), .A2(n13720), .ZN(n13290) );
  OAI21_X1 U10302 ( .B1(n11363), .B2(n7931), .A(n7929), .ZN(n11845) );
  NOR2_X1 U10303 ( .A1(n11363), .A2(n7936), .ZN(n11662) );
  OR2_X1 U10304 ( .A1(n8247), .A2(n11851), .ZN(n7935) );
  NAND2_X1 U10305 ( .A1(n13016), .A2(n7938), .ZN(n13010) );
  NAND2_X1 U10306 ( .A1(n15964), .A2(n7938), .ZN(n10902) );
  NAND2_X1 U10308 ( .A1(n12858), .A2(n7948), .ZN(n7945) );
  NAND2_X1 U10309 ( .A1(n8066), .A2(n7952), .ZN(n8123) );
  NAND3_X1 U10310 ( .A1(n8120), .A2(n8064), .A3(n7954), .ZN(n7953) );
  NAND3_X1 U10311 ( .A1(n7964), .A2(n7965), .A3(n7962), .ZN(n7961) );
  OAI211_X1 U10312 ( .C1(n13650), .C2(n7975), .A(n7973), .B(n7971), .ZN(n12882) );
  NAND2_X1 U10313 ( .A1(n13650), .A2(n7972), .ZN(n7971) );
  AND2_X1 U10314 ( .A1(n12926), .A2(n12868), .ZN(n7972) );
  OAI21_X1 U10315 ( .B1(n12926), .B2(n7977), .A(n7974), .ZN(n7973) );
  OAI21_X1 U10316 ( .B1(n12926), .B2(n12868), .A(n7977), .ZN(n7974) );
  NAND2_X1 U10317 ( .A1(n13651), .A2(n12868), .ZN(n13638) );
  NAND2_X2 U10318 ( .A1(n9507), .A2(n7176), .ZN(n9793) );
  NAND2_X1 U10319 ( .A1(n13462), .A2(n15972), .ZN(n13014) );
  NAND2_X1 U10320 ( .A1(n9433), .A2(n11551), .ZN(n10482) );
  OAI211_X1 U10321 ( .C1(n13671), .C2(n15988), .A(n13670), .B(n13669), .ZN(
        n13854) );
  INV_X1 U10322 ( .A(n8919), .ZN(n8610) );
  OR2_X1 U10323 ( .A1(n10657), .A2(n9793), .ZN(n9615) );
  AND2_X1 U10324 ( .A1(n12447), .A2(n14890), .ZN(n12448) );
  NAND2_X1 U10325 ( .A1(n8615), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8595) );
  AOI21_X1 U10326 ( .B1(n16013), .B2(n13855), .A(n13854), .ZN(n13931) );
  INV_X1 U10327 ( .A(n15751), .ZN(n10950) );
  OR2_X1 U10328 ( .A1(n15220), .A2(n9295), .ZN(n9302) );
  OR2_X1 U10329 ( .A1(n15262), .A2(n9295), .ZN(n9242) );
  INV_X1 U10330 ( .A(n15469), .ZN(n15161) );
  NAND4_X4 U10331 ( .A1(n8867), .A2(n8866), .A3(n8865), .A4(n8864), .ZN(n15751) );
  OR2_X1 U10332 ( .A1(n8863), .A2(n8862), .ZN(n8865) );
  NAND2_X1 U10333 ( .A1(n15467), .A2(n8002), .ZN(n15566) );
  NAND2_X1 U10334 ( .A1(n15343), .A2(n15327), .ZN(n15318) );
  INV_X1 U10335 ( .A(n15205), .ZN(n15203) );
  NAND2_X1 U10336 ( .A1(n15454), .A2(n15835), .ZN(n15455) );
  XNOR2_X1 U10337 ( .A(n15155), .B(n15148), .ZN(n15149) );
  NAND2_X1 U10338 ( .A1(n10173), .A2(n10172), .ZN(n10183) );
  NAND2_X2 U10339 ( .A1(n12699), .A2(n12698), .ZN(n15330) );
  XNOR2_X1 U10340 ( .A(n15982), .B(n8332), .ZN(n8161) );
  NAND2_X1 U10341 ( .A1(n10401), .A2(n10378), .ZN(n10402) );
  NAND2_X2 U10342 ( .A1(n8843), .A2(n6542), .ZN(n8898) );
  OAI211_X2 U10343 ( .C1(n7252), .C2(n10521), .A(n8223), .B(n8222), .ZN(n15959) );
  XNOR2_X1 U10344 ( .A(n14349), .B(n14348), .ZN(n14350) );
  INV_X1 U10345 ( .A(n13255), .ZN(n8128) );
  INV_X1 U10346 ( .A(n14586), .ZN(n9705) );
  NOR3_X1 U10347 ( .A1(n9388), .A2(n12011), .A3(n11755), .ZN(n7978) );
  AND2_X1 U10348 ( .A1(n12571), .A2(n12437), .ZN(n7980) );
  AND2_X1 U10349 ( .A1(n12721), .A2(n12720), .ZN(n7981) );
  OR2_X1 U10350 ( .A1(n13422), .A2(n6960), .ZN(n7984) );
  OR2_X1 U10351 ( .A1(n15162), .A2(n15181), .ZN(n7985) );
  OR2_X1 U10352 ( .A1(n15161), .A2(n15213), .ZN(n7986) );
  AND2_X1 U10353 ( .A1(n13185), .A2(n13184), .ZN(n7987) );
  AND2_X1 U10354 ( .A1(n12811), .A2(n12810), .ZN(n7989) );
  AND2_X1 U10355 ( .A1(n10360), .A2(n10351), .ZN(n7991) );
  INV_X1 U10356 ( .A(n14444), .ZN(n9843) );
  AND3_X1 U10357 ( .A1(n9367), .A2(n9342), .A3(n9371), .ZN(n7992) );
  INV_X1 U10358 ( .A(n14197), .ZN(n14169) );
  NAND2_X1 U10359 ( .A1(n9205), .A2(n9204), .ZN(n15002) );
  INV_X1 U10360 ( .A(n15002), .ZN(n12727) );
  INV_X1 U10361 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n8607) );
  INV_X1 U10362 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n8698) );
  INV_X1 U10363 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n8594) );
  INV_X1 U10364 ( .A(n12979), .ZN(n13045) );
  INV_X1 U10365 ( .A(P3_B_REG_SCAN_IN), .ZN(n8086) );
  OR2_X1 U10366 ( .A1(n8232), .A2(n12059), .ZN(n7993) );
  AND2_X1 U10367 ( .A1(n13330), .A2(n13454), .ZN(n7995) );
  AND2_X1 U10368 ( .A1(n12962), .A2(n13599), .ZN(n7996) );
  OR2_X1 U10369 ( .A1(n15355), .A2(n12719), .ZN(n7999) );
  AND2_X1 U10370 ( .A1(n10873), .A2(n10872), .ZN(n8000) );
  INV_X1 U10371 ( .A(n14695), .ZN(n14401) );
  AND4_X1 U10372 ( .A1(n10319), .A2(n10318), .A3(n10317), .A4(n10316), .ZN(
        n8001) );
  AND2_X1 U10373 ( .A1(n9855), .A2(n9854), .ZN(n14634) );
  INV_X1 U10374 ( .A(n14634), .ZN(n14657) );
  AND2_X1 U10375 ( .A1(n15466), .A2(n15465), .ZN(n8002) );
  AND2_X1 U10376 ( .A1(n14552), .A2(n14563), .ZN(n8003) );
  OAI21_X1 U10377 ( .B1(n10183), .B2(n10176), .A(n10175), .ZN(n10186) );
  OAI21_X1 U10378 ( .B1(n8961), .B2(n8960), .A(n8959), .ZN(n8970) );
  INV_X1 U10379 ( .A(n8984), .ZN(n8985) );
  OAI22_X1 U10380 ( .A1(n12366), .A2(n10340), .B1(n12329), .B2(n10339), .ZN(
        n10212) );
  INV_X1 U10381 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9417) );
  NOR2_X1 U10382 ( .A1(n9151), .A2(SI_18_), .ZN(n8650) );
  INV_X1 U10383 ( .A(n13198), .ZN(n13199) );
  NAND2_X1 U10384 ( .A1(n13189), .A2(n8869), .ZN(n10873) );
  INV_X1 U10385 ( .A(n15334), .ZN(n12720) );
  OR2_X1 U10386 ( .A1(n8175), .A2(n7338), .ZN(n8158) );
  INV_X1 U10387 ( .A(n15967), .ZN(n10901) );
  MUX2_X1 U10388 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9443), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n9444) );
  NAND2_X1 U10389 ( .A1(n13200), .A2(n13199), .ZN(n13201) );
  INV_X1 U10390 ( .A(n9179), .ZN(n8748) );
  INV_X1 U10391 ( .A(n9093), .ZN(n8747) );
  INV_X1 U10392 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n8971) );
  NAND2_X1 U10393 ( .A1(n15488), .A2(n12731), .ZN(n12732) );
  NAND2_X1 U10394 ( .A1(n11505), .A2(n11504), .ZN(n15428) );
  INV_X1 U10395 ( .A(n13498), .ZN(n13488) );
  INV_X1 U10396 ( .A(n13448), .ZN(n13655) );
  INV_X1 U10397 ( .A(n10907), .ZN(n12976) );
  INV_X1 U10398 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n8010) );
  AND2_X1 U10399 ( .A1(n9898), .A2(n15902), .ZN(n10490) );
  INV_X1 U10400 ( .A(n12349), .ZN(n10443) );
  INV_X1 U10401 ( .A(n10377), .ZN(n10378) );
  INV_X1 U10402 ( .A(n9716), .ZN(n9879) );
  OR2_X1 U10403 ( .A1(n9235), .A2(n14862), .ZN(n9250) );
  NAND2_X1 U10404 ( .A1(n10987), .A2(n10989), .ZN(n10990) );
  OR2_X1 U10405 ( .A1(n13206), .A2(n13205), .ZN(n13207) );
  NAND2_X1 U10406 ( .A1(n8749), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9235) );
  INV_X1 U10407 ( .A(n11908), .ZN(n13233) );
  INV_X1 U10408 ( .A(n9293), .ZN(n8751) );
  NAND2_X1 U10409 ( .A1(n8750), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U10410 ( .A1(n8748), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n9199) );
  INV_X1 U10411 ( .A(n15462), .ZN(n15162) );
  NAND2_X1 U10412 ( .A1(n7829), .A2(n15009), .ZN(n12711) );
  NAND2_X1 U10413 ( .A1(n8625), .A2(n10580), .ZN(n8772) );
  OR2_X1 U10414 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n10833), .ZN(n10834) );
  INV_X1 U10415 ( .A(n13829), .ZN(n13284) );
  INV_X1 U10416 ( .A(n11848), .ZN(n13303) );
  INV_X1 U10417 ( .A(n13455), .ZN(n13407) );
  INV_X1 U10418 ( .A(n13430), .ZN(n13441) );
  NAND2_X1 U10419 ( .A1(n12261), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8177) );
  OR2_X1 U10420 ( .A1(n11157), .A2(n11141), .ZN(n11148) );
  INV_X1 U10421 ( .A(n13091), .ZN(n12893) );
  AND2_X1 U10422 ( .A1(n13016), .A2(n13015), .ZN(n10907) );
  AND2_X1 U10423 ( .A1(n10451), .A2(n10448), .ZN(n12333) );
  INV_X1 U10424 ( .A(n12657), .ZN(n10462) );
  INV_X1 U10425 ( .A(n10405), .ZN(n10485) );
  AND2_X1 U10426 ( .A1(n15914), .A2(n10491), .ZN(n11682) );
  INV_X1 U10427 ( .A(n15894), .ZN(n14306) );
  INV_X1 U10428 ( .A(n14428), .ZN(n14423) );
  INV_X1 U10429 ( .A(n14203), .ZN(n14594) );
  OR2_X1 U10430 ( .A1(n11022), .A2(n9478), .ZN(n14636) );
  INV_X1 U10431 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9904) );
  INV_X1 U10432 ( .A(n10994), .ZN(n10995) );
  NOR2_X1 U10433 ( .A1(n13240), .A2(n14994), .ZN(n13241) );
  OR2_X1 U10434 ( .A1(n9199), .A2(n14879), .ZN(n9216) );
  XNOR2_X1 U10435 ( .A(n13228), .B(n11908), .ZN(n13230) );
  INV_X1 U10436 ( .A(n9273), .ZN(n8887) );
  INV_X1 U10437 ( .A(n15152), .ZN(n15148) );
  NAND2_X1 U10438 ( .A1(n15201), .A2(n15200), .ZN(n15205) );
  NAND2_X1 U10439 ( .A1(n12709), .A2(n12736), .ZN(n12710) );
  INV_X1 U10440 ( .A(n12714), .ZN(n15376) );
  NAND2_X1 U10441 ( .A1(n8991), .A2(n9333), .ZN(n8997) );
  INV_X1 U10442 ( .A(n10870), .ZN(n15742) );
  OAI21_X1 U10443 ( .B1(n8590), .B2(n13446), .A(n8589), .ZN(n8591) );
  AND2_X1 U10444 ( .A1(n8571), .A2(n10912), .ZN(n13430) );
  NOR2_X1 U10445 ( .A1(n15997), .A2(n15956), .ZN(n13837) );
  AND2_X1 U10446 ( .A1(n13911), .A2(n16007), .ZN(n13902) );
  AND2_X1 U10447 ( .A1(n11376), .A2(n11375), .ZN(n11395) );
  INV_X1 U10448 ( .A(n13997), .ZN(n13981) );
  OR2_X1 U10449 ( .A1(n15969), .A2(n16013), .ZN(n16007) );
  AND2_X1 U10450 ( .A1(n8535), .A2(n8534), .ZN(n11387) );
  INV_X1 U10452 ( .A(n14823), .ZN(n14151) );
  INV_X1 U10453 ( .A(n14173), .ZN(n14189) );
  AND3_X1 U10454 ( .A1(n9725), .A2(n9724), .A3(n9723), .ZN(n14563) );
  AND2_X1 U10455 ( .A1(n11047), .A2(n11046), .ZN(n15894) );
  INV_X1 U10456 ( .A(n14330), .ZN(n15892) );
  INV_X1 U10457 ( .A(n10392), .ZN(n14561) );
  INV_X1 U10458 ( .A(n14636), .ZN(n14652) );
  INV_X1 U10459 ( .A(n10391), .ZN(n12504) );
  INV_X1 U10460 ( .A(n15932), .ZN(n12350) );
  INV_X1 U10461 ( .A(n15917), .ZN(n12114) );
  INV_X1 U10462 ( .A(n14781), .ZN(n14682) );
  INV_X1 U10463 ( .A(n15910), .ZN(n12371) );
  INV_X1 U10464 ( .A(n14774), .ZN(n15929) );
  INV_X1 U10465 ( .A(n15931), .ZN(n14770) );
  AND2_X1 U10466 ( .A1(n9897), .A2(n9896), .ZN(n15902) );
  NAND2_X1 U10467 ( .A1(n13265), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9458) );
  AND2_X1 U10468 ( .A1(n10997), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14928) );
  AND2_X1 U10469 ( .A1(n10974), .A2(n15813), .ZN(n14992) );
  OR2_X1 U10470 ( .A1(n14900), .A2(n9295), .ZN(n9278) );
  INV_X1 U10471 ( .A(n15102), .ZN(n15723) );
  INV_X1 U10472 ( .A(n15142), .ZN(n15724) );
  INV_X1 U10473 ( .A(n15754), .ZN(n15829) );
  INV_X1 U10474 ( .A(n15835), .ZN(n15801) );
  AND2_X1 U10475 ( .A1(n10957), .A2(n10532), .ZN(n10955) );
  AND2_X1 U10476 ( .A1(n11157), .A2(n11156), .ZN(n15945) );
  INV_X1 U10477 ( .A(n10163), .ZN(n10164) );
  INV_X1 U10478 ( .A(n13437), .ZN(n13413) );
  AND2_X1 U10479 ( .A1(n12945), .A2(n12267), .ZN(n12958) );
  INV_X1 U10480 ( .A(n13773), .ZN(n13801) );
  INV_X1 U10481 ( .A(n13463), .ZN(n13461) );
  INV_X1 U10482 ( .A(n13615), .ZN(n13586) );
  INV_X1 U10483 ( .A(n15958), .ZN(n13825) );
  INV_X1 U10484 ( .A(n13837), .ZN(n13807) );
  NAND3_X1 U10485 ( .A1(n11396), .A2(n11395), .A3(n11394), .ZN(n16023) );
  AND2_X1 U10486 ( .A1(n10921), .A2(n10920), .ZN(n16018) );
  INV_X1 U10487 ( .A(SI_10_), .ZN(n10578) );
  INV_X1 U10488 ( .A(SI_4_), .ZN(n10501) );
  INV_X1 U10489 ( .A(n14700), .ZN(n14415) );
  OR2_X1 U10490 ( .A1(n14147), .A2(n14638), .ZN(n14184) );
  NAND2_X1 U10491 ( .A1(n10486), .A2(n10479), .ZN(n14154) );
  INV_X1 U10492 ( .A(n10407), .ZN(n10408) );
  INV_X1 U10493 ( .A(n14089), .ZN(n14576) );
  INV_X1 U10494 ( .A(n14066), .ZN(n14653) );
  NAND2_X1 U10495 ( .A1(n14645), .A2(n11977), .ZN(n14664) );
  AND2_X1 U10496 ( .A1(n14554), .A2(n11986), .ZN(n14669) );
  INV_X1 U10497 ( .A(n15944), .ZN(n15941) );
  INV_X1 U10498 ( .A(n10367), .ZN(n14788) );
  INV_X1 U10499 ( .A(n14818), .ZN(n15938) );
  NAND2_X1 U10500 ( .A1(n14818), .A2(n14770), .ZN(n14822) );
  INV_X1 U10501 ( .A(n15907), .ZN(n15908) );
  XNOR2_X1 U10502 ( .A(n9873), .B(n9872), .ZN(n12225) );
  INV_X1 U10503 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10769) );
  OR2_X1 U10504 ( .A1(n9412), .A2(n10644), .ZN(n9413) );
  NAND2_X1 U10505 ( .A1(n9330), .A2(n9329), .ZN(n15181) );
  INV_X1 U10506 ( .A(n15321), .ZN(n15359) );
  INV_X1 U10507 ( .A(n15383), .ZN(n15423) );
  OR2_X1 U10508 ( .A1(n10969), .A2(n10968), .ZN(n15836) );
  INV_X1 U10509 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10775) );
  INV_X1 U10510 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10651) );
  NAND2_X1 U10511 ( .A1(n8010), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8011) );
  NAND2_X1 U10512 ( .A1(n10583), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8013) );
  XNOR2_X1 U10513 ( .A(n10618), .B(P1_DATAO_REG_8__SCAN_IN), .ZN(n8248) );
  INV_X1 U10514 ( .A(n8248), .ZN(n8015) );
  NAND2_X1 U10515 ( .A1(n10618), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8016) );
  NAND2_X1 U10516 ( .A1(n8281), .A2(n8280), .ZN(n8018) );
  NAND2_X1 U10517 ( .A1(n10655), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8017) );
  NAND2_X1 U10518 ( .A1(n8301), .A2(n8300), .ZN(n8020) );
  NAND2_X1 U10519 ( .A1(n7257), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8019) );
  XNOR2_X1 U10520 ( .A(n7199), .B(P1_DATAO_REG_12__SCAN_IN), .ZN(n8313) );
  INV_X1 U10521 ( .A(n8313), .ZN(n8021) );
  NAND2_X1 U10522 ( .A1(n7199), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8022) );
  INV_X1 U10523 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10778) );
  NAND2_X1 U10524 ( .A1(n10778), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8023) );
  INV_X1 U10525 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10648) );
  NOR2_X1 U10526 ( .A1(n10648), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n8024) );
  INV_X1 U10527 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10777) );
  AOI22_X1 U10528 ( .A1(n8024), .A2(n8023), .B1(P1_DATAO_REG_14__SCAN_IN), 
        .B2(n10777), .ZN(n8025) );
  XNOR2_X1 U10529 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n8359) );
  INV_X1 U10530 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n8026) );
  NAND2_X1 U10531 ( .A1(n8026), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8027) );
  XNOR2_X1 U10532 ( .A(n10769), .B(P2_DATAO_REG_16__SCAN_IN), .ZN(n8379) );
  INV_X1 U10533 ( .A(n8379), .ZN(n8028) );
  INV_X1 U10534 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10771) );
  NAND2_X1 U10535 ( .A1(n10771), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8029) );
  XNOR2_X1 U10536 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .ZN(n8386) );
  INV_X1 U10537 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11004) );
  XNOR2_X1 U10538 ( .A(n11004), .B(P2_DATAO_REG_18__SCAN_IN), .ZN(n8402) );
  INV_X1 U10539 ( .A(n8402), .ZN(n8030) );
  NAND2_X1 U10540 ( .A1(n8403), .A2(n8030), .ZN(n8032) );
  INV_X1 U10541 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11006) );
  NAND2_X1 U10542 ( .A1(n11006), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8031) );
  INV_X1 U10543 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11347) );
  XNOR2_X1 U10544 ( .A(n11347), .B(P1_DATAO_REG_19__SCAN_IN), .ZN(n8419) );
  INV_X1 U10545 ( .A(n8419), .ZN(n8033) );
  NAND2_X1 U10546 ( .A1(n11347), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8034) );
  INV_X1 U10547 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11552) );
  NAND2_X1 U10548 ( .A1(n11552), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8038) );
  INV_X1 U10549 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11311) );
  NAND2_X1 U10550 ( .A1(n11311), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8036) );
  AND2_X1 U10551 ( .A1(n8038), .A2(n8036), .ZN(n8037) );
  INV_X1 U10552 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n12825) );
  AND2_X1 U10553 ( .A1(n12825), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8039) );
  INV_X1 U10554 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12749) );
  AOI22_X1 U10555 ( .A1(n8039), .A2(n8038), .B1(P1_DATAO_REG_21__SCAN_IN), 
        .B2(n12749), .ZN(n8040) );
  INV_X1 U10556 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11726) );
  NAND2_X1 U10557 ( .A1(n11726), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8043) );
  INV_X1 U10558 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8658) );
  NAND2_X1 U10559 ( .A1(n8658), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8042) );
  NAND2_X1 U10560 ( .A1(n8043), .A2(n8042), .ZN(n8461) );
  INV_X1 U10561 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8660) );
  NAND2_X1 U10562 ( .A1(n8660), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8045) );
  INV_X1 U10563 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n9232) );
  NAND2_X1 U10564 ( .A1(n9232), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8044) );
  AND2_X1 U10565 ( .A1(n8045), .A2(n8044), .ZN(n8474) );
  INV_X1 U10566 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12221) );
  NAND2_X1 U10567 ( .A1(n8488), .A2(n12221), .ZN(n8048) );
  INV_X1 U10568 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12223) );
  INV_X1 U10569 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12479) );
  NAND2_X1 U10570 ( .A1(n12479), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8050) );
  INV_X1 U10571 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12482) );
  NAND2_X1 U10572 ( .A1(n12482), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8049) );
  NAND2_X1 U10573 ( .A1(n8050), .A2(n8049), .ZN(n8501) );
  INV_X1 U10574 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n12485) );
  INV_X1 U10575 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n12483) );
  XNOR2_X1 U10576 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n8051) );
  XNOR2_X1 U10577 ( .A(n12827), .B(n8051), .ZN(n12394) );
  NOR2_X1 U10578 ( .A1(P3_IR_REG_26__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), 
        .ZN(n8058) );
  XNOR2_X2 U10579 ( .A(n8065), .B(n8120), .ZN(n12879) );
  INV_X1 U10580 ( .A(SI_27_), .ZN(n12395) );
  OR2_X1 U10581 ( .A1(n7252), .A2(n12395), .ZN(n8070) );
  INV_X1 U10582 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8073) );
  NAND2_X1 U10583 ( .A1(n8102), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8077) );
  MUX2_X1 U10584 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8077), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8078) );
  INV_X1 U10585 ( .A(n8328), .ZN(n8556) );
  NAND2_X1 U10586 ( .A1(n8072), .A2(n8079), .ZN(n8555) );
  OR2_X1 U10587 ( .A1(n8555), .A2(P3_IR_REG_23__SCAN_IN), .ZN(n8081) );
  XNOR2_X1 U10588 ( .A(P3_IR_REG_24__SCAN_IN), .B(P3_IR_REG_31__SCAN_IN), .ZN(
        n8080) );
  INV_X1 U10589 ( .A(n8555), .ZN(n8084) );
  INV_X1 U10590 ( .A(n8315), .ZN(n8083) );
  NAND3_X1 U10591 ( .A1(n8084), .A2(n8083), .A3(n8082), .ZN(n8088) );
  NAND2_X1 U10592 ( .A1(n8088), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8087) );
  XNOR2_X1 U10593 ( .A(n8087), .B(P3_IR_REG_25__SCAN_IN), .ZN(n8563) );
  INV_X1 U10594 ( .A(n8563), .ZN(n8091) );
  OAI21_X1 U10595 ( .B1(n8088), .B2(P3_IR_REG_25__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8090) );
  INV_X1 U10596 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8089) );
  XNOR2_X1 U10597 ( .A(n8090), .B(n8089), .ZN(n12288) );
  AOI21_X1 U10598 ( .B1(n8092), .B2(n8091), .A(n12288), .ZN(n8532) );
  INV_X1 U10599 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n8093) );
  NAND2_X1 U10600 ( .A1(n8532), .A2(n8093), .ZN(n8096) );
  INV_X1 U10601 ( .A(n8094), .ZN(n11814) );
  NAND2_X1 U10602 ( .A1(n12288), .A2(n11814), .ZN(n8095) );
  INV_X1 U10603 ( .A(n8098), .ZN(n8099) );
  NAND2_X1 U10604 ( .A1(n8099), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8100) );
  MUX2_X1 U10605 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8100), .S(
        P3_IR_REG_19__SCAN_IN), .Z(n8101) );
  XNOR2_X1 U10606 ( .A(n13927), .B(n12911), .ZN(n12918) );
  INV_X1 U10607 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n8107) );
  INV_X1 U10608 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8108) );
  INV_X1 U10609 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n8110) );
  INV_X1 U10610 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8112) );
  INV_X1 U10611 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n8114) );
  INV_X1 U10612 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n9957) );
  INV_X1 U10613 ( .A(n8523), .ZN(n8118) );
  INV_X1 U10614 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8117) );
  NAND2_X1 U10615 ( .A1(n8523), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8119) );
  NAND2_X1 U10616 ( .A1(n8572), .A2(n8119), .ZN(n13659) );
  INV_X1 U10617 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8121) );
  INV_X1 U10618 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n14002) );
  NAND2_X1 U10619 ( .A1(n8123), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8124) );
  INV_X1 U10620 ( .A(n8125), .ZN(n14001) );
  INV_X1 U10621 ( .A(n14008), .ZN(n8127) );
  NAND2_X1 U10622 ( .A1(n13659), .A2(n6551), .ZN(n8133) );
  INV_X1 U10623 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n13851) );
  AND2_X4 U10624 ( .A1(n13255), .A2(n14008), .ZN(n12261) );
  NAND2_X1 U10625 ( .A1(n12261), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8130) );
  NAND2_X1 U10626 ( .A1(n12939), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8129) );
  OAI211_X1 U10627 ( .C1(n13851), .C2(n12264), .A(n8130), .B(n8129), .ZN(n8131) );
  INV_X1 U10628 ( .A(n8131), .ZN(n8132) );
  NOR2_X1 U10629 ( .A1(n12918), .A2(n13666), .ZN(n12914) );
  AOI21_X1 U10630 ( .B1(n12918), .B2(n13666), .A(n12914), .ZN(n8531) );
  XNOR2_X1 U10631 ( .A(n8135), .B(n8134), .ZN(n10503) );
  OR2_X1 U10632 ( .A1(n12950), .A2(n10503), .ZN(n8143) );
  OR2_X1 U10633 ( .A1(n12951), .A2(SI_5_), .ZN(n8142) );
  INV_X1 U10634 ( .A(n8202), .ZN(n8138) );
  INV_X1 U10635 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8137) );
  NAND2_X1 U10636 ( .A1(n8138), .A2(n8137), .ZN(n8220) );
  NAND2_X1 U10637 ( .A1(n8220), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8140) );
  INV_X1 U10638 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8139) );
  XNOR2_X1 U10639 ( .A(n8140), .B(n8139), .ZN(n11217) );
  NAND2_X1 U10640 ( .A1(n6538), .A2(n11217), .ZN(n8141) );
  XNOR2_X1 U10641 ( .A(n8332), .B(n16012), .ZN(n8217) );
  NAND2_X1 U10642 ( .A1(n8209), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8144) );
  NAND2_X1 U10643 ( .A1(n8224), .A2(n8144), .ZN(n11416) );
  NAND2_X1 U10644 ( .A1(n6549), .A2(n11416), .ZN(n8149) );
  NAND2_X1 U10645 ( .A1(n12938), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8148) );
  OR2_X1 U10646 ( .A1(n6548), .A2(n7583), .ZN(n8147) );
  INV_X1 U10647 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n8145) );
  OR2_X1 U10648 ( .A1(n6545), .A2(n8145), .ZN(n8146) );
  INV_X1 U10649 ( .A(SI_1_), .ZN(n10517) );
  OR2_X1 U10650 ( .A1(n12951), .A2(n10517), .ZN(n8155) );
  NAND2_X1 U10651 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n8150) );
  XNOR2_X1 U10652 ( .A(n8168), .B(n8152), .ZN(n10516) );
  NAND2_X1 U10653 ( .A1(n12261), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8157) );
  NAND2_X1 U10654 ( .A1(n8174), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8156) );
  NOR2_X1 U10655 ( .A1(n8161), .A2(n8170), .ZN(n8172) );
  NOR3_X1 U10656 ( .A1(n10860), .A2(n8332), .A3(n15982), .ZN(n8162) );
  NOR2_X1 U10657 ( .A1(n8172), .A2(n8162), .ZN(n10863) );
  NAND2_X1 U10658 ( .A1(n12261), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8166) );
  NAND2_X1 U10659 ( .A1(n8174), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8165) );
  NAND2_X1 U10660 ( .A1(n12938), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8164) );
  INV_X1 U10661 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11149) );
  OR2_X1 U10662 ( .A1(n6547), .A2(n11149), .ZN(n8163) );
  NAND4_X1 U10663 ( .A1(n8166), .A2(n8165), .A3(n8164), .A4(n8163), .ZN(n13464) );
  INV_X1 U10664 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8845) );
  NAND2_X1 U10665 ( .A1(n8845), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8167) );
  AND2_X1 U10666 ( .A1(n8168), .A2(n8167), .ZN(n8169) );
  INV_X1 U10667 ( .A(SI_0_), .ZN(n8844) );
  MUX2_X1 U10668 ( .A(n8169), .B(n8844), .S(n6542), .Z(n10499) );
  MUX2_X1 U10669 ( .A(n11165), .B(n10499), .S(n8136), .Z(n11399) );
  INV_X1 U10670 ( .A(n11399), .ZN(n12677) );
  INV_X1 U10671 ( .A(n10904), .ZN(n15986) );
  NAND2_X1 U10672 ( .A1(n15980), .A2(n13008), .ZN(n10899) );
  NAND2_X1 U10673 ( .A1(n10899), .A2(n8332), .ZN(n8171) );
  NAND3_X1 U10674 ( .A1(n10863), .A2(n15986), .A3(n8171), .ZN(n10862) );
  INV_X1 U10675 ( .A(n8172), .ZN(n8173) );
  NAND2_X1 U10676 ( .A1(n10862), .A2(n8173), .ZN(n10854) );
  NAND2_X1 U10677 ( .A1(n8174), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8179) );
  NAND2_X1 U10678 ( .A1(n12938), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8178) );
  INV_X1 U10679 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15979) );
  OR2_X1 U10680 ( .A1(n6547), .A2(n15979), .ZN(n8176) );
  XNOR2_X1 U10681 ( .A(n10900), .B(n8332), .ZN(n8195) );
  XNOR2_X1 U10682 ( .A(n13462), .B(n8195), .ZN(n10855) );
  NAND2_X1 U10683 ( .A1(n10854), .A2(n10855), .ZN(n10853) );
  OR2_X1 U10684 ( .A1(n12951), .A2(SI_3_), .ZN(n8188) );
  XNOR2_X1 U10685 ( .A(n8183), .B(n8182), .ZN(n10507) );
  OR2_X1 U10686 ( .A1(n12950), .A2(n10507), .ZN(n8187) );
  NAND2_X1 U10687 ( .A1(n8253), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8185) );
  INV_X1 U10688 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8184) );
  NAND2_X1 U10689 ( .A1(n6538), .A2(n11185), .ZN(n8186) );
  XNOR2_X1 U10690 ( .A(n8332), .B(n10929), .ZN(n8197) );
  NAND2_X1 U10691 ( .A1(n6549), .A2(n8189), .ZN(n8194) );
  NAND2_X1 U10692 ( .A1(n12938), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8193) );
  INV_X1 U10693 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n8190) );
  OR2_X1 U10694 ( .A1(n6545), .A2(n8190), .ZN(n8192) );
  INV_X1 U10695 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11130) );
  OR2_X1 U10696 ( .A1(n6548), .A2(n11130), .ZN(n8191) );
  XNOR2_X1 U10697 ( .A(n8197), .B(n10901), .ZN(n10925) );
  NAND2_X1 U10698 ( .A1(n8195), .A2(n15991), .ZN(n10926) );
  INV_X1 U10699 ( .A(n8197), .ZN(n8198) );
  XNOR2_X1 U10700 ( .A(n8201), .B(n8200), .ZN(n10500) );
  OR2_X1 U10701 ( .A1(n12950), .A2(n10500), .ZN(n8207) );
  OR2_X1 U10702 ( .A1(n12951), .A2(SI_4_), .ZN(n8206) );
  NAND2_X1 U10703 ( .A1(n8202), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8203) );
  MUX2_X1 U10704 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8203), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n8204) );
  NAND2_X1 U10705 ( .A1(n6537), .A2(n11302), .ZN(n8205) );
  XNOR2_X1 U10706 ( .A(n8332), .B(n16006), .ZN(n8215) );
  NAND2_X1 U10707 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8208) );
  NAND2_X1 U10708 ( .A1(n8209), .A2(n8208), .ZN(n11460) );
  NAND2_X1 U10709 ( .A1(n6549), .A2(n11460), .ZN(n8214) );
  NAND2_X1 U10710 ( .A1(n12938), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8213) );
  INV_X1 U10711 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11459) );
  OR2_X1 U10712 ( .A1(n6548), .A2(n11459), .ZN(n8212) );
  INV_X1 U10713 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n8210) );
  NAND2_X1 U10714 ( .A1(n8215), .A2(n11408), .ZN(n8216) );
  OAI21_X1 U10715 ( .B1(n8215), .B2(n11408), .A(n8216), .ZN(n11104) );
  XNOR2_X1 U10716 ( .A(n8217), .B(n11664), .ZN(n11364) );
  INV_X1 U10717 ( .A(SI_6_), .ZN(n10521) );
  XNOR2_X1 U10718 ( .A(n10527), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8218) );
  XNOR2_X1 U10719 ( .A(n8219), .B(n8218), .ZN(n10522) );
  OR2_X1 U10720 ( .A1(n10522), .A2(n12950), .ZN(n8223) );
  XNOR2_X2 U10721 ( .A(n8221), .B(P3_IR_REG_6__SCAN_IN), .ZN(n11258) );
  NAND2_X1 U10722 ( .A1(n6538), .A2(n11258), .ZN(n8222) );
  XNOR2_X1 U10723 ( .A(n8332), .B(n11667), .ZN(n8231) );
  NAND2_X1 U10724 ( .A1(n8224), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8225) );
  NAND2_X1 U10725 ( .A1(n8240), .A2(n8225), .ZN(n15957) );
  NAND2_X1 U10726 ( .A1(n8174), .A2(n15957), .ZN(n8230) );
  NAND2_X1 U10727 ( .A1(n12938), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8229) );
  INV_X1 U10728 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n8226) );
  OR2_X1 U10729 ( .A1(n6545), .A2(n8226), .ZN(n8228) );
  INV_X1 U10730 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n15962) );
  XNOR2_X1 U10731 ( .A(n8231), .B(n12059), .ZN(n11661) );
  INV_X1 U10732 ( .A(n8231), .ZN(n8232) );
  XNOR2_X1 U10733 ( .A(n8234), .B(n8233), .ZN(n10577) );
  NAND2_X1 U10734 ( .A1(n10577), .A2(n12935), .ZN(n8239) );
  INV_X1 U10735 ( .A(SI_7_), .ZN(n10576) );
  OAI21_X1 U10736 ( .B1(n8235), .B2(P3_IR_REG_6__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8237) );
  INV_X1 U10737 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8236) );
  XNOR2_X1 U10738 ( .A(n8237), .B(n8236), .ZN(n11327) );
  AOI22_X1 U10739 ( .A1(n7065), .A2(n10576), .B1(n6538), .B2(n11327), .ZN(
        n8238) );
  XNOR2_X1 U10740 ( .A(n8332), .B(n15950), .ZN(n8247) );
  NAND2_X1 U10741 ( .A1(n8240), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8241) );
  NAND2_X1 U10742 ( .A1(n8257), .A2(n8241), .ZN(n15949) );
  NAND2_X1 U10743 ( .A1(n6549), .A2(n15949), .ZN(n8246) );
  NAND2_X1 U10744 ( .A1(n12938), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8245) );
  OR2_X1 U10745 ( .A1(n6548), .A2(n7586), .ZN(n8244) );
  INV_X1 U10746 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n8242) );
  OR2_X1 U10747 ( .A1(n6545), .A2(n8242), .ZN(n8243) );
  XNOR2_X1 U10748 ( .A(n8247), .B(n11851), .ZN(n12063) );
  XNOR2_X1 U10749 ( .A(n8249), .B(n8248), .ZN(n10518) );
  NAND2_X1 U10750 ( .A1(n10518), .A2(n12935), .ZN(n8256) );
  INV_X1 U10751 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8250) );
  OR2_X1 U10752 ( .A1(n8253), .A2(n8252), .ZN(n8267) );
  NAND2_X1 U10753 ( .A1(n8267), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8254) );
  XNOR2_X1 U10754 ( .A(n8254), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11464) );
  AOI22_X1 U10755 ( .A1(n7065), .A2(SI_8_), .B1(n6538), .B2(n11464), .ZN(n8255) );
  XNOR2_X1 U10756 ( .A(n11800), .B(n8332), .ZN(n8264) );
  NAND2_X1 U10757 ( .A1(n12939), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8263) );
  NAND2_X1 U10758 ( .A1(n8257), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8258) );
  NAND2_X1 U10759 ( .A1(n8273), .A2(n8258), .ZN(n11846) );
  NAND2_X1 U10760 ( .A1(n6549), .A2(n11846), .ZN(n8262) );
  NAND2_X1 U10761 ( .A1(n12938), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8261) );
  INV_X1 U10762 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n8259) );
  OR2_X1 U10763 ( .A1(n6545), .A2(n8259), .ZN(n8260) );
  NAND4_X1 U10764 ( .A1(n8263), .A2(n8262), .A3(n8261), .A4(n8260), .ZN(n13456) );
  XNOR2_X1 U10765 ( .A(n8264), .B(n12198), .ZN(n11844) );
  XNOR2_X1 U10766 ( .A(n8266), .B(n8265), .ZN(n10515) );
  NAND2_X1 U10767 ( .A1(n10515), .A2(n12935), .ZN(n8272) );
  INV_X1 U10768 ( .A(SI_9_), .ZN(n10514) );
  INV_X1 U10769 ( .A(n8267), .ZN(n8269) );
  INV_X1 U10770 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8268) );
  NAND2_X1 U10771 ( .A1(n8269), .A2(n8268), .ZN(n8282) );
  NAND2_X1 U10772 ( .A1(n8282), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8270) );
  INV_X1 U10773 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8283) );
  XNOR2_X1 U10774 ( .A(n8270), .B(n8283), .ZN(n11483) );
  AOI22_X1 U10775 ( .A1(n7065), .A2(n10514), .B1(n6538), .B2(n11483), .ZN(
        n8271) );
  NAND2_X1 U10776 ( .A1(n8272), .A2(n8271), .ZN(n12203) );
  XNOR2_X1 U10777 ( .A(n12203), .B(n8332), .ZN(n8296) );
  NAND2_X1 U10778 ( .A1(n12939), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8279) );
  NAND2_X1 U10779 ( .A1(n8273), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n8274) );
  NAND2_X1 U10780 ( .A1(n8289), .A2(n8274), .ZN(n12200) );
  NAND2_X1 U10781 ( .A1(n6551), .A2(n12200), .ZN(n8278) );
  NAND2_X1 U10782 ( .A1(n12938), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8277) );
  INV_X1 U10783 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n8275) );
  OR2_X1 U10784 ( .A1(n6545), .A2(n8275), .ZN(n8276) );
  NAND4_X1 U10785 ( .A1(n8279), .A2(n8278), .A3(n8277), .A4(n8276), .ZN(n11848) );
  XNOR2_X1 U10786 ( .A(n8296), .B(n13303), .ZN(n12194) );
  XNOR2_X1 U10787 ( .A(n8281), .B(n8280), .ZN(n10579) );
  NAND2_X1 U10788 ( .A1(n10579), .A2(n12935), .ZN(n8288) );
  INV_X1 U10789 ( .A(n8282), .ZN(n8284) );
  NAND2_X1 U10790 ( .A1(n8284), .A2(n8283), .ZN(n8302) );
  NAND2_X1 U10791 ( .A1(n8302), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8286) );
  INV_X1 U10792 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8285) );
  XNOR2_X1 U10793 ( .A(n8286), .B(n8285), .ZN(n11885) );
  AOI22_X1 U10794 ( .A1(n7065), .A2(n10578), .B1(n6538), .B2(n11885), .ZN(
        n8287) );
  XNOR2_X1 U10795 ( .A(n13308), .B(n8332), .ZN(n8299) );
  NAND2_X1 U10796 ( .A1(n12939), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8295) );
  NAND2_X1 U10797 ( .A1(n8289), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8290) );
  NAND2_X1 U10798 ( .A1(n8307), .A2(n8290), .ZN(n13305) );
  NAND2_X1 U10799 ( .A1(n6551), .A2(n13305), .ZN(n8294) );
  NAND2_X1 U10800 ( .A1(n12938), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8293) );
  INV_X1 U10801 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n8291) );
  OR2_X1 U10802 ( .A1(n6545), .A2(n8291), .ZN(n8292) );
  XNOR2_X1 U10803 ( .A(n8299), .B(n13407), .ZN(n13299) );
  INV_X1 U10804 ( .A(n8296), .ZN(n8297) );
  NAND2_X1 U10805 ( .A1(n8297), .A2(n13303), .ZN(n13296) );
  AND2_X1 U10806 ( .A1(n13299), .A2(n13296), .ZN(n8298) );
  XNOR2_X1 U10807 ( .A(n8301), .B(n8300), .ZN(n10581) );
  NAND2_X1 U10808 ( .A1(n10581), .A2(n12935), .ZN(n8306) );
  INV_X1 U10809 ( .A(SI_11_), .ZN(n10580) );
  OAI21_X1 U10810 ( .B1(n8302), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8303) );
  MUX2_X1 U10811 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8303), .S(
        P3_IR_REG_11__SCAN_IN), .Z(n8304) );
  NAND2_X1 U10812 ( .A1(n8304), .A2(n8315), .ZN(n12145) );
  AOI22_X1 U10813 ( .A1(n7065), .A2(n10580), .B1(n6538), .B2(n12145), .ZN(
        n8305) );
  NAND2_X1 U10814 ( .A1(n8306), .A2(n8305), .ZN(n13408) );
  XNOR2_X1 U10815 ( .A(n13408), .B(n8332), .ZN(n13330) );
  NAND2_X1 U10816 ( .A1(n12939), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8312) );
  NAND2_X1 U10817 ( .A1(n8307), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8308) );
  NAND2_X1 U10818 ( .A1(n6605), .A2(n8308), .ZN(n13411) );
  NAND2_X1 U10819 ( .A1(n6549), .A2(n13411), .ZN(n8311) );
  NAND2_X1 U10820 ( .A1(n12938), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8310) );
  INV_X1 U10821 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n9979) );
  OR2_X1 U10822 ( .A1(n6545), .A2(n9979), .ZN(n8309) );
  NAND4_X1 U10823 ( .A1(n8312), .A2(n8311), .A3(n8310), .A4(n8309), .ZN(n13454) );
  XNOR2_X1 U10824 ( .A(n8314), .B(n8313), .ZN(n10638) );
  NAND2_X1 U10825 ( .A1(n10638), .A2(n12935), .ZN(n8318) );
  NAND2_X1 U10826 ( .A1(n8315), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8316) );
  XNOR2_X1 U10827 ( .A(n8316), .B(P3_IR_REG_12__SCAN_IN), .ZN(n13475) );
  AOI22_X1 U10828 ( .A1(n7065), .A2(SI_12_), .B1(n6538), .B2(n13475), .ZN(
        n8317) );
  XNOR2_X1 U10829 ( .A(n13344), .B(n8332), .ZN(n8325) );
  NAND2_X1 U10830 ( .A1(n6605), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8319) );
  NAND2_X1 U10831 ( .A1(n8333), .A2(n8319), .ZN(n13338) );
  NAND2_X1 U10832 ( .A1(n6551), .A2(n13338), .ZN(n8324) );
  NAND2_X1 U10833 ( .A1(n12938), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8323) );
  INV_X1 U10834 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12495) );
  OR2_X1 U10835 ( .A1(n6547), .A2(n12495), .ZN(n8322) );
  INV_X1 U10836 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n8320) );
  OR2_X1 U10837 ( .A1(n6545), .A2(n8320), .ZN(n8321) );
  NAND2_X1 U10838 ( .A1(n8325), .A2(n13388), .ZN(n13328) );
  OAI21_X1 U10839 ( .B1(n13330), .B2(n13454), .A(n13328), .ZN(n8327) );
  INV_X1 U10840 ( .A(n8325), .ZN(n8326) );
  INV_X1 U10841 ( .A(n13388), .ZN(n13453) );
  NAND2_X1 U10842 ( .A1(n8326), .A2(n13453), .ZN(n13329) );
  XNOR2_X1 U10843 ( .A(n8342), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8341) );
  XNOR2_X1 U10844 ( .A(n8341), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n10660) );
  NAND2_X1 U10845 ( .A1(n10660), .A2(n12935), .ZN(n8331) );
  INV_X1 U10846 ( .A(SI_13_), .ZN(n10659) );
  OR2_X1 U10847 ( .A1(n8328), .A2(n8121), .ZN(n8329) );
  INV_X1 U10848 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8347) );
  XNOR2_X1 U10849 ( .A(n8329), .B(n8347), .ZN(n13486) );
  AOI22_X1 U10850 ( .A1(n7065), .A2(n10659), .B1(n6538), .B2(n13486), .ZN(
        n8330) );
  XNOR2_X1 U10851 ( .A(n13389), .B(n12911), .ZN(n13384) );
  NAND2_X1 U10852 ( .A1(n8333), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8334) );
  NAND2_X1 U10853 ( .A1(n8351), .A2(n8334), .ZN(n13392) );
  NAND2_X1 U10854 ( .A1(n13392), .A2(n8174), .ZN(n8338) );
  NAND2_X1 U10855 ( .A1(n12939), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8337) );
  INV_X1 U10856 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n12533) );
  OR2_X1 U10857 ( .A1(n6545), .A2(n12533), .ZN(n8336) );
  NAND2_X1 U10858 ( .A1(n12938), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8335) );
  NAND2_X1 U10859 ( .A1(n13384), .A2(n13284), .ZN(n8340) );
  NOR2_X1 U10860 ( .A1(n13384), .A2(n13284), .ZN(n8339) );
  NAND2_X1 U10861 ( .A1(n8341), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8344) );
  NAND2_X1 U10862 ( .A1(n8342), .A2(n10651), .ZN(n8343) );
  NAND2_X1 U10863 ( .A1(n8344), .A2(n8343), .ZN(n8346) );
  XNOR2_X1 U10864 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8345) );
  XNOR2_X1 U10865 ( .A(n8346), .B(n8345), .ZN(n10664) );
  NAND2_X1 U10866 ( .A1(n10664), .A2(n12935), .ZN(n8350) );
  INV_X1 U10867 ( .A(SI_14_), .ZN(n10663) );
  AND2_X1 U10868 ( .A1(n8328), .A2(n8347), .ZN(n8362) );
  OR2_X1 U10869 ( .A1(n8362), .A2(n8121), .ZN(n8348) );
  INV_X1 U10870 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8361) );
  XNOR2_X1 U10871 ( .A(n8348), .B(n8361), .ZN(n13508) );
  AOI22_X1 U10872 ( .A1(n7065), .A2(n10663), .B1(n6538), .B2(n13508), .ZN(
        n8349) );
  XNOR2_X1 U10873 ( .A(n13996), .B(n8332), .ZN(n8358) );
  INV_X1 U10874 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13901) );
  NAND2_X1 U10875 ( .A1(n8351), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8352) );
  NAND2_X1 U10876 ( .A1(n8368), .A2(n8352), .ZN(n13823) );
  NAND2_X1 U10877 ( .A1(n13823), .A2(n6551), .ZN(n8356) );
  NAND2_X1 U10878 ( .A1(n12939), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8354) );
  INV_X1 U10879 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13991) );
  OR2_X1 U10880 ( .A1(n6545), .A2(n13991), .ZN(n8353) );
  AND2_X1 U10881 ( .A1(n8354), .A2(n8353), .ZN(n8355) );
  XNOR2_X1 U10882 ( .A(n8358), .B(n13811), .ZN(n13281) );
  INV_X1 U10883 ( .A(n13281), .ZN(n8357) );
  NOR2_X1 U10884 ( .A1(n8358), .A2(n13452), .ZN(n13434) );
  XNOR2_X1 U10885 ( .A(n8360), .B(n8359), .ZN(n10662) );
  NAND2_X1 U10886 ( .A1(n10662), .A2(n12935), .ZN(n8367) );
  INV_X1 U10887 ( .A(SI_15_), .ZN(n10661) );
  NAND2_X1 U10888 ( .A1(n8362), .A2(n8361), .ZN(n8364) );
  NAND2_X1 U10889 ( .A1(n8364), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8363) );
  MUX2_X1 U10890 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8363), .S(
        P3_IR_REG_15__SCAN_IN), .Z(n8365) );
  OR2_X1 U10891 ( .A1(n8364), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n8388) );
  NAND2_X1 U10892 ( .A1(n8365), .A2(n8388), .ZN(n13534) );
  AOI22_X1 U10893 ( .A1(n7065), .A2(n10661), .B1(n13534), .B2(n6538), .ZN(
        n8366) );
  XNOR2_X1 U10894 ( .A(n13817), .B(n8332), .ZN(n8372) );
  INV_X1 U10895 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13898) );
  NAND2_X1 U10896 ( .A1(n8368), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8369) );
  NAND2_X1 U10897 ( .A1(n8374), .A2(n8369), .ZN(n13815) );
  NAND2_X1 U10898 ( .A1(n13815), .A2(n6551), .ZN(n8371) );
  AOI22_X1 U10899 ( .A1(n12939), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n12261), 
        .B2(P3_REG0_REG_15__SCAN_IN), .ZN(n8370) );
  XNOR2_X1 U10900 ( .A(n8372), .B(n13831), .ZN(n13433) );
  NAND2_X1 U10901 ( .A1(n8372), .A2(n13831), .ZN(n8373) );
  NAND2_X1 U10902 ( .A1(n8374), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8375) );
  NAND2_X1 U10903 ( .A1(n8394), .A2(n8375), .ZN(n13804) );
  NAND2_X1 U10904 ( .A1(n13804), .A2(n6551), .ZN(n8378) );
  AOI22_X1 U10905 ( .A1(n12939), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n12261), 
        .B2(P3_REG0_REG_16__SCAN_IN), .ZN(n8377) );
  NAND2_X1 U10906 ( .A1(n12938), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8376) );
  XNOR2_X1 U10907 ( .A(n8380), .B(n8379), .ZN(n10742) );
  NAND2_X1 U10908 ( .A1(n10742), .A2(n12935), .ZN(n8383) );
  NAND2_X1 U10909 ( .A1(n8388), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8381) );
  XNOR2_X1 U10910 ( .A(n8381), .B(P3_IR_REG_16__SCAN_IN), .ZN(n13556) );
  AOI22_X1 U10911 ( .A1(n6538), .A2(n13556), .B1(n7065), .B2(SI_16_), .ZN(
        n8382) );
  XNOR2_X1 U10912 ( .A(n13980), .B(n8332), .ZN(n8384) );
  XOR2_X1 U10913 ( .A(n13812), .B(n8384), .Z(n13359) );
  INV_X1 U10914 ( .A(n8384), .ZN(n8385) );
  INV_X1 U10915 ( .A(n13812), .ZN(n13788) );
  XNOR2_X1 U10916 ( .A(n8387), .B(n8386), .ZN(n10767) );
  NAND2_X1 U10917 ( .A1(n10767), .A2(n12935), .ZN(n8393) );
  INV_X1 U10918 ( .A(n8388), .ZN(n8389) );
  INV_X1 U10919 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n9924) );
  NAND2_X1 U10920 ( .A1(n8389), .A2(n9924), .ZN(n8404) );
  NAND2_X1 U10921 ( .A1(n8404), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8391) );
  INV_X1 U10922 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8390) );
  XNOR2_X1 U10923 ( .A(n8391), .B(n8390), .ZN(n13581) );
  INV_X1 U10924 ( .A(SI_17_), .ZN(n10766) );
  AOI22_X1 U10925 ( .A1(n13581), .A2(n6538), .B1(n7065), .B2(n10766), .ZN(
        n8392) );
  XNOR2_X1 U10926 ( .A(n13974), .B(n8332), .ZN(n8399) );
  NAND2_X1 U10927 ( .A1(n8394), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8395) );
  NAND2_X1 U10928 ( .A1(n8409), .A2(n8395), .ZN(n13792) );
  INV_X1 U10929 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13889) );
  NAND2_X1 U10930 ( .A1(n12261), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8397) );
  NAND2_X1 U10931 ( .A1(n12939), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8396) );
  OAI211_X1 U10932 ( .C1(n13889), .C2(n12264), .A(n8397), .B(n8396), .ZN(n8398) );
  NAND2_X1 U10933 ( .A1(n8399), .A2(n13773), .ZN(n13366) );
  INV_X1 U10934 ( .A(n8399), .ZN(n8400) );
  NAND2_X1 U10935 ( .A1(n8400), .A2(n13801), .ZN(n13367) );
  NAND2_X1 U10936 ( .A1(n8401), .A2(n13367), .ZN(n13417) );
  XNOR2_X1 U10937 ( .A(n8403), .B(n8402), .ZN(n10780) );
  NAND2_X1 U10938 ( .A1(n10780), .A2(n12935), .ZN(n8408) );
  OAI21_X1 U10939 ( .B1(n8404), .B2(P3_IR_REG_17__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8405) );
  XNOR2_X1 U10940 ( .A(n8405), .B(P3_IR_REG_18__SCAN_IN), .ZN(n13607) );
  INV_X1 U10941 ( .A(SI_18_), .ZN(n10781) );
  NOR2_X1 U10942 ( .A1(n7252), .A2(n10781), .ZN(n8406) );
  AOI21_X1 U10943 ( .B1(n13607), .B2(n6538), .A(n8406), .ZN(n8407) );
  XNOR2_X1 U10944 ( .A(n13782), .B(n8332), .ZN(n8416) );
  NAND2_X1 U10945 ( .A1(n8409), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8410) );
  NAND2_X1 U10946 ( .A1(n8423), .A2(n8410), .ZN(n13774) );
  NAND2_X1 U10947 ( .A1(n13774), .A2(n6551), .ZN(n8415) );
  INV_X1 U10948 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13887) );
  NAND2_X1 U10949 ( .A1(n12261), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8412) );
  NAND2_X1 U10950 ( .A1(n12939), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8411) );
  OAI211_X1 U10951 ( .C1(n12264), .C2(n13887), .A(n8412), .B(n8411), .ZN(n8413) );
  INV_X1 U10952 ( .A(n8413), .ZN(n8414) );
  XNOR2_X1 U10953 ( .A(n8416), .B(n13789), .ZN(n13416) );
  INV_X1 U10954 ( .A(n8416), .ZN(n8417) );
  NAND2_X1 U10955 ( .A1(n8417), .A2(n13789), .ZN(n8418) );
  XNOR2_X1 U10956 ( .A(n8420), .B(n8419), .ZN(n10965) );
  NAND2_X1 U10957 ( .A1(n10965), .A2(n12935), .ZN(n8422) );
  INV_X1 U10958 ( .A(n13599), .ZN(n13616) );
  AOI22_X1 U10959 ( .A1(n7065), .A2(SI_19_), .B1(n13616), .B2(n6538), .ZN(
        n8421) );
  XNOR2_X1 U10960 ( .A(n13964), .B(n8332), .ZN(n8430) );
  NAND2_X1 U10961 ( .A1(n8423), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8424) );
  NAND2_X1 U10962 ( .A1(n8435), .A2(n8424), .ZN(n13764) );
  NAND2_X1 U10963 ( .A1(n13764), .A2(n6551), .ZN(n8429) );
  INV_X1 U10964 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13880) );
  NAND2_X1 U10965 ( .A1(n12261), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8426) );
  NAND2_X1 U10966 ( .A1(n12939), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8425) );
  OAI211_X1 U10967 ( .C1(n13880), .C2(n12264), .A(n8426), .B(n8425), .ZN(n8427) );
  INV_X1 U10968 ( .A(n8427), .ZN(n8428) );
  XNOR2_X1 U10969 ( .A(n8430), .B(n13743), .ZN(n13310) );
  INV_X1 U10970 ( .A(n8430), .ZN(n8431) );
  NAND2_X1 U10971 ( .A1(n8431), .A2(n13743), .ZN(n8432) );
  XNOR2_X1 U10972 ( .A(n8443), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n11488) );
  NAND2_X1 U10973 ( .A1(n11488), .A2(n12935), .ZN(n8434) );
  INV_X1 U10974 ( .A(SI_20_), .ZN(n11490) );
  OR2_X1 U10975 ( .A1(n7252), .A2(n11490), .ZN(n8433) );
  XNOR2_X1 U10976 ( .A(n13958), .B(n8332), .ZN(n8442) );
  NAND2_X1 U10977 ( .A1(n8435), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8436) );
  NAND2_X1 U10978 ( .A1(n8451), .A2(n8436), .ZN(n13747) );
  NAND2_X1 U10979 ( .A1(n13747), .A2(n6551), .ZN(n8441) );
  INV_X1 U10980 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13877) );
  NAND2_X1 U10981 ( .A1(n12939), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8438) );
  NAND2_X1 U10982 ( .A1(n12261), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8437) );
  OAI211_X1 U10983 ( .C1(n13877), .C2(n12264), .A(n8438), .B(n8437), .ZN(n8439) );
  INV_X1 U10984 ( .A(n8439), .ZN(n8440) );
  NOR2_X1 U10985 ( .A1(n8442), .A2(n13760), .ZN(n13377) );
  NAND2_X1 U10986 ( .A1(n8443), .A2(n12825), .ZN(n8446) );
  NAND2_X1 U10987 ( .A1(n8444), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8445) );
  NAND2_X1 U10988 ( .A1(n8446), .A2(n8445), .ZN(n8448) );
  XNOR2_X1 U10989 ( .A(n11552), .B(P2_DATAO_REG_21__SCAN_IN), .ZN(n8447) );
  XNOR2_X1 U10990 ( .A(n8448), .B(n8447), .ZN(n11627) );
  NAND2_X1 U10991 ( .A1(n11627), .A2(n12935), .ZN(n8450) );
  INV_X1 U10992 ( .A(SI_21_), .ZN(n11629) );
  OR2_X1 U10993 ( .A1(n7252), .A2(n11629), .ZN(n8449) );
  NAND2_X1 U10994 ( .A1(n8451), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8452) );
  NAND2_X1 U10995 ( .A1(n8467), .A2(n8452), .ZN(n13321) );
  NAND2_X1 U10996 ( .A1(n13321), .A2(n6551), .ZN(n8457) );
  INV_X1 U10997 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n13732) );
  NAND2_X1 U10998 ( .A1(n12938), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8454) );
  NAND2_X1 U10999 ( .A1(n12261), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8453) );
  OAI211_X1 U11000 ( .C1(n6547), .C2(n13732), .A(n8454), .B(n8453), .ZN(n8455)
         );
  INV_X1 U11001 ( .A(n8455), .ZN(n8456) );
  AOI21_X1 U11002 ( .B1(n8458), .B2(n13744), .A(n8459), .ZN(n13319) );
  INV_X1 U11003 ( .A(n8459), .ZN(n8460) );
  NAND2_X1 U11004 ( .A1(n8462), .A2(n8461), .ZN(n8463) );
  NAND2_X1 U11005 ( .A1(n8464), .A2(n8463), .ZN(n11213) );
  NAND2_X1 U11006 ( .A1(n11213), .A2(n12935), .ZN(n8466) );
  OR2_X1 U11007 ( .A1(n7252), .A2(n7230), .ZN(n8465) );
  XNOR2_X1 U11008 ( .A(n13948), .B(n8332), .ZN(n10152) );
  NAND2_X1 U11009 ( .A1(n8467), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8468) );
  NAND2_X1 U11010 ( .A1(n8480), .A2(n8468), .ZN(n13723) );
  NAND2_X1 U11011 ( .A1(n13723), .A2(n6551), .ZN(n8473) );
  INV_X1 U11012 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n13722) );
  NAND2_X1 U11013 ( .A1(n12938), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8470) );
  NAND2_X1 U11014 ( .A1(n12261), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8469) );
  OAI211_X1 U11015 ( .C1(n6548), .C2(n13722), .A(n8470), .B(n8469), .ZN(n8471)
         );
  INV_X1 U11016 ( .A(n8471), .ZN(n8472) );
  OR2_X1 U11017 ( .A1(n8475), .A2(n8474), .ZN(n8476) );
  NAND2_X1 U11018 ( .A1(n8477), .A2(n8476), .ZN(n11613) );
  NAND2_X1 U11019 ( .A1(n11613), .A2(n12935), .ZN(n8479) );
  INV_X1 U11020 ( .A(SI_23_), .ZN(n11615) );
  OR2_X1 U11021 ( .A1(n7252), .A2(n11615), .ZN(n8478) );
  XNOR2_X1 U11022 ( .A(n13710), .B(n8332), .ZN(n10156) );
  NAND2_X1 U11023 ( .A1(n8480), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8481) );
  NAND2_X1 U11024 ( .A1(n8491), .A2(n8481), .ZN(n13711) );
  NAND2_X1 U11025 ( .A1(n13711), .A2(n6551), .ZN(n8486) );
  INV_X1 U11026 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13868) );
  NAND2_X1 U11027 ( .A1(n12939), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8483) );
  NAND2_X1 U11028 ( .A1(n12261), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8482) );
  OAI211_X1 U11029 ( .C1(n13868), .C2(n12264), .A(n8483), .B(n8482), .ZN(n8484) );
  INV_X1 U11030 ( .A(n8484), .ZN(n8485) );
  INV_X1 U11031 ( .A(n13720), .ZN(n13693) );
  AOI22_X1 U11032 ( .A1(n10156), .A2(n13693), .B1(n13731), .B2(n10152), .ZN(
        n8487) );
  INV_X1 U11033 ( .A(n10156), .ZN(n8499) );
  XNOR2_X1 U11034 ( .A(n8488), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n11811) );
  NAND2_X1 U11035 ( .A1(n11811), .A2(n12935), .ZN(n8490) );
  INV_X1 U11036 ( .A(SI_24_), .ZN(n11812) );
  OR2_X1 U11037 ( .A1(n7252), .A2(n11812), .ZN(n8489) );
  XNOR2_X1 U11038 ( .A(n12898), .B(n8332), .ZN(n8498) );
  NAND2_X1 U11039 ( .A1(n8491), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8492) );
  NAND2_X1 U11040 ( .A1(n8507), .A2(n8492), .ZN(n13696) );
  NAND2_X1 U11041 ( .A1(n13696), .A2(n6551), .ZN(n8497) );
  INV_X1 U11042 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13864) );
  NAND2_X1 U11043 ( .A1(n12939), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8494) );
  NAND2_X1 U11044 ( .A1(n12261), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8493) );
  OAI211_X1 U11045 ( .C1(n13864), .C2(n12264), .A(n8494), .B(n8493), .ZN(n8495) );
  INV_X1 U11046 ( .A(n8495), .ZN(n8496) );
  NAND2_X1 U11047 ( .A1(n8498), .A2(n13704), .ZN(n13348) );
  OAI21_X1 U11048 ( .B1(n8498), .B2(n13704), .A(n13348), .ZN(n10158) );
  AOI21_X1 U11049 ( .B1(n8499), .B2(n13720), .A(n10158), .ZN(n8500) );
  NAND2_X1 U11050 ( .A1(n8502), .A2(n8501), .ZN(n8503) );
  NAND2_X1 U11051 ( .A1(n8504), .A2(n8503), .ZN(n11983) );
  NAND2_X1 U11052 ( .A1(n11983), .A2(n12935), .ZN(n8506) );
  INV_X1 U11053 ( .A(SI_25_), .ZN(n11985) );
  OR2_X1 U11054 ( .A1(n7252), .A2(n11985), .ZN(n8505) );
  XNOR2_X1 U11055 ( .A(n13119), .B(n12911), .ZN(n8514) );
  NAND2_X1 U11056 ( .A1(n8507), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8508) );
  NAND2_X1 U11057 ( .A1(n8521), .A2(n8508), .ZN(n13685) );
  NAND2_X1 U11058 ( .A1(n13685), .A2(n6551), .ZN(n8513) );
  INV_X1 U11059 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13860) );
  NAND2_X1 U11060 ( .A1(n12939), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8510) );
  NAND2_X1 U11061 ( .A1(n12261), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8509) );
  OAI211_X1 U11062 ( .C1(n13860), .C2(n12264), .A(n8510), .B(n8509), .ZN(n8511) );
  INV_X1 U11063 ( .A(n8511), .ZN(n8512) );
  NOR2_X1 U11064 ( .A1(n8514), .A2(n13665), .ZN(n8516) );
  AOI21_X1 U11065 ( .B1(n8514), .B2(n13665), .A(n8516), .ZN(n13349) );
  NAND2_X1 U11066 ( .A1(n8515), .A2(n13349), .ZN(n13351) );
  INV_X1 U11067 ( .A(n8516), .ZN(n8517) );
  NAND2_X1 U11068 ( .A1(n13351), .A2(n8517), .ZN(n13424) );
  XNOR2_X1 U11069 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .ZN(n8518) );
  OR2_X1 U11070 ( .A1(n7252), .A2(n12286), .ZN(n8520) );
  XNOR2_X1 U11071 ( .A(n13422), .B(n12911), .ZN(n8527) );
  NAND2_X1 U11072 ( .A1(n8521), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8522) );
  INV_X1 U11073 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13856) );
  NAND2_X1 U11074 ( .A1(n12939), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8525) );
  NAND2_X1 U11075 ( .A1(n12261), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8524) );
  OAI211_X1 U11076 ( .C1(n13856), .C2(n12264), .A(n8525), .B(n8524), .ZN(n8526) );
  NOR2_X1 U11077 ( .A1(n8527), .A2(n6960), .ZN(n8528) );
  AOI21_X1 U11078 ( .B1(n8527), .B2(n6960), .A(n8528), .ZN(n13425) );
  NAND2_X1 U11079 ( .A1(n13424), .A2(n13425), .ZN(n13423) );
  INV_X1 U11080 ( .A(n8528), .ZN(n8529) );
  NAND2_X1 U11081 ( .A1(n13423), .A2(n8529), .ZN(n8530) );
  INV_X1 U11082 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8533) );
  NAND2_X1 U11083 ( .A1(n8532), .A2(n8533), .ZN(n8535) );
  NAND2_X1 U11084 ( .A1(n12288), .A2(n8091), .ZN(n8534) );
  NOR4_X1 U11085 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_27__SCAN_IN), .ZN(n8544) );
  NOR4_X1 U11086 ( .A1(P3_D_REG_24__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n8543) );
  OR4_X1 U11087 ( .A1(P3_D_REG_22__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_17__SCAN_IN), .A4(P3_D_REG_25__SCAN_IN), .ZN(n8541) );
  NOR4_X1 U11088 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n8539) );
  NOR4_X1 U11089 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_11__SCAN_IN), .ZN(n8538) );
  NOR4_X1 U11090 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8537) );
  NOR4_X1 U11091 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n8536) );
  NAND4_X1 U11092 ( .A1(n8539), .A2(n8538), .A3(n8537), .A4(n8536), .ZN(n8540)
         );
  NOR4_X1 U11093 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_2__SCAN_IN), .A3(
        n8541), .A4(n8540), .ZN(n8542) );
  NAND3_X1 U11094 ( .A1(n8544), .A2(n8543), .A3(n8542), .ZN(n8545) );
  NAND2_X1 U11095 ( .A1(n8532), .A2(n8545), .ZN(n11373) );
  NAND3_X1 U11096 ( .A1(n8097), .A2(n11387), .A3(n11373), .ZN(n10914) );
  INV_X1 U11097 ( .A(n10914), .ZN(n10919) );
  NOR2_X1 U11098 ( .A1(n8546), .A2(n10908), .ZN(n11390) );
  OAI21_X1 U11099 ( .B1(n8547), .B2(P3_IR_REG_21__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8548) );
  XNOR2_X1 U11100 ( .A(n11390), .B(n6543), .ZN(n8550) );
  NOR2_X1 U11101 ( .A1(n8546), .A2(n13616), .ZN(n8549) );
  OR2_X1 U11102 ( .A1(n6543), .A2(n8546), .ZN(n15981) );
  NAND3_X1 U11103 ( .A1(n10919), .A2(n10933), .A3(n15981), .ZN(n8554) );
  NAND2_X1 U11104 ( .A1(n11372), .A2(n11373), .ZN(n8551) );
  NOR2_X1 U11105 ( .A1(n8551), .A2(n11387), .ZN(n10912) );
  NAND2_X1 U11106 ( .A1(n6543), .A2(n13616), .ZN(n11389) );
  OR2_X1 U11107 ( .A1(n11389), .A2(n12995), .ZN(n10915) );
  INV_X1 U11108 ( .A(n10915), .ZN(n8552) );
  NAND2_X1 U11109 ( .A1(n10912), .A2(n8552), .ZN(n8553) );
  NAND2_X1 U11110 ( .A1(n8554), .A2(n8553), .ZN(n8565) );
  OR2_X1 U11111 ( .A1(n8556), .A2(n8555), .ZN(n8558) );
  NAND2_X1 U11112 ( .A1(n8558), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8557) );
  MUX2_X1 U11113 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8557), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n8562) );
  INV_X1 U11114 ( .A(n8558), .ZN(n8560) );
  NAND2_X1 U11115 ( .A1(n8560), .A2(n8559), .ZN(n8561) );
  NAND2_X1 U11116 ( .A1(n8562), .A2(n8561), .ZN(n11139) );
  NAND2_X1 U11117 ( .A1(n11139), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10584) );
  INV_X1 U11118 ( .A(n10584), .ZN(n10512) );
  NAND2_X1 U11119 ( .A1(n8563), .A2(n8094), .ZN(n8564) );
  OR2_X1 U11120 ( .A1(n12288), .A2(n8564), .ZN(n10411) );
  NAND2_X1 U11121 ( .A1(n10512), .A2(n10411), .ZN(n11140) );
  INV_X1 U11122 ( .A(n11140), .ZN(n11374) );
  INV_X1 U11123 ( .A(n13927), .ZN(n8590) );
  NOR2_X1 U11124 ( .A1(n15981), .A2(n11140), .ZN(n8566) );
  NAND2_X1 U11125 ( .A1(n10919), .A2(n8566), .ZN(n8568) );
  AND2_X1 U11126 ( .A1(n11492), .A2(n13616), .ZN(n15983) );
  NAND2_X1 U11127 ( .A1(n11374), .A2(n15983), .ZN(n8567) );
  NAND2_X1 U11128 ( .A1(n13146), .A2(n8546), .ZN(n8579) );
  INV_X1 U11129 ( .A(n12879), .ZN(n13142) );
  INV_X1 U11130 ( .A(n13576), .ZN(n13600) );
  NAND2_X1 U11131 ( .A1(n13142), .A2(n13600), .ZN(n11147) );
  NAND2_X1 U11132 ( .A1(n8136), .A2(n11147), .ZN(n10909) );
  INV_X1 U11133 ( .A(n10909), .ZN(n8569) );
  NOR2_X1 U11134 ( .A1(n11140), .A2(n7391), .ZN(n8580) );
  INV_X1 U11135 ( .A(n8580), .ZN(n8570) );
  NOR2_X1 U11136 ( .A1(n15992), .A2(n8570), .ZN(n8571) );
  NAND2_X1 U11137 ( .A1(n8572), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U11138 ( .A1(n13625), .A2(n8573), .ZN(n13645) );
  NAND2_X1 U11139 ( .A1(n13645), .A2(n6551), .ZN(n8578) );
  INV_X1 U11140 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13848) );
  NAND2_X1 U11141 ( .A1(n12939), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8575) );
  NAND2_X1 U11142 ( .A1(n12261), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8574) );
  OAI211_X1 U11143 ( .C1(n13848), .C2(n12264), .A(n8575), .B(n8574), .ZN(n8576) );
  INV_X1 U11144 ( .A(n8576), .ZN(n8577) );
  NAND2_X1 U11145 ( .A1(n13101), .A2(n8580), .ZN(n10917) );
  NOR2_X1 U11146 ( .A1(n10917), .A2(n10909), .ZN(n13143) );
  NAND2_X1 U11147 ( .A1(n13143), .A2(n10912), .ZN(n13428) );
  NAND2_X1 U11148 ( .A1(n10933), .A2(n10914), .ZN(n8583) );
  OAI211_X1 U11149 ( .C1(n13124), .C2(n13139), .A(n10411), .B(n11139), .ZN(
        n8581) );
  INV_X1 U11150 ( .A(n8581), .ZN(n8582) );
  OAI211_X1 U11151 ( .C1(n10912), .C2(n10915), .A(n8583), .B(n8582), .ZN(n8584) );
  NAND2_X1 U11152 ( .A1(n8584), .A2(P3_STATE_REG_SCAN_IN), .ZN(n8586) );
  OR2_X1 U11153 ( .A1(n10912), .A2(n10917), .ZN(n8585) );
  AOI22_X1 U11154 ( .A1(n13659), .A2(n13443), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n8587) );
  OAI21_X1 U11155 ( .B1(n13654), .B2(n13428), .A(n8587), .ZN(n8588) );
  AOI21_X1 U11156 ( .B1(n13430), .B2(n13448), .A(n8588), .ZN(n8589) );
  INV_X1 U11157 ( .A(n8591), .ZN(n8592) );
  INV_X1 U11158 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10572) );
  MUX2_X1 U11159 ( .A(n10572), .B(n8593), .S(n8615), .Z(n8600) );
  INV_X1 U11160 ( .A(SI_2_), .ZN(n10506) );
  NAND2_X1 U11161 ( .A1(n8600), .A2(n10506), .ZN(n8877) );
  INV_X1 U11162 ( .A(n8598), .ZN(n8596) );
  INV_X1 U11163 ( .A(n8874), .ZN(n8599) );
  NAND2_X1 U11164 ( .A1(n8599), .A2(n8877), .ZN(n8602) );
  INV_X1 U11165 ( .A(n8600), .ZN(n8601) );
  NAND2_X1 U11166 ( .A1(n8601), .A2(SI_2_), .ZN(n8876) );
  MUX2_X1 U11167 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n8615), .Z(n8604) );
  NAND2_X1 U11168 ( .A1(n8604), .A2(SI_3_), .ZN(n8917) );
  OAI21_X1 U11169 ( .B1(n8604), .B2(SI_3_), .A(n8917), .ZN(n8894) );
  INV_X1 U11170 ( .A(n8894), .ZN(n8605) );
  NAND2_X1 U11171 ( .A1(n8609), .A2(SI_4_), .ZN(n8942) );
  NAND3_X1 U11172 ( .A1(n8918), .A2(n8917), .A3(n8942), .ZN(n8613) );
  NAND2_X1 U11173 ( .A1(n6541), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8606) );
  OAI21_X1 U11174 ( .B1(n8608), .B2(SI_5_), .A(n8611), .ZN(n8944) );
  MUX2_X1 U11175 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n8615), .Z(n8616) );
  OAI21_X1 U11176 ( .B1(n8616), .B2(SI_7_), .A(n8618), .ZN(n8831) );
  MUX2_X1 U11177 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n6541), .Z(n8619) );
  INV_X1 U11178 ( .A(n8620), .ZN(n8807) );
  MUX2_X1 U11179 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n6541), .Z(n8622) );
  INV_X1 U11180 ( .A(n8978), .ZN(n8623) );
  INV_X1 U11181 ( .A(n8626), .ZN(n8625) );
  INV_X1 U11182 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10658) );
  XNOR2_X1 U11183 ( .A(n8626), .B(SI_11_), .ZN(n9014) );
  INV_X1 U11184 ( .A(n8630), .ZN(n8631) );
  NAND2_X1 U11185 ( .A1(n8631), .A2(n10639), .ZN(n8632) );
  MUX2_X1 U11186 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n7176), .Z(n8633) );
  MUX2_X1 U11187 ( .A(n10777), .B(n10778), .S(n7176), .Z(n9046) );
  NAND2_X1 U11188 ( .A1(n9046), .A2(n10663), .ZN(n9114) );
  MUX2_X1 U11189 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n6542), .Z(n8637) );
  INV_X1 U11190 ( .A(n8637), .ZN(n8636) );
  XNOR2_X1 U11191 ( .A(n8637), .B(SI_15_), .ZN(n9065) );
  NOR2_X1 U11192 ( .A1(n9046), .A2(n10663), .ZN(n8638) );
  INV_X1 U11193 ( .A(n9116), .ZN(n8640) );
  MUX2_X1 U11194 ( .A(n10771), .B(n10769), .S(n7176), .Z(n8642) );
  INV_X1 U11195 ( .A(SI_16_), .ZN(n10743) );
  NAND2_X1 U11196 ( .A1(n8642), .A2(n10743), .ZN(n9098) );
  INV_X1 U11197 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10773) );
  MUX2_X1 U11198 ( .A(n10775), .B(n10773), .S(n6542), .Z(n8644) );
  NAND2_X1 U11199 ( .A1(n8644), .A2(n10766), .ZN(n8643) );
  AND2_X1 U11200 ( .A1(n9098), .A2(n8643), .ZN(n8646) );
  INV_X1 U11201 ( .A(n8643), .ZN(n8645) );
  XNOR2_X1 U11202 ( .A(n8644), .B(SI_17_), .ZN(n9100) );
  MUX2_X1 U11203 ( .A(n11006), .B(n11004), .S(n7176), .Z(n9078) );
  MUX2_X1 U11204 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n7176), .Z(n8648) );
  NAND2_X1 U11205 ( .A1(n8648), .A2(SI_19_), .ZN(n8649) );
  OAI21_X1 U11206 ( .B1(n10781), .B2(n9078), .A(n8649), .ZN(n8647) );
  INV_X1 U11207 ( .A(n9078), .ZN(n9151) );
  INV_X1 U11208 ( .A(SI_19_), .ZN(n10967) );
  INV_X1 U11209 ( .A(n8648), .ZN(n9152) );
  MUX2_X1 U11210 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n6542), .Z(n8654) );
  MUX2_X1 U11211 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n7176), .Z(n9188) );
  NOR2_X1 U11212 ( .A1(n9188), .A2(SI_20_), .ZN(n8652) );
  INV_X1 U11213 ( .A(n8653), .ZN(n9209) );
  NAND3_X1 U11214 ( .A1(n9209), .A2(n9188), .A3(SI_20_), .ZN(n8655) );
  NAND2_X1 U11215 ( .A1(n8654), .A2(SI_21_), .ZN(n9208) );
  MUX2_X1 U11216 ( .A(n8658), .B(n11726), .S(n7176), .Z(n9759) );
  MUX2_X1 U11217 ( .A(n9232), .B(n8660), .S(n6542), .Z(n8661) );
  MUX2_X1 U11218 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n7176), .Z(n9259) );
  MUX2_X1 U11219 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n7176), .Z(n8664) );
  MUX2_X1 U11220 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n7176), .Z(n8665) );
  NAND2_X1 U11221 ( .A1(n8665), .A2(SI_26_), .ZN(n8666) );
  OAI21_X1 U11222 ( .B1(n8665), .B2(SI_26_), .A(n8666), .ZN(n9286) );
  MUX2_X1 U11223 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n7176), .Z(n9312) );
  INV_X1 U11224 ( .A(n9312), .ZN(n8667) );
  NAND2_X1 U11225 ( .A1(n8667), .A2(n12395), .ZN(n8668) );
  NAND2_X1 U11226 ( .A1(n9312), .A2(SI_27_), .ZN(n8669) );
  MUX2_X1 U11227 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n7176), .Z(n8671) );
  INV_X1 U11228 ( .A(n8671), .ZN(n8672) );
  INV_X1 U11229 ( .A(SI_28_), .ZN(n12865) );
  NAND2_X1 U11230 ( .A1(n8672), .A2(n12865), .ZN(n8673) );
  INV_X1 U11231 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15593) );
  INV_X1 U11232 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14827) );
  MUX2_X1 U11233 ( .A(n15593), .B(n14827), .S(n6542), .Z(n8674) );
  INV_X1 U11234 ( .A(SI_29_), .ZN(n14007) );
  NAND2_X1 U11235 ( .A1(n8674), .A2(n14007), .ZN(n8675) );
  INV_X1 U11236 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13277) );
  INV_X1 U11237 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13280) );
  MUX2_X1 U11238 ( .A(n13277), .B(n13280), .S(n7176), .Z(n8676) );
  XNOR2_X1 U11239 ( .A(n8676), .B(SI_30_), .ZN(n8726) );
  INV_X1 U11240 ( .A(n8676), .ZN(n8677) );
  MUX2_X1 U11241 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7176), .Z(n8678) );
  XNOR2_X1 U11242 ( .A(n8678), .B(SI_31_), .ZN(n8679) );
  NAND3_X1 U11243 ( .A1(n8709), .A2(n8705), .A3(n7238), .ZN(n8682) );
  NOR2_X1 U11244 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n8685) );
  NOR2_X1 U11245 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n8688) );
  INV_X1 U11246 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8691) );
  INV_X1 U11247 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8692) );
  XNOR2_X2 U11248 ( .A(n8693), .B(n8692), .ZN(n8855) );
  NAND2_X1 U11249 ( .A1(n6603), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8694) );
  NAND2_X1 U11250 ( .A1(n15583), .A2(n9333), .ZN(n8697) );
  INV_X1 U11251 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9955) );
  OR2_X1 U11252 ( .A1(n8898), .A2(n9955), .ZN(n8696) );
  INV_X1 U11253 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10123) );
  AND2_X2 U11254 ( .A1(n13276), .A2(n15591), .ZN(n8906) );
  NAND2_X1 U11255 ( .A1(n9296), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8704) );
  INV_X1 U11256 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n8701) );
  OR2_X1 U11257 ( .A1(n9308), .A2(n8701), .ZN(n8703) );
  INV_X1 U11258 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n10020) );
  OR2_X1 U11259 ( .A1(n7213), .A2(n10020), .ZN(n8702) );
  AND3_X1 U11260 ( .A1(n8704), .A2(n8703), .A3(n8702), .ZN(n14996) );
  XNOR2_X1 U11261 ( .A(n15152), .B(n14996), .ZN(n9397) );
  NAND3_X1 U11262 ( .A1(n8710), .A2(n8709), .A3(n9918), .ZN(n8711) );
  OR2_X1 U11263 ( .A1(n10871), .A2(n6539), .ZN(n11751) );
  NAND2_X1 U11264 ( .A1(n9067), .A2(n8717), .ZN(n9366) );
  INV_X1 U11265 ( .A(n10807), .ZN(n8718) );
  NAND2_X1 U11266 ( .A1(n8720), .A2(n15598), .ZN(n10944) );
  NAND2_X1 U11267 ( .A1(n8718), .A2(n10944), .ZN(n8719) );
  NAND2_X1 U11268 ( .A1(n11751), .A2(n8719), .ZN(n9404) );
  NOR2_X1 U11269 ( .A1(n9397), .A2(n9404), .ZN(n9359) );
  INV_X1 U11270 ( .A(n8720), .ZN(n10808) );
  NAND2_X1 U11271 ( .A1(n15598), .A2(n15392), .ZN(n10790) );
  NAND2_X1 U11272 ( .A1(n10788), .A2(n15748), .ZN(n8721) );
  NAND2_X1 U11273 ( .A1(n10790), .A2(n8721), .ZN(n8731) );
  INV_X1 U11274 ( .A(n8722), .ZN(n8730) );
  NAND2_X1 U11275 ( .A1(n8720), .A2(n8730), .ZN(n10793) );
  INV_X1 U11276 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8725) );
  NAND2_X1 U11277 ( .A1(n9296), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8724) );
  INV_X1 U11278 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n15156) );
  OR2_X1 U11279 ( .A1(n7213), .A2(n15156), .ZN(n8723) );
  OAI211_X1 U11280 ( .C1(n9308), .C2(n8725), .A(n8724), .B(n8723), .ZN(n15177)
         );
  INV_X1 U11281 ( .A(n15177), .ZN(n8735) );
  AOI21_X1 U11282 ( .B1(n14996), .B2(n8733), .A(n8735), .ZN(n8734) );
  NAND2_X1 U11283 ( .A1(n13275), .A2(n9333), .ZN(n8729) );
  OR2_X1 U11284 ( .A1(n8898), .A2(n13277), .ZN(n8728) );
  NAND2_X1 U11285 ( .A1(n8731), .A2(n8730), .ZN(n8732) );
  MUX2_X1 U11286 ( .A(n8734), .B(n15159), .S(n9076), .Z(n9348) );
  INV_X4 U11287 ( .A(n9076), .ZN(n9344) );
  OR2_X1 U11288 ( .A1(n9131), .A2(n14996), .ZN(n8737) );
  AOI21_X1 U11289 ( .B1(n8737), .B2(n8736), .A(n8735), .ZN(n8738) );
  AOI21_X1 U11290 ( .B1(n15159), .B2(n9344), .A(n8738), .ZN(n9347) );
  NAND2_X1 U11291 ( .A1(n9348), .A2(n9347), .ZN(n9363) );
  NAND2_X1 U11292 ( .A1(n9359), .A2(n9363), .ZN(n9351) );
  INV_X1 U11293 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8998) );
  AND2_X1 U11294 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_REG3_REG_11__SCAN_IN), 
        .ZN(n8742) );
  NAND2_X1 U11295 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_REG3_REG_16__SCAN_IN), 
        .ZN(n8746) );
  INV_X1 U11296 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9158) );
  OR2_X2 U11297 ( .A1(n9159), .A2(n9158), .ZN(n9179) );
  INV_X1 U11298 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14879) );
  INV_X1 U11299 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14862) );
  INV_X1 U11300 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9249) );
  OR2_X2 U11301 ( .A1(n9250), .A2(n9249), .ZN(n9270) );
  NAND2_X1 U11302 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n8752) );
  OR2_X2 U11303 ( .A1(n9321), .A2(n8752), .ZN(n15176) );
  INV_X1 U11304 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9985) );
  NAND2_X1 U11305 ( .A1(n9296), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U11306 ( .A1(n9252), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8754) );
  OAI211_X1 U11307 ( .C1(n9985), .C2(n9308), .A(n8755), .B(n8754), .ZN(n8756)
         );
  INV_X1 U11308 ( .A(n8756), .ZN(n8757) );
  OAI21_X1 U11309 ( .B1(n15176), .B2(n9295), .A(n8757), .ZN(n14997) );
  INV_X1 U11310 ( .A(n14997), .ZN(n8762) );
  NAND2_X1 U11311 ( .A1(n14825), .A2(n9333), .ZN(n8761) );
  OR2_X1 U11312 ( .A1(n8898), .A2(n15593), .ZN(n8760) );
  INV_X1 U11313 ( .A(n15175), .ZN(n15451) );
  MUX2_X1 U11314 ( .A(n8762), .B(n15451), .S(n9131), .Z(n9339) );
  MUX2_X1 U11315 ( .A(n14997), .B(n15175), .S(n9020), .Z(n9338) );
  NAND2_X1 U11316 ( .A1(n9339), .A2(n9338), .ZN(n9349) );
  NAND2_X1 U11317 ( .A1(n9351), .A2(n9349), .ZN(n9358) );
  NAND2_X1 U11318 ( .A1(n9296), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8768) );
  INV_X1 U11319 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n12541) );
  OR2_X1 U11320 ( .A1(n9308), .A2(n12541), .ZN(n8767) );
  INV_X1 U11321 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n11073) );
  INV_X1 U11322 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n8763) );
  OAI21_X1 U11323 ( .B1(n9007), .B2(n11073), .A(n8763), .ZN(n8764) );
  NAND2_X1 U11324 ( .A1(n9029), .A2(n8764), .ZN(n14893) );
  OR2_X1 U11325 ( .A1(n9295), .A2(n14893), .ZN(n8766) );
  INV_X1 U11326 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n12386) );
  OR2_X1 U11327 ( .A1(n7213), .A2(n12386), .ZN(n8765) );
  NAND4_X1 U11328 ( .A1(n8768), .A2(n8767), .A3(n8766), .A4(n8765), .ZN(n15010) );
  NAND2_X1 U11329 ( .A1(n8987), .A2(n8769), .ZN(n8771) );
  NAND2_X1 U11330 ( .A1(n8771), .A2(n8770), .ZN(n8773) );
  NAND2_X1 U11331 ( .A1(n8773), .A2(n8772), .ZN(n8774) );
  NAND2_X1 U11332 ( .A1(n10646), .A2(n9333), .ZN(n8786) );
  INV_X1 U11333 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8775) );
  INV_X1 U11334 ( .A(n8792), .ZN(n8777) );
  INV_X1 U11335 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8776) );
  NAND2_X1 U11336 ( .A1(n8777), .A2(n8776), .ZN(n8833) );
  INV_X1 U11337 ( .A(n8833), .ZN(n8779) );
  INV_X1 U11338 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n8778) );
  NAND2_X1 U11339 ( .A1(n8779), .A2(n8778), .ZN(n8811) );
  OR2_X1 U11340 ( .A1(n8781), .A2(n15585), .ZN(n8782) );
  NAND2_X1 U11341 ( .A1(n8993), .A2(n8782), .ZN(n9017) );
  INV_X1 U11342 ( .A(n9017), .ZN(n8783) );
  NAND2_X1 U11343 ( .A1(n8783), .A2(n9016), .ZN(n8784) );
  NAND2_X1 U11344 ( .A1(n8784), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9040) );
  XNOR2_X1 U11345 ( .A(n9040), .B(P1_IR_REG_12__SCAN_IN), .ZN(n15710) );
  AOI22_X1 U11346 ( .A1(n9154), .A2(n15710), .B1(n9155), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n8785) );
  MUX2_X1 U11347 ( .A(n15010), .B(n12605), .S(n9131), .Z(n9028) );
  NAND2_X1 U11348 ( .A1(n8788), .A2(n8787), .ZN(n8791) );
  NAND2_X1 U11349 ( .A1(n8791), .A2(n8830), .ZN(n10570) );
  OR2_X1 U11350 ( .A1(n10570), .A2(n8897), .ZN(n8795) );
  NAND2_X1 U11351 ( .A1(n8792), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8793) );
  XNOR2_X1 U11352 ( .A(n8793), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10709) );
  AOI22_X1 U11353 ( .A1(n9155), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9154), .B2(
        n10709), .ZN(n8794) );
  NAND2_X1 U11354 ( .A1(n9324), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8802) );
  INV_X1 U11355 ( .A(n8906), .ZN(n9327) );
  INV_X1 U11356 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n8796) );
  OR2_X1 U11357 ( .A1(n9327), .A2(n8796), .ZN(n8801) );
  INV_X1 U11358 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n8797) );
  NAND2_X1 U11359 ( .A1(n8937), .A2(n8797), .ZN(n8798) );
  NAND2_X1 U11360 ( .A1(n8822), .A2(n8798), .ZN(n11791) );
  OR2_X1 U11361 ( .A1(n9295), .A2(n11791), .ZN(n8800) );
  INV_X1 U11362 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10690) );
  OR2_X1 U11363 ( .A1(n9273), .A2(n10690), .ZN(n8799) );
  MUX2_X1 U11364 ( .A(n15731), .B(n15016), .S(n9076), .Z(n8953) );
  INV_X1 U11365 ( .A(n8953), .ZN(n8804) );
  INV_X1 U11366 ( .A(n15731), .ZN(n11797) );
  MUX2_X1 U11367 ( .A(n11797), .B(n14839), .S(n9131), .Z(n8954) );
  INV_X1 U11368 ( .A(n8954), .ZN(n8803) );
  NAND2_X1 U11369 ( .A1(n8806), .A2(n8805), .ZN(n8808) );
  NAND2_X1 U11370 ( .A1(n8808), .A2(n8807), .ZN(n8810) );
  NAND2_X1 U11371 ( .A1(n10617), .A2(n9333), .ZN(n8814) );
  NAND2_X1 U11372 ( .A1(n8811), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8812) );
  XNOR2_X1 U11373 ( .A(n8812), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10751) );
  AOI22_X1 U11374 ( .A1(n9155), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9154), .B2(
        n10751), .ZN(n8813) );
  INV_X1 U11375 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10746) );
  OR2_X1 U11376 ( .A1(n9308), .A2(n10746), .ZN(n8820) );
  NAND2_X1 U11377 ( .A1(n8906), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8819) );
  NAND2_X1 U11378 ( .A1(n9252), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n8818) );
  INV_X1 U11379 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n8815) );
  NAND2_X1 U11380 ( .A1(n8824), .A2(n8815), .ZN(n8816) );
  NAND2_X1 U11381 ( .A1(n8972), .A2(n8816), .ZN(n11951) );
  OR2_X1 U11382 ( .A1(n9295), .A2(n11951), .ZN(n8817) );
  NAND4_X1 U11383 ( .A1(n8820), .A2(n8819), .A3(n8818), .A4(n8817), .ZN(n15014) );
  NAND2_X1 U11384 ( .A1(n9296), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n8828) );
  INV_X1 U11385 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10692) );
  OR2_X1 U11386 ( .A1(n9273), .A2(n10692), .ZN(n8827) );
  INV_X1 U11387 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n8821) );
  NAND2_X1 U11388 ( .A1(n8822), .A2(n8821), .ZN(n8823) );
  NAND2_X1 U11389 ( .A1(n8824), .A2(n8823), .ZN(n14843) );
  OR2_X1 U11390 ( .A1(n9295), .A2(n14843), .ZN(n8826) );
  INV_X1 U11391 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10671) );
  OR2_X1 U11392 ( .A1(n9308), .A2(n10671), .ZN(n8825) );
  XNOR2_X1 U11393 ( .A(n8832), .B(n8831), .ZN(n10582) );
  NAND2_X1 U11394 ( .A1(n10582), .A2(n9333), .ZN(n8836) );
  NAND2_X1 U11395 ( .A1(n8833), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8834) );
  XNOR2_X1 U11396 ( .A(n8834), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10691) );
  AOI22_X1 U11397 ( .A1(n9155), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9154), .B2(
        n10691), .ZN(n8835) );
  INV_X1 U11398 ( .A(n15812), .ZN(n11761) );
  INV_X1 U11399 ( .A(n11955), .ZN(n15015) );
  MUX2_X1 U11400 ( .A(n15015), .B(n15812), .S(n9131), .Z(n8962) );
  NAND2_X1 U11401 ( .A1(n8963), .A2(n8962), .ZN(n8837) );
  AND2_X1 U11402 ( .A1(n11959), .A2(n8837), .ZN(n8958) );
  NAND2_X1 U11403 ( .A1(n8906), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8842) );
  INV_X1 U11404 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n15673) );
  OR2_X1 U11405 ( .A1(n8863), .A2(n15673), .ZN(n8841) );
  INV_X1 U11406 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11443) );
  OR2_X1 U11407 ( .A1(n9295), .A2(n11443), .ZN(n8840) );
  INV_X1 U11408 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n8838) );
  OR2_X1 U11409 ( .A1(n9273), .A2(n8838), .ZN(n8839) );
  AND4_X2 U11410 ( .A1(n8842), .A2(n8841), .A3(n8840), .A4(n8839), .ZN(n15749)
         );
  NOR2_X1 U11411 ( .A1(n6542), .A2(n8844), .ZN(n8846) );
  XNOR2_X1 U11412 ( .A(n8846), .B(n8845), .ZN(n15600) );
  OAI21_X2 U11413 ( .B1(n10642), .B2(n8858), .A(n8847), .ZN(n8869) );
  NAND2_X1 U11414 ( .A1(n8874), .A2(n8848), .ZN(n8852) );
  INV_X1 U11415 ( .A(n8852), .ZN(n8849) );
  NAND2_X1 U11416 ( .A1(n8849), .A2(n8850), .ZN(n8875) );
  INV_X1 U11417 ( .A(n8850), .ZN(n8851) );
  NAND2_X1 U11418 ( .A1(n8852), .A2(n8851), .ZN(n8853) );
  NAND2_X1 U11419 ( .A1(n8875), .A2(n8853), .ZN(n10573) );
  NOR2_X1 U11420 ( .A1(n10573), .A2(n6542), .ZN(n8854) );
  INV_X1 U11421 ( .A(n8855), .ZN(n10676) );
  INV_X1 U11422 ( .A(n15674), .ZN(n15150) );
  AND2_X1 U11423 ( .A1(n7176), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8856) );
  INV_X1 U11424 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n8858) );
  INV_X1 U11425 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n8857) );
  INV_X1 U11426 ( .A(n10678), .ZN(n15023) );
  NAND3_X1 U11427 ( .A1(n8855), .A2(n15023), .A3(n15674), .ZN(n8859) );
  INV_X1 U11428 ( .A(n9295), .ZN(n8886) );
  NAND2_X1 U11429 ( .A1(n8906), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n8866) );
  INV_X1 U11430 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n8862) );
  NAND2_X1 U11431 ( .A1(n11501), .A2(n15751), .ZN(n9384) );
  NAND2_X1 U11432 ( .A1(n8868), .A2(n9384), .ZN(n11505) );
  INV_X1 U11433 ( .A(n8869), .ZN(n11502) );
  NAND2_X1 U11434 ( .A1(n11502), .A2(n15749), .ZN(n8870) );
  INV_X1 U11435 ( .A(n15749), .ZN(n15753) );
  NAND2_X1 U11436 ( .A1(n8870), .A2(n15738), .ZN(n11447) );
  NAND2_X1 U11437 ( .A1(n11447), .A2(n6953), .ZN(n8871) );
  OR2_X2 U11438 ( .A1(n15751), .A2(n11501), .ZN(n11504) );
  MUX2_X1 U11439 ( .A(n11504), .B(n9384), .S(n9131), .Z(n8872) );
  NAND2_X1 U11440 ( .A1(n8875), .A2(n8874), .ZN(n8879) );
  AND2_X1 U11441 ( .A1(n8877), .A2(n8876), .ZN(n8878) );
  XNOR2_X1 U11442 ( .A(n8879), .B(n8878), .ZN(n10624) );
  OR2_X1 U11443 ( .A1(n10624), .A2(n8897), .ZN(n8885) );
  OR2_X1 U11444 ( .A1(n8898), .A2(n10572), .ZN(n8884) );
  INV_X1 U11445 ( .A(n8880), .ZN(n8882) );
  INV_X1 U11446 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8881) );
  NAND2_X1 U11447 ( .A1(n8882), .A2(n8881), .ZN(n8899) );
  INV_X1 U11448 ( .A(n10683), .ZN(n10889) );
  NAND2_X1 U11449 ( .A1(n9154), .A2(n10889), .ZN(n8883) );
  NAND2_X1 U11450 ( .A1(n8886), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n8891) );
  NAND2_X1 U11451 ( .A1(n8906), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8890) );
  NAND2_X1 U11452 ( .A1(n9324), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8889) );
  NAND2_X1 U11453 ( .A1(n8887), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n8888) );
  MUX2_X1 U11454 ( .A(n9383), .B(n11506), .S(n9131), .Z(n8892) );
  NAND2_X1 U11455 ( .A1(n8893), .A2(n8892), .ZN(n8913) );
  NAND2_X1 U11456 ( .A1(n8895), .A2(n8894), .ZN(n8896) );
  NAND2_X1 U11457 ( .A1(n8896), .A2(n8918), .ZN(n10630) );
  OR2_X1 U11458 ( .A1(n8897), .A2(n10630), .ZN(n8905) );
  INV_X1 U11459 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10575) );
  OR2_X1 U11460 ( .A1(n8898), .A2(n10575), .ZN(n8904) );
  NAND2_X1 U11461 ( .A1(n8899), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8900) );
  MUX2_X1 U11462 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8900), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n8902) );
  INV_X1 U11463 ( .A(n8925), .ZN(n8901) );
  NAND2_X1 U11464 ( .A1(n9154), .A2(n15040), .ZN(n8903) );
  NAND2_X1 U11465 ( .A1(n9324), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8910) );
  NAND2_X1 U11466 ( .A1(n8906), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8909) );
  OR2_X1 U11467 ( .A1(n9295), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8907) );
  NAND2_X1 U11468 ( .A1(n11541), .A2(n15425), .ZN(n8914) );
  NAND2_X1 U11469 ( .A1(n15786), .A2(n11498), .ZN(n11507) );
  MUX2_X1 U11470 ( .A(n10985), .B(n15780), .S(n9131), .Z(n8911) );
  NAND2_X1 U11471 ( .A1(n15780), .A2(n10985), .ZN(n11496) );
  NAND2_X1 U11472 ( .A1(n8911), .A2(n11496), .ZN(n8912) );
  NAND3_X1 U11473 ( .A1(n8913), .A2(n11539), .A3(n8912), .ZN(n8916) );
  MUX2_X1 U11474 ( .A(n8914), .B(n11507), .S(n9344), .Z(n8915) );
  NAND2_X1 U11475 ( .A1(n8916), .A2(n8915), .ZN(n8952) );
  AND2_X1 U11476 ( .A1(n8918), .A2(n8917), .ZN(n8920) );
  NAND2_X1 U11477 ( .A1(n8942), .A2(n8919), .ZN(n8921) );
  NAND2_X1 U11478 ( .A1(n8920), .A2(n8921), .ZN(n8924) );
  INV_X1 U11479 ( .A(n8920), .ZN(n8923) );
  INV_X1 U11480 ( .A(n8921), .ZN(n8922) );
  NAND2_X1 U11481 ( .A1(n8923), .A2(n8922), .ZN(n8943) );
  OR2_X1 U11482 ( .A1(n10626), .A2(n8897), .ZN(n8928) );
  INV_X1 U11483 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n15585) );
  AOI22_X1 U11484 ( .A1(n9155), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n9154), .B2(
        n15684), .ZN(n8927) );
  NAND2_X1 U11485 ( .A1(n9324), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8932) );
  NAND2_X1 U11486 ( .A1(n9296), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n8931) );
  NAND2_X1 U11487 ( .A1(n9252), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n8930) );
  XNOR2_X1 U11488 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n11357) );
  OR2_X1 U11489 ( .A1(n9295), .A2(n11357), .ZN(n8929) );
  MUX2_X1 U11490 ( .A(n11525), .B(n15018), .S(n9020), .Z(n8951) );
  NAND2_X1 U11491 ( .A1(n9296), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8941) );
  NAND2_X1 U11492 ( .A1(n9252), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n8940) );
  INV_X1 U11493 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8935) );
  NAND2_X1 U11494 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n8934) );
  NAND2_X1 U11495 ( .A1(n8935), .A2(n8934), .ZN(n8936) );
  NAND2_X1 U11496 ( .A1(n8937), .A2(n8936), .ZN(n11653) );
  OR2_X1 U11497 ( .A1(n9295), .A2(n11653), .ZN(n8939) );
  INV_X1 U11498 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10669) );
  OR2_X1 U11499 ( .A1(n9308), .A2(n10669), .ZN(n8938) );
  NAND4_X1 U11500 ( .A1(n8941), .A2(n8940), .A3(n8939), .A4(n8938), .ZN(n15017) );
  INV_X1 U11501 ( .A(n15017), .ZN(n11711) );
  NAND2_X1 U11502 ( .A1(n8943), .A2(n8942), .ZN(n8945) );
  XNOR2_X1 U11503 ( .A(n8944), .B(n8945), .ZN(n10569) );
  NAND2_X1 U11504 ( .A1(n10569), .A2(n9333), .ZN(n8949) );
  NAND2_X1 U11505 ( .A1(n8946), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8947) );
  XNOR2_X1 U11506 ( .A(n8947), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10688) );
  AOI22_X1 U11507 ( .A1(n9155), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9154), .B2(
        n10688), .ZN(n8948) );
  INV_X1 U11508 ( .A(n11742), .ZN(n11534) );
  MUX2_X1 U11509 ( .A(n11711), .B(n11534), .S(n9076), .Z(n8956) );
  MUX2_X1 U11510 ( .A(n15017), .B(n11742), .S(n9131), .Z(n8955) );
  OAI22_X1 U11511 ( .A1(n8952), .A2(n8951), .B1(n8956), .B2(n8955), .ZN(n8961)
         );
  INV_X1 U11512 ( .A(n15018), .ZN(n11524) );
  MUX2_X1 U11513 ( .A(n11521), .B(n11524), .S(n9131), .Z(n8950) );
  AOI21_X1 U11514 ( .B1(n8952), .B2(n8951), .A(n8950), .ZN(n8960) );
  AOI22_X1 U11515 ( .A1(n8956), .A2(n8955), .B1(n8954), .B2(n8953), .ZN(n8957)
         );
  INV_X1 U11516 ( .A(n8962), .ZN(n8965) );
  INV_X1 U11517 ( .A(n8963), .ZN(n8964) );
  NAND3_X1 U11518 ( .A1(n11959), .A2(n8965), .A3(n8964), .ZN(n8969) );
  AND2_X1 U11519 ( .A1(n9131), .A2(n15014), .ZN(n8967) );
  OAI21_X1 U11520 ( .B1(n15014), .B2(n9344), .A(n12001), .ZN(n8966) );
  OAI21_X1 U11521 ( .B1(n8967), .B2(n12001), .A(n8966), .ZN(n8968) );
  NAND2_X1 U11522 ( .A1(n9296), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8977) );
  INV_X1 U11523 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n12017) );
  OR2_X1 U11524 ( .A1(n7213), .A2(n12017), .ZN(n8976) );
  NAND2_X1 U11525 ( .A1(n8972), .A2(n8971), .ZN(n8973) );
  NAND2_X1 U11526 ( .A1(n8999), .A2(n8973), .ZN(n12643) );
  OR2_X1 U11527 ( .A1(n9295), .A2(n12643), .ZN(n8975) );
  INV_X1 U11528 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n11068) );
  OR2_X1 U11529 ( .A1(n9308), .A2(n11068), .ZN(n8974) );
  INV_X1 U11530 ( .A(n12432), .ZN(n15013) );
  NAND2_X1 U11531 ( .A1(n10621), .A2(n9333), .ZN(n8981) );
  XNOR2_X1 U11532 ( .A(n8993), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10752) );
  AOI22_X1 U11533 ( .A1(n9155), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9154), .B2(
        n10752), .ZN(n8980) );
  NAND2_X2 U11534 ( .A1(n8981), .A2(n8980), .ZN(n12655) );
  MUX2_X1 U11535 ( .A(n15013), .B(n12655), .S(n9076), .Z(n8984) );
  MUX2_X1 U11536 ( .A(n15013), .B(n12655), .S(n9344), .Z(n8982) );
  INV_X1 U11537 ( .A(n8983), .ZN(n8986) );
  NAND2_X1 U11538 ( .A1(n8987), .A2(SI_10_), .ZN(n9012) );
  NAND2_X1 U11539 ( .A1(n8989), .A2(n8988), .ZN(n8990) );
  INV_X1 U11540 ( .A(n10657), .ZN(n8991) );
  INV_X1 U11541 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8992) );
  NAND2_X1 U11542 ( .A1(n8993), .A2(n8992), .ZN(n8994) );
  NAND2_X1 U11543 ( .A1(n8994), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8995) );
  XNOR2_X1 U11544 ( .A(n8995), .B(P1_IR_REG_10__SCAN_IN), .ZN(n15054) );
  AOI22_X1 U11545 ( .A1(n9155), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n9154), 
        .B2(n15054), .ZN(n8996) );
  NAND2_X1 U11546 ( .A1(n9296), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n9004) );
  NAND2_X1 U11547 ( .A1(n9252), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9003) );
  NAND2_X1 U11548 ( .A1(n9324), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9002) );
  NAND2_X1 U11549 ( .A1(n8999), .A2(n8998), .ZN(n9000) );
  NAND2_X1 U11550 ( .A1(n9007), .A2(n9000), .ZN(n12576) );
  OR2_X1 U11551 ( .A1(n9295), .A2(n12576), .ZN(n9001) );
  NAND4_X1 U11552 ( .A1(n9004), .A2(n9003), .A3(n9002), .A4(n9001), .ZN(n15012) );
  MUX2_X1 U11553 ( .A(n12426), .B(n15012), .S(n9076), .Z(n9006) );
  INV_X1 U11554 ( .A(n15012), .ZN(n12170) );
  INV_X1 U11555 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11766) );
  OR2_X1 U11556 ( .A1(n9308), .A2(n11766), .ZN(n9011) );
  NAND2_X1 U11557 ( .A1(n9296), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n9010) );
  NAND2_X1 U11558 ( .A1(n9252), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9009) );
  XNOR2_X1 U11559 ( .A(n9007), .B(n11073), .ZN(n14956) );
  OR2_X1 U11560 ( .A1(n9295), .A2(n14956), .ZN(n9008) );
  NAND4_X1 U11561 ( .A1(n9011), .A2(n9010), .A3(n9009), .A4(n9008), .ZN(n15011) );
  NAND2_X1 U11562 ( .A1(n9013), .A2(n9012), .ZN(n9015) );
  XNOR2_X1 U11563 ( .A(n9014), .B(n9015), .ZN(n10761) );
  NAND2_X1 U11564 ( .A1(n10761), .A2(n9333), .ZN(n9019) );
  XNOR2_X1 U11565 ( .A(n9017), .B(n9016), .ZN(n11771) );
  AOI22_X1 U11566 ( .A1(n9155), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9154), 
        .B2(n11771), .ZN(n9018) );
  MUX2_X1 U11567 ( .A(n15011), .B(n15559), .S(n9020), .Z(n9023) );
  MUX2_X1 U11568 ( .A(n15011), .B(n15559), .S(n9344), .Z(n9021) );
  NAND2_X1 U11569 ( .A1(n9027), .A2(n9028), .ZN(n9025) );
  MUX2_X1 U11570 ( .A(n15010), .B(n12605), .S(n9076), .Z(n9024) );
  NAND2_X1 U11571 ( .A1(n9025), .A2(n9024), .ZN(n9026) );
  NAND2_X1 U11572 ( .A1(n8906), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n9034) );
  INV_X1 U11573 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10108) );
  OR2_X1 U11574 ( .A1(n9308), .A2(n10108), .ZN(n9033) );
  NAND2_X1 U11575 ( .A1(n9252), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9032) );
  INV_X1 U11576 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n11775) );
  NAND2_X1 U11577 ( .A1(n9029), .A2(n11775), .ZN(n9030) );
  NAND2_X1 U11578 ( .A1(n9057), .A2(n9030), .ZN(n12614) );
  OR2_X1 U11579 ( .A1(n9295), .A2(n12614), .ZN(n9031) );
  NAND4_X1 U11580 ( .A1(n9034), .A2(n9033), .A3(n9032), .A4(n9031), .ZN(n15009) );
  NAND2_X1 U11581 ( .A1(n9036), .A2(n9035), .ZN(n9037) );
  NAND2_X1 U11582 ( .A1(n9038), .A2(n9037), .ZN(n10650) );
  OR2_X1 U11583 ( .A1(n10650), .A2(n8897), .ZN(n9044) );
  INV_X1 U11584 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9039) );
  NAND2_X1 U11585 ( .A1(n9040), .A2(n9039), .ZN(n9041) );
  NAND2_X1 U11586 ( .A1(n9041), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9050) );
  XNOR2_X1 U11587 ( .A(n9050), .B(P1_IR_REG_13__SCAN_IN), .ZN(n15066) );
  NOR2_X1 U11588 ( .A1(n8898), .A2(n10651), .ZN(n9042) );
  AOI21_X1 U11589 ( .B1(n15066), .B2(n9154), .A(n9042), .ZN(n9043) );
  MUX2_X1 U11590 ( .A(n15009), .B(n15553), .S(n9020), .Z(n9141) );
  NAND2_X1 U11591 ( .A1(n9115), .A2(SI_14_), .ZN(n9063) );
  INV_X1 U11592 ( .A(n9046), .ZN(n9045) );
  NAND2_X1 U11593 ( .A1(n9047), .A2(n9046), .ZN(n9048) );
  NAND2_X1 U11594 ( .A1(n10776), .A2(n9333), .ZN(n9054) );
  INV_X1 U11595 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9049) );
  NAND2_X1 U11596 ( .A1(n9050), .A2(n9049), .ZN(n9051) );
  NAND2_X1 U11597 ( .A1(n9051), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9052) );
  XNOR2_X1 U11598 ( .A(n9052), .B(P1_IR_REG_14__SCAN_IN), .ZN(n15081) );
  AOI22_X1 U11599 ( .A1(n15081), .A2(n9154), .B1(n9155), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n9053) );
  INV_X1 U11600 ( .A(n9055), .ZN(n9071) );
  INV_X1 U11601 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9056) );
  NAND2_X1 U11602 ( .A1(n9057), .A2(n9056), .ZN(n9058) );
  AND2_X1 U11603 ( .A1(n9071), .A2(n9058), .ZN(n15416) );
  NAND2_X1 U11604 ( .A1(n15416), .A2(n9323), .ZN(n9062) );
  NAND2_X1 U11605 ( .A1(n9296), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9061) );
  NAND2_X1 U11606 ( .A1(n9252), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9060) );
  INV_X1 U11607 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n15064) );
  OR2_X1 U11608 ( .A1(n9308), .A2(n15064), .ZN(n9059) );
  NAND4_X1 U11609 ( .A1(n9062), .A2(n9061), .A3(n9060), .A4(n9059), .ZN(n15008) );
  AND2_X1 U11610 ( .A1(n15419), .A2(n15008), .ZN(n12713) );
  INV_X1 U11611 ( .A(n15008), .ZN(n12622) );
  NAND2_X1 U11612 ( .A1(n15548), .A2(n12622), .ZN(n12716) );
  INV_X1 U11613 ( .A(n15009), .ZN(n15410) );
  OR2_X1 U11614 ( .A1(n9067), .A2(n15585), .ZN(n9068) );
  XNOR2_X1 U11615 ( .A(n9068), .B(P1_IR_REG_15__SCAN_IN), .ZN(n15721) );
  AOI22_X1 U11616 ( .A1(n9155), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9154), 
        .B2(n15721), .ZN(n9069) );
  INV_X1 U11617 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9070) );
  NAND2_X1 U11618 ( .A1(n9071), .A2(n9070), .ZN(n9072) );
  NAND2_X1 U11619 ( .A1(n9108), .A2(n9072), .ZN(n15394) );
  OR2_X1 U11620 ( .A1(n15394), .A2(n9295), .ZN(n9075) );
  AOI22_X1 U11621 ( .A1(n9324), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n9296), .B2(
        P1_REG0_REG_15__SCAN_IN), .ZN(n9074) );
  NAND2_X1 U11622 ( .A1(n9252), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n9073) );
  AND4_X1 U11623 ( .A1(n15408), .A2(n15410), .A3(n9076), .A4(n15370), .ZN(
        n9077) );
  OAI21_X1 U11624 ( .B1(n9140), .B2(n9141), .A(n9077), .ZN(n9144) );
  XNOR2_X1 U11625 ( .A(n9149), .B(SI_18_), .ZN(n9148) );
  XNOR2_X1 U11626 ( .A(n9148), .B(n9078), .ZN(n11003) );
  NAND2_X1 U11627 ( .A1(n11003), .A2(n9333), .ZN(n9082) );
  NAND2_X1 U11628 ( .A1(n9079), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9080) );
  XNOR2_X1 U11629 ( .A(n9080), .B(P1_IR_REG_18__SCAN_IN), .ZN(n15137) );
  AOI22_X1 U11630 ( .A1(n9155), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9154), 
        .B2(n15137), .ZN(n9081) );
  INV_X1 U11631 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n15116) );
  NAND2_X1 U11632 ( .A1(n9093), .A2(n15116), .ZN(n9083) );
  NAND2_X1 U11633 ( .A1(n9159), .A2(n9083), .ZN(n15346) );
  OR2_X1 U11634 ( .A1(n15346), .A2(n9295), .ZN(n9088) );
  INV_X1 U11635 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n15125) );
  NAND2_X1 U11636 ( .A1(n9296), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n9085) );
  INV_X1 U11637 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n15347) );
  OR2_X1 U11638 ( .A1(n7213), .A2(n15347), .ZN(n9084) );
  OAI211_X1 U11639 ( .C1(n9308), .C2(n15125), .A(n9085), .B(n9084), .ZN(n9086)
         );
  INV_X1 U11640 ( .A(n9086), .ZN(n9087) );
  XNOR2_X1 U11641 ( .A(n14965), .B(n15321), .ZN(n15334) );
  INV_X1 U11642 ( .A(n15370), .ZN(n9089) );
  NAND2_X1 U11643 ( .A1(n9089), .A2(n9020), .ZN(n9134) );
  AND2_X1 U11644 ( .A1(n15408), .A2(n12717), .ZN(n9090) );
  NOR2_X1 U11645 ( .A1(n15553), .A2(n9020), .ZN(n9142) );
  NAND2_X1 U11646 ( .A1(n9141), .A2(n9142), .ZN(n9137) );
  INV_X1 U11647 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9092) );
  INV_X1 U11648 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9091) );
  OAI21_X1 U11649 ( .B1(n9108), .B2(n9092), .A(n9091), .ZN(n9094) );
  AND2_X1 U11650 ( .A1(n9094), .A2(n9093), .ZN(n15364) );
  NAND2_X1 U11651 ( .A1(n15364), .A2(n9323), .ZN(n9097) );
  AOI22_X1 U11652 ( .A1(n9324), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n9296), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n9096) );
  INV_X1 U11653 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n15107) );
  OR2_X1 U11654 ( .A1(n7213), .A2(n15107), .ZN(n9095) );
  INV_X1 U11655 ( .A(n15340), .ZN(n15005) );
  NAND2_X1 U11656 ( .A1(n15005), .A2(n9344), .ZN(n9107) );
  NAND2_X1 U11657 ( .A1(n15340), .A2(n9076), .ZN(n9106) );
  NAND2_X1 U11658 ( .A1(n9099), .A2(n9098), .ZN(n9101) );
  XNOR2_X1 U11659 ( .A(n9101), .B(n9100), .ZN(n10772) );
  NAND2_X1 U11660 ( .A1(n10772), .A2(n9333), .ZN(n9105) );
  NAND2_X1 U11661 ( .A1(n9124), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9102) );
  MUX2_X1 U11662 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9102), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n9103) );
  NAND2_X1 U11663 ( .A1(n9103), .A2(n9079), .ZN(n15120) );
  INV_X1 U11664 ( .A(n15120), .ZN(n15123) );
  AOI22_X1 U11665 ( .A1(n9155), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9154), 
        .B2(n15123), .ZN(n9104) );
  MUX2_X1 U11666 ( .A(n9107), .B(n9106), .S(n15531), .Z(n9170) );
  XNOR2_X1 U11667 ( .A(n9108), .B(P1_REG3_REG_16__SCAN_IN), .ZN(n15379) );
  NAND2_X1 U11668 ( .A1(n15379), .A2(n9323), .ZN(n9113) );
  INV_X1 U11669 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10016) );
  NAND2_X1 U11670 ( .A1(n9324), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9110) );
  NAND2_X1 U11671 ( .A1(n9252), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9109) );
  OAI211_X1 U11672 ( .C1(n9327), .C2(n10016), .A(n9110), .B(n9109), .ZN(n9111)
         );
  INV_X1 U11673 ( .A(n9111), .ZN(n9112) );
  NAND2_X1 U11674 ( .A1(n9113), .A2(n9112), .ZN(n15006) );
  NAND2_X1 U11675 ( .A1(n9115), .A2(n9114), .ZN(n9117) );
  NAND2_X1 U11676 ( .A1(n9117), .A2(n9116), .ZN(n9119) );
  NAND2_X1 U11677 ( .A1(n9119), .A2(n9118), .ZN(n9121) );
  XNOR2_X1 U11678 ( .A(n9121), .B(n9120), .ZN(n10768) );
  NAND2_X1 U11679 ( .A1(n10768), .A2(n9333), .ZN(n9127) );
  NAND2_X1 U11680 ( .A1(n9122), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9123) );
  MUX2_X1 U11681 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9123), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n9125) );
  AND2_X1 U11682 ( .A1(n9125), .A2(n9124), .ZN(n15101) );
  AOI22_X1 U11683 ( .A1(n9155), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9154), 
        .B2(n15101), .ZN(n9126) );
  MUX2_X1 U11684 ( .A(n15006), .B(n15537), .S(n9076), .Z(n9168) );
  NAND2_X1 U11685 ( .A1(n15537), .A2(n9344), .ZN(n9145) );
  NAND2_X1 U11686 ( .A1(n9076), .A2(n15006), .ZN(n9167) );
  NAND3_X1 U11687 ( .A1(n9168), .A2(n9145), .A3(n9167), .ZN(n9128) );
  AND2_X1 U11688 ( .A1(n9170), .A2(n9128), .ZN(n9136) );
  NAND2_X1 U11689 ( .A1(n12716), .A2(n9076), .ZN(n9129) );
  NAND2_X1 U11690 ( .A1(n12717), .A2(n9129), .ZN(n9130) );
  OAI21_X1 U11691 ( .B1(n12717), .B2(n9344), .A(n9130), .ZN(n9133) );
  NAND3_X1 U11692 ( .A1(n15369), .A2(n15370), .A3(n9131), .ZN(n9132) );
  NAND3_X1 U11693 ( .A1(n9134), .A2(n9133), .A3(n9132), .ZN(n9135) );
  INV_X1 U11694 ( .A(n9138), .ZN(n9143) );
  AND2_X1 U11695 ( .A1(n15345), .A2(n15359), .ZN(n12722) );
  AND2_X1 U11696 ( .A1(n14965), .A2(n15321), .ZN(n9171) );
  NOR2_X1 U11697 ( .A1(n15531), .A2(n15005), .ZN(n12697) );
  OAI21_X1 U11698 ( .B1(n9168), .B2(n9145), .A(n15357), .ZN(n9146) );
  NAND2_X1 U11699 ( .A1(n9146), .A2(n9170), .ZN(n9147) );
  OR3_X1 U11700 ( .A1(n12722), .A2(n9171), .A3(n9147), .ZN(n9166) );
  INV_X1 U11701 ( .A(n9149), .ZN(n9150) );
  XNOR2_X1 U11702 ( .A(n9152), .B(SI_19_), .ZN(n9153) );
  NAND2_X1 U11703 ( .A1(n11346), .A2(n9333), .ZN(n9157) );
  AOI22_X1 U11704 ( .A1(n9155), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n15748), 
        .B2(n9154), .ZN(n9156) );
  NAND2_X1 U11705 ( .A1(n9159), .A2(n9158), .ZN(n9160) );
  AND2_X1 U11706 ( .A1(n9179), .A2(n9160), .ZN(n15323) );
  NAND2_X1 U11707 ( .A1(n15323), .A2(n9323), .ZN(n9165) );
  INV_X1 U11708 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n15140) );
  NAND2_X1 U11709 ( .A1(n9324), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n9162) );
  NAND2_X1 U11710 ( .A1(n8906), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9161) );
  OAI211_X1 U11711 ( .C1(n15140), .C2(n7213), .A(n9162), .B(n9161), .ZN(n9163)
         );
  INV_X1 U11712 ( .A(n9163), .ZN(n9164) );
  OR2_X1 U11713 ( .A1(n15519), .A2(n15341), .ZN(n9382) );
  NOR2_X1 U11714 ( .A1(n9168), .A2(n9167), .ZN(n9169) );
  AND2_X1 U11715 ( .A1(n9170), .A2(n9169), .ZN(n9172) );
  INV_X1 U11716 ( .A(n9171), .ZN(n9173) );
  AOI22_X1 U11717 ( .A1(n12722), .A2(n9076), .B1(n9172), .B2(n9173), .ZN(n9176) );
  NAND2_X1 U11718 ( .A1(n15519), .A2(n15341), .ZN(n12725) );
  NAND2_X1 U11719 ( .A1(n12725), .A2(n9173), .ZN(n9174) );
  NAND2_X1 U11720 ( .A1(n9174), .A2(n9344), .ZN(n9175) );
  MUX2_X1 U11721 ( .A(n12725), .B(n9382), .S(n9344), .Z(n9177) );
  INV_X1 U11722 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9178) );
  NAND2_X1 U11723 ( .A1(n9179), .A2(n9178), .ZN(n9180) );
  NAND2_X1 U11724 ( .A1(n9199), .A2(n9180), .ZN(n15306) );
  OR2_X1 U11725 ( .A1(n15306), .A2(n9295), .ZN(n9185) );
  INV_X1 U11726 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n15310) );
  NAND2_X1 U11727 ( .A1(n9324), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n9182) );
  NAND2_X1 U11728 ( .A1(n9296), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9181) );
  OAI211_X1 U11729 ( .C1(n15310), .C2(n7213), .A(n9182), .B(n9181), .ZN(n9183)
         );
  INV_X1 U11730 ( .A(n9183), .ZN(n9184) );
  NAND2_X1 U11731 ( .A1(n9185), .A2(n9184), .ZN(n15003) );
  INV_X1 U11732 ( .A(n15003), .ZN(n15322) );
  OR2_X1 U11733 ( .A1(n9186), .A2(n11490), .ZN(n9206) );
  NAND2_X1 U11734 ( .A1(n9186), .A2(n11490), .ZN(n9187) );
  NAND2_X1 U11735 ( .A1(n9206), .A2(n9187), .ZN(n9190) );
  INV_X1 U11736 ( .A(n9188), .ZN(n9189) );
  NAND2_X1 U11737 ( .A1(n9190), .A2(n9189), .ZN(n9191) );
  OR2_X1 U11738 ( .A1(n8898), .A2(n12825), .ZN(n9192) );
  MUX2_X1 U11739 ( .A(n15322), .B(n15512), .S(n9344), .Z(n9195) );
  MUX2_X1 U11740 ( .A(n15305), .B(n15003), .S(n9344), .Z(n9194) );
  NAND2_X1 U11741 ( .A1(n9196), .A2(n9195), .ZN(n9197) );
  NAND2_X1 U11742 ( .A1(n9199), .A2(n14879), .ZN(n9200) );
  AND2_X1 U11743 ( .A1(n9216), .A2(n9200), .ZN(n15293) );
  NAND2_X1 U11744 ( .A1(n15293), .A2(n9323), .ZN(n9205) );
  INV_X1 U11745 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n15287) );
  NAND2_X1 U11746 ( .A1(n9324), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n9202) );
  NAND2_X1 U11747 ( .A1(n9296), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9201) );
  OAI211_X1 U11748 ( .C1(n15287), .C2(n7213), .A(n9202), .B(n9201), .ZN(n9203)
         );
  INV_X1 U11749 ( .A(n9203), .ZN(n9204) );
  NAND2_X1 U11750 ( .A1(n9207), .A2(n9206), .ZN(n9211) );
  NAND2_X1 U11751 ( .A1(n9209), .A2(n9208), .ZN(n9210) );
  NAND2_X1 U11752 ( .A1(n11550), .A2(n9333), .ZN(n9213) );
  OR2_X1 U11753 ( .A1(n8898), .A2(n12749), .ZN(n9212) );
  MUX2_X1 U11755 ( .A(n15002), .B(n15507), .S(n9076), .Z(n9215) );
  MUX2_X1 U11756 ( .A(n15002), .B(n15507), .S(n9344), .Z(n9214) );
  INV_X1 U11757 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14945) );
  NAND2_X1 U11758 ( .A1(n9216), .A2(n14945), .ZN(n9217) );
  NAND2_X1 U11759 ( .A1(n9235), .A2(n9217), .ZN(n15272) );
  OR2_X1 U11760 ( .A1(n15272), .A2(n9295), .ZN(n9222) );
  INV_X1 U11761 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n10135) );
  NAND2_X1 U11762 ( .A1(n9296), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9219) );
  NAND2_X1 U11763 ( .A1(n9252), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9218) );
  OAI211_X1 U11764 ( .C1(n10135), .C2(n9308), .A(n9219), .B(n9218), .ZN(n9220)
         );
  INV_X1 U11765 ( .A(n9220), .ZN(n9221) );
  INV_X1 U11766 ( .A(n13194), .ZN(n15001) );
  OR2_X1 U11767 ( .A1(n9760), .A2(n7176), .ZN(n9223) );
  INV_X1 U11768 ( .A(n15277), .ZN(n15500) );
  MUX2_X1 U11769 ( .A(n15001), .B(n15500), .S(n9344), .Z(n9226) );
  NAND2_X1 U11770 ( .A1(n9227), .A2(n9226), .ZN(n9225) );
  MUX2_X1 U11771 ( .A(n15500), .B(n15001), .S(n9344), .Z(n9224) );
  NAND2_X1 U11772 ( .A1(n9225), .A2(n9224), .ZN(n9228) );
  XNOR2_X1 U11773 ( .A(n9229), .B(SI_23_), .ZN(n9230) );
  XNOR2_X1 U11774 ( .A(n9231), .B(n9230), .ZN(n11734) );
  NAND2_X1 U11775 ( .A1(n11734), .A2(n9333), .ZN(n9234) );
  OR2_X1 U11776 ( .A1(n8898), .A2(n9232), .ZN(n9233) );
  NAND2_X1 U11777 ( .A1(n9235), .A2(n14862), .ZN(n9236) );
  NAND2_X1 U11778 ( .A1(n9250), .A2(n9236), .ZN(n15262) );
  INV_X1 U11779 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9239) );
  NAND2_X1 U11780 ( .A1(n9252), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9238) );
  NAND2_X1 U11781 ( .A1(n9296), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9237) );
  OAI211_X1 U11782 ( .C1(n9308), .C2(n9239), .A(n9238), .B(n9237), .ZN(n9240)
         );
  INV_X1 U11783 ( .A(n9240), .ZN(n9241) );
  AND2_X2 U11784 ( .A1(n9242), .A2(n9241), .ZN(n15274) );
  MUX2_X1 U11785 ( .A(n15265), .B(n15000), .S(n9344), .Z(n9243) );
  NAND2_X1 U11786 ( .A1(n9244), .A2(n9243), .ZN(n9246) );
  MUX2_X1 U11787 ( .A(n15000), .B(n15265), .S(n9344), .Z(n9245) );
  NAND2_X1 U11788 ( .A1(n9246), .A2(n9245), .ZN(n9247) );
  NAND2_X1 U11789 ( .A1(n9250), .A2(n9249), .ZN(n9251) );
  NAND2_X1 U11790 ( .A1(n15252), .A2(n9323), .ZN(n9258) );
  INV_X1 U11791 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9255) );
  NAND2_X1 U11792 ( .A1(n9296), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9254) );
  NAND2_X1 U11793 ( .A1(n9252), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9253) );
  OAI211_X1 U11794 ( .C1(n9255), .C2(n9308), .A(n9254), .B(n9253), .ZN(n9256)
         );
  INV_X1 U11795 ( .A(n9256), .ZN(n9257) );
  NAND2_X2 U11796 ( .A1(n9258), .A2(n9257), .ZN(n14999) );
  INV_X1 U11797 ( .A(n9259), .ZN(n9260) );
  NAND2_X1 U11798 ( .A1(n9261), .A2(n9260), .ZN(n9262) );
  OR2_X1 U11799 ( .A1(n8898), .A2(n12221), .ZN(n9264) );
  MUX2_X1 U11800 ( .A(n14999), .B(n15488), .S(n9344), .Z(n9268) );
  MUX2_X1 U11801 ( .A(n15488), .B(n14999), .S(n9344), .Z(n9266) );
  INV_X1 U11802 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9269) );
  NAND2_X1 U11803 ( .A1(n9270), .A2(n9269), .ZN(n9271) );
  NAND2_X1 U11804 ( .A1(n9293), .A2(n9271), .ZN(n14900) );
  INV_X1 U11805 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9984) );
  NAND2_X1 U11806 ( .A1(n9324), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n9275) );
  INV_X1 U11807 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9272) );
  OR2_X1 U11808 ( .A1(n7213), .A2(n9272), .ZN(n9274) );
  OAI211_X1 U11809 ( .C1(n9327), .C2(n9984), .A(n9275), .B(n9274), .ZN(n9276)
         );
  INV_X1 U11810 ( .A(n9276), .ZN(n9277) );
  NAND2_X2 U11811 ( .A1(n9278), .A2(n9277), .ZN(n15212) );
  OR2_X1 U11812 ( .A1(n8898), .A2(n12482), .ZN(n9281) );
  MUX2_X1 U11813 ( .A(n15212), .B(n15482), .S(n9020), .Z(n9285) );
  MUX2_X1 U11814 ( .A(n15212), .B(n15482), .S(n9344), .Z(n9283) );
  NAND2_X1 U11815 ( .A1(n9287), .A2(n9286), .ZN(n9288) );
  OR2_X1 U11816 ( .A1(n8898), .A2(n12485), .ZN(n9290) );
  INV_X1 U11817 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9292) );
  NAND2_X1 U11818 ( .A1(n9293), .A2(n9292), .ZN(n9294) );
  NAND2_X1 U11819 ( .A1(n9321), .A2(n9294), .ZN(n15220) );
  INV_X1 U11820 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9299) );
  NAND2_X1 U11821 ( .A1(n9252), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9298) );
  NAND2_X1 U11822 ( .A1(n9296), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9297) );
  OAI211_X1 U11823 ( .C1(n9308), .C2(n9299), .A(n9298), .B(n9297), .ZN(n9300)
         );
  INV_X1 U11824 ( .A(n9300), .ZN(n9301) );
  MUX2_X1 U11825 ( .A(n15222), .B(n14998), .S(n9020), .Z(n9304) );
  MUX2_X1 U11826 ( .A(n15222), .B(n14998), .S(n9344), .Z(n9303) );
  XNOR2_X1 U11827 ( .A(n9321), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n14854) );
  NAND2_X1 U11828 ( .A1(n14854), .A2(n9323), .ZN(n9311) );
  INV_X1 U11829 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9307) );
  NAND2_X1 U11830 ( .A1(n9252), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9306) );
  NAND2_X1 U11831 ( .A1(n8906), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9305) );
  OAI211_X1 U11832 ( .C1(n9308), .C2(n9307), .A(n9306), .B(n9305), .ZN(n9309)
         );
  INV_X1 U11833 ( .A(n9309), .ZN(n9310) );
  XNOR2_X1 U11834 ( .A(n9312), .B(SI_27_), .ZN(n9313) );
  INV_X1 U11835 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15596) );
  OR2_X1 U11836 ( .A1(n8898), .A2(n15596), .ZN(n9315) );
  MUX2_X1 U11837 ( .A(n15213), .B(n15469), .S(n9076), .Z(n9319) );
  MUX2_X1 U11838 ( .A(n15213), .B(n15469), .S(n9344), .Z(n9317) );
  INV_X1 U11839 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n14851) );
  INV_X1 U11840 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9320) );
  OAI21_X1 U11841 ( .B1(n9321), .B2(n14851), .A(n9320), .ZN(n9322) );
  NAND2_X1 U11842 ( .A1(n15192), .A2(n9323), .ZN(n9330) );
  INV_X1 U11843 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n10032) );
  NAND2_X1 U11844 ( .A1(n9324), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n9326) );
  NAND2_X1 U11845 ( .A1(n9252), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9325) );
  OAI211_X1 U11846 ( .C1(n9327), .C2(n10032), .A(n9326), .B(n9325), .ZN(n9328)
         );
  INV_X1 U11847 ( .A(n9328), .ZN(n9329) );
  INV_X1 U11848 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n13259) );
  OR2_X1 U11849 ( .A1(n8898), .A2(n13259), .ZN(n9334) );
  MUX2_X1 U11850 ( .A(n15181), .B(n15462), .S(n9344), .Z(n9337) );
  MUX2_X1 U11851 ( .A(n15181), .B(n15462), .S(n9076), .Z(n9336) );
  INV_X1 U11852 ( .A(n9338), .ZN(n9341) );
  INV_X1 U11853 ( .A(n9339), .ZN(n9340) );
  AND2_X1 U11854 ( .A1(n9341), .A2(n9340), .ZN(n9353) );
  NAND2_X1 U11855 ( .A1(n9366), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9343) );
  XNOR2_X1 U11856 ( .A(n9343), .B(n9342), .ZN(n10956) );
  OR2_X1 U11857 ( .A1(n10956), .A2(P1_U3086), .ZN(n10644) );
  NAND2_X1 U11858 ( .A1(n15152), .A2(n14996), .ZN(n9346) );
  OR2_X1 U11859 ( .A1(n15152), .A2(n14996), .ZN(n9345) );
  OR2_X1 U11860 ( .A1(n8720), .A2(n8722), .ZN(n11441) );
  AND2_X1 U11861 ( .A1(n9404), .A2(n11441), .ZN(n9401) );
  NAND2_X1 U11862 ( .A1(n9405), .A2(n9401), .ZN(n9364) );
  NOR2_X1 U11863 ( .A1(n9348), .A2(n9347), .ZN(n9360) );
  NOR2_X1 U11864 ( .A1(n9352), .A2(n9349), .ZN(n9350) );
  AOI211_X1 U11865 ( .C1(n9353), .C2(n9351), .A(n10644), .B(n9350), .ZN(n9356)
         );
  INV_X1 U11866 ( .A(n9352), .ZN(n9355) );
  INV_X1 U11867 ( .A(n9353), .ZN(n9354) );
  INV_X1 U11868 ( .A(n9359), .ZN(n9362) );
  INV_X1 U11869 ( .A(n9360), .ZN(n9361) );
  OAI22_X1 U11870 ( .A1(n9364), .A2(n9363), .B1(n9362), .B2(n9361), .ZN(n9380)
         );
  INV_X1 U11871 ( .A(n10644), .ZN(n11736) );
  INV_X1 U11872 ( .A(P1_B_REG_SCAN_IN), .ZN(n9365) );
  AOI21_X1 U11873 ( .B1(n10788), .B2(n11736), .A(n9365), .ZN(n9379) );
  AND2_X1 U11874 ( .A1(n8722), .A2(n6539), .ZN(n10941) );
  OR2_X1 U11875 ( .A1(n10941), .A2(n10944), .ZN(n10958) );
  OAI21_X1 U11876 ( .B1(n9370), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9368) );
  MUX2_X1 U11877 ( .A(n9368), .B(P1_IR_REG_31__SCAN_IN), .S(n9367), .Z(n9369)
         );
  NAND2_X1 U11878 ( .A1(n9369), .A2(n9373), .ZN(n12480) );
  INV_X1 U11879 ( .A(n12480), .ZN(n9377) );
  MUX2_X1 U11880 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9374), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n9375) );
  NAND2_X1 U11881 ( .A1(n9375), .A2(n6603), .ZN(n12487) );
  NOR2_X1 U11882 ( .A1(n12222), .A2(n12487), .ZN(n9376) );
  AND2_X1 U11883 ( .A1(n10956), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10532) );
  INV_X1 U11884 ( .A(n10944), .ZN(n10789) );
  NAND3_X1 U11885 ( .A1(n11438), .A2(n15150), .A3(n15426), .ZN(n9378) );
  AOI22_X1 U11886 ( .A1(n9380), .A2(n11736), .B1(n9379), .B2(n9378), .ZN(n9414) );
  INV_X1 U11887 ( .A(n15168), .ZN(n15164) );
  INV_X1 U11888 ( .A(n15204), .ZN(n15202) );
  INV_X1 U11889 ( .A(n12736), .ZN(n12739) );
  NAND2_X1 U11890 ( .A1(n15265), .A2(n15274), .ZN(n12730) );
  OR2_X1 U11891 ( .A1(n15265), .A2(n15274), .ZN(n9381) );
  NAND2_X1 U11892 ( .A1(n12730), .A2(n9381), .ZN(n15259) );
  INV_X1 U11893 ( .A(n15289), .ZN(n15284) );
  XNOR2_X1 U11894 ( .A(n15277), .B(n13194), .ZN(n12729) );
  NAND2_X1 U11895 ( .A1(n9382), .A2(n12725), .ZN(n15317) );
  INV_X1 U11896 ( .A(n15317), .ZN(n15329) );
  NAND2_X1 U11897 ( .A1(n15370), .A2(n12717), .ZN(n12694) );
  INV_X1 U11898 ( .A(n12694), .ZN(n15396) );
  XNOR2_X1 U11899 ( .A(n15559), .B(n15011), .ZN(n12160) );
  INV_X1 U11900 ( .A(n12160), .ZN(n12173) );
  XNOR2_X1 U11901 ( .A(n12605), .B(n15010), .ZN(n12382) );
  INV_X1 U11902 ( .A(n12382), .ZN(n12377) );
  XNOR2_X1 U11903 ( .A(n15553), .B(n15009), .ZN(n12610) );
  INV_X1 U11904 ( .A(n15750), .ZN(n9385) );
  NAND4_X1 U11905 ( .A1(n15429), .A2(n11539), .A3(n9385), .A4(n11447), .ZN(
        n9386) );
  XNOR2_X1 U11906 ( .A(n11521), .B(n15018), .ZN(n11509) );
  NOR2_X1 U11907 ( .A1(n9386), .A2(n11509), .ZN(n9387) );
  XNOR2_X1 U11908 ( .A(n15731), .B(n15016), .ZN(n11713) );
  NAND4_X1 U11909 ( .A1(n11959), .A2(n9387), .A3(n11709), .A4(n11713), .ZN(
        n9388) );
  XNOR2_X1 U11910 ( .A(n12655), .B(n12432), .ZN(n12011) );
  XNOR2_X1 U11911 ( .A(n15812), .B(n11955), .ZN(n11755) );
  XNOR2_X1 U11912 ( .A(n12426), .B(n15012), .ZN(n12026) );
  NAND3_X1 U11913 ( .A1(n12610), .A2(n7978), .A3(n12026), .ZN(n9389) );
  NOR4_X1 U11914 ( .A1(n15405), .A2(n12173), .A3(n12377), .A4(n9389), .ZN(
        n9390) );
  XNOR2_X1 U11915 ( .A(n15537), .B(n15006), .ZN(n12714) );
  AND4_X1 U11916 ( .A1(n15396), .A2(n9390), .A3(n12714), .A4(n15357), .ZN(
        n9391) );
  AND2_X1 U11917 ( .A1(n15299), .A2(n9391), .ZN(n9392) );
  NAND4_X1 U11918 ( .A1(n12729), .A2(n15329), .A3(n9392), .A4(n12720), .ZN(
        n9393) );
  NOR3_X1 U11919 ( .A1(n15259), .A2(n15284), .A3(n9393), .ZN(n9395) );
  XNOR2_X2 U11920 ( .A(n15488), .B(n14999), .ZN(n15244) );
  NAND4_X1 U11921 ( .A1(n12734), .A2(n9395), .A3(n15235), .A4(n15244), .ZN(
        n9396) );
  NOR4_X1 U11922 ( .A1(n15164), .A2(n15202), .A3(n12739), .A4(n9396), .ZN(
        n9399) );
  INV_X1 U11923 ( .A(n9397), .ZN(n9403) );
  XOR2_X1 U11924 ( .A(n15177), .B(n15447), .Z(n9398) );
  NAND3_X1 U11925 ( .A1(n9399), .A2(n9403), .A3(n9398), .ZN(n9400) );
  XNOR2_X1 U11926 ( .A(n9400), .B(n15748), .ZN(n9411) );
  INV_X1 U11927 ( .A(n11441), .ZN(n9410) );
  INV_X1 U11928 ( .A(n9401), .ZN(n9402) );
  NOR2_X1 U11929 ( .A1(n9403), .A2(n9402), .ZN(n9408) );
  INV_X1 U11930 ( .A(n9404), .ZN(n9407) );
  INV_X1 U11931 ( .A(n9405), .ZN(n9406) );
  MUX2_X1 U11932 ( .A(n9408), .B(n9407), .S(n9406), .Z(n9409) );
  AOI21_X1 U11933 ( .B1(n9411), .B2(n9410), .A(n9409), .ZN(n9412) );
  NAND3_X1 U11934 ( .A1(n9415), .A2(n9414), .A3(n9413), .ZN(P1_U3242) );
  NOR2_X4 U11935 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n9481) );
  INV_X1 U11936 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9426) );
  NAND2_X1 U11937 ( .A1(n9428), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9424) );
  XNOR2_X2 U11938 ( .A(n9427), .B(n9426), .ZN(n9853) );
  INV_X1 U11939 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n9429) );
  NOR2_X1 U11940 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .ZN(n9436) );
  INV_X1 U11941 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n9440) );
  INV_X1 U11942 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9437) );
  INV_X1 U11943 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n9453) );
  AND2_X2 U11944 ( .A1(n9507), .A2(n7219), .ZN(n9678) );
  NAND2_X1 U11945 ( .A1(n10336), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9445) );
  INV_X1 U11946 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n14145) );
  INV_X1 U11947 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11607) );
  INV_X1 U11948 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n11694) );
  INV_X1 U11949 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9711) );
  NAND2_X1 U11950 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_23__SCAN_IN), 
        .ZN(n9452) );
  INV_X1 U11951 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n14098) );
  XNOR2_X1 U11952 ( .A(n9808), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n14385) );
  INV_X1 U11953 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n9454) );
  AND2_X1 U11954 ( .A1(n9454), .A2(n9453), .ZN(n9456) );
  NAND2_X1 U11955 ( .A1(n14385), .A2(n7527), .ZN(n9466) );
  INV_X1 U11956 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n10014) );
  NAND2_X1 U11957 ( .A1(n10328), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9463) );
  NAND2_X1 U11958 ( .A1(n10321), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9462) );
  OAI211_X1 U11959 ( .C1(n10014), .C2(n9861), .A(n9463), .B(n9462), .ZN(n9464)
         );
  INV_X1 U11960 ( .A(n9464), .ZN(n9465) );
  NAND2_X1 U11961 ( .A1(n10336), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9467) );
  INV_X1 U11962 ( .A(n14705), .ZN(n14103) );
  INV_X1 U11963 ( .A(n9469), .ZN(n9785) );
  NAND2_X1 U11964 ( .A1(n9774), .A2(n14098), .ZN(n9470) );
  NAND2_X1 U11965 ( .A1(n9785), .A2(n9470), .ZN(n14430) );
  OR2_X1 U11966 ( .A1(n14430), .A2(n9517), .ZN(n9475) );
  INV_X1 U11967 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n14431) );
  NAND2_X1 U11968 ( .A1(n10321), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9472) );
  NAND2_X1 U11969 ( .A1(n10329), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n9471) );
  OAI211_X1 U11970 ( .C1(n14431), .C2(n10325), .A(n9472), .B(n9471), .ZN(n9473) );
  INV_X1 U11971 ( .A(n9473), .ZN(n9474) );
  NAND2_X1 U11972 ( .A1(n9475), .A2(n9474), .ZN(n14198) );
  INV_X1 U11973 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9476) );
  INV_X1 U11974 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9477) );
  INV_X1 U11975 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n11029) );
  NOR2_X1 U11976 ( .A1(n6542), .A2(n10525), .ZN(n9485) );
  NOR2_X1 U11977 ( .A1(n10573), .A2(n8069), .ZN(n9479) );
  NAND2_X1 U11978 ( .A1(n9507), .A2(n9479), .ZN(n9489) );
  NAND2_X1 U11979 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9480) );
  MUX2_X1 U11980 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9480), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n9483) );
  NAND2_X1 U11981 ( .A1(n9483), .A2(n9482), .ZN(n14220) );
  INV_X1 U11982 ( .A(n14220), .ZN(n11007) );
  INV_X1 U11983 ( .A(n9484), .ZN(n11026) );
  AOI21_X1 U11984 ( .B1(n9478), .B2(n9487), .A(n9486), .ZN(n9488) );
  INV_X1 U11985 ( .A(n12091), .ZN(n9496) );
  NAND2_X1 U11986 ( .A1(n10321), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n9493) );
  INV_X1 U11987 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n12669) );
  OR2_X1 U11988 ( .A1(n9861), .A2(n12669), .ZN(n9492) );
  INV_X1 U11989 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n12673) );
  OR2_X1 U11990 ( .A1(n9517), .A2(n12673), .ZN(n9491) );
  INV_X1 U11991 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n12668) );
  OR2_X1 U11992 ( .A1(n10325), .A2(n12668), .ZN(n9490) );
  INV_X1 U11993 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n14222) );
  NAND2_X1 U11994 ( .A1(n6542), .A2(SI_0_), .ZN(n9495) );
  XNOR2_X1 U11995 ( .A(n9494), .B(n9495), .ZN(n14834) );
  MUX2_X1 U11996 ( .A(n14222), .B(n14834), .S(n9507), .Z(n10414) );
  INV_X1 U11997 ( .A(n10414), .ZN(n13267) );
  NAND2_X1 U11998 ( .A1(n10168), .A2(n13267), .ZN(n12089) );
  NAND2_X1 U11999 ( .A1(n13274), .A2(n12688), .ZN(n9501) );
  NAND2_X1 U12000 ( .A1(n12093), .A2(n9501), .ZN(n12103) );
  NAND2_X1 U12001 ( .A1(n10321), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n9506) );
  INV_X1 U12002 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n12117) );
  OR2_X1 U12003 ( .A1(n9517), .A2(n12117), .ZN(n9505) );
  INV_X1 U12004 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9502) );
  OR2_X1 U12005 ( .A1(n9861), .A2(n9502), .ZN(n9504) );
  INV_X1 U12006 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n11028) );
  OR2_X1 U12007 ( .A1(n10325), .A2(n11028), .ZN(n9503) );
  NAND2_X1 U12008 ( .A1(n9678), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n9513) );
  MUX2_X1 U12009 ( .A(n9693), .B(n9508), .S(P2_IR_REG_2__SCAN_IN), .Z(n9511)
         );
  OAI211_X1 U12010 ( .C1(n9793), .C2(n10624), .A(n9513), .B(n9512), .ZN(n9864)
         );
  NAND2_X1 U12011 ( .A1(n9678), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n9516) );
  NAND2_X1 U12012 ( .A1(n9510), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9514) );
  MUX2_X1 U12013 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9514), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n9515) );
  OR2_X1 U12014 ( .A1(n9510), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n9546) );
  AND2_X1 U12015 ( .A1(n9515), .A2(n9546), .ZN(n15855) );
  NAND2_X1 U12016 ( .A1(n10321), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n9522) );
  OR2_X1 U12017 ( .A1(n9517), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9521) );
  INV_X1 U12018 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9518) );
  OR2_X1 U12019 ( .A1(n9861), .A2(n9518), .ZN(n9520) );
  INV_X1 U12020 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11033) );
  OR2_X1 U12021 ( .A1(n10325), .A2(n11033), .ZN(n9519) );
  NAND2_X1 U12022 ( .A1(n12103), .A2(n9523), .ZN(n9527) );
  NAND2_X1 U12023 ( .A1(n12085), .A2(n15917), .ZN(n12248) );
  NAND2_X1 U12024 ( .A1(n12248), .A2(n14214), .ZN(n9525) );
  AND2_X1 U12025 ( .A1(n12085), .A2(n12104), .ZN(n9524) );
  AOI22_X1 U12026 ( .A1(n9525), .A2(n12407), .B1(n9524), .B2(n15917), .ZN(
        n9526) );
  NAND2_X1 U12027 ( .A1(n9527), .A2(n9526), .ZN(n11988) );
  NAND2_X1 U12028 ( .A1(n10328), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9533) );
  INV_X1 U12029 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9528) );
  OR2_X1 U12030 ( .A1(n6793), .A2(n9528), .ZN(n9532) );
  OAI21_X1 U12031 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n9539), .ZN(n14105) );
  OR2_X1 U12032 ( .A1(n9517), .A2(n14105), .ZN(n9531) );
  INV_X1 U12033 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9529) );
  OR2_X1 U12034 ( .A1(n9861), .A2(n9529), .ZN(n9530) );
  NAND2_X1 U12035 ( .A1(n10336), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n9536) );
  NAND2_X1 U12036 ( .A1(n9546), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9534) );
  XNOR2_X1 U12037 ( .A(n9534), .B(P2_IR_REG_4__SCAN_IN), .ZN(n14246) );
  NAND2_X1 U12038 ( .A1(n9727), .A2(n14246), .ZN(n9535) );
  OAI211_X1 U12039 ( .C1(n9793), .C2(n10626), .A(n9536), .B(n9535), .ZN(n14107) );
  XNOR2_X1 U12040 ( .A(n14213), .B(n14107), .ZN(n10383) );
  INV_X1 U12041 ( .A(n10383), .ZN(n11992) );
  NAND2_X1 U12042 ( .A1(n11988), .A2(n11992), .ZN(n11987) );
  NAND2_X1 U12043 ( .A1(n12179), .A2(n15924), .ZN(n9537) );
  NAND2_X1 U12044 ( .A1(n10321), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9545) );
  INV_X1 U12045 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n12185) );
  OR2_X1 U12046 ( .A1(n10325), .A2(n12185), .ZN(n9544) );
  INV_X1 U12047 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9538) );
  NAND2_X1 U12048 ( .A1(n9539), .A2(n9538), .ZN(n9540) );
  NAND2_X1 U12049 ( .A1(n9571), .A2(n9540), .ZN(n12188) );
  OR2_X1 U12050 ( .A1(n9517), .A2(n12188), .ZN(n9543) );
  INV_X1 U12051 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9541) );
  OR2_X1 U12052 ( .A1(n9861), .A2(n9541), .ZN(n9542) );
  INV_X1 U12053 ( .A(n9546), .ZN(n9548) );
  INV_X1 U12054 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n9547) );
  NAND2_X1 U12055 ( .A1(n9548), .A2(n9547), .ZN(n9550) );
  NAND2_X1 U12056 ( .A1(n9550), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9549) );
  MUX2_X1 U12057 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9549), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n9553) );
  INV_X1 U12058 ( .A(n9550), .ZN(n9552) );
  NAND2_X1 U12059 ( .A1(n9552), .A2(n9551), .ZN(n9566) );
  AOI22_X1 U12060 ( .A1(n10336), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9727), 
        .B2(n15869), .ZN(n9555) );
  NAND2_X1 U12061 ( .A1(n10569), .A2(n10335), .ZN(n9554) );
  XNOR2_X1 U12062 ( .A(n14212), .B(n12315), .ZN(n10386) );
  INV_X1 U12063 ( .A(n10386), .ZN(n12181) );
  NAND2_X1 U12064 ( .A1(n14104), .A2(n12412), .ZN(n9556) );
  NAND2_X1 U12065 ( .A1(n12177), .A2(n9556), .ZN(n11967) );
  NAND2_X1 U12066 ( .A1(n10328), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9561) );
  INV_X1 U12067 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9557) );
  OR2_X1 U12068 ( .A1(n6793), .A2(n9557), .ZN(n9560) );
  INV_X1 U12069 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9570) );
  XNOR2_X1 U12070 ( .A(n9571), .B(n9570), .ZN(n12352) );
  OR2_X1 U12071 ( .A1(n9517), .A2(n12352), .ZN(n9559) );
  OR2_X1 U12072 ( .A1(n9861), .A2(n15942), .ZN(n9558) );
  NAND4_X1 U12073 ( .A1(n9561), .A2(n9560), .A3(n9559), .A4(n9558), .ZN(n14211) );
  NAND2_X1 U12074 ( .A1(n9566), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9562) );
  XNOR2_X1 U12075 ( .A(n9562), .B(P2_IR_REG_6__SCAN_IN), .ZN(n14260) );
  AOI22_X1 U12076 ( .A1(n10336), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9727), 
        .B2(n14260), .ZN(n9564) );
  OR2_X1 U12077 ( .A1(n10570), .A2(n9793), .ZN(n9563) );
  NAND2_X1 U12078 ( .A1(n12336), .A2(n15932), .ZN(n9565) );
  NAND2_X1 U12079 ( .A1(n10582), .A2(n10335), .ZN(n9569) );
  OAI21_X1 U12080 ( .B1(n9566), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9567) );
  XNOR2_X1 U12081 ( .A(n9567), .B(P2_IR_REG_7__SCAN_IN), .ZN(n14272) );
  AOI22_X1 U12082 ( .A1(n10336), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9727), 
        .B2(n14272), .ZN(n9568) );
  NAND2_X1 U12083 ( .A1(n10328), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9576) );
  INV_X1 U12084 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n12397) );
  OR2_X1 U12085 ( .A1(n6793), .A2(n12397), .ZN(n9575) );
  INV_X1 U12086 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n12339) );
  OAI21_X1 U12087 ( .B1(n9571), .B2(n9570), .A(n12339), .ZN(n9572) );
  NAND2_X1 U12088 ( .A1(n9572), .A2(n9584), .ZN(n12345) );
  OR2_X1 U12089 ( .A1(n9517), .A2(n12345), .ZN(n9574) );
  INV_X1 U12090 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n11014) );
  OR2_X1 U12091 ( .A1(n9861), .A2(n11014), .ZN(n9573) );
  AND2_X1 U12092 ( .A1(n12398), .A2(n12548), .ZN(n12317) );
  NAND2_X1 U12093 ( .A1(n10617), .A2(n10335), .ZN(n9582) );
  NAND2_X1 U12094 ( .A1(n9577), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9578) );
  MUX2_X1 U12095 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9578), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n9580) );
  INV_X1 U12096 ( .A(n9577), .ZN(n9626) );
  INV_X1 U12097 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n9579) );
  NAND2_X1 U12098 ( .A1(n9626), .A2(n9579), .ZN(n9609) );
  NAND2_X1 U12099 ( .A1(n9580), .A2(n9609), .ZN(n11059) );
  INV_X1 U12100 ( .A(n11059), .ZN(n11042) );
  AOI22_X1 U12101 ( .A1(n10336), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n9727), 
        .B2(n11042), .ZN(n9581) );
  NAND2_X1 U12102 ( .A1(n10328), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9590) );
  INV_X1 U12103 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n12402) );
  OR2_X1 U12104 ( .A1(n6793), .A2(n12402), .ZN(n9589) );
  INV_X1 U12105 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9583) );
  NAND2_X1 U12106 ( .A1(n9584), .A2(n9583), .ZN(n9585) );
  NAND2_X1 U12107 ( .A1(n9599), .A2(n9585), .ZN(n12358) );
  OR2_X1 U12108 ( .A1(n9517), .A2(n12358), .ZN(n9588) );
  INV_X1 U12109 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9586) );
  OR2_X1 U12110 ( .A1(n9861), .A2(n9586), .ZN(n9587) );
  NAND4_X1 U12111 ( .A1(n9590), .A2(n9589), .A3(n9588), .A4(n9587), .ZN(n14209) );
  NOR2_X1 U12112 ( .A1(n12331), .A2(n14209), .ZN(n9591) );
  OAI21_X1 U12113 ( .B1(n12398), .B2(n12548), .A(n12471), .ZN(n9593) );
  NOR2_X1 U12114 ( .A1(n12471), .A2(n12548), .ZN(n9592) );
  AOI22_X1 U12115 ( .A1(n9593), .A2(n12331), .B1(n12342), .B2(n9592), .ZN(
        n12273) );
  NAND2_X1 U12116 ( .A1(n10621), .A2(n10335), .ZN(n9596) );
  NAND2_X1 U12117 ( .A1(n9609), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9594) );
  XNOR2_X1 U12118 ( .A(n9594), .B(P2_IR_REG_9__SCAN_IN), .ZN(n11094) );
  AOI22_X1 U12119 ( .A1(n10336), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n9727), 
        .B2(n11094), .ZN(n9595) );
  NAND2_X1 U12120 ( .A1(n10328), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n9604) );
  INV_X1 U12121 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9597) );
  OR2_X1 U12122 ( .A1(n6793), .A2(n9597), .ZN(n9603) );
  NAND2_X1 U12123 ( .A1(n9599), .A2(n9598), .ZN(n9600) );
  NAND2_X1 U12124 ( .A1(n9617), .A2(n9600), .ZN(n12465) );
  OR2_X1 U12125 ( .A1(n9517), .A2(n12465), .ZN(n9602) );
  INV_X1 U12126 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10030) );
  OR2_X1 U12127 ( .A1(n9861), .A2(n10030), .ZN(n9601) );
  OR2_X1 U12128 ( .A1(n12366), .A2(n12329), .ZN(n9605) );
  AND2_X1 U12129 ( .A1(n12273), .A2(n9605), .ZN(n9608) );
  INV_X1 U12130 ( .A(n9605), .ZN(n9606) );
  XNOR2_X1 U12131 ( .A(n12468), .B(n12329), .ZN(n10388) );
  INV_X1 U12132 ( .A(n9609), .ZN(n9610) );
  INV_X1 U12133 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9921) );
  NAND2_X1 U12134 ( .A1(n9610), .A2(n9921), .ZN(n9612) );
  NAND2_X1 U12135 ( .A1(n9612), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9611) );
  MUX2_X1 U12136 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9611), .S(
        P2_IR_REG_10__SCAN_IN), .Z(n9613) );
  OR2_X1 U12137 ( .A1(n9612), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n9623) );
  AOI22_X1 U12138 ( .A1(n10336), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n9727), 
        .B2(n11114), .ZN(n9614) );
  NAND2_X1 U12139 ( .A1(n10328), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9622) );
  INV_X1 U12140 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n12517) );
  OR2_X1 U12141 ( .A1(n6793), .A2(n12517), .ZN(n9621) );
  INV_X1 U12142 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9616) );
  NAND2_X1 U12143 ( .A1(n9617), .A2(n9616), .ZN(n9618) );
  NAND2_X1 U12144 ( .A1(n9630), .A2(n9618), .ZN(n12243) );
  OR2_X1 U12145 ( .A1(n9517), .A2(n12243), .ZN(n9620) );
  INV_X1 U12146 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n12520) );
  OR2_X1 U12147 ( .A1(n9861), .A2(n12520), .ZN(n9619) );
  NAND4_X1 U12148 ( .A1(n9622), .A2(n9621), .A3(n9620), .A4(n9619), .ZN(n14207) );
  NAND2_X1 U12149 ( .A1(n10761), .A2(n10335), .ZN(n9629) );
  NAND2_X1 U12150 ( .A1(n9623), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9624) );
  MUX2_X1 U12151 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9624), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n9627) );
  NAND2_X1 U12152 ( .A1(n9626), .A2(n9625), .ZN(n9650) );
  NAND2_X1 U12153 ( .A1(n9627), .A2(n9650), .ZN(n11601) );
  INV_X1 U12154 ( .A(n11601), .ZN(n11594) );
  AOI22_X1 U12155 ( .A1(n10336), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n9727), 
        .B2(n11594), .ZN(n9628) );
  AND2_X2 U12156 ( .A1(n9629), .A2(n9628), .ZN(n14823) );
  NAND2_X1 U12157 ( .A1(n10328), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n9635) );
  INV_X1 U12158 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n14820) );
  OR2_X1 U12159 ( .A1(n6793), .A2(n14820), .ZN(n9634) );
  NAND2_X1 U12160 ( .A1(n9630), .A2(n14145), .ZN(n9631) );
  NAND2_X1 U12161 ( .A1(n9641), .A2(n9631), .ZN(n14148) );
  OR2_X1 U12162 ( .A1(n9517), .A2(n14148), .ZN(n9633) );
  INV_X1 U12163 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n14779) );
  OR2_X1 U12164 ( .A1(n9861), .A2(n14779), .ZN(n9632) );
  OR2_X1 U12165 ( .A1(n14823), .A2(n14066), .ZN(n14665) );
  NAND2_X1 U12166 ( .A1(n10646), .A2(n10335), .ZN(n9638) );
  NAND2_X1 U12167 ( .A1(n9650), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9636) );
  XNOR2_X1 U12168 ( .A(n9636), .B(P2_IR_REG_12__SCAN_IN), .ZN(n15895) );
  AOI22_X1 U12169 ( .A1(n10336), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n9727), 
        .B2(n15895), .ZN(n9637) );
  INV_X1 U12170 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9905) );
  OR2_X1 U12171 ( .A1(n6793), .A2(n9905), .ZN(n9646) );
  INV_X1 U12172 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n9639) );
  OR2_X1 U12173 ( .A1(n10325), .A2(n9639), .ZN(n9645) );
  INV_X1 U12174 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9640) );
  NAND2_X1 U12175 ( .A1(n9641), .A2(n9640), .ZN(n9642) );
  NAND2_X1 U12176 ( .A1(n9656), .A2(n9642), .ZN(n14660) );
  OR2_X1 U12177 ( .A1(n9517), .A2(n14660), .ZN(n9644) );
  INV_X1 U12178 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11595) );
  OR2_X1 U12179 ( .A1(n9861), .A2(n11595), .ZN(n9643) );
  NAND4_X1 U12180 ( .A1(n9646), .A2(n9645), .A3(n9644), .A4(n9643), .ZN(n14206) );
  NAND2_X1 U12181 ( .A1(n14769), .A2(n14206), .ZN(n10389) );
  NAND2_X1 U12182 ( .A1(n14665), .A2(n10389), .ZN(n9648) );
  NOR2_X1 U12183 ( .A1(n12242), .A2(n14207), .ZN(n12498) );
  AOI21_X1 U12184 ( .B1(n14823), .B2(n14066), .A(n12498), .ZN(n9647) );
  OR2_X1 U12185 ( .A1(n14769), .A2(n14206), .ZN(n10390) );
  OAI21_X1 U12186 ( .B1(n9648), .B2(n9647), .A(n10390), .ZN(n9649) );
  INV_X1 U12187 ( .A(n9649), .ZN(n14621) );
  OR2_X1 U12188 ( .A1(n10650), .A2(n9793), .ZN(n9655) );
  INV_X1 U12189 ( .A(n9650), .ZN(n9652) );
  NAND2_X1 U12190 ( .A1(n9652), .A2(n9651), .ZN(n9662) );
  NAND2_X1 U12191 ( .A1(n9662), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9653) );
  XNOR2_X1 U12192 ( .A(n9653), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U12193 ( .A1(n10336), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n9727), 
        .B2(n11698), .ZN(n9654) );
  NAND2_X1 U12194 ( .A1(n10321), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n9661) );
  INV_X1 U12195 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n14644) );
  OR2_X1 U12196 ( .A1(n10325), .A2(n14644), .ZN(n9660) );
  NAND2_X1 U12197 ( .A1(n9656), .A2(n11607), .ZN(n9657) );
  NAND2_X1 U12198 ( .A1(n9666), .A2(n9657), .ZN(n14643) );
  OR2_X1 U12199 ( .A1(n9517), .A2(n14643), .ZN(n9659) );
  INV_X1 U12200 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n14766) );
  OR2_X1 U12201 ( .A1(n9861), .A2(n14766), .ZN(n9658) );
  NAND2_X1 U12202 ( .A1(n14816), .A2(n14205), .ZN(n14623) );
  NAND2_X1 U12203 ( .A1(n10776), .A2(n10335), .ZN(n9665) );
  OAI21_X1 U12204 ( .B1(n9662), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9663) );
  XNOR2_X1 U12205 ( .A(n9663), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11940) );
  AOI22_X1 U12206 ( .A1(n10336), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n9727), 
        .B2(n11940), .ZN(n9664) );
  AND2_X2 U12207 ( .A1(n9665), .A2(n9664), .ZN(n14620) );
  NAND2_X1 U12208 ( .A1(n10321), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n9672) );
  INV_X1 U12209 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11701) );
  OR2_X1 U12210 ( .A1(n9861), .A2(n11701), .ZN(n9671) );
  NAND2_X1 U12211 ( .A1(n9666), .A2(n11694), .ZN(n9667) );
  NAND2_X1 U12212 ( .A1(n9681), .A2(n9667), .ZN(n14617) );
  OR2_X1 U12213 ( .A1(n9517), .A2(n14617), .ZN(n9670) );
  INV_X1 U12214 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n9668) );
  OR2_X1 U12215 ( .A1(n10325), .A2(n9668), .ZN(n9669) );
  NAND2_X1 U12216 ( .A1(n14620), .A2(n14637), .ZN(n9688) );
  AND2_X1 U12217 ( .A1(n14623), .A2(n9688), .ZN(n9673) );
  AND2_X1 U12218 ( .A1(n14621), .A2(n9673), .ZN(n9676) );
  INV_X1 U12219 ( .A(n9673), .ZN(n9675) );
  NAND2_X1 U12220 ( .A1(n14641), .A2(n14205), .ZN(n9828) );
  OR2_X1 U12221 ( .A1(n14641), .A2(n14205), .ZN(n9674) );
  NAND2_X1 U12222 ( .A1(n9828), .A2(n9674), .ZN(n14632) );
  OR2_X1 U12223 ( .A1(n6746), .A2(n9693), .ZN(n9677) );
  XNOR2_X1 U12224 ( .A(n9677), .B(P2_IR_REG_15__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U12225 ( .A1(n9678), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n9727), 
        .B2(n12210), .ZN(n9679) );
  NAND2_X1 U12226 ( .A1(n10328), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n9687) );
  INV_X1 U12227 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9680) );
  OR2_X1 U12228 ( .A1(n6793), .A2(n9680), .ZN(n9686) );
  INV_X1 U12229 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n14183) );
  NAND2_X1 U12230 ( .A1(n9681), .A2(n14183), .ZN(n9682) );
  NAND2_X1 U12231 ( .A1(n9699), .A2(n9682), .ZN(n14602) );
  OR2_X1 U12232 ( .A1(n9517), .A2(n14602), .ZN(n9685) );
  INV_X1 U12233 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9683) );
  OR2_X1 U12234 ( .A1(n9861), .A2(n9683), .ZN(n9684) );
  INV_X1 U12235 ( .A(n14609), .ZN(n14592) );
  INV_X1 U12236 ( .A(n9688), .ZN(n9689) );
  AND2_X1 U12237 ( .A1(n14592), .A2(n14606), .ZN(n9690) );
  NAND2_X1 U12238 ( .A1(n14605), .A2(n14089), .ZN(n9691) );
  NAND2_X1 U12239 ( .A1(n10768), .A2(n10335), .ZN(n9697) );
  OR2_X1 U12240 ( .A1(n9694), .A2(n9693), .ZN(n9695) );
  XNOR2_X1 U12241 ( .A(n9695), .B(P2_IR_REG_16__SCAN_IN), .ZN(n14291) );
  AOI22_X1 U12242 ( .A1(n10336), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n9727), 
        .B2(n14291), .ZN(n9696) );
  INV_X1 U12244 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9698) );
  NAND2_X1 U12245 ( .A1(n9699), .A2(n9698), .ZN(n9700) );
  NAND2_X1 U12246 ( .A1(n9712), .A2(n9700), .ZN(n14572) );
  OR2_X1 U12247 ( .A1(n14572), .A2(n9517), .ZN(n9704) );
  NAND2_X1 U12248 ( .A1(n10321), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n9703) );
  NAND2_X1 U12249 ( .A1(n10329), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n9702) );
  INV_X1 U12250 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n14583) );
  OR2_X1 U12251 ( .A1(n10325), .A2(n14583), .ZN(n9701) );
  NAND4_X1 U12252 ( .A1(n9704), .A2(n9703), .A3(n9702), .A4(n9701), .ZN(n14203) );
  XNOR2_X1 U12253 ( .A(n14580), .B(n14203), .ZN(n14586) );
  NAND2_X1 U12254 ( .A1(n14580), .A2(n14203), .ZN(n9706) );
  NAND2_X1 U12255 ( .A1(n10772), .A2(n10335), .ZN(n9710) );
  NAND2_X1 U12256 ( .A1(n9707), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9708) );
  XNOR2_X1 U12257 ( .A(n9708), .B(P2_IR_REG_17__SCAN_IN), .ZN(n14309) );
  AOI22_X1 U12258 ( .A1(n10336), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n9727), 
        .B2(n14309), .ZN(n9709) );
  NAND2_X1 U12259 ( .A1(n9712), .A2(n9711), .ZN(n9713) );
  NAND2_X1 U12260 ( .A1(n9721), .A2(n9713), .ZN(n14567) );
  AOI22_X1 U12261 ( .A1(n10321), .A2(P2_REG0_REG_17__SCAN_IN), .B1(n10328), 
        .B2(P2_REG2_REG_17__SCAN_IN), .ZN(n9715) );
  NAND2_X1 U12262 ( .A1(n10329), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n9714) );
  OAI211_X1 U12263 ( .C1(n14567), .C2(n9517), .A(n9715), .B(n9714), .ZN(n14575) );
  XNOR2_X1 U12264 ( .A(n14566), .B(n14575), .ZN(n10392) );
  INV_X1 U12265 ( .A(n14537), .ZN(n9726) );
  NAND2_X1 U12266 ( .A1(n11003), .A2(n10335), .ZN(n9720) );
  NAND2_X1 U12267 ( .A1(n9879), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9717) );
  MUX2_X1 U12268 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9717), .S(
        P2_IR_REG_18__SCAN_IN), .Z(n9718) );
  AND2_X1 U12269 ( .A1(n9718), .A2(n9431), .ZN(n14312) );
  AOI22_X1 U12270 ( .A1(n10336), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n9727), 
        .B2(n14312), .ZN(n9719) );
  INV_X2 U12272 ( .A(n14552), .ZN(n14737) );
  NAND2_X1 U12273 ( .A1(n9721), .A2(n6860), .ZN(n9722) );
  NAND2_X1 U12274 ( .A1(n9748), .A2(n9722), .ZN(n14549) );
  OR2_X1 U12275 ( .A1(n14549), .A2(n9517), .ZN(n9725) );
  AOI22_X1 U12276 ( .A1(n10321), .A2(P2_REG0_REG_18__SCAN_IN), .B1(n10328), 
        .B2(P2_REG2_REG_18__SCAN_IN), .ZN(n9724) );
  NAND2_X1 U12277 ( .A1(n10329), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n9723) );
  NAND2_X1 U12278 ( .A1(n14737), .A2(n14563), .ZN(n9837) );
  NAND2_X1 U12279 ( .A1(n14505), .A2(n9837), .ZN(n14503) );
  AOI22_X1 U12280 ( .A1(n10336), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n11860), 
        .B2(n9727), .ZN(n9728) );
  XNOR2_X1 U12281 ( .A(n9748), .B(P2_REG3_REG_19__SCAN_IN), .ZN(n14528) );
  NAND2_X1 U12282 ( .A1(n14528), .A2(n7527), .ZN(n9735) );
  INV_X1 U12283 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9732) );
  NAND2_X1 U12284 ( .A1(n10328), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n9731) );
  NAND2_X1 U12285 ( .A1(n10321), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n9730) );
  OAI211_X1 U12286 ( .C1(n9732), .C2(n9861), .A(n9731), .B(n9730), .ZN(n9733)
         );
  INV_X1 U12287 ( .A(n9733), .ZN(n9734) );
  NAND2_X1 U12288 ( .A1(n9735), .A2(n9734), .ZN(n14201) );
  XNOR2_X1 U12289 ( .A(n14732), .B(n14201), .ZN(n14522) );
  INV_X1 U12290 ( .A(n14522), .ZN(n14532) );
  NAND2_X1 U12291 ( .A1(n14732), .A2(n14201), .ZN(n9736) );
  NAND2_X1 U12292 ( .A1(n11550), .A2(n10335), .ZN(n9738) );
  NAND2_X1 U12293 ( .A1(n10336), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9737) );
  INV_X1 U12295 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9740) );
  NAND2_X1 U12296 ( .A1(n9749), .A2(n9740), .ZN(n9741) );
  NAND2_X1 U12297 ( .A1(n9773), .A2(n9741), .ZN(n14492) );
  INV_X1 U12298 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n14723) );
  NAND2_X1 U12299 ( .A1(n10321), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9743) );
  NAND2_X1 U12300 ( .A1(n10328), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9742) );
  OAI211_X1 U12301 ( .C1(n14723), .C2(n9861), .A(n9743), .B(n9742), .ZN(n9744)
         );
  INV_X1 U12302 ( .A(n9744), .ZN(n9745) );
  NAND2_X1 U12303 ( .A1(n10336), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9746) );
  INV_X1 U12304 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n14034) );
  INV_X1 U12305 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n14122) );
  OAI21_X1 U12306 ( .B1(n9748), .B2(n14034), .A(n14122), .ZN(n9750) );
  AND2_X1 U12307 ( .A1(n9750), .A2(n9749), .ZN(n14516) );
  NAND2_X1 U12308 ( .A1(n14516), .A2(n7527), .ZN(n9755) );
  INV_X1 U12309 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n14801) );
  NAND2_X1 U12310 ( .A1(n10328), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n9752) );
  NAND2_X1 U12311 ( .A1(n10329), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n9751) );
  OAI211_X1 U12312 ( .C1(n6793), .C2(n14801), .A(n9752), .B(n9751), .ZN(n9753)
         );
  INV_X1 U12313 ( .A(n9753), .ZN(n9754) );
  NAND2_X1 U12314 ( .A1(n9755), .A2(n9754), .ZN(n14484) );
  INV_X1 U12315 ( .A(n14491), .ZN(n14799) );
  OAI21_X1 U12316 ( .B1(n14515), .B2(n14484), .A(n14200), .ZN(n9757) );
  INV_X1 U12317 ( .A(n14515), .ZN(n14803) );
  NOR2_X1 U12318 ( .A1(n14200), .A2(n14484), .ZN(n9756) );
  AOI22_X1 U12319 ( .A1(n14799), .A2(n9757), .B1(n14803), .B2(n9756), .ZN(
        n9758) );
  NAND2_X1 U12320 ( .A1(n9760), .A2(n9759), .ZN(n9761) );
  AND2_X1 U12321 ( .A1(n9762), .A2(n9761), .ZN(n11724) );
  NAND2_X1 U12322 ( .A1(n11724), .A2(n10335), .ZN(n9764) );
  NAND2_X1 U12323 ( .A1(n10336), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9763) );
  XNOR2_X1 U12324 ( .A(n9773), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n14475) );
  NAND2_X1 U12325 ( .A1(n14475), .A2(n7527), .ZN(n9769) );
  INV_X1 U12326 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9969) );
  NAND2_X1 U12327 ( .A1(n10328), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n9766) );
  NAND2_X1 U12328 ( .A1(n10329), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n9765) );
  OAI211_X1 U12329 ( .C1(n6793), .C2(n9969), .A(n9766), .B(n9765), .ZN(n9767)
         );
  INV_X1 U12330 ( .A(n9767), .ZN(n9768) );
  NAND2_X1 U12331 ( .A1(n9769), .A2(n9768), .ZN(n14485) );
  INV_X1 U12332 ( .A(n14485), .ZN(n14056) );
  XNOR2_X1 U12333 ( .A(n12751), .B(n14056), .ZN(n14470) );
  INV_X1 U12334 ( .A(n14470), .ZN(n14464) );
  NAND2_X1 U12335 ( .A1(n12751), .A2(n14485), .ZN(n9770) );
  NAND2_X1 U12336 ( .A1(n14467), .A2(n9770), .ZN(n14460) );
  NAND2_X1 U12337 ( .A1(n11734), .A2(n10335), .ZN(n9772) );
  NAND2_X1 U12338 ( .A1(n10336), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n9771) );
  INV_X1 U12339 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n14135) );
  INV_X1 U12340 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n14024) );
  OAI21_X1 U12341 ( .B1(n9773), .B2(n14135), .A(n14024), .ZN(n9775) );
  NAND2_X1 U12342 ( .A1(n9775), .A2(n9774), .ZN(n14454) );
  OR2_X1 U12343 ( .A1(n14454), .A2(n9517), .ZN(n9781) );
  INV_X1 U12344 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9778) );
  NAND2_X1 U12345 ( .A1(n10328), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n9777) );
  NAND2_X1 U12346 ( .A1(n10321), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n9776) );
  OAI211_X1 U12347 ( .C1(n9778), .C2(n9861), .A(n9777), .B(n9776), .ZN(n9779)
         );
  INV_X1 U12348 ( .A(n9779), .ZN(n9780) );
  NAND2_X1 U12349 ( .A1(n9781), .A2(n9780), .ZN(n14199) );
  XNOR2_X1 U12350 ( .A(n14710), .B(n14199), .ZN(n14446) );
  INV_X1 U12351 ( .A(n14446), .ZN(n14459) );
  NAND2_X1 U12352 ( .A1(n14460), .A2(n14459), .ZN(n14458) );
  INV_X1 U12353 ( .A(n14710), .ZN(n14457) );
  INV_X1 U12354 ( .A(n14199), .ZN(n12795) );
  NAND2_X1 U12355 ( .A1(n14458), .A2(n7990), .ZN(n14429) );
  NAND2_X1 U12356 ( .A1(n12477), .A2(n10335), .ZN(n9783) );
  NAND2_X1 U12357 ( .A1(n10336), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9782) );
  INV_X1 U12358 ( .A(n9784), .ZN(n9796) );
  INV_X1 U12359 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n14081) );
  NAND2_X1 U12360 ( .A1(n9785), .A2(n14081), .ZN(n9786) );
  NAND2_X1 U12361 ( .A1(n14413), .A2(n7527), .ZN(n9791) );
  INV_X1 U12362 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9972) );
  NAND2_X1 U12363 ( .A1(n10321), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9788) );
  NAND2_X1 U12364 ( .A1(n10328), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9787) );
  OAI211_X1 U12365 ( .C1(n9861), .C2(n9972), .A(n9788), .B(n9787), .ZN(n9789)
         );
  INV_X1 U12366 ( .A(n9789), .ZN(n9790) );
  NAND2_X1 U12367 ( .A1(n14700), .A2(n14197), .ZN(n9792) );
  NAND2_X1 U12368 ( .A1(n10336), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9794) );
  INV_X1 U12369 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9795) );
  NAND2_X1 U12370 ( .A1(n9796), .A2(n9795), .ZN(n9797) );
  NAND2_X1 U12371 ( .A1(n9808), .A2(n9797), .ZN(n14167) );
  INV_X1 U12372 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9800) );
  NAND2_X1 U12373 ( .A1(n10328), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n9799) );
  NAND2_X1 U12374 ( .A1(n10321), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n9798) );
  OAI211_X1 U12375 ( .C1(n9800), .C2(n9861), .A(n9799), .B(n9798), .ZN(n9801)
         );
  INV_X1 U12376 ( .A(n9801), .ZN(n9802) );
  NAND2_X1 U12377 ( .A1(n10336), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9805) );
  INV_X1 U12378 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n12820) );
  INV_X1 U12379 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9807) );
  OAI21_X1 U12380 ( .B1(n9808), .B2(n12820), .A(n9807), .ZN(n9809) );
  NAND2_X1 U12381 ( .A1(n14366), .A2(n7527), .ZN(n9814) );
  NAND2_X1 U12382 ( .A1(n10321), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9811) );
  NAND2_X1 U12383 ( .A1(n10328), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9810) );
  OAI211_X1 U12384 ( .C1(n9904), .C2(n9861), .A(n9811), .B(n9810), .ZN(n9812)
         );
  INV_X1 U12385 ( .A(n9812), .ZN(n9813) );
  INV_X1 U12386 ( .A(n10168), .ZN(n12086) );
  NAND2_X1 U12387 ( .A1(n12086), .A2(n13267), .ZN(n10381) );
  INV_X1 U12388 ( .A(n10381), .ZN(n12084) );
  NAND2_X1 U12389 ( .A1(n13274), .A2(n12099), .ZN(n12105) );
  NAND2_X1 U12390 ( .A1(n12107), .A2(n12105), .ZN(n9816) );
  XNOR2_X1 U12391 ( .A(n14215), .B(n9864), .ZN(n12102) );
  NAND2_X1 U12392 ( .A1(n9816), .A2(n12102), .ZN(n12109) );
  NAND2_X1 U12393 ( .A1(n12085), .A2(n12114), .ZN(n9817) );
  NAND2_X1 U12394 ( .A1(n12109), .A2(n9817), .ZN(n12254) );
  NAND2_X1 U12395 ( .A1(n12179), .A2(n14107), .ZN(n12180) );
  NAND2_X1 U12396 ( .A1(n14104), .A2(n12315), .ZN(n11970) );
  NAND2_X1 U12397 ( .A1(n12336), .A2(n12350), .ZN(n9818) );
  NAND2_X1 U12398 ( .A1(n12398), .A2(n14210), .ZN(n9819) );
  OR2_X1 U12399 ( .A1(n12398), .A2(n14210), .ZN(n9820) );
  XNOR2_X1 U12400 ( .A(n12331), .B(n14209), .ZN(n12319) );
  INV_X1 U12401 ( .A(n12319), .ZN(n12327) );
  OR2_X1 U12402 ( .A1(n12331), .A2(n12471), .ZN(n9822) );
  INV_X1 U12403 ( .A(n10388), .ZN(n12275) );
  INV_X1 U12404 ( .A(n12329), .ZN(n14208) );
  NAND2_X1 U12405 ( .A1(n12366), .A2(n14208), .ZN(n12234) );
  NAND2_X1 U12406 ( .A1(n9865), .A2(n14207), .ZN(n9824) );
  XNOR2_X1 U12407 ( .A(n14151), .B(n14653), .ZN(n10391) );
  INV_X1 U12408 ( .A(n14206), .ZN(n14635) );
  AND2_X1 U12409 ( .A1(n14769), .A2(n14635), .ZN(n9826) );
  OR2_X1 U12410 ( .A1(n14769), .A2(n14635), .ZN(n9827) );
  INV_X1 U12411 ( .A(n14637), .ZN(n14204) );
  NAND2_X1 U12412 ( .A1(n14620), .A2(n14204), .ZN(n9829) );
  NAND2_X1 U12413 ( .A1(n14759), .A2(n14637), .ZN(n9830) );
  NAND2_X1 U12414 ( .A1(n14605), .A2(n14576), .ZN(n9832) );
  NAND2_X1 U12415 ( .A1(n14580), .A2(n14594), .ZN(n9833) );
  OR2_X1 U12416 ( .A1(n14580), .A2(n14594), .ZN(n9834) );
  INV_X1 U12417 ( .A(n14201), .ZN(n14539) );
  NAND2_X1 U12418 ( .A1(n14732), .A2(n14539), .ZN(n14507) );
  INV_X1 U12419 ( .A(n14575), .ZN(n14538) );
  NAND2_X1 U12420 ( .A1(n14566), .A2(n14538), .ZN(n14541) );
  AND3_X1 U12421 ( .A1(n14507), .A2(n9837), .A3(n14541), .ZN(n9841) );
  INV_X1 U12422 ( .A(n14566), .ZN(n14809) );
  NAND3_X1 U12423 ( .A1(n9837), .A2(n14809), .A3(n14575), .ZN(n9835) );
  NAND3_X1 U12424 ( .A1(n9835), .A2(n14539), .A3(n14505), .ZN(n9836) );
  NAND2_X1 U12425 ( .A1(n9836), .A2(n14530), .ZN(n9839) );
  NAND4_X1 U12426 ( .A1(n9837), .A2(n14809), .A3(n14201), .A4(n14575), .ZN(
        n9838) );
  OAI211_X1 U12427 ( .C1(n14539), .C2(n14505), .A(n9839), .B(n9838), .ZN(n9840) );
  NOR2_X1 U12428 ( .A1(n14716), .A2(n14485), .ZN(n14444) );
  INV_X1 U12429 ( .A(n14484), .ZN(n14057) );
  NAND2_X1 U12430 ( .A1(n14515), .A2(n14057), .ZN(n14468) );
  OAI21_X1 U12431 ( .B1(n14799), .B2(n14200), .A(n14468), .ZN(n14443) );
  INV_X1 U12432 ( .A(n14443), .ZN(n9842) );
  NAND2_X1 U12433 ( .A1(n9843), .A2(n9842), .ZN(n9851) );
  AOI21_X1 U12434 ( .B1(n14803), .B2(n14484), .A(n14200), .ZN(n9844) );
  OR2_X1 U12435 ( .A1(n9844), .A2(n14491), .ZN(n9847) );
  NAND2_X1 U12436 ( .A1(n14200), .A2(n14484), .ZN(n9845) );
  OR2_X1 U12437 ( .A1(n14515), .A2(n9845), .ZN(n9846) );
  OAI211_X1 U12438 ( .C1(n12751), .C2(n14056), .A(n9847), .B(n9846), .ZN(n9848) );
  INV_X1 U12439 ( .A(n9848), .ZN(n14442) );
  OAI21_X1 U12440 ( .B1(n14444), .B2(n14442), .A(n14446), .ZN(n9849) );
  INV_X1 U12441 ( .A(n9849), .ZN(n9850) );
  OAI21_X1 U12442 ( .B1(n14441), .B2(n9851), .A(n9850), .ZN(n9852) );
  OR2_X1 U12443 ( .A1(n9433), .A2(n14332), .ZN(n9855) );
  INV_X1 U12444 ( .A(n9853), .ZN(n10382) );
  NAND2_X1 U12445 ( .A1(n10382), .A2(n10375), .ZN(n9854) );
  AOI21_X1 U12446 ( .B1(n9857), .B2(n9856), .A(n14634), .ZN(n9863) );
  INV_X1 U12447 ( .A(n9433), .ZN(n10333) );
  NAND2_X1 U12448 ( .A1(n10333), .A2(n10375), .ZN(n11022) );
  INV_X1 U12449 ( .A(n9858), .ZN(n14361) );
  INV_X1 U12450 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9994) );
  NAND2_X1 U12451 ( .A1(n10321), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9860) );
  NAND2_X1 U12452 ( .A1(n10328), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9859) );
  OAI211_X1 U12453 ( .C1(n9994), .C2(n9861), .A(n9860), .B(n9859), .ZN(n9862)
         );
  AOI21_X1 U12454 ( .B1(n14361), .B2(n7527), .A(n9862), .ZN(n10379) );
  OAI22_X1 U12455 ( .A1(n7884), .A2(n14636), .B1(n10379), .B2(n14638), .ZN(
        n14045) );
  NAND2_X1 U12456 ( .A1(n9853), .A2(n14332), .ZN(n10405) );
  NAND2_X1 U12457 ( .A1(n12113), .A2(n15917), .ZN(n12251) );
  NAND2_X1 U12458 ( .A1(n11996), .A2(n15924), .ZN(n12187) );
  INV_X1 U12459 ( .A(n9867), .ZN(n14639) );
  NOR2_X4 U12460 ( .A1(n14564), .A2(n14737), .ZN(n14548) );
  NOR2_X4 U12461 ( .A1(n14452), .A2(n14705), .ZN(n14436) );
  NAND2_X1 U12462 ( .A1(n14369), .A2(n14383), .ZN(n9868) );
  NAND2_X1 U12463 ( .A1(n9868), .A2(n10450), .ZN(n9869) );
  NOR2_X1 U12464 ( .A1(n14359), .A2(n9869), .ZN(n14370) );
  AOI21_X1 U12465 ( .B1(n14770), .B2(n14369), .A(n14370), .ZN(n9870) );
  INV_X1 U12466 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9872) );
  NAND2_X1 U12467 ( .A1(n9874), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9875) );
  MUX2_X1 U12468 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9875), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n9877) );
  NAND2_X1 U12469 ( .A1(n9877), .A2(n9876), .ZN(n12484) );
  OAI21_X1 U12470 ( .B1(n9879), .B2(n9878), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9880) );
  MUX2_X1 U12471 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9880), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n9881) );
  NAND2_X1 U12472 ( .A1(n9881), .A2(n9874), .ZN(n12478) );
  OR2_X1 U12473 ( .A1(n9883), .A2(n9882), .ZN(n9884) );
  NAND2_X1 U12474 ( .A1(n9885), .A2(n9884), .ZN(n11020) );
  OR2_X1 U12475 ( .A1(n11022), .A2(n10485), .ZN(n10491) );
  NOR4_X1 U12476 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n9894) );
  INV_X1 U12477 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n15904) );
  INV_X1 U12478 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n15905) );
  INV_X1 U12479 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n15906) );
  INV_X1 U12480 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n15903) );
  NAND4_X1 U12481 ( .A1(n15904), .A2(n15905), .A3(n15906), .A4(n15903), .ZN(
        n9891) );
  NOR4_X1 U12482 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n9889) );
  NOR4_X1 U12483 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n9888) );
  NOR4_X1 U12484 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9887) );
  NOR4_X1 U12485 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n9886) );
  NAND4_X1 U12486 ( .A1(n9889), .A2(n9888), .A3(n9887), .A4(n9886), .ZN(n9890)
         );
  NOR4_X1 U12487 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n9891), .A4(n9890), .ZN(n9893) );
  NOR4_X1 U12488 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n9892) );
  NAND3_X1 U12489 ( .A1(n9894), .A2(n9893), .A3(n9892), .ZN(n9898) );
  XNOR2_X1 U12490 ( .A(n12225), .B(P2_B_REG_SCAN_IN), .ZN(n9895) );
  NAND2_X1 U12491 ( .A1(n12478), .A2(n9895), .ZN(n9897) );
  INV_X1 U12492 ( .A(n12484), .ZN(n9896) );
  NAND2_X1 U12493 ( .A1(n11682), .A2(n10478), .ZN(n11858) );
  INV_X1 U12494 ( .A(n11866), .ZN(n10400) );
  INV_X1 U12495 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15912) );
  NAND2_X1 U12496 ( .A1(n15902), .A2(n15912), .ZN(n9900) );
  NAND2_X1 U12497 ( .A1(n12478), .A2(n12484), .ZN(n9899) );
  NAND2_X1 U12498 ( .A1(n9900), .A2(n9899), .ZN(n15913) );
  NAND2_X1 U12499 ( .A1(n10488), .A2(n15913), .ZN(n9901) );
  OR2_X1 U12500 ( .A1(n11858), .A2(n9901), .ZN(n12372) );
  NAND2_X1 U12501 ( .A1(n12225), .A2(n12484), .ZN(n9903) );
  INV_X1 U12502 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15909) );
  NAND2_X1 U12503 ( .A1(n15902), .A2(n15909), .ZN(n9902) );
  NOR2_X4 U12504 ( .A1(n12372), .A2(n15910), .ZN(n15944) );
  NOR4_X1 U12505 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .A3(P2_REG2_REG_17__SCAN_IN), .A4(n10030), .ZN(n9909) );
  INV_X1 U12506 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n15840) );
  NOR4_X1 U12507 ( .A1(P3_REG0_REG_31__SCAN_IN), .A2(n9905), .A3(n11029), .A4(
        n15840), .ZN(n9908) );
  NOR4_X1 U12508 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .A3(P1_REG0_REG_16__SCAN_IN), .A4(P1_REG1_REG_6__SCAN_IN), .ZN(n9907)
         );
  NOR4_X1 U12509 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_REG1_REG_15__SCAN_IN), 
        .A3(P2_REG1_REG_23__SCAN_IN), .A4(P1_REG2_REG_2__SCAN_IN), .ZN(n9906)
         );
  NAND4_X1 U12510 ( .A1(n9909), .A2(n9908), .A3(n9907), .A4(n9906), .ZN(n9917)
         );
  INV_X1 U12511 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n9960) );
  AND4_X1 U12512 ( .A1(P3_REG0_REG_5__SCAN_IN), .A2(P1_REG1_REG_22__SCAN_IN), 
        .A3(P1_REG2_REG_21__SCAN_IN), .A4(n7530), .ZN(n9911) );
  AND4_X1 U12513 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(n10661), .A3(n13277), .A4(
        n9994), .ZN(n9910) );
  NAND4_X1 U12514 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_REG0_REG_6__SCAN_IN), 
        .A3(n9911), .A4(n9910), .ZN(n9916) );
  NOR4_X1 U12515 ( .A1(P1_REG0_REG_25__SCAN_IN), .A2(P1_IR_REG_30__SCAN_IN), 
        .A3(P2_REG2_REG_31__SCAN_IN), .A4(P3_ADDR_REG_12__SCAN_IN), .ZN(n9914)
         );
  NOR4_X1 U12516 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P1_REG1_REG_1__SCAN_IN), .A4(P1_ADDR_REG_12__SCAN_IN), .ZN(n9913)
         );
  NOR4_X1 U12517 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(P2_REG2_REG_16__SCAN_IN), 
        .A3(n10032), .A4(n14945), .ZN(n9912) );
  NAND4_X1 U12518 ( .A1(P2_REG0_REG_6__SCAN_IN), .A2(n9914), .A3(n9913), .A4(
        n9912), .ZN(n9915) );
  NOR4_X1 U12519 ( .A1(n9918), .A2(n9917), .A3(n9916), .A4(n9915), .ZN(n9919)
         );
  NAND2_X1 U12520 ( .A1(n9919), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n9920) );
  INV_X1 U12521 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n15769) );
  NOR4_X1 U12522 ( .A1(n9920), .A2(n15769), .A3(P3_DATAO_REG_12__SCAN_IN), 
        .A4(P2_D_REG_5__SCAN_IN), .ZN(n9934) );
  NAND4_X1 U12523 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P1_DATAO_REG_1__SCAN_IN), .A4(P2_REG0_REG_4__SCAN_IN), .ZN(n9923) );
  NAND2_X1 U12524 ( .A1(n9921), .A2(n6818), .ZN(n9922) );
  NOR4_X1 U12525 ( .A1(n9923), .A2(n9922), .A3(P2_IR_REG_22__SCAN_IN), .A4(
        P2_REG0_REG_20__SCAN_IN), .ZN(n9933) );
  NAND4_X1 U12526 ( .A1(n10639), .A2(SI_10_), .A3(P1_REG1_REG_12__SCAN_IN), 
        .A4(P1_REG0_REG_17__SCAN_IN), .ZN(n9928) );
  NAND4_X1 U12527 ( .A1(n9924), .A2(P3_IR_REG_17__SCAN_IN), .A3(
        P3_IR_REG_28__SCAN_IN), .A4(P3_REG3_REG_16__SCAN_IN), .ZN(n9927) );
  NAND4_X1 U12528 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P3_REG0_REG_10__SCAN_IN), 
        .A3(P3_REG3_REG_3__SCAN_IN), .A4(P3_REG2_REG_22__SCAN_IN), .ZN(n9926)
         );
  OR4_X1 U12529 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(SI_6_), .A3(SI_2_), .A4(
        P1_IR_REG_31__SCAN_IN), .ZN(n9925) );
  NOR4_X1 U12530 ( .A1(n9928), .A2(n9927), .A3(n9926), .A4(n9925), .ZN(n9932)
         );
  NAND4_X1 U12531 ( .A1(P3_REG0_REG_11__SCAN_IN), .A2(P3_DATAO_REG_13__SCAN_IN), .A3(n10769), .A4(n7897), .ZN(n9930) );
  INV_X1 U12532 ( .A(P1_WR_REG_SCAN_IN), .ZN(n9982) );
  NAND4_X1 U12533 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(SI_8_), .A3(
        P1_REG1_REG_29__SCAN_IN), .A4(n9982), .ZN(n9929) );
  NOR2_X1 U12534 ( .A1(n9930), .A2(n9929), .ZN(n9931) );
  NAND4_X1 U12535 ( .A1(n9934), .A2(n9933), .A3(n9932), .A4(n9931), .ZN(n9945)
         );
  INV_X1 U12536 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n11307) );
  NAND4_X1 U12537 ( .A1(P2_REG1_REG_25__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), 
        .A3(P2_REG0_REG_22__SCAN_IN), .A4(n11307), .ZN(n9935) );
  NOR3_X1 U12538 ( .A1(P3_REG1_REG_25__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .A3(n9935), .ZN(n9936) );
  NAND3_X1 U12539 ( .A1(P3_REG2_REG_21__SCAN_IN), .A2(n9936), .A3(n11812), 
        .ZN(n9944) );
  NOR4_X1 U12540 ( .A1(P3_REG3_REG_25__SCAN_IN), .A2(P2_DATAO_REG_29__SCAN_IN), 
        .A3(P2_D_REG_21__SCAN_IN), .A4(n9955), .ZN(n9940) );
  NOR4_X1 U12541 ( .A1(P2_REG0_REG_30__SCAN_IN), .A2(P3_REG1_REG_17__SCAN_IN), 
        .A3(P1_REG2_REG_20__SCAN_IN), .A4(n10967), .ZN(n9939) );
  INV_X1 U12542 ( .A(SI_26_), .ZN(n12286) );
  NOR4_X1 U12543 ( .A1(P2_REG1_REG_27__SCAN_IN), .A2(P3_REG0_REG_13__SCAN_IN), 
        .A3(P2_REG1_REG_4__SCAN_IN), .A4(n12286), .ZN(n9938) );
  NOR4_X1 U12544 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P1_REG2_REG_25__SCAN_IN), .A4(n10743), .ZN(n9937) );
  NAND4_X1 U12545 ( .A1(n9940), .A2(n9939), .A3(n9938), .A4(n9937), .ZN(n9943)
         );
  NOR4_X1 U12546 ( .A1(P1_RD_REG_SCAN_IN), .A2(P2_RD_REG_SCAN_IN), .A3(
        P1_ADDR_REG_4__SCAN_IN), .A4(P2_ADDR_REG_5__SCAN_IN), .ZN(n9941) );
  NAND4_X1 U12547 ( .A1(SI_1_), .A2(P2_REG2_REG_24__SCAN_IN), .A3(n9941), .A4(
        n12223), .ZN(n9942) );
  NOR4_X1 U12548 ( .A1(n9945), .A2(n9944), .A3(n9943), .A4(n9942), .ZN(n9949)
         );
  NOR4_X1 U12549 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P3_DATAO_REG_9__SCAN_IN), 
        .A3(P1_ADDR_REG_14__SCAN_IN), .A4(n10108), .ZN(n9948) );
  INV_X1 U12550 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n12883) );
  INV_X1 U12551 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15825) );
  NOR4_X1 U12552 ( .A1(P3_REG0_REG_14__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), 
        .A3(n12883), .A4(n15825), .ZN(n9947) );
  NOR4_X1 U12553 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), 
        .A3(P1_IR_REG_8__SCAN_IN), .A4(n15903), .ZN(n9946) );
  NAND4_X1 U12554 ( .A1(n9949), .A2(n9948), .A3(n9947), .A4(n9946), .ZN(n9953)
         );
  INV_X1 U12555 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n15767) );
  NOR4_X1 U12556 ( .A1(P3_REG2_REG_29__SCAN_IN), .A2(P2_ADDR_REG_16__SCAN_IN), 
        .A3(n15767), .A4(n12017), .ZN(n9951) );
  INV_X1 U12557 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15765) );
  NOR4_X1 U12558 ( .A1(P1_REG2_REG_31__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), 
        .A3(n15765), .A4(n10671), .ZN(n9950) );
  NAND2_X1 U12559 ( .A1(n9951), .A2(n9950), .ZN(n9952) );
  OAI21_X1 U12560 ( .B1(n9953), .B2(n9952), .A(keyinput125), .ZN(n10148) );
  INV_X1 U12561 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n15020) );
  AOI22_X1 U12562 ( .A1(n9955), .A2(keyinput88), .B1(keyinput38), .B2(n15593), 
        .ZN(n9954) );
  OAI221_X1 U12563 ( .B1(n9955), .B2(keyinput88), .C1(n15593), .C2(keyinput38), 
        .A(n9954), .ZN(n9966) );
  AOI22_X1 U12564 ( .A1(n15310), .A2(keyinput35), .B1(n9957), .B2(keyinput61), 
        .ZN(n9956) );
  OAI221_X1 U12565 ( .B1(n15310), .B2(keyinput35), .C1(n9957), .C2(keyinput61), 
        .A(n9956), .ZN(n9965) );
  INV_X1 U12566 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9959) );
  AOI22_X1 U12567 ( .A1(n9960), .A2(keyinput66), .B1(keyinput15), .B2(n9959), 
        .ZN(n9958) );
  OAI221_X1 U12568 ( .B1(n9960), .B2(keyinput66), .C1(n9959), .C2(keyinput15), 
        .A(n9958), .ZN(n9964) );
  INV_X1 U12569 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n9962) );
  AOI22_X1 U12570 ( .A1(n15904), .A2(keyinput81), .B1(n9962), .B2(keyinput33), 
        .ZN(n9961) );
  OAI221_X1 U12571 ( .B1(n15904), .B2(keyinput81), .C1(n9962), .C2(keyinput33), 
        .A(n9961), .ZN(n9963) );
  NOR4_X1 U12572 ( .A1(n9966), .A2(n9965), .A3(n9964), .A4(n9963), .ZN(n10002)
         );
  AOI22_X1 U12573 ( .A1(n13732), .A2(keyinput117), .B1(keyinput97), .B2(n11307), .ZN(n9967) );
  OAI221_X1 U12574 ( .B1(n13732), .B2(keyinput117), .C1(n11307), .C2(
        keyinput97), .A(n9967), .ZN(n9976) );
  AOI22_X1 U12575 ( .A1(n9969), .A2(keyinput109), .B1(n13860), .B2(keyinput62), 
        .ZN(n9968) );
  OAI221_X1 U12576 ( .B1(n9969), .B2(keyinput109), .C1(n13860), .C2(keyinput62), .A(n9968), .ZN(n9975) );
  INV_X1 U12577 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n15052) );
  INV_X1 U12578 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10600) );
  AOI22_X1 U12579 ( .A1(n15052), .A2(keyinput29), .B1(n10600), .B2(keyinput114), .ZN(n9970) );
  OAI221_X1 U12580 ( .B1(n15052), .B2(keyinput29), .C1(n10600), .C2(
        keyinput114), .A(n9970), .ZN(n9974) );
  AOI22_X1 U12581 ( .A1(n9972), .A2(keyinput126), .B1(n7897), .B2(keyinput108), 
        .ZN(n9971) );
  OAI221_X1 U12582 ( .B1(n9972), .B2(keyinput126), .C1(n7897), .C2(keyinput108), .A(n9971), .ZN(n9973) );
  NOR4_X1 U12583 ( .A1(n9976), .A2(n9975), .A3(n9974), .A4(n9973), .ZN(n10001)
         );
  INV_X1 U12584 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n9978) );
  AOI22_X1 U12585 ( .A1(n9979), .A2(keyinput92), .B1(keyinput70), .B2(n9978), 
        .ZN(n9977) );
  OAI221_X1 U12586 ( .B1(n9979), .B2(keyinput92), .C1(n9978), .C2(keyinput70), 
        .A(n9977), .ZN(n9989) );
  INV_X1 U12587 ( .A(SI_8_), .ZN(n10519) );
  AOI22_X1 U12588 ( .A1(n10769), .A2(keyinput90), .B1(keyinput56), .B2(n10519), 
        .ZN(n9980) );
  OAI221_X1 U12589 ( .B1(n10769), .B2(keyinput90), .C1(n10519), .C2(keyinput56), .A(n9980), .ZN(n9988) );
  AOI22_X1 U12590 ( .A1(n11701), .A2(keyinput64), .B1(keyinput19), .B2(n9982), 
        .ZN(n9981) );
  OAI221_X1 U12591 ( .B1(n11701), .B2(keyinput64), .C1(n9982), .C2(keyinput19), 
        .A(n9981), .ZN(n9987) );
  AOI22_X1 U12592 ( .A1(n9985), .A2(keyinput20), .B1(keyinput7), .B2(n9984), 
        .ZN(n9983) );
  OAI221_X1 U12593 ( .B1(n9985), .B2(keyinput20), .C1(n9984), .C2(keyinput7), 
        .A(n9983), .ZN(n9986) );
  NOR4_X1 U12594 ( .A1(n9989), .A2(n9988), .A3(n9987), .A4(n9986), .ZN(n10000)
         );
  INV_X1 U12595 ( .A(keyinput6), .ZN(n10066) );
  INV_X1 U12596 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15880) );
  XOR2_X1 U12597 ( .A(n15880), .B(keyinput110), .Z(n9990) );
  OAI21_X1 U12598 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n10066), .A(n9990), .ZN(
        n9998) );
  AOI22_X1 U12599 ( .A1(n12223), .A2(keyinput106), .B1(keyinput23), .B2(n14431), .ZN(n9991) );
  OAI221_X1 U12600 ( .B1(n12223), .B2(keyinput106), .C1(n14431), .C2(
        keyinput23), .A(n9991), .ZN(n9997) );
  AOI22_X1 U12601 ( .A1(n10661), .A2(keyinput24), .B1(keyinput113), .B2(n9872), 
        .ZN(n9992) );
  OAI221_X1 U12602 ( .B1(n10661), .B2(keyinput24), .C1(n9872), .C2(keyinput113), .A(n9992), .ZN(n9996) );
  AOI22_X1 U12603 ( .A1(n13277), .A2(keyinput43), .B1(keyinput104), .B2(n9994), 
        .ZN(n9993) );
  OAI221_X1 U12604 ( .B1(n13277), .B2(keyinput43), .C1(n9994), .C2(keyinput104), .A(n9993), .ZN(n9995) );
  NOR4_X1 U12605 ( .A1(n9998), .A2(n9997), .A3(n9996), .A4(n9995), .ZN(n9999)
         );
  NAND4_X1 U12606 ( .A1(n10002), .A2(n10001), .A3(n10000), .A4(n9999), .ZN(
        n10147) );
  AOI22_X1 U12607 ( .A1(n13991), .A2(keyinput14), .B1(keyinput40), .B2(n15825), 
        .ZN(n10003) );
  OAI221_X1 U12608 ( .B1(n13991), .B2(keyinput14), .C1(n15825), .C2(keyinput40), .A(n10003), .ZN(n10008) );
  INV_X1 U12609 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n12910) );
  INV_X1 U12610 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n15715) );
  AOI22_X1 U12611 ( .A1(n12910), .A2(keyinput55), .B1(keyinput49), .B2(n15715), 
        .ZN(n10004) );
  OAI221_X1 U12612 ( .B1(n12910), .B2(keyinput55), .C1(n15715), .C2(keyinput49), .A(n10004), .ZN(n10007) );
  INV_X1 U12613 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12942) );
  AOI22_X1 U12614 ( .A1(n13722), .A2(keyinput32), .B1(keyinput5), .B2(n12942), 
        .ZN(n10005) );
  OAI221_X1 U12615 ( .B1(n13722), .B2(keyinput32), .C1(n12942), .C2(keyinput5), 
        .A(n10005), .ZN(n10006) );
  NOR3_X1 U12616 ( .A1(n10008), .A2(n10007), .A3(n10006), .ZN(n10027) );
  INV_X1 U12617 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n15856) );
  AOI22_X1 U12618 ( .A1(n8862), .A2(keyinput124), .B1(n15856), .B2(keyinput18), 
        .ZN(n10009) );
  OAI221_X1 U12619 ( .B1(n8862), .B2(keyinput124), .C1(n15856), .C2(keyinput18), .A(n10009), .ZN(n10012) );
  AOI22_X1 U12620 ( .A1(n12533), .A2(keyinput118), .B1(n12286), .B2(keyinput50), .ZN(n10010) );
  OAI221_X1 U12621 ( .B1(n12533), .B2(keyinput118), .C1(n12286), .C2(
        keyinput50), .A(n10010), .ZN(n10011) );
  NOR2_X1 U12622 ( .A1(n10012), .A2(n10011), .ZN(n10026) );
  AOI22_X1 U12623 ( .A1(n10014), .A2(keyinput93), .B1(keyinput73), .B2(n9529), 
        .ZN(n10013) );
  OAI221_X1 U12624 ( .B1(n10014), .B2(keyinput93), .C1(n9529), .C2(keyinput73), 
        .A(n10013), .ZN(n10018) );
  INV_X1 U12625 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n11723) );
  AOI22_X1 U12626 ( .A1(n10016), .A2(keyinput10), .B1(keyinput45), .B2(n11723), 
        .ZN(n10015) );
  OAI221_X1 U12627 ( .B1(n10016), .B2(keyinput10), .C1(n11723), .C2(keyinput45), .A(n10015), .ZN(n10017) );
  NOR2_X1 U12628 ( .A1(n10018), .A2(n10017), .ZN(n10025) );
  AOI22_X1 U12629 ( .A1(n10020), .A2(keyinput76), .B1(keyinput84), .B2(n15765), 
        .ZN(n10019) );
  OAI221_X1 U12630 ( .B1(n10020), .B2(keyinput76), .C1(n15765), .C2(keyinput84), .A(n10019), .ZN(n10023) );
  AOI22_X1 U12631 ( .A1(n12541), .A2(keyinput27), .B1(keyinput13), .B2(n15769), 
        .ZN(n10021) );
  OAI221_X1 U12632 ( .B1(n12541), .B2(keyinput27), .C1(n15769), .C2(keyinput13), .A(n10021), .ZN(n10022) );
  NOR2_X1 U12633 ( .A1(n10023), .A2(n10022), .ZN(n10024) );
  NAND4_X1 U12634 ( .A1(n10027), .A2(n10026), .A3(n10025), .A4(n10024), .ZN(
        n10064) );
  AOI22_X1 U12635 ( .A1(n9272), .A2(keyinput122), .B1(n15905), .B2(keyinput22), 
        .ZN(n10028) );
  OAI221_X1 U12636 ( .B1(n9272), .B2(keyinput122), .C1(n15905), .C2(keyinput22), .A(n10028), .ZN(n10035) );
  INV_X1 U12637 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n11740) );
  AOI22_X1 U12638 ( .A1(n10030), .A2(keyinput63), .B1(n11740), .B2(keyinput41), 
        .ZN(n10029) );
  OAI221_X1 U12639 ( .B1(n10030), .B2(keyinput63), .C1(n11740), .C2(keyinput41), .A(n10029), .ZN(n10034) );
  AOI22_X1 U12640 ( .A1(n10032), .A2(keyinput85), .B1(n10651), .B2(keyinput74), 
        .ZN(n10031) );
  OAI221_X1 U12641 ( .B1(n10032), .B2(keyinput85), .C1(n10651), .C2(keyinput74), .A(n10031), .ZN(n10033) );
  NOR3_X1 U12642 ( .A1(n10035), .A2(n10034), .A3(n10033), .ZN(n10062) );
  INV_X1 U12643 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15768) );
  AOI22_X1 U12644 ( .A1(n15768), .A2(keyinput1), .B1(n11812), .B2(keyinput72), 
        .ZN(n10036) );
  OAI221_X1 U12645 ( .B1(n15768), .B2(keyinput1), .C1(n11812), .C2(keyinput72), 
        .A(n10036), .ZN(n10053) );
  XNOR2_X1 U12646 ( .A(SI_2_), .B(keyinput26), .ZN(n10040) );
  XNOR2_X1 U12647 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput47), .ZN(n10039) );
  XNOR2_X1 U12648 ( .A(P2_IR_REG_9__SCAN_IN), .B(keyinput9), .ZN(n10038) );
  XNOR2_X1 U12649 ( .A(P3_REG0_REG_10__SCAN_IN), .B(keyinput4), .ZN(n10037) );
  AND4_X1 U12650 ( .A1(n10040), .A2(n10039), .A3(n10038), .A4(n10037), .ZN(
        n10046) );
  XNOR2_X1 U12651 ( .A(keyinput68), .B(n8226), .ZN(n10042) );
  XNOR2_X1 U12652 ( .A(keyinput115), .B(n7125), .ZN(n10041) );
  NOR2_X1 U12653 ( .A1(n10042), .A2(n10041), .ZN(n10045) );
  XNOR2_X1 U12654 ( .A(P3_IR_REG_28__SCAN_IN), .B(keyinput0), .ZN(n10044) );
  XNOR2_X1 U12655 ( .A(P3_IR_REG_17__SCAN_IN), .B(keyinput8), .ZN(n10043) );
  NAND4_X1 U12656 ( .A1(n10046), .A2(n10045), .A3(n10044), .A4(n10043), .ZN(
        n10052) );
  XNOR2_X1 U12657 ( .A(keyinput89), .B(P2_REG0_REG_6__SCAN_IN), .ZN(n10050) );
  XNOR2_X1 U12658 ( .A(keyinput67), .B(P2_REG0_REG_4__SCAN_IN), .ZN(n10049) );
  XNOR2_X1 U12659 ( .A(keyinput98), .B(P3_DATAO_REG_12__SCAN_IN), .ZN(n10048)
         );
  XNOR2_X1 U12660 ( .A(keyinput52), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n10047) );
  NAND4_X1 U12661 ( .A1(n10050), .A2(n10049), .A3(n10048), .A4(n10047), .ZN(
        n10051) );
  NOR3_X1 U12662 ( .A1(n10053), .A2(n10052), .A3(n10051), .ZN(n10061) );
  INV_X1 U12663 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n10055) );
  AOI22_X1 U12664 ( .A1(n15903), .A2(keyinput16), .B1(keyinput103), .B2(n10055), .ZN(n10054) );
  OAI221_X1 U12665 ( .B1(n15903), .B2(keyinput16), .C1(n10055), .C2(
        keyinput103), .A(n10054), .ZN(n10059) );
  INV_X1 U12666 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n15766) );
  INV_X1 U12667 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10057) );
  AOI22_X1 U12668 ( .A1(n15766), .A2(keyinput96), .B1(n10057), .B2(keyinput2), 
        .ZN(n10056) );
  OAI221_X1 U12669 ( .B1(n15766), .B2(keyinput96), .C1(n10057), .C2(keyinput2), 
        .A(n10056), .ZN(n10058) );
  NOR2_X1 U12670 ( .A1(n10059), .A2(n10058), .ZN(n10060) );
  NAND3_X1 U12671 ( .A1(n10062), .A2(n10061), .A3(n10060), .ZN(n10063) );
  OR2_X1 U12672 ( .A1(n10064), .A2(n10063), .ZN(n10121) );
  INV_X1 U12673 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n10764) );
  INV_X1 U12674 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15614) );
  AOI22_X1 U12675 ( .A1(n10764), .A2(keyinput53), .B1(keyinput60), .B2(n15614), 
        .ZN(n10065) );
  OAI221_X1 U12676 ( .B1(n10764), .B2(keyinput53), .C1(n15614), .C2(keyinput60), .A(n10065), .ZN(n10072) );
  XNOR2_X1 U12677 ( .A(SI_1_), .B(keyinput36), .ZN(n10070) );
  XNOR2_X1 U12678 ( .A(keyinput11), .B(P2_D_REG_5__SCAN_IN), .ZN(n10069) );
  NAND2_X1 U12679 ( .A1(keyinput125), .A2(n15020), .ZN(n10068) );
  NAND2_X1 U12680 ( .A1(n10066), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n10067) );
  NAND4_X1 U12681 ( .A1(n10070), .A2(n10069), .A3(n10068), .A4(n10067), .ZN(
        n10071) );
  NOR2_X1 U12682 ( .A1(n10072), .A2(n10071), .ZN(n10106) );
  XNOR2_X1 U12683 ( .A(SI_16_), .B(keyinput101), .ZN(n10076) );
  XNOR2_X1 U12684 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(keyinput28), .ZN(n10075) );
  XNOR2_X1 U12685 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput86), .ZN(n10074) );
  XNOR2_X1 U12686 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput80), .ZN(n10073) );
  NAND4_X1 U12687 ( .A1(n10076), .A2(n10075), .A3(n10074), .A4(n10073), .ZN(
        n10082) );
  XNOR2_X1 U12688 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput99), .ZN(n10080)
         );
  XNOR2_X1 U12689 ( .A(P2_REG1_REG_23__SCAN_IN), .B(keyinput44), .ZN(n10079)
         );
  XNOR2_X1 U12690 ( .A(P2_REG0_REG_12__SCAN_IN), .B(keyinput116), .ZN(n10078)
         );
  XNOR2_X1 U12691 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput105), .ZN(n10077)
         );
  NAND4_X1 U12692 ( .A1(n10080), .A2(n10079), .A3(n10078), .A4(n10077), .ZN(
        n10081) );
  NOR2_X1 U12693 ( .A1(n10082), .A2(n10081), .ZN(n10105) );
  XNOR2_X1 U12694 ( .A(P2_REG3_REG_24__SCAN_IN), .B(keyinput91), .ZN(n10086)
         );
  XNOR2_X1 U12695 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput31), .ZN(n10085)
         );
  XNOR2_X1 U12696 ( .A(P3_IR_REG_9__SCAN_IN), .B(keyinput69), .ZN(n10084) );
  XNOR2_X1 U12697 ( .A(P3_IR_REG_6__SCAN_IN), .B(keyinput54), .ZN(n10083) );
  NAND4_X1 U12698 ( .A1(n10086), .A2(n10085), .A3(n10084), .A4(n10083), .ZN(
        n10092) );
  XNOR2_X1 U12699 ( .A(P3_REG0_REG_29__SCAN_IN), .B(keyinput37), .ZN(n10090)
         );
  XNOR2_X1 U12700 ( .A(P3_IR_REG_21__SCAN_IN), .B(keyinput102), .ZN(n10089) );
  XNOR2_X1 U12701 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput121), .ZN(n10088) );
  XNOR2_X1 U12702 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput127), .ZN(n10087) );
  NAND4_X1 U12703 ( .A1(n10090), .A2(n10089), .A3(n10088), .A4(n10087), .ZN(
        n10091) );
  NOR2_X1 U12704 ( .A1(n10092), .A2(n10091), .ZN(n10104) );
  XNOR2_X1 U12705 ( .A(SI_10_), .B(keyinput107), .ZN(n10096) );
  XNOR2_X1 U12706 ( .A(SI_12_), .B(keyinput111), .ZN(n10095) );
  XNOR2_X1 U12707 ( .A(P3_REG3_REG_3__SCAN_IN), .B(keyinput78), .ZN(n10094) );
  XNOR2_X1 U12708 ( .A(P3_IR_REG_16__SCAN_IN), .B(keyinput83), .ZN(n10093) );
  NAND4_X1 U12709 ( .A1(n10096), .A2(n10095), .A3(n10094), .A4(n10093), .ZN(
        n10102) );
  XNOR2_X1 U12710 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput71), .ZN(n10100) );
  XNOR2_X1 U12711 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput77), .ZN(n10099) );
  XNOR2_X1 U12712 ( .A(SI_6_), .B(keyinput51), .ZN(n10098) );
  XNOR2_X1 U12713 ( .A(P1_REG0_REG_17__SCAN_IN), .B(keyinput65), .ZN(n10097)
         );
  NAND4_X1 U12714 ( .A1(n10100), .A2(n10099), .A3(n10098), .A4(n10097), .ZN(
        n10101) );
  NOR2_X1 U12715 ( .A1(n10102), .A2(n10101), .ZN(n10103) );
  AND4_X1 U12716 ( .A1(n10106), .A2(n10105), .A3(n10104), .A4(n10103), .ZN(
        n10119) );
  AOI22_X1 U12717 ( .A1(n7127), .A2(keyinput79), .B1(keyinput48), .B2(n10108), 
        .ZN(n10107) );
  OAI221_X1 U12718 ( .B1(n7127), .B2(keyinput79), .C1(n10108), .C2(keyinput48), 
        .A(n10107), .ZN(n10112) );
  AOI22_X1 U12719 ( .A1(n14583), .A2(keyinput57), .B1(keyinput12), .B2(n14945), 
        .ZN(n10109) );
  OAI221_X1 U12720 ( .B1(n14583), .B2(keyinput57), .C1(n14945), .C2(keyinput12), .A(n10109), .ZN(n10111) );
  INV_X1 U12721 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10612) );
  XNOR2_X1 U12722 ( .A(n10612), .B(keyinput25), .ZN(n10110) );
  NOR3_X1 U12723 ( .A1(n10112), .A2(n10111), .A3(n10110), .ZN(n10118) );
  INV_X1 U12724 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10682) );
  AOI22_X1 U12725 ( .A1(n13898), .A2(keyinput39), .B1(keyinput119), .B2(n10682), .ZN(n10113) );
  OAI221_X1 U12726 ( .B1(n13898), .B2(keyinput39), .C1(n10682), .C2(
        keyinput119), .A(n10113), .ZN(n10116) );
  AOI22_X1 U12727 ( .A1(n11029), .A2(keyinput123), .B1(keyinput94), .B2(n15840), .ZN(n10114) );
  OAI221_X1 U12728 ( .B1(n11029), .B2(keyinput123), .C1(n15840), .C2(
        keyinput94), .A(n10114), .ZN(n10115) );
  NOR2_X1 U12729 ( .A1(n10116), .A2(n10115), .ZN(n10117) );
  NAND3_X1 U12730 ( .A1(n10119), .A2(n10118), .A3(n10117), .ZN(n10120) );
  NOR2_X1 U12731 ( .A1(n10121), .A2(n10120), .ZN(n10145) );
  INV_X1 U12732 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n10324) );
  AOI22_X1 U12733 ( .A1(n10123), .A2(keyinput21), .B1(keyinput58), .B2(n10324), 
        .ZN(n10122) );
  OAI221_X1 U12734 ( .B1(n10123), .B2(keyinput21), .C1(n10324), .C2(keyinput58), .A(n10122), .ZN(n10133) );
  INV_X1 U12735 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n10126) );
  INV_X1 U12736 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n10125) );
  AOI22_X1 U12737 ( .A1(n10126), .A2(keyinput75), .B1(n10125), .B2(keyinput42), 
        .ZN(n10124) );
  OAI221_X1 U12738 ( .B1(n10126), .B2(keyinput75), .C1(n10125), .C2(keyinput42), .A(n10124), .ZN(n10132) );
  AOI22_X1 U12739 ( .A1(n15767), .A2(keyinput112), .B1(keyinput46), .B2(n12017), .ZN(n10127) );
  OAI221_X1 U12740 ( .B1(n15767), .B2(keyinput112), .C1(n12017), .C2(
        keyinput46), .A(n10127), .ZN(n10131) );
  INV_X1 U12741 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n10129) );
  AOI22_X1 U12742 ( .A1(n10129), .A2(keyinput34), .B1(n14801), .B2(keyinput87), 
        .ZN(n10128) );
  OAI221_X1 U12743 ( .B1(n10129), .B2(keyinput34), .C1(n14801), .C2(keyinput87), .A(n10128), .ZN(n10130) );
  NOR4_X1 U12744 ( .A1(n10133), .A2(n10132), .A3(n10131), .A4(n10130), .ZN(
        n10144) );
  AOI22_X1 U12745 ( .A1(n8145), .A2(keyinput30), .B1(keyinput95), .B2(n10135), 
        .ZN(n10134) );
  OAI221_X1 U12746 ( .B1(n8145), .B2(keyinput30), .C1(n10135), .C2(keyinput95), 
        .A(n10134), .ZN(n10142) );
  AOI22_X1 U12747 ( .A1(n12479), .A2(keyinput17), .B1(keyinput100), .B2(n7530), 
        .ZN(n10136) );
  OAI221_X1 U12748 ( .B1(n12479), .B2(keyinput17), .C1(n7530), .C2(keyinput100), .A(n10136), .ZN(n10141) );
  INV_X1 U12749 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n10332) );
  AOI22_X1 U12750 ( .A1(n13889), .A2(keyinput120), .B1(keyinput82), .B2(n10332), .ZN(n10137) );
  OAI221_X1 U12751 ( .B1(n13889), .B2(keyinput120), .C1(n10332), .C2(
        keyinput82), .A(n10137), .ZN(n10140) );
  AOI22_X1 U12752 ( .A1(n15287), .A2(keyinput3), .B1(n10967), .B2(keyinput59), 
        .ZN(n10138) );
  OAI221_X1 U12753 ( .B1(n15287), .B2(keyinput3), .C1(n10967), .C2(keyinput59), 
        .A(n10138), .ZN(n10139) );
  NOR4_X1 U12754 ( .A1(n10142), .A2(n10141), .A3(n10140), .A4(n10139), .ZN(
        n10143) );
  NAND3_X1 U12755 ( .A1(n10145), .A2(n10144), .A3(n10143), .ZN(n10146) );
  AOI211_X1 U12756 ( .C1(n10148), .C2(P1_REG3_REG_1__SCAN_IN), .A(n10147), .B(
        n10146), .ZN(n10149) );
  INV_X1 U12757 ( .A(n10153), .ZN(n10151) );
  INV_X1 U12758 ( .A(n10152), .ZN(n10150) );
  NAND2_X1 U12759 ( .A1(n10151), .A2(n10150), .ZN(n10154) );
  NAND2_X1 U12760 ( .A1(n10153), .A2(n10152), .ZN(n10155) );
  NAND2_X1 U12761 ( .A1(n10157), .A2(n10156), .ZN(n10159) );
  NAND2_X1 U12762 ( .A1(n6641), .A2(n10159), .ZN(n13288) );
  INV_X1 U12763 ( .A(n12898), .ZN(n13941) );
  AOI22_X1 U12764 ( .A1(n13696), .A2(n13443), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10160) );
  OAI21_X1 U12765 ( .B1(n13693), .B2(n13428), .A(n10160), .ZN(n10161) );
  AOI21_X1 U12766 ( .B1(n13430), .B2(n13665), .A(n10161), .ZN(n10162) );
  OAI21_X1 U12767 ( .B1(n13941), .B2(n13446), .A(n10162), .ZN(n10163) );
  NAND2_X1 U12768 ( .A1(n10165), .A2(n10164), .ZN(P3_U3169) );
  NAND2_X1 U12769 ( .A1(n10240), .A2(n10414), .ZN(n10167) );
  NAND2_X1 U12770 ( .A1(n6685), .A2(n10167), .ZN(n10169) );
  NAND2_X1 U12771 ( .A1(n10168), .A2(n10414), .ZN(n13266) );
  NAND2_X1 U12772 ( .A1(n13266), .A2(n11861), .ZN(n10170) );
  NAND2_X1 U12773 ( .A1(n10169), .A2(n10170), .ZN(n10173) );
  INV_X1 U12774 ( .A(n10170), .ZN(n10171) );
  NAND3_X1 U12775 ( .A1(n10171), .A2(n11860), .A3(n9433), .ZN(n10172) );
  NAND2_X1 U12776 ( .A1(n10194), .A2(n14216), .ZN(n10182) );
  NAND2_X1 U12777 ( .A1(n10340), .A2(n12099), .ZN(n10181) );
  AND2_X1 U12778 ( .A1(n10182), .A2(n10181), .ZN(n10176) );
  NAND2_X1 U12779 ( .A1(n10240), .A2(n14216), .ZN(n10174) );
  OAI21_X1 U12780 ( .B1(n10232), .B2(n12688), .A(n10174), .ZN(n10175) );
  NAND2_X1 U12781 ( .A1(n10340), .A2(n14215), .ZN(n10177) );
  NAND2_X1 U12782 ( .A1(n10178), .A2(n10177), .ZN(n10187) );
  OR2_X1 U12783 ( .A1(n10240), .A2(n12085), .ZN(n10180) );
  NAND2_X1 U12784 ( .A1(n10340), .A2(n12114), .ZN(n10179) );
  NAND2_X1 U12785 ( .A1(n10183), .A2(n10176), .ZN(n10184) );
  NAND3_X1 U12786 ( .A1(n10186), .A2(n10185), .A3(n10184), .ZN(n10191) );
  INV_X1 U12787 ( .A(n10187), .ZN(n10189) );
  NAND2_X1 U12788 ( .A1(n10189), .A2(n10188), .ZN(n10190) );
  NAND2_X1 U12789 ( .A1(n10191), .A2(n10190), .ZN(n10196) );
  OR2_X1 U12790 ( .A1(n10232), .A2(n12104), .ZN(n10193) );
  OR2_X1 U12791 ( .A1(n10232), .A2(n15924), .ZN(n10198) );
  NAND2_X1 U12792 ( .A1(n10232), .A2(n14213), .ZN(n10197) );
  NAND2_X1 U12793 ( .A1(n10198), .A2(n10197), .ZN(n10200) );
  AOI22_X1 U12794 ( .A1(n10339), .A2(n14213), .B1(n14107), .B2(n10340), .ZN(
        n10199) );
  OR2_X1 U12795 ( .A1(n10232), .A2(n14104), .ZN(n10201) );
  NAND2_X1 U12796 ( .A1(n10232), .A2(n14212), .ZN(n10202) );
  OAI21_X1 U12797 ( .B1(n10232), .B2(n12412), .A(n10202), .ZN(n10203) );
  OR2_X1 U12798 ( .A1(n10240), .A2(n15932), .ZN(n10205) );
  NAND2_X1 U12799 ( .A1(n10232), .A2(n14211), .ZN(n10204) );
  AOI22_X1 U12800 ( .A1(n10194), .A2(n14211), .B1(n12350), .B2(n10340), .ZN(
        n10206) );
  OAI22_X1 U12801 ( .A1(n12398), .A2(n10339), .B1(n10232), .B2(n12548), .ZN(
        n10209) );
  AOI22_X1 U12802 ( .A1(n10345), .A2(n12342), .B1(n14210), .B2(n10232), .ZN(
        n10207) );
  AOI22_X1 U12803 ( .A1(n12331), .A2(n10345), .B1(n14209), .B2(n10340), .ZN(
        n10211) );
  OAI22_X1 U12804 ( .A1(n12554), .A2(n10339), .B1(n12471), .B2(n10240), .ZN(
        n10210) );
  OAI22_X1 U12805 ( .A1(n12366), .A2(n10339), .B1(n12329), .B2(n10232), .ZN(
        n10214) );
  AOI22_X1 U12806 ( .A1(n12242), .A2(n10345), .B1(n14207), .B2(n10232), .ZN(
        n10216) );
  INV_X1 U12807 ( .A(n14207), .ZN(n10461) );
  OAI22_X1 U12808 ( .A1(n9865), .A2(n10339), .B1(n10461), .B2(n10240), .ZN(
        n10215) );
  OAI22_X1 U12809 ( .A1(n14823), .A2(n10339), .B1(n14066), .B2(n10232), .ZN(
        n10219) );
  OAI22_X1 U12810 ( .A1(n14823), .A2(n10340), .B1(n14066), .B2(n10339), .ZN(
        n10220) );
  AOI22_X1 U12811 ( .A1(n14769), .A2(n10345), .B1(n14206), .B2(n10232), .ZN(
        n10223) );
  AOI22_X1 U12812 ( .A1(n14769), .A2(n10232), .B1(n10345), .B2(n14206), .ZN(
        n10221) );
  INV_X1 U12813 ( .A(n10221), .ZN(n10222) );
  OAI22_X1 U12814 ( .A1(n14816), .A2(n10339), .B1(n14205), .B2(n10232), .ZN(
        n10226) );
  OAI22_X1 U12815 ( .A1(n14816), .A2(n10240), .B1(n14205), .B2(n10339), .ZN(
        n10225) );
  INV_X1 U12816 ( .A(n10226), .ZN(n10227) );
  OAI22_X1 U12817 ( .A1(n14620), .A2(n10340), .B1(n14637), .B2(n10345), .ZN(
        n10228) );
  OAI22_X1 U12818 ( .A1(n14620), .A2(n10339), .B1(n14637), .B2(n10232), .ZN(
        n10229) );
  OAI22_X1 U12819 ( .A1(n14605), .A2(n10339), .B1(n14089), .B2(n10240), .ZN(
        n10230) );
  OAI22_X1 U12820 ( .A1(n14605), .A2(n10340), .B1(n14089), .B2(n10339), .ZN(
        n10231) );
  AOI22_X1 U12821 ( .A1(n14580), .A2(n10345), .B1(n14203), .B2(n10232), .ZN(
        n10234) );
  OAI22_X1 U12822 ( .A1(n7627), .A2(n10339), .B1(n14594), .B2(n10232), .ZN(
        n10233) );
  NAND2_X1 U12823 ( .A1(n10235), .A2(n10234), .ZN(n10236) );
  AOI22_X1 U12824 ( .A1(n14566), .A2(n10240), .B1(n10345), .B2(n14575), .ZN(
        n10237) );
  AOI22_X1 U12825 ( .A1(n14566), .A2(n10339), .B1(n14575), .B2(n10340), .ZN(
        n10238) );
  INV_X1 U12826 ( .A(n14563), .ZN(n14202) );
  AOI22_X1 U12827 ( .A1(n14737), .A2(n10232), .B1(n10345), .B2(n14202), .ZN(
        n10270) );
  OAI22_X1 U12828 ( .A1(n14552), .A2(n10240), .B1(n14563), .B2(n10339), .ZN(
        n10269) );
  AND2_X1 U12829 ( .A1(n14484), .A2(n10339), .ZN(n10241) );
  AOI21_X1 U12830 ( .B1(n14515), .B2(n10232), .A(n10241), .ZN(n10308) );
  NAND2_X1 U12831 ( .A1(n14515), .A2(n10339), .ZN(n10243) );
  NAND2_X1 U12832 ( .A1(n14484), .A2(n10232), .ZN(n10242) );
  NAND2_X1 U12833 ( .A1(n10243), .A2(n10242), .ZN(n10307) );
  AND2_X1 U12834 ( .A1(n14196), .A2(n10339), .ZN(n10244) );
  AOI21_X1 U12835 ( .B1(n14695), .B2(n10232), .A(n10244), .ZN(n10289) );
  NAND2_X1 U12836 ( .A1(n14196), .A2(n10232), .ZN(n10245) );
  NAND2_X1 U12837 ( .A1(n10246), .A2(n10245), .ZN(n10288) );
  AND2_X1 U12838 ( .A1(n14197), .A2(n10345), .ZN(n10247) );
  AOI21_X1 U12839 ( .B1(n14700), .B2(n10232), .A(n10247), .ZN(n10285) );
  NAND2_X1 U12840 ( .A1(n14700), .A2(n10339), .ZN(n10249) );
  NAND2_X1 U12841 ( .A1(n14197), .A2(n10232), .ZN(n10248) );
  NAND2_X1 U12842 ( .A1(n10249), .A2(n10248), .ZN(n10284) );
  NAND2_X1 U12843 ( .A1(n10285), .A2(n10284), .ZN(n10250) );
  AND2_X1 U12844 ( .A1(n14198), .A2(n10345), .ZN(n10251) );
  AOI21_X1 U12845 ( .B1(n14705), .B2(n10232), .A(n10251), .ZN(n10276) );
  NAND2_X1 U12846 ( .A1(n14705), .A2(n10339), .ZN(n10253) );
  NAND2_X1 U12847 ( .A1(n14198), .A2(n10232), .ZN(n10252) );
  NAND2_X1 U12848 ( .A1(n10253), .A2(n10252), .ZN(n10275) );
  AND2_X1 U12849 ( .A1(n14199), .A2(n10345), .ZN(n10254) );
  AOI21_X1 U12850 ( .B1(n14710), .B2(n10232), .A(n10254), .ZN(n10280) );
  NAND2_X1 U12851 ( .A1(n14710), .A2(n10345), .ZN(n10256) );
  NAND2_X1 U12852 ( .A1(n14199), .A2(n10232), .ZN(n10255) );
  NAND2_X1 U12853 ( .A1(n10256), .A2(n10255), .ZN(n10279) );
  NAND2_X1 U12854 ( .A1(n10280), .A2(n10279), .ZN(n10257) );
  INV_X1 U12855 ( .A(n10300), .ZN(n10262) );
  AND2_X1 U12856 ( .A1(n14485), .A2(n10345), .ZN(n10258) );
  AOI21_X1 U12857 ( .B1(n12751), .B2(n10232), .A(n10258), .ZN(n10299) );
  NAND2_X1 U12858 ( .A1(n12751), .A2(n10339), .ZN(n10260) );
  NAND2_X1 U12859 ( .A1(n14485), .A2(n10232), .ZN(n10259) );
  NAND2_X1 U12860 ( .A1(n10260), .A2(n10259), .ZN(n10298) );
  NAND2_X1 U12861 ( .A1(n10299), .A2(n10298), .ZN(n10261) );
  AND2_X1 U12862 ( .A1(n14200), .A2(n10339), .ZN(n10263) );
  AOI21_X1 U12863 ( .B1(n14491), .B2(n10232), .A(n10263), .ZN(n10313) );
  NAND2_X1 U12864 ( .A1(n14491), .A2(n10345), .ZN(n10265) );
  NAND2_X1 U12865 ( .A1(n14200), .A2(n10232), .ZN(n10264) );
  NAND2_X1 U12866 ( .A1(n10265), .A2(n10264), .ZN(n10312) );
  AND2_X1 U12867 ( .A1(n14201), .A2(n10240), .ZN(n10266) );
  AOI21_X1 U12868 ( .B1(n14732), .B2(n10345), .A(n10266), .ZN(n10304) );
  NAND2_X1 U12869 ( .A1(n14732), .A2(n10232), .ZN(n10268) );
  NAND2_X1 U12870 ( .A1(n14201), .A2(n10339), .ZN(n10267) );
  NAND2_X1 U12871 ( .A1(n10268), .A2(n10267), .ZN(n10303) );
  OAI22_X1 U12872 ( .A1(n10304), .A2(n10303), .B1(n7466), .B2(n7467), .ZN(
        n10271) );
  AND2_X1 U12873 ( .A1(n14195), .A2(n10240), .ZN(n10272) );
  AOI21_X1 U12874 ( .B1(n14690), .B2(n10345), .A(n10272), .ZN(n10349) );
  NAND2_X1 U12875 ( .A1(n14690), .A2(n10340), .ZN(n10274) );
  NAND2_X1 U12876 ( .A1(n14195), .A2(n10339), .ZN(n10273) );
  NAND2_X1 U12877 ( .A1(n10274), .A2(n10273), .ZN(n10348) );
  INV_X1 U12878 ( .A(n10275), .ZN(n10278) );
  INV_X1 U12879 ( .A(n10276), .ZN(n10277) );
  NAND2_X1 U12880 ( .A1(n10278), .A2(n10277), .ZN(n10296) );
  INV_X1 U12881 ( .A(n10279), .ZN(n10282) );
  INV_X1 U12882 ( .A(n10280), .ZN(n10281) );
  NAND3_X1 U12883 ( .A1(n10283), .A2(n10282), .A3(n10281), .ZN(n10295) );
  INV_X1 U12884 ( .A(n10284), .ZN(n10287) );
  INV_X1 U12885 ( .A(n10285), .ZN(n10286) );
  AND2_X1 U12886 ( .A1(n10287), .A2(n10286), .ZN(n10292) );
  INV_X1 U12887 ( .A(n10288), .ZN(n10291) );
  INV_X1 U12888 ( .A(n10289), .ZN(n10290) );
  AOI22_X1 U12889 ( .A1(n10293), .A2(n10292), .B1(n10291), .B2(n10290), .ZN(
        n10294) );
  OAI211_X1 U12890 ( .C1(n10297), .C2(n10296), .A(n10295), .B(n10294), .ZN(
        n10302) );
  NOR3_X1 U12891 ( .A1(n10300), .A2(n10299), .A3(n10298), .ZN(n10301) );
  AOI211_X1 U12892 ( .C1(n10349), .C2(n10348), .A(n10302), .B(n10301), .ZN(
        n10319) );
  NAND3_X1 U12893 ( .A1(n10305), .A2(n10304), .A3(n10303), .ZN(n10318) );
  INV_X1 U12894 ( .A(n10306), .ZN(n10311) );
  INV_X1 U12895 ( .A(n10307), .ZN(n10310) );
  INV_X1 U12896 ( .A(n10308), .ZN(n10309) );
  NAND3_X1 U12897 ( .A1(n10311), .A2(n10310), .A3(n10309), .ZN(n10317) );
  INV_X1 U12898 ( .A(n10312), .ZN(n10315) );
  INV_X1 U12899 ( .A(n10313), .ZN(n10314) );
  NAND3_X1 U12900 ( .A1(n6591), .A2(n10315), .A3(n10314), .ZN(n10316) );
  NAND2_X1 U12901 ( .A1(n10336), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n10320) );
  NAND2_X1 U12902 ( .A1(n10329), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n10323) );
  NAND2_X1 U12903 ( .A1(n10321), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n10322) );
  OAI211_X1 U12904 ( .C1(n10325), .C2(n10324), .A(n10323), .B(n10322), .ZN(
        n14193) );
  AOI22_X1 U12905 ( .A1(n10367), .A2(n10340), .B1(n10339), .B2(n14193), .ZN(
        n10342) );
  NAND2_X1 U12906 ( .A1(n10336), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n10326) );
  NAND2_X1 U12907 ( .A1(n10328), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n10331) );
  NAND2_X1 U12908 ( .A1(n10329), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n10330) );
  OAI211_X1 U12909 ( .C1(n6793), .C2(n10332), .A(n10331), .B(n10330), .ZN(
        n14351) );
  NAND2_X1 U12910 ( .A1(n10240), .A2(n14193), .ZN(n10369) );
  NAND2_X1 U12911 ( .A1(n10333), .A2(n11866), .ZN(n10373) );
  NAND4_X1 U12912 ( .A1(n10369), .A2(n10375), .A3(n10373), .A4(n10405), .ZN(
        n10334) );
  AOI22_X1 U12913 ( .A1(n14681), .A2(n10345), .B1(n14351), .B2(n10334), .ZN(
        n10363) );
  INV_X1 U12914 ( .A(n10363), .ZN(n10341) );
  AOI22_X1 U12915 ( .A1(n14681), .A2(n10232), .B1(n10345), .B2(n14351), .ZN(
        n10362) );
  NAND2_X1 U12916 ( .A1(n14825), .A2(n10335), .ZN(n10338) );
  NAND2_X1 U12917 ( .A1(n10336), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n10337) );
  INV_X1 U12918 ( .A(n10379), .ZN(n14194) );
  AOI22_X1 U12919 ( .A1(n10380), .A2(n10240), .B1(n10345), .B2(n14194), .ZN(
        n10358) );
  OAI22_X1 U12920 ( .A1(n14686), .A2(n10340), .B1(n10379), .B2(n10339), .ZN(
        n10359) );
  INV_X1 U12921 ( .A(n10343), .ZN(n10360) );
  AND2_X1 U12922 ( .A1(n14355), .A2(n10240), .ZN(n10344) );
  AOI21_X1 U12923 ( .B1(n14369), .B2(n10345), .A(n10344), .ZN(n10355) );
  NAND2_X1 U12924 ( .A1(n14369), .A2(n10240), .ZN(n10347) );
  NAND2_X1 U12925 ( .A1(n14355), .A2(n10339), .ZN(n10346) );
  NAND2_X1 U12926 ( .A1(n10347), .A2(n10346), .ZN(n10354) );
  OAI22_X1 U12927 ( .A1(n10355), .A2(n10354), .B1(n10349), .B2(n10348), .ZN(
        n10350) );
  INV_X1 U12928 ( .A(n10350), .ZN(n10351) );
  NAND2_X1 U12929 ( .A1(n10352), .A2(n7991), .ZN(n10366) );
  INV_X1 U12930 ( .A(n10354), .ZN(n10357) );
  INV_X1 U12931 ( .A(n10355), .ZN(n10356) );
  OAI22_X1 U12932 ( .A1(n10359), .A2(n10358), .B1(n10357), .B2(n10356), .ZN(
        n10361) );
  INV_X1 U12933 ( .A(n10362), .ZN(n10364) );
  OAI211_X1 U12934 ( .C1(n14788), .C2(n10240), .A(n10369), .B(n10368), .ZN(
        n10370) );
  AOI211_X1 U12935 ( .C1(n10375), .C2(n14332), .A(n10485), .B(n10371), .ZN(
        n10372) );
  NOR2_X1 U12936 ( .A1(n9853), .A2(n14332), .ZN(n10376) );
  INV_X1 U12937 ( .A(n10373), .ZN(n10374) );
  AOI21_X1 U12938 ( .B1(n10376), .B2(n10375), .A(n10374), .ZN(n10377) );
  XNOR2_X1 U12939 ( .A(n14515), .B(n14057), .ZN(n14508) );
  AND2_X1 U12940 ( .A1(n10381), .A2(n13266), .ZN(n14784) );
  NAND2_X1 U12941 ( .A1(n10383), .A2(n12091), .ZN(n10384) );
  NOR3_X1 U12942 ( .A1(n10385), .A2(n11971), .A3(n10384), .ZN(n10387) );
  XNOR2_X1 U12943 ( .A(n12342), .B(n14210), .ZN(n12125) );
  NAND2_X1 U12944 ( .A1(n10390), .A2(n10389), .ZN(n14668) );
  NOR4_X1 U12945 ( .A1(n14470), .A2(n14508), .A3(n14503), .A4(n10393), .ZN(
        n10394) );
  XNOR2_X1 U12946 ( .A(n14491), .B(n14200), .ZN(n14488) );
  NAND4_X1 U12947 ( .A1(n10394), .A2(n14446), .A3(n14522), .A4(n14488), .ZN(
        n10395) );
  NOR4_X1 U12948 ( .A1(n14403), .A2(n14417), .A3(n14428), .A4(n10395), .ZN(
        n10397) );
  NAND2_X1 U12949 ( .A1(n10404), .A2(n6782), .ZN(n10409) );
  INV_X1 U12950 ( .A(P2_B_REG_SCAN_IN), .ZN(n12902) );
  INV_X1 U12951 ( .A(n15914), .ZN(n15911) );
  AOI211_X1 U12952 ( .C1(n6782), .C2(n9433), .A(n12902), .B(n10406), .ZN(
        n10407) );
  NAND2_X1 U12953 ( .A1(n10409), .A2(n10408), .ZN(P2_U3328) );
  INV_X1 U12954 ( .A(n10532), .ZN(n10619) );
  NOR2_X2 U12955 ( .A1(n10957), .A2(n10619), .ZN(P1_U4016) );
  NAND2_X1 U12956 ( .A1(n11020), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10410) );
  OR2_X2 U12957 ( .A1(n11021), .A2(n10410), .ZN(n14217) );
  INV_X1 U12958 ( .A(n14217), .ZN(P2_U3947) );
  NOR2_X1 U12959 ( .A1(n10411), .A2(n10584), .ZN(P3_U3897) );
  INV_X1 U12960 ( .A(n11861), .ZN(n10412) );
  XNOR2_X1 U12961 ( .A(n10419), .B(n10417), .ZN(n11680) );
  NAND2_X1 U12962 ( .A1(n10413), .A2(n10414), .ZN(n10416) );
  NAND2_X1 U12963 ( .A1(n10415), .A2(n13267), .ZN(n13269) );
  INV_X1 U12964 ( .A(n10417), .ZN(n10418) );
  NAND2_X1 U12965 ( .A1(n10419), .A2(n10418), .ZN(n10420) );
  XNOR2_X1 U12966 ( .A(n10413), .B(n15917), .ZN(n10424) );
  NOR2_X1 U12967 ( .A1(n10450), .A2(n12085), .ZN(n10422) );
  XNOR2_X1 U12968 ( .A(n10424), .B(n10422), .ZN(n11687) );
  NAND2_X1 U12969 ( .A1(n11688), .A2(n11687), .ZN(n10426) );
  INV_X1 U12970 ( .A(n10422), .ZN(n10423) );
  NAND2_X1 U12971 ( .A1(n10424), .A2(n10423), .ZN(n10425) );
  NOR2_X1 U12972 ( .A1(n10450), .A2(n12104), .ZN(n10428) );
  NAND2_X1 U12973 ( .A1(n10427), .A2(n10428), .ZN(n10431) );
  INV_X1 U12974 ( .A(n10427), .ZN(n14112) );
  INV_X1 U12975 ( .A(n10428), .ZN(n10429) );
  NAND2_X1 U12976 ( .A1(n14112), .A2(n10429), .ZN(n10430) );
  NAND2_X1 U12977 ( .A1(n10431), .A2(n10430), .ZN(n11675) );
  XNOR2_X1 U12978 ( .A(n10413), .B(n15924), .ZN(n12047) );
  NOR2_X1 U12979 ( .A1(n10450), .A2(n12179), .ZN(n10432) );
  XNOR2_X1 U12980 ( .A(n12047), .B(n10432), .ZN(n14111) );
  INV_X1 U12981 ( .A(n10432), .ZN(n10433) );
  NAND2_X1 U12982 ( .A1(n12047), .A2(n10433), .ZN(n10434) );
  XNOR2_X1 U12983 ( .A(n10413), .B(n12412), .ZN(n10437) );
  NOR2_X1 U12984 ( .A1(n10450), .A2(n14104), .ZN(n10435) );
  XNOR2_X1 U12985 ( .A(n10437), .B(n10435), .ZN(n12049) );
  INV_X1 U12986 ( .A(n10435), .ZN(n10436) );
  NAND2_X1 U12987 ( .A1(n10437), .A2(n10436), .ZN(n10438) );
  XNOR2_X1 U12988 ( .A(n10413), .B(n12350), .ZN(n10439) );
  NOR2_X1 U12989 ( .A1(n10450), .A2(n12336), .ZN(n10440) );
  NAND2_X1 U12990 ( .A1(n10439), .A2(n10440), .ZN(n10444) );
  INV_X1 U12991 ( .A(n10439), .ZN(n12335) );
  INV_X1 U12992 ( .A(n10440), .ZN(n10441) );
  NAND2_X1 U12993 ( .A1(n12335), .A2(n10441), .ZN(n10442) );
  NAND2_X1 U12994 ( .A1(n10444), .A2(n10442), .ZN(n12349) );
  XNOR2_X1 U12995 ( .A(n10413), .B(n12342), .ZN(n10445) );
  NOR2_X1 U12996 ( .A1(n10450), .A2(n12548), .ZN(n10446) );
  NAND2_X1 U12997 ( .A1(n10445), .A2(n10446), .ZN(n10451) );
  INV_X1 U12998 ( .A(n10445), .ZN(n12547) );
  INV_X1 U12999 ( .A(n10446), .ZN(n10447) );
  NAND2_X1 U13000 ( .A1(n12547), .A2(n10447), .ZN(n10448) );
  XNOR2_X1 U13001 ( .A(n10413), .B(n12331), .ZN(n10453) );
  OR2_X1 U13002 ( .A1(n10450), .A2(n12471), .ZN(n10454) );
  XNOR2_X1 U13003 ( .A(n10453), .B(n10454), .ZN(n12560) );
  AND2_X1 U13004 ( .A1(n12560), .A2(n10451), .ZN(n10452) );
  INV_X1 U13005 ( .A(n10453), .ZN(n12470) );
  NAND2_X1 U13006 ( .A1(n12470), .A2(n10454), .ZN(n10455) );
  NAND2_X1 U13007 ( .A1(n12555), .A2(n10455), .ZN(n10456) );
  XNOR2_X1 U13008 ( .A(n12366), .B(n10413), .ZN(n10459) );
  NOR2_X1 U13009 ( .A1(n10450), .A2(n12329), .ZN(n10457) );
  XNOR2_X1 U13010 ( .A(n10459), .B(n10457), .ZN(n12469) );
  INV_X1 U13011 ( .A(n10457), .ZN(n10458) );
  NAND2_X1 U13012 ( .A1(n10459), .A2(n10458), .ZN(n10460) );
  XNOR2_X1 U13013 ( .A(n12242), .B(n10413), .ZN(n10464) );
  NOR2_X1 U13014 ( .A1(n10450), .A2(n10461), .ZN(n10463) );
  XNOR2_X1 U13015 ( .A(n10464), .B(n10463), .ZN(n12657) );
  NAND2_X1 U13016 ( .A1(n10464), .A2(n10463), .ZN(n10465) );
  XNOR2_X1 U13017 ( .A(n14823), .B(n10413), .ZN(n10466) );
  OR2_X1 U13018 ( .A1(n10450), .A2(n14066), .ZN(n10467) );
  NAND2_X1 U13019 ( .A1(n10466), .A2(n10467), .ZN(n14142) );
  INV_X1 U13020 ( .A(n10466), .ZN(n10469) );
  INV_X1 U13021 ( .A(n10467), .ZN(n10468) );
  NAND2_X1 U13022 ( .A1(n10469), .A2(n10468), .ZN(n14141) );
  XNOR2_X1 U13023 ( .A(n14769), .B(n12750), .ZN(n10471) );
  OR2_X1 U13024 ( .A1(n10450), .A2(n14635), .ZN(n10472) );
  NAND2_X1 U13025 ( .A1(n10471), .A2(n10472), .ZN(n14062) );
  INV_X1 U13026 ( .A(n10471), .ZN(n10474) );
  INV_X1 U13027 ( .A(n10472), .ZN(n10473) );
  NAND2_X1 U13028 ( .A1(n10474), .A2(n10473), .ZN(n14063) );
  INV_X1 U13029 ( .A(n12760), .ZN(n10481) );
  XNOR2_X1 U13030 ( .A(n14816), .B(n10413), .ZN(n14010) );
  INV_X1 U13031 ( .A(n14010), .ZN(n10476) );
  OR2_X1 U13032 ( .A1(n10450), .A2(n14205), .ZN(n10477) );
  INV_X1 U13033 ( .A(n10477), .ZN(n10475) );
  NAND2_X1 U13034 ( .A1(n10476), .A2(n10475), .ZN(n12832) );
  NAND2_X1 U13035 ( .A1(n14010), .A2(n10477), .ZN(n12755) );
  NAND2_X1 U13036 ( .A1(n12832), .A2(n12755), .ZN(n10480) );
  NOR2_X1 U13037 ( .A1(n15910), .A2(n15913), .ZN(n10487) );
  AND2_X1 U13038 ( .A1(n15931), .A2(n11022), .ZN(n10479) );
  AOI211_X1 U13039 ( .C1(n10481), .C2(n10480), .A(n14154), .B(n14012), .ZN(
        n10497) );
  NOR2_X1 U13040 ( .A1(n10482), .A2(n9853), .ZN(n11977) );
  NAND2_X1 U13041 ( .A1(n10486), .A2(n11977), .ZN(n10484) );
  INV_X1 U13042 ( .A(n10488), .ZN(n10483) );
  NOR2_X1 U13043 ( .A1(n14173), .A2(n14816), .ZN(n10496) );
  NAND2_X1 U13044 ( .A1(n10486), .A2(n10485), .ZN(n14147) );
  OAI22_X1 U13045 ( .A1(n14184), .A2(n14637), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11607), .ZN(n10495) );
  INV_X1 U13046 ( .A(n10487), .ZN(n10489) );
  OAI21_X1 U13047 ( .B1(n10490), .B2(n10489), .A(n10488), .ZN(n11683) );
  NAND3_X1 U13048 ( .A1(n11683), .A2(n10492), .A3(n10491), .ZN(n10493) );
  OAI22_X1 U13049 ( .A1(n14643), .A2(n14186), .B1(n14185), .B2(n14635), .ZN(
        n10494) );
  OR4_X1 U13050 ( .A1(n10497), .A2(n10496), .A3(n10495), .A4(n10494), .ZN(
        P2_U3206) );
  NAND2_X1 U13051 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_STATE_REG_SCAN_IN), .ZN(
        n10498) );
  OAI21_X1 U13052 ( .B1(n10499), .B2(P3_STATE_REG_SCAN_IN), .A(n10498), .ZN(
        P3_U3295) );
  NOR2_X1 U13053 ( .A1(n6542), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13999) );
  INV_X1 U13054 ( .A(n10500), .ZN(n10502) );
  OAI222_X1 U13055 ( .A1(n11302), .A2(P3_U3151), .B1(n13257), .B2(n10502), 
        .C1(n10501), .C2(n14006), .ZN(P3_U3291) );
  INV_X1 U13056 ( .A(n10503), .ZN(n10505) );
  INV_X1 U13057 ( .A(SI_5_), .ZN(n10504) );
  OAI222_X1 U13058 ( .A1(n11217), .A2(P3_U3151), .B1(n13257), .B2(n10505), 
        .C1(n10504), .C2(n14006), .ZN(P3_U3290) );
  OAI222_X1 U13059 ( .A1(n11280), .A2(P3_U3151), .B1(n13257), .B2(n6785), .C1(
        n10506), .C2(n14006), .ZN(P3_U3293) );
  INV_X1 U13060 ( .A(n10507), .ZN(n10509) );
  INV_X1 U13061 ( .A(SI_3_), .ZN(n10508) );
  OAI222_X1 U13062 ( .A1(n11185), .A2(P3_U3151), .B1(n13257), .B2(n10509), 
        .C1(n10508), .C2(n14006), .ZN(P3_U3292) );
  NAND2_X1 U13063 ( .A1(n11387), .A2(n10512), .ZN(n10510) );
  OAI21_X1 U13064 ( .B1(n10512), .B2(n8533), .A(n10510), .ZN(P3_U3377) );
  NAND2_X1 U13065 ( .A1(n8097), .A2(n10512), .ZN(n10511) );
  OAI21_X1 U13066 ( .B1(n10512), .B2(n8093), .A(n10511), .ZN(P3_U3376) );
  INV_X1 U13067 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10513) );
  INV_X1 U13068 ( .A(n15684), .ZN(n15698) );
  OAI222_X1 U13069 ( .A1(n15597), .A2(n10513), .B1(n15595), .B2(n10626), .C1(
        n15698), .C2(P1_U3086), .ZN(P1_U3351) );
  OAI222_X1 U13070 ( .A1(n13257), .A2(n10515), .B1(n14006), .B2(n10514), .C1(
        n11483), .C2(P3_U3151), .ZN(P3_U3286) );
  OAI222_X1 U13071 ( .A1(P3_U3151), .A2(n11183), .B1(n14006), .B2(n10517), 
        .C1(n13257), .C2(n10516), .ZN(P3_U3294) );
  INV_X1 U13072 ( .A(n10518), .ZN(n10520) );
  INV_X1 U13073 ( .A(n11464), .ZN(n11467) );
  OAI222_X1 U13074 ( .A1(n13257), .A2(n10520), .B1(n14006), .B2(n10519), .C1(
        n11467), .C2(P3_U3151), .ZN(P3_U3287) );
  INV_X1 U13075 ( .A(n11258), .ZN(n11221) );
  OAI222_X1 U13076 ( .A1(n11221), .A2(P3_U3151), .B1(n13257), .B2(n10522), 
        .C1(n10521), .C2(n14006), .ZN(P3_U3289) );
  NAND2_X1 U13077 ( .A1(n6542), .A2(P2_U3088), .ZN(n12909) );
  NOR2_X1 U13078 ( .A1(n6542), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14830) );
  INV_X1 U13079 ( .A(n14830), .ZN(n14826) );
  OAI222_X1 U13080 ( .A1(P2_U3088), .A2(n14220), .B1(n12909), .B2(n10573), 
        .C1(n10525), .C2(n14826), .ZN(P2_U3326) );
  INV_X1 U13081 ( .A(n14260), .ZN(n10526) );
  OAI222_X1 U13082 ( .A1(n14826), .A2(n10527), .B1(n12909), .B2(n10570), .C1(
        n10526), .C2(P2_U3088), .ZN(P2_U3321) );
  NAND2_X1 U13083 ( .A1(n12480), .A2(P1_B_REG_SCAN_IN), .ZN(n10529) );
  INV_X1 U13084 ( .A(n12222), .ZN(n10528) );
  MUX2_X1 U13085 ( .A(n10529), .B(P1_B_REG_SCAN_IN), .S(n10528), .Z(n10530) );
  INV_X1 U13086 ( .A(n10530), .ZN(n10531) );
  NOR2_X1 U13087 ( .A1(n10531), .A2(n12487), .ZN(n10806) );
  INV_X1 U13088 ( .A(n10806), .ZN(n10810) );
  NAND2_X1 U13089 ( .A1(n10810), .A2(n10955), .ZN(n15771) );
  INV_X1 U13090 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10534) );
  NAND2_X1 U13091 ( .A1(n12480), .A2(n12487), .ZN(n10795) );
  INV_X1 U13092 ( .A(n10795), .ZN(n10533) );
  AOI22_X1 U13093 ( .A1(n15771), .A2(n10534), .B1(n10533), .B2(n10532), .ZN(
        P1_U3446) );
  INV_X1 U13094 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n15021) );
  NAND2_X1 U13095 ( .A1(n15021), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n10535) );
  NAND2_X1 U13096 ( .A1(n10554), .A2(n10535), .ZN(n10559) );
  NAND2_X1 U13097 ( .A1(n10536), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n10539) );
  INV_X1 U13098 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10537) );
  NAND2_X1 U13099 ( .A1(n10537), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n10538) );
  NAND2_X1 U13100 ( .A1(n10540), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n10541) );
  INV_X1 U13101 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n15035) );
  INV_X1 U13102 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n15704) );
  NAND2_X1 U13103 ( .A1(n15704), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n10543) );
  INV_X1 U13104 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n11285) );
  NAND2_X1 U13105 ( .A1(n11285), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n10542) );
  AND2_X1 U13106 ( .A1(n10543), .A2(n10542), .ZN(n10547) );
  NAND2_X1 U13107 ( .A1(n10548), .A2(n10547), .ZN(n10550) );
  INV_X1 U13108 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n11194) );
  INV_X1 U13109 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10544) );
  OR2_X1 U13110 ( .A1(n10545), .A2(n10544), .ZN(n10546) );
  NAND2_X1 U13111 ( .A1(n10550), .A2(n10549), .ZN(n10568) );
  INV_X1 U13112 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10551) );
  XNOR2_X1 U13113 ( .A(n10568), .B(n10551), .ZN(n15604) );
  OAI21_X1 U13114 ( .B1(n10553), .B2(n15035), .A(n10552), .ZN(n10567) );
  NAND2_X1 U13115 ( .A1(n10556), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n10557) );
  XNOR2_X1 U13116 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P3_ADDR_REG_0__SCAN_IN), 
        .ZN(n15601) );
  INV_X1 U13117 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15602) );
  NOR2_X1 U13118 ( .A1(n15601), .A2(n15602), .ZN(n16030) );
  OR2_X1 U13119 ( .A1(n10559), .A2(n10558), .ZN(n10560) );
  NAND2_X1 U13120 ( .A1(n10561), .A2(n10560), .ZN(n10563) );
  INV_X1 U13121 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n15670) );
  NAND2_X1 U13122 ( .A1(n15668), .A2(n15670), .ZN(n10566) );
  INV_X1 U13123 ( .A(n10562), .ZN(n10565) );
  INV_X1 U13124 ( .A(n10563), .ZN(n10564) );
  NAND2_X1 U13125 ( .A1(n10565), .A2(n10564), .ZN(n15669) );
  INV_X1 U13126 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n16027) );
  OAI21_X1 U13127 ( .B1(n6783), .B2(n15880), .A(n10813), .ZN(SUB_1596_U58) );
  INV_X1 U13128 ( .A(n10569), .ZN(n10628) );
  INV_X1 U13129 ( .A(n10688), .ZN(n10731) );
  OAI222_X1 U13130 ( .A1(n15597), .A2(n8607), .B1(n15595), .B2(n10628), .C1(
        P1_U3086), .C2(n10731), .ZN(P1_U3350) );
  INV_X1 U13131 ( .A(n10709), .ZN(n10670) );
  OAI222_X1 U13132 ( .A1(n15597), .A2(n10571), .B1(n15595), .B2(n10570), .C1(
        n10670), .C2(P1_U3086), .ZN(P1_U3349) );
  OAI222_X1 U13133 ( .A1(n15597), .A2(n10572), .B1(n15595), .B2(n10624), .C1(
        P1_U3086), .C2(n10683), .ZN(P1_U3353) );
  OAI222_X1 U13134 ( .A1(n15597), .A2(n8594), .B1(n15595), .B2(n10573), .C1(
        n10678), .C2(P1_U3086), .ZN(P1_U3354) );
  INV_X1 U13135 ( .A(n15040), .ZN(n10574) );
  OAI222_X1 U13136 ( .A1(n15597), .A2(n10575), .B1(n15595), .B2(n10630), .C1(
        n10574), .C2(P1_U3086), .ZN(P1_U3352) );
  OAI222_X1 U13137 ( .A1(n13257), .A2(n10577), .B1(n14006), .B2(n10576), .C1(
        n11327), .C2(P3_U3151), .ZN(P3_U3288) );
  OAI222_X1 U13138 ( .A1(n13257), .A2(n10579), .B1(n14006), .B2(n10578), .C1(
        n11885), .C2(P3_U3151), .ZN(P3_U3285) );
  OAI222_X1 U13139 ( .A1(n13257), .A2(n10581), .B1(n14006), .B2(n10580), .C1(
        n12145), .C2(P3_U3151), .ZN(P3_U3284) );
  INV_X1 U13140 ( .A(n10582), .ZN(n10636) );
  INV_X1 U13141 ( .A(n10691), .ZN(n10718) );
  OAI222_X1 U13142 ( .A1(n15597), .A2(n10583), .B1(n15595), .B2(n10636), .C1(
        P1_U3086), .C2(n10718), .ZN(P1_U3348) );
  NOR2_X1 U13143 ( .A1(n8532), .A2(n10584), .ZN(n10586) );
  INV_X1 U13144 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10585) );
  NOR2_X1 U13145 ( .A1(n10615), .A2(n10585), .ZN(P3_U3246) );
  CLKBUF_X1 U13146 ( .A(n10586), .Z(n10615) );
  INV_X1 U13147 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10587) );
  NOR2_X1 U13148 ( .A1(n10615), .A2(n10587), .ZN(P3_U3237) );
  INV_X1 U13149 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10588) );
  NOR2_X1 U13150 ( .A1(n10615), .A2(n10588), .ZN(P3_U3236) );
  INV_X1 U13151 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10589) );
  NOR2_X1 U13152 ( .A1(n10586), .A2(n10589), .ZN(P3_U3247) );
  INV_X1 U13153 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10590) );
  NOR2_X1 U13154 ( .A1(n10615), .A2(n10590), .ZN(P3_U3234) );
  INV_X1 U13155 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10591) );
  NOR2_X1 U13156 ( .A1(n10615), .A2(n10591), .ZN(P3_U3244) );
  INV_X1 U13157 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10592) );
  NOR2_X1 U13158 ( .A1(n10615), .A2(n10592), .ZN(P3_U3245) );
  INV_X1 U13159 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10593) );
  NOR2_X1 U13160 ( .A1(n10615), .A2(n10593), .ZN(P3_U3242) );
  INV_X1 U13161 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10594) );
  NOR2_X1 U13162 ( .A1(n10615), .A2(n10594), .ZN(P3_U3241) );
  INV_X1 U13163 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10595) );
  NOR2_X1 U13164 ( .A1(n10586), .A2(n10595), .ZN(P3_U3248) );
  INV_X1 U13165 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10596) );
  NOR2_X1 U13166 ( .A1(n10615), .A2(n10596), .ZN(P3_U3239) );
  INV_X1 U13167 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10597) );
  NOR2_X1 U13168 ( .A1(n10615), .A2(n10597), .ZN(P3_U3238) );
  INV_X1 U13169 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10598) );
  NOR2_X1 U13170 ( .A1(n10615), .A2(n10598), .ZN(P3_U3235) );
  INV_X1 U13171 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10599) );
  NOR2_X1 U13172 ( .A1(n10586), .A2(n10599), .ZN(P3_U3250) );
  NOR2_X1 U13173 ( .A1(n10586), .A2(n10600), .ZN(P3_U3257) );
  INV_X1 U13174 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10601) );
  NOR2_X1 U13175 ( .A1(n10615), .A2(n10601), .ZN(P3_U3258) );
  INV_X1 U13176 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10602) );
  NOR2_X1 U13177 ( .A1(n10586), .A2(n10602), .ZN(P3_U3259) );
  INV_X1 U13178 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10603) );
  NOR2_X1 U13179 ( .A1(n10615), .A2(n10603), .ZN(P3_U3260) );
  INV_X1 U13180 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10604) );
  NOR2_X1 U13181 ( .A1(n10586), .A2(n10604), .ZN(P3_U3261) );
  INV_X1 U13182 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10605) );
  NOR2_X1 U13183 ( .A1(n10615), .A2(n10605), .ZN(P3_U3262) );
  INV_X1 U13184 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10606) );
  NOR2_X1 U13185 ( .A1(n10586), .A2(n10606), .ZN(P3_U3263) );
  INV_X1 U13186 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10607) );
  NOR2_X1 U13187 ( .A1(n10586), .A2(n10607), .ZN(P3_U3256) );
  INV_X1 U13188 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10608) );
  NOR2_X1 U13189 ( .A1(n10586), .A2(n10608), .ZN(P3_U3255) );
  INV_X1 U13190 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10609) );
  NOR2_X1 U13191 ( .A1(n10586), .A2(n10609), .ZN(P3_U3249) );
  INV_X1 U13192 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10610) );
  NOR2_X1 U13193 ( .A1(n10586), .A2(n10610), .ZN(P3_U3253) );
  INV_X1 U13194 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10611) );
  NOR2_X1 U13195 ( .A1(n10615), .A2(n10611), .ZN(P3_U3251) );
  NOR2_X1 U13196 ( .A1(n10615), .A2(n10612), .ZN(P3_U3243) );
  INV_X1 U13197 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10613) );
  NOR2_X1 U13198 ( .A1(n10615), .A2(n10613), .ZN(P3_U3252) );
  INV_X1 U13199 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10614) );
  NOR2_X1 U13200 ( .A1(n10615), .A2(n10614), .ZN(P3_U3240) );
  INV_X1 U13201 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10616) );
  NOR2_X1 U13202 ( .A1(n10615), .A2(n10616), .ZN(P3_U3254) );
  INV_X1 U13203 ( .A(n10617), .ZN(n10633) );
  INV_X1 U13204 ( .A(n10751), .ZN(n10747) );
  OAI222_X1 U13205 ( .A1(n15597), .A2(n10618), .B1(n15595), .B2(n10633), .C1(
        n10747), .C2(P1_U3086), .ZN(P1_U3347) );
  INV_X1 U13206 ( .A(n15771), .ZN(n15770) );
  NAND2_X1 U13207 ( .A1(n12222), .A2(n12487), .ZN(n10809) );
  OAI22_X1 U13208 ( .A1(n15770), .A2(P1_D_REG_0__SCAN_IN), .B1(n10809), .B2(
        n10619), .ZN(n10620) );
  INV_X1 U13209 ( .A(n10620), .ZN(P1_U3445) );
  INV_X1 U13210 ( .A(n10621), .ZN(n10631) );
  INV_X1 U13211 ( .A(n10752), .ZN(n11075) );
  OAI222_X1 U13212 ( .A1(n15597), .A2(n10622), .B1(n15595), .B2(n10631), .C1(
        P1_U3086), .C2(n11075), .ZN(P1_U3346) );
  INV_X1 U13213 ( .A(n12909), .ZN(n13261) );
  INV_X1 U13214 ( .A(n13261), .ZN(n14832) );
  AOI22_X1 U13215 ( .A1(n14231), .A2(P2_STATE_REG_SCAN_IN), .B1(n14830), .B2(
        P1_DATAO_REG_2__SCAN_IN), .ZN(n10623) );
  OAI21_X1 U13216 ( .B1(n10624), .B2(n14832), .A(n10623), .ZN(P2_U3325) );
  AOI22_X1 U13217 ( .A1(n14246), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n14830), .ZN(n10625) );
  OAI21_X1 U13218 ( .B1(n10626), .B2(n14832), .A(n10625), .ZN(P2_U3323) );
  AOI22_X1 U13219 ( .A1(n15869), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n14830), .ZN(n10627) );
  OAI21_X1 U13220 ( .B1(n10628), .B2(n14832), .A(n10627), .ZN(P2_U3322) );
  AOI22_X1 U13221 ( .A1(n15855), .A2(P2_STATE_REG_SCAN_IN), .B1(n14830), .B2(
        P1_DATAO_REG_3__SCAN_IN), .ZN(n10629) );
  OAI21_X1 U13222 ( .B1(n10630), .B2(n14832), .A(n10629), .ZN(P2_U3324) );
  INV_X1 U13223 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10632) );
  INV_X1 U13224 ( .A(n11094), .ZN(n11049) );
  OAI222_X1 U13225 ( .A1(n14826), .A2(n10632), .B1(n14832), .B2(n10631), .C1(
        P2_U3088), .C2(n11049), .ZN(P2_U3318) );
  INV_X1 U13226 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10634) );
  OAI222_X1 U13227 ( .A1(n14826), .A2(n10634), .B1(n14832), .B2(n10633), .C1(
        n11059), .C2(P2_U3088), .ZN(P2_U3319) );
  INV_X1 U13228 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10637) );
  INV_X1 U13229 ( .A(n14272), .ZN(n10635) );
  OAI222_X1 U13230 ( .A1(n14826), .A2(n10637), .B1(n14832), .B2(n10636), .C1(
        P2_U3088), .C2(n10635), .ZN(P2_U3320) );
  INV_X1 U13231 ( .A(n10638), .ZN(n10640) );
  INV_X1 U13232 ( .A(n13475), .ZN(n13467) );
  OAI222_X1 U13233 ( .A1(n13257), .A2(n10640), .B1(n13467), .B2(P3_U3151), 
        .C1(n10639), .C2(n14006), .ZN(P3_U3283) );
  INV_X1 U13234 ( .A(n10956), .ZN(n10641) );
  OR2_X1 U13235 ( .A1(n10944), .A2(n10641), .ZN(n10643) );
  AND2_X1 U13236 ( .A1(n10643), .A2(n10642), .ZN(n10675) );
  INV_X1 U13237 ( .A(n10675), .ZN(n10645) );
  INV_X1 U13238 ( .A(n10955), .ZN(n11439) );
  NAND2_X1 U13239 ( .A1(n11439), .A2(n10644), .ZN(n10674) );
  AND2_X1 U13240 ( .A1(n10645), .A2(n10674), .ZN(n15680) );
  NOR2_X1 U13241 ( .A1(n15680), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U13242 ( .A(n10646), .ZN(n10653) );
  INV_X1 U13243 ( .A(n15597), .ZN(n15588) );
  AOI22_X1 U13244 ( .A1(n15710), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n15588), .ZN(n10647) );
  OAI21_X1 U13245 ( .B1(n10653), .B2(n15595), .A(n10647), .ZN(P1_U3343) );
  INV_X1 U13246 ( .A(n11698), .ZN(n10649) );
  OAI222_X1 U13247 ( .A1(P2_U3088), .A2(n10649), .B1(n12909), .B2(n10650), 
        .C1(n10648), .C2(n14826), .ZN(P2_U3314) );
  INV_X1 U13248 ( .A(n15066), .ZN(n15072) );
  OAI222_X1 U13249 ( .A1(n15597), .A2(n10651), .B1(n15595), .B2(n10650), .C1(
        n15072), .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U13250 ( .A(n15895), .ZN(n10654) );
  INV_X1 U13251 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10652) );
  OAI222_X1 U13252 ( .A1(P2_U3088), .A2(n10654), .B1(n12909), .B2(n10653), 
        .C1(n10652), .C2(n14826), .ZN(P2_U3315) );
  INV_X1 U13253 ( .A(n15054), .ZN(n11069) );
  OAI222_X1 U13254 ( .A1(n15597), .A2(n10655), .B1(n15595), .B2(n10657), .C1(
        n11069), .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U13255 ( .A(n11114), .ZN(n10656) );
  OAI222_X1 U13256 ( .A1(n14826), .A2(n10658), .B1(n14832), .B2(n10657), .C1(
        n10656), .C2(P2_U3088), .ZN(P2_U3317) );
  OAI222_X1 U13257 ( .A1(n13257), .A2(n10660), .B1(n14006), .B2(n10659), .C1(
        n13486), .C2(P3_U3151), .ZN(P3_U3282) );
  OAI222_X1 U13258 ( .A1(n13257), .A2(n10662), .B1(n13534), .B2(P3_U3151), 
        .C1(n14006), .C2(n10661), .ZN(P3_U3280) );
  OAI222_X1 U13259 ( .A1(n13257), .A2(n10664), .B1(n14006), .B2(n10663), .C1(
        n13508), .C2(P3_U3151), .ZN(P3_U3281) );
  MUX2_X1 U13260 ( .A(n10746), .B(P1_REG1_REG_8__SCAN_IN), .S(n10751), .Z(
        n10673) );
  INV_X1 U13261 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10668) );
  AND2_X1 U13262 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n15025) );
  NAND2_X1 U13263 ( .A1(n15026), .A2(n15025), .ZN(n15024) );
  NAND2_X1 U13264 ( .A1(n15023), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10665) );
  NAND2_X1 U13265 ( .A1(n15024), .A2(n10665), .ZN(n10884) );
  MUX2_X1 U13266 ( .A(n15840), .B(P1_REG1_REG_2__SCAN_IN), .S(n10683), .Z(
        n10885) );
  NAND2_X1 U13267 ( .A1(n10884), .A2(n10885), .ZN(n10883) );
  NAND2_X1 U13268 ( .A1(n10889), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n10666) );
  NAND2_X1 U13269 ( .A1(n10883), .A2(n10666), .ZN(n15038) );
  INV_X1 U13270 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n15842) );
  MUX2_X1 U13271 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n15842), .S(n15040), .Z(
        n15039) );
  NAND2_X1 U13272 ( .A1(n15040), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n15692) );
  NAND2_X1 U13273 ( .A1(n15691), .A2(n15692), .ZN(n10667) );
  MUX2_X1 U13274 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10668), .S(n15684), .Z(
        n15690) );
  NAND2_X1 U13275 ( .A1(n10667), .A2(n15690), .ZN(n15695) );
  OAI21_X1 U13276 ( .B1(n10668), .B2(n15698), .A(n15695), .ZN(n10729) );
  XNOR2_X1 U13277 ( .A(n10688), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n10730) );
  MUX2_X1 U13278 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n11723), .S(n10709), .Z(
        n10711) );
  MUX2_X1 U13279 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n10671), .S(n10691), .Z(
        n10722) );
  OAI21_X1 U13280 ( .B1(n10671), .B2(n10718), .A(n10721), .ZN(n10672) );
  AOI21_X1 U13281 ( .B1(n10673), .B2(n10672), .A(n10745), .ZN(n10702) );
  NAND2_X1 U13282 ( .A1(n10675), .A2(n10674), .ZN(n15683) );
  OR2_X1 U13283 ( .A1(n15683), .A2(n15150), .ZN(n15102) );
  OR2_X1 U13284 ( .A1(n15683), .A2(n10676), .ZN(n15699) );
  INV_X1 U13285 ( .A(n15699), .ZN(n15720) );
  INV_X1 U13286 ( .A(n15680), .ZN(n15728) );
  INV_X1 U13287 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10837) );
  NAND2_X1 U13288 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11929) );
  OAI21_X1 U13289 ( .B1(n15728), .B2(n10837), .A(n11929), .ZN(n10677) );
  AOI21_X1 U13290 ( .B1(n10751), .B2(n15720), .A(n10677), .ZN(n10701) );
  INV_X1 U13291 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10679) );
  AND2_X1 U13292 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n10680) );
  NAND2_X1 U13293 ( .A1(n15029), .A2(n10680), .ZN(n15028) );
  NAND2_X1 U13294 ( .A1(n15023), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10681) );
  NAND2_X1 U13295 ( .A1(n15028), .A2(n10681), .ZN(n10886) );
  MUX2_X1 U13296 ( .A(n10682), .B(P1_REG2_REG_2__SCAN_IN), .S(n10683), .Z(
        n10887) );
  NAND2_X1 U13297 ( .A1(n10886), .A2(n10887), .ZN(n15042) );
  NAND2_X1 U13298 ( .A1(n10889), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n15041) );
  NAND2_X1 U13299 ( .A1(n15042), .A2(n15041), .ZN(n10685) );
  MUX2_X1 U13300 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n7249), .S(n15040), .Z(
        n10684) );
  NAND2_X1 U13301 ( .A1(n10685), .A2(n10684), .ZN(n15687) );
  NAND2_X1 U13302 ( .A1(n15040), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n15686) );
  NAND2_X1 U13303 ( .A1(n15687), .A2(n15686), .ZN(n10687) );
  INV_X1 U13304 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11514) );
  MUX2_X1 U13305 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n11514), .S(n15684), .Z(
        n10686) );
  NAND2_X1 U13306 ( .A1(n15684), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10736) );
  INV_X1 U13307 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10689) );
  MUX2_X1 U13308 ( .A(n10689), .B(P1_REG2_REG_5__SCAN_IN), .S(n10688), .Z(
        n10735) );
  NOR2_X1 U13309 ( .A1(n10731), .A2(n10689), .ZN(n10704) );
  MUX2_X1 U13310 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10690), .S(n10709), .Z(
        n10703) );
  NAND2_X1 U13311 ( .A1(n10709), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10715) );
  MUX2_X1 U13312 ( .A(n10692), .B(P1_REG2_REG_7__SCAN_IN), .S(n10691), .Z(
        n10714) );
  NOR2_X1 U13313 ( .A1(n10718), .A2(n10692), .ZN(n10697) );
  INV_X1 U13314 ( .A(n10697), .ZN(n10695) );
  INV_X1 U13315 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10693) );
  MUX2_X1 U13316 ( .A(n10693), .B(P1_REG2_REG_8__SCAN_IN), .S(n10751), .Z(
        n10694) );
  NAND2_X1 U13317 ( .A1(n10695), .A2(n10694), .ZN(n10699) );
  MUX2_X1 U13318 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10693), .S(n10751), .Z(
        n10696) );
  OAI21_X1 U13319 ( .B1(n10727), .B2(n10697), .A(n10696), .ZN(n10755) );
  OR2_X1 U13320 ( .A1(n15674), .A2(n8855), .ZN(n10698) );
  OR2_X1 U13321 ( .A1(n15683), .A2(n10698), .ZN(n15142) );
  OAI211_X1 U13322 ( .C1(n10727), .C2(n10699), .A(n10755), .B(n15724), .ZN(
        n10700) );
  OAI211_X1 U13323 ( .C1(n10702), .C2(n15102), .A(n10701), .B(n10700), .ZN(
        P1_U3251) );
  INV_X1 U13324 ( .A(n10716), .ZN(n10706) );
  NOR3_X1 U13325 ( .A1(n10734), .A2(n10704), .A3(n10703), .ZN(n10705) );
  NOR3_X1 U13326 ( .A1(n15142), .A2(n10706), .A3(n10705), .ZN(n10708) );
  INV_X1 U13327 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10825) );
  NAND2_X1 U13328 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n11792) );
  OAI21_X1 U13329 ( .B1(n15728), .B2(n10825), .A(n11792), .ZN(n10707) );
  AOI211_X1 U13330 ( .C1(n15720), .C2(n10709), .A(n10708), .B(n10707), .ZN(
        n10713) );
  OAI211_X1 U13331 ( .C1(n10711), .C2(n6784), .A(n15723), .B(n10710), .ZN(
        n10712) );
  NAND2_X1 U13332 ( .A1(n10713), .A2(n10712), .ZN(P1_U3249) );
  NAND3_X1 U13333 ( .A1(n10716), .A2(n10715), .A3(n10714), .ZN(n10717) );
  NAND2_X1 U13334 ( .A1(n15724), .A2(n10717), .ZN(n10726) );
  NOR2_X1 U13335 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8821), .ZN(n10720) );
  NOR2_X1 U13336 ( .A1(n15699), .A2(n10718), .ZN(n10719) );
  AOI211_X1 U13337 ( .C1(n15680), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n10720), .B(
        n10719), .ZN(n10725) );
  OAI211_X1 U13338 ( .C1(n10723), .C2(n10722), .A(n10721), .B(n15723), .ZN(
        n10724) );
  OAI211_X1 U13339 ( .C1(n10727), .C2(n10726), .A(n10725), .B(n10724), .ZN(
        P1_U3250) );
  AOI21_X1 U13340 ( .B1(n10730), .B2(n10729), .A(n10728), .ZN(n10741) );
  AND2_X1 U13341 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10733) );
  NOR2_X1 U13342 ( .A1(n15699), .A2(n10731), .ZN(n10732) );
  AOI211_X1 U13343 ( .C1(n15680), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n10733), .B(
        n10732), .ZN(n10740) );
  INV_X1 U13344 ( .A(n10734), .ZN(n10738) );
  NAND3_X1 U13345 ( .A1(n15689), .A2(n10736), .A3(n10735), .ZN(n10737) );
  NAND3_X1 U13346 ( .A1(n15724), .A2(n10738), .A3(n10737), .ZN(n10739) );
  OAI211_X1 U13347 ( .C1(n10741), .C2(n15102), .A(n10740), .B(n10739), .ZN(
        P1_U3248) );
  INV_X1 U13348 ( .A(n10742), .ZN(n10744) );
  INV_X1 U13349 ( .A(n13556), .ZN(n13569) );
  OAI222_X1 U13350 ( .A1(n13257), .A2(n10744), .B1(n13569), .B2(P3_U3151), 
        .C1(n10743), .C2(n14006), .ZN(P3_U3279) );
  MUX2_X1 U13351 ( .A(n11068), .B(P1_REG1_REG_9__SCAN_IN), .S(n10752), .Z(
        n10749) );
  AOI21_X1 U13352 ( .B1(n10749), .B2(n10748), .A(n11067), .ZN(n10760) );
  INV_X1 U13353 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n11320) );
  NAND2_X1 U13354 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n12645) );
  OAI21_X1 U13355 ( .B1(n15728), .B2(n11320), .A(n12645), .ZN(n10750) );
  AOI21_X1 U13356 ( .B1(n10752), .B2(n15720), .A(n10750), .ZN(n10759) );
  NAND2_X1 U13357 ( .A1(n10751), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10754) );
  MUX2_X1 U13358 ( .A(n12017), .B(P1_REG2_REG_9__SCAN_IN), .S(n10752), .Z(
        n10753) );
  AOI21_X1 U13359 ( .B1(n10755), .B2(n10754), .A(n10753), .ZN(n15060) );
  INV_X1 U13360 ( .A(n15060), .ZN(n10757) );
  NAND3_X1 U13361 ( .A1(n10755), .A2(n10754), .A3(n10753), .ZN(n10756) );
  NAND3_X1 U13362 ( .A1(n10757), .A2(n15724), .A3(n10756), .ZN(n10758) );
  OAI211_X1 U13363 ( .C1(n10760), .C2(n15102), .A(n10759), .B(n10758), .ZN(
        P1_U3252) );
  INV_X1 U13364 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10762) );
  INV_X1 U13365 ( .A(n10761), .ZN(n10765) );
  OAI222_X1 U13366 ( .A1(n14826), .A2(n10762), .B1(n14832), .B2(n10765), .C1(
        P2_U3088), .C2(n11601), .ZN(P2_U3316) );
  NAND2_X1 U13367 ( .A1(n11848), .A2(n13461), .ZN(n10763) );
  OAI21_X1 U13368 ( .B1(n13461), .B2(n10764), .A(n10763), .ZN(P3_U3500) );
  INV_X1 U13369 ( .A(n11771), .ZN(n11767) );
  OAI222_X1 U13370 ( .A1(n7257), .A2(n15597), .B1(P1_U3086), .B2(n11767), .C1(
        n15595), .C2(n10765), .ZN(P1_U3344) );
  OAI222_X1 U13371 ( .A1(n13257), .A2(n10767), .B1(n14006), .B2(n10766), .C1(
        n13581), .C2(P3_U3151), .ZN(P3_U3278) );
  INV_X1 U13372 ( .A(n14291), .ZN(n12208) );
  INV_X1 U13373 ( .A(n10768), .ZN(n10770) );
  OAI222_X1 U13374 ( .A1(P2_U3088), .A2(n12208), .B1(n12909), .B2(n10770), 
        .C1(n10769), .C2(n14826), .ZN(P2_U3311) );
  INV_X1 U13375 ( .A(n15101), .ZN(n15106) );
  OAI222_X1 U13376 ( .A1(n15597), .A2(n10771), .B1(n15595), .B2(n10770), .C1(
        n15106), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U13377 ( .A(n14309), .ZN(n14289) );
  INV_X1 U13378 ( .A(n10772), .ZN(n10774) );
  OAI222_X1 U13379 ( .A1(P2_U3088), .A2(n14289), .B1(n12909), .B2(n10774), 
        .C1(n10773), .C2(n14826), .ZN(P2_U3310) );
  OAI222_X1 U13380 ( .A1(n15597), .A2(n10775), .B1(n15595), .B2(n10774), .C1(
        n15120), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U13381 ( .A(n10776), .ZN(n10779) );
  INV_X1 U13382 ( .A(n15081), .ZN(n15087) );
  OAI222_X1 U13383 ( .A1(n15597), .A2(n10777), .B1(n15595), .B2(n10779), .C1(
        n15087), .C2(P1_U3086), .ZN(P1_U3341) );
  INV_X1 U13384 ( .A(n11940), .ZN(n11695) );
  OAI222_X1 U13385 ( .A1(P2_U3088), .A2(n11695), .B1(n12909), .B2(n10779), 
        .C1(n10778), .C2(n14826), .ZN(P2_U3313) );
  INV_X1 U13386 ( .A(n10780), .ZN(n10782) );
  INV_X1 U13387 ( .A(n13607), .ZN(n13585) );
  OAI222_X1 U13388 ( .A1(n13257), .A2(n10782), .B1(n14006), .B2(n10781), .C1(
        n13585), .C2(P3_U3151), .ZN(P3_U3277) );
  INV_X1 U13389 ( .A(n10783), .ZN(n10851) );
  AOI22_X1 U13390 ( .A1(n15721), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n15588), .ZN(n10784) );
  OAI21_X1 U13391 ( .B1(n10851), .B2(n15595), .A(n10784), .ZN(P1_U3340) );
  INV_X1 U13392 ( .A(n15980), .ZN(n13006) );
  NAND2_X1 U13393 ( .A1(n13464), .A2(n11399), .ZN(n13000) );
  AND2_X1 U13394 ( .A1(n13006), .A2(n13000), .ZN(n12972) );
  NOR2_X1 U13395 ( .A1(n13443), .A2(P3_U3151), .ZN(n10869) );
  INV_X1 U13396 ( .A(n10869), .ZN(n10785) );
  NAND2_X1 U13397 ( .A1(n10785), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10787) );
  INV_X1 U13398 ( .A(n13446), .ZN(n13400) );
  AOI22_X1 U13399 ( .A1(n13400), .A2(n12677), .B1(n13430), .B2(n8170), .ZN(
        n10786) );
  OAI211_X1 U13400 ( .C1(n12972), .C2(n13413), .A(n10787), .B(n10786), .ZN(
        P3_U3172) );
  AND2_X1 U13401 ( .A1(n10808), .A2(n10788), .ZN(n10943) );
  NOR2_X1 U13402 ( .A1(n15411), .A2(n10950), .ZN(n11445) );
  OR2_X1 U13403 ( .A1(n10871), .A2(n10790), .ZN(n10791) );
  AND2_X1 U13404 ( .A1(n11908), .A2(n10791), .ZN(n11446) );
  NAND2_X1 U13405 ( .A1(n11446), .A2(n6539), .ZN(n15433) );
  NAND2_X1 U13406 ( .A1(n10807), .A2(n15748), .ZN(n15815) );
  NAND2_X1 U13407 ( .A1(n15433), .A2(n15815), .ZN(n15835) );
  NAND2_X1 U13408 ( .A1(n15598), .A2(n15748), .ZN(n10792) );
  NAND2_X1 U13409 ( .A1(n10793), .A2(n10792), .ZN(n15754) );
  AOI21_X1 U13410 ( .B1(n15801), .B2(n15829), .A(n11447), .ZN(n10794) );
  AOI211_X1 U13411 ( .C1(n10943), .C2(n8869), .A(n11445), .B(n10794), .ZN(
        n10970) );
  OAI21_X1 U13412 ( .B1(n10810), .B2(P1_D_REG_1__SCAN_IN), .A(n10795), .ZN(
        n10940) );
  NOR4_X1 U13413 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n10804) );
  NOR4_X1 U13414 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n10803) );
  NAND4_X1 U13415 ( .A1(n15765), .A2(n15769), .A3(n15766), .A4(n15768), .ZN(
        n10801) );
  NOR4_X1 U13416 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n10799) );
  NOR4_X1 U13417 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n10798) );
  NOR4_X1 U13418 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n10797) );
  NOR4_X1 U13419 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n10796) );
  NAND4_X1 U13420 ( .A1(n10799), .A2(n10798), .A3(n10797), .A4(n10796), .ZN(
        n10800) );
  NOR4_X1 U13421 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        n10801), .A4(n10800), .ZN(n10802) );
  NAND3_X1 U13422 ( .A1(n10804), .A2(n10803), .A3(n10802), .ZN(n10805) );
  NAND2_X1 U13423 ( .A1(n10806), .A2(n10805), .ZN(n11435) );
  NAND2_X1 U13424 ( .A1(n10870), .A2(n15748), .ZN(n11440) );
  NAND4_X1 U13425 ( .A1(n11438), .A2(n10940), .A3(n11435), .A4(n11440), .ZN(
        n10969) );
  OAI21_X1 U13426 ( .B1(n10810), .B2(P1_D_REG_0__SCAN_IN), .A(n10809), .ZN(
        n11436) );
  NAND2_X1 U13427 ( .A1(n15848), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10811) );
  OAI21_X1 U13428 ( .B1(n10970), .B2(n15848), .A(n10811), .ZN(P1_U3528) );
  NAND2_X1 U13429 ( .A1(n10813), .A2(n10812), .ZN(n10818) );
  NAND2_X1 U13430 ( .A1(n10814), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n10815) );
  NAND2_X1 U13431 ( .A1(n10816), .A2(n10815), .ZN(n10824) );
  XNOR2_X1 U13432 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n10817) );
  XNOR2_X1 U13433 ( .A(n10824), .B(n10817), .ZN(n15606) );
  INV_X1 U13434 ( .A(n10818), .ZN(n10819) );
  NAND2_X1 U13435 ( .A1(n10819), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n10820) );
  INV_X1 U13436 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10821) );
  INV_X1 U13437 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n10822) );
  NAND2_X1 U13438 ( .A1(n10822), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n10823) );
  NAND2_X1 U13439 ( .A1(n10824), .A2(n10823), .ZN(n10827) );
  NAND2_X1 U13440 ( .A1(n10825), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n10826) );
  NAND2_X1 U13441 ( .A1(n10827), .A2(n10826), .ZN(n10833) );
  XNOR2_X1 U13442 ( .A(n10833), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n10832) );
  XNOR2_X1 U13443 ( .A(n10832), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15608) );
  NAND2_X1 U13444 ( .A1(n10828), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n10829) );
  INV_X1 U13445 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10831) );
  INV_X1 U13446 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n10836) );
  NAND2_X1 U13447 ( .A1(n10836), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n10846) );
  NAND2_X1 U13448 ( .A1(n10837), .A2(P3_ADDR_REG_8__SCAN_IN), .ZN(n10838) );
  AND2_X1 U13449 ( .A1(n10846), .A2(n10838), .ZN(n10844) );
  XNOR2_X1 U13450 ( .A(n10845), .B(n10844), .ZN(n10839) );
  NAND2_X1 U13451 ( .A1(n15609), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n10843) );
  INV_X1 U13452 ( .A(n10839), .ZN(n10840) );
  NAND2_X1 U13453 ( .A1(n10841), .A2(n10840), .ZN(n10842) );
  NAND2_X1 U13454 ( .A1(n10845), .A2(n10844), .ZN(n10847) );
  NAND2_X1 U13455 ( .A1(n10847), .A2(n10846), .ZN(n11319) );
  INV_X1 U13456 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n10848) );
  XNOR2_X1 U13457 ( .A(n10848), .B(P1_ADDR_REG_9__SCAN_IN), .ZN(n11318) );
  INV_X1 U13458 ( .A(n11318), .ZN(n10849) );
  XNOR2_X1 U13459 ( .A(n11319), .B(n10849), .ZN(n11315) );
  INV_X1 U13460 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n11312) );
  XNOR2_X1 U13461 ( .A(n11315), .B(n11312), .ZN(n10850) );
  XNOR2_X1 U13462 ( .A(n11314), .B(n10850), .ZN(SUB_1596_U54) );
  INV_X1 U13463 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10852) );
  INV_X1 U13464 ( .A(n12210), .ZN(n11943) );
  OAI222_X1 U13465 ( .A1(n14826), .A2(n10852), .B1(n12909), .B2(n10851), .C1(
        P2_U3088), .C2(n11943), .ZN(P2_U3312) );
  INV_X1 U13466 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n11266) );
  OAI21_X1 U13467 ( .B1(n10855), .B2(n10854), .A(n10853), .ZN(n10856) );
  NAND2_X1 U13468 ( .A1(n10856), .A2(n13437), .ZN(n10859) );
  OAI22_X1 U13469 ( .A1(n13441), .A2(n15967), .B1(n13428), .B2(n10860), .ZN(
        n10857) );
  AOI21_X1 U13470 ( .B1(n10900), .B2(n13400), .A(n10857), .ZN(n10858) );
  OAI211_X1 U13471 ( .C1(n10869), .C2(n11266), .A(n10859), .B(n10858), .ZN(
        P3_U3177) );
  NAND2_X1 U13472 ( .A1(n10866), .A2(n10860), .ZN(n13007) );
  AND2_X2 U13473 ( .A1(n13008), .A2(n13007), .ZN(n10905) );
  INV_X1 U13474 ( .A(n10905), .ZN(n13004) );
  NAND3_X1 U13475 ( .A1(n13004), .A2(n13006), .A3(n8332), .ZN(n10861) );
  OAI211_X1 U13476 ( .C1(n10863), .C2(n15986), .A(n10862), .B(n10861), .ZN(
        n10864) );
  NAND2_X1 U13477 ( .A1(n10864), .A2(n13437), .ZN(n10868) );
  INV_X1 U13478 ( .A(n13464), .ZN(n15989) );
  OAI22_X1 U13479 ( .A1(n13441), .A2(n15991), .B1(n13428), .B2(n15989), .ZN(
        n10865) );
  AOI21_X1 U13480 ( .B1(n10866), .B2(n13400), .A(n10865), .ZN(n10867) );
  OAI211_X1 U13481 ( .C1(n10869), .C2(n10057), .A(n10868), .B(n10867), .ZN(
        P3_U3162) );
  NAND2_X1 U13482 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n15027) );
  NAND2_X1 U13483 ( .A1(n10875), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n10872) );
  NAND2_X1 U13484 ( .A1(n10875), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10878) );
  NAND2_X1 U13485 ( .A1(n8869), .A2(n10876), .ZN(n10877) );
  OAI211_X1 U13486 ( .C1(n15749), .C2(n13224), .A(n10878), .B(n10877), .ZN(
        n10947) );
  NAND2_X1 U13487 ( .A1(n10879), .A2(n10947), .ZN(n10949) );
  OAI21_X1 U13488 ( .B1(n10879), .B2(n10947), .A(n10949), .ZN(n10973) );
  MUX2_X1 U13489 ( .A(n15027), .B(n10973), .S(n15674), .Z(n10880) );
  NOR2_X1 U13490 ( .A1(n10880), .A2(n8855), .ZN(n10882) );
  NOR2_X1 U13491 ( .A1(n15674), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10881) );
  NOR2_X1 U13492 ( .A1(n8855), .A2(n10881), .ZN(n15675) );
  NOR2_X1 U13493 ( .A1(n15675), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n15672) );
  NOR3_X1 U13494 ( .A1(n10882), .A2(n15672), .A3(n15019), .ZN(n15701) );
  OAI211_X1 U13495 ( .C1(n10885), .C2(n10884), .A(n15723), .B(n10883), .ZN(
        n10893) );
  OAI211_X1 U13496 ( .C1(n10887), .C2(n10886), .A(n15724), .B(n15042), .ZN(
        n10892) );
  NOR2_X1 U13497 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11307), .ZN(n10888) );
  AOI21_X1 U13498 ( .B1(n15680), .B2(P1_ADDR_REG_2__SCAN_IN), .A(n10888), .ZN(
        n10891) );
  NAND2_X1 U13499 ( .A1(n15720), .A2(n10889), .ZN(n10890) );
  NAND4_X1 U13500 ( .A1(n10893), .A2(n10892), .A3(n10891), .A4(n10890), .ZN(
        n10894) );
  OR2_X1 U13501 ( .A1(n15701), .A2(n10894), .ZN(P1_U3245) );
  AND2_X1 U13502 ( .A1(n15981), .A2(n13139), .ZN(n10895) );
  NAND2_X1 U13503 ( .A1(n10933), .A2(n10895), .ZN(n10897) );
  AND2_X1 U13504 ( .A1(n10908), .A2(n13599), .ZN(n10896) );
  NAND2_X1 U13505 ( .A1(n6543), .A2(n10896), .ZN(n11371) );
  NAND2_X1 U13506 ( .A1(n10897), .A2(n11371), .ZN(n15969) );
  INV_X1 U13507 ( .A(n6543), .ZN(n10898) );
  AND2_X1 U13508 ( .A1(n10898), .A2(n15983), .ZN(n16013) );
  NAND2_X1 U13509 ( .A1(n10899), .A2(n13007), .ZN(n15966) );
  NAND2_X1 U13510 ( .A1(n15967), .A2(n10929), .ZN(n13016) );
  INV_X1 U13511 ( .A(n10929), .ZN(n11553) );
  NAND2_X1 U13512 ( .A1(n10901), .A2(n11553), .ZN(n13015) );
  OAI21_X1 U13513 ( .B1(n10902), .B2(n10907), .A(n11402), .ZN(n11385) );
  NAND2_X1 U13514 ( .A1(n10860), .A2(n15982), .ZN(n10903) );
  AND2_X1 U13515 ( .A1(n15991), .A2(n15972), .ZN(n10906) );
  NAND2_X1 U13516 ( .A1(n11406), .A2(n12976), .ZN(n11455) );
  OAI211_X1 U13517 ( .C1(n11406), .C2(n12976), .A(n11455), .B(n13833), .ZN(
        n10911) );
  INV_X1 U13518 ( .A(n11408), .ZN(n13460) );
  AOI22_X1 U13519 ( .A1(n13830), .A2(n13460), .B1(n13462), .B2(n13828), .ZN(
        n10910) );
  NAND2_X1 U13520 ( .A1(n10911), .A2(n10910), .ZN(n11382) );
  AOI21_X1 U13521 ( .B1(n16007), .B2(n11385), .A(n11382), .ZN(n11556) );
  NAND2_X1 U13522 ( .A1(n10933), .A2(n10912), .ZN(n10913) );
  OAI21_X1 U13523 ( .B1(n10915), .B2(n10914), .A(n10913), .ZN(n10916) );
  NAND2_X1 U13524 ( .A1(n10916), .A2(n11374), .ZN(n10921) );
  INV_X1 U13525 ( .A(n10917), .ZN(n10918) );
  NAND2_X1 U13526 ( .A1(n10919), .A2(n10918), .ZN(n10920) );
  INV_X2 U13527 ( .A(n16018), .ZN(n16017) );
  OAI22_X1 U13528 ( .A1(n11553), .A2(n13997), .B1(n16017), .B2(n8190), .ZN(
        n10922) );
  INV_X1 U13529 ( .A(n10922), .ZN(n10923) );
  OAI21_X1 U13530 ( .B1(n11556), .B2(n16018), .A(n10923), .ZN(P3_U3399) );
  NAND2_X1 U13531 ( .A1(n10924), .A2(n13437), .ZN(n10932) );
  AOI21_X1 U13532 ( .B1(n10853), .B2(n10926), .A(n10925), .ZN(n10931) );
  OAI22_X1 U13533 ( .A1(n13441), .A2(n11408), .B1(n13428), .B2(n15991), .ZN(
        n10928) );
  MUX2_X1 U13534 ( .A(n13443), .B(P3_U3151), .S(P3_REG3_REG_3__SCAN_IN), .Z(
        n10927) );
  AOI211_X1 U13535 ( .C1(n10929), .C2(n13400), .A(n10928), .B(n10927), .ZN(
        n10930) );
  OAI21_X1 U13536 ( .B1(n10932), .B2(n10931), .A(n10930), .ZN(P3_U3158) );
  AOI21_X1 U13537 ( .B1(n10933), .B2(n15981), .A(n13833), .ZN(n10934) );
  OR2_X1 U13538 ( .A1(n12972), .A2(n10934), .ZN(n10936) );
  NAND2_X1 U13539 ( .A1(n8170), .A2(n13830), .ZN(n10935) );
  NAND2_X1 U13540 ( .A1(n10936), .A2(n10935), .ZN(n12676) );
  INV_X1 U13541 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10937) );
  NOR2_X1 U13542 ( .A1(n16017), .A2(n10937), .ZN(n10938) );
  AOI21_X1 U13543 ( .B1(n16017), .B2(n12676), .A(n10938), .ZN(n10939) );
  OAI21_X1 U13544 ( .B1(n11399), .B2(n13997), .A(n10939), .ZN(P3_U3390) );
  INV_X1 U13545 ( .A(n11436), .ZN(n10968) );
  INV_X1 U13546 ( .A(n10940), .ZN(n11437) );
  AND3_X1 U13547 ( .A1(n10968), .A2(n11437), .A3(n11435), .ZN(n10953) );
  INV_X1 U13548 ( .A(n10941), .ZN(n10942) );
  NAND2_X1 U13549 ( .A1(n10944), .A2(n10955), .ZN(n10945) );
  NOR2_X1 U13550 ( .A1(n15813), .A2(n10945), .ZN(n10946) );
  NAND2_X1 U13551 ( .A1(n10953), .A2(n10946), .ZN(n14994) );
  OR2_X1 U13552 ( .A1(n10947), .A2(n13233), .ZN(n10948) );
  NAND2_X1 U13553 ( .A1(n10949), .A2(n10948), .ZN(n10978) );
  OR2_X1 U13554 ( .A1(n13223), .A2(n10950), .ZN(n10952) );
  INV_X1 U13555 ( .A(n11501), .ZN(n15744) );
  NAND2_X1 U13556 ( .A1(n13189), .A2(n15744), .ZN(n10951) );
  NAND2_X1 U13557 ( .A1(n10952), .A2(n10951), .ZN(n10979) );
  XNOR2_X1 U13558 ( .A(n10981), .B(n10979), .ZN(n10977) );
  XOR2_X1 U13559 ( .A(n10978), .B(n10977), .Z(n10964) );
  NAND2_X1 U13560 ( .A1(n10953), .A2(n11438), .ZN(n14989) );
  OR2_X1 U13561 ( .A1(n14989), .A2(n15411), .ZN(n14921) );
  INV_X1 U13562 ( .A(n14921), .ZN(n14983) );
  INV_X1 U13563 ( .A(n10953), .ZN(n10954) );
  NAND2_X1 U13564 ( .A1(n10954), .A2(n11440), .ZN(n10960) );
  AND2_X1 U13565 ( .A1(n10960), .A2(n10955), .ZN(n10974) );
  INV_X1 U13566 ( .A(n10974), .ZN(n14980) );
  NAND2_X1 U13567 ( .A1(n15744), .A2(n15813), .ZN(n15773) );
  INV_X1 U13568 ( .A(n15426), .ZN(n15758) );
  OR2_X1 U13569 ( .A1(n14989), .A2(n15758), .ZN(n14971) );
  OAI22_X1 U13570 ( .A1(n14980), .A2(n15773), .B1(n14971), .B2(n15749), .ZN(
        n10962) );
  AND3_X1 U13571 ( .A1(n10958), .A2(n10957), .A3(n10956), .ZN(n10959) );
  NAND2_X1 U13572 ( .A1(n10960), .A2(n10959), .ZN(n10997) );
  NOR2_X1 U13573 ( .A1(n10997), .A2(P1_U3086), .ZN(n11306) );
  NOR2_X1 U13574 ( .A1(n11306), .A2(n15020), .ZN(n10961) );
  AOI211_X1 U13575 ( .C1(n14983), .C2(n15745), .A(n10962), .B(n10961), .ZN(
        n10963) );
  OAI21_X1 U13576 ( .B1(n14994), .B2(n10964), .A(n10963), .ZN(P1_U3222) );
  INV_X1 U13577 ( .A(n10965), .ZN(n10966) );
  OAI222_X1 U13578 ( .A1(n13599), .A2(P3_U3151), .B1(n14006), .B2(n10967), 
        .C1(n13257), .C2(n10966), .ZN(P3_U3276) );
  INV_X2 U13579 ( .A(n15836), .ZN(n15838) );
  INV_X1 U13580 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10972) );
  OR2_X1 U13581 ( .A1(n10970), .A2(n15836), .ZN(n10971) );
  OAI21_X1 U13582 ( .B1(n15838), .B2(n10972), .A(n10971), .ZN(P1_U3459) );
  AOI22_X1 U13583 ( .A1(n14983), .A2(n15751), .B1(n10973), .B2(n14969), .ZN(
        n10976) );
  NAND2_X1 U13584 ( .A1(n14992), .A2(n8869), .ZN(n10975) );
  OAI211_X1 U13585 ( .C1(n11306), .C2(n11443), .A(n10976), .B(n10975), .ZN(
        P1_U3232) );
  INV_X1 U13586 ( .A(n14992), .ZN(n14963) );
  INV_X1 U13587 ( .A(n10979), .ZN(n10980) );
  NAND2_X1 U13588 ( .A1(n10981), .A2(n10980), .ZN(n10982) );
  NAND2_X1 U13589 ( .A1(n13189), .A2(n15745), .ZN(n10983) );
  OAI21_X1 U13590 ( .B1(n15780), .B2(n13195), .A(n10983), .ZN(n10984) );
  XNOR2_X1 U13591 ( .A(n10984), .B(n13233), .ZN(n10987) );
  OR2_X1 U13592 ( .A1(n13223), .A2(n10985), .ZN(n10986) );
  OAI21_X1 U13593 ( .B1(n15780), .B2(n13224), .A(n10986), .ZN(n10988) );
  XNOR2_X1 U13594 ( .A(n10987), .B(n10988), .ZN(n11304) );
  XNOR2_X1 U13595 ( .A(n10992), .B(n11908), .ZN(n11349) );
  OAI22_X1 U13596 ( .A1(n13223), .A2(n11498), .B1(n11541), .B2(n13224), .ZN(
        n11348) );
  XNOR2_X1 U13597 ( .A(n11349), .B(n11348), .ZN(n10994) );
  AOI21_X1 U13598 ( .B1(n10993), .B2(n10994), .A(n14994), .ZN(n10996) );
  NAND2_X1 U13599 ( .A1(n10996), .A2(n11351), .ZN(n11002) );
  INV_X1 U13600 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n15034) );
  NAND2_X1 U13601 ( .A1(n15746), .A2(n15018), .ZN(n10999) );
  NAND2_X1 U13602 ( .A1(n15426), .A2(n15745), .ZN(n10998) );
  AND2_X1 U13603 ( .A1(n10999), .A2(n10998), .ZN(n11546) );
  OAI22_X1 U13604 ( .A1(n14989), .A2(n11546), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15034), .ZN(n11000) );
  AOI21_X1 U13605 ( .B1(n14928), .B2(n15034), .A(n11000), .ZN(n11001) );
  OAI211_X1 U13606 ( .C1(n11541), .C2(n14963), .A(n11002), .B(n11001), .ZN(
        P1_U3218) );
  INV_X1 U13607 ( .A(n14312), .ZN(n14305) );
  INV_X1 U13608 ( .A(n11003), .ZN(n11005) );
  OAI222_X1 U13609 ( .A1(P2_U3088), .A2(n14305), .B1(n12909), .B2(n11005), 
        .C1(n11004), .C2(n14826), .ZN(P2_U3309) );
  INV_X1 U13610 ( .A(n15137), .ZN(n15131) );
  OAI222_X1 U13611 ( .A1(n15597), .A2(n11006), .B1(n15595), .B2(n11005), .C1(
        n15131), .C2(P1_U3086), .ZN(P1_U3337) );
  XNOR2_X1 U13612 ( .A(n11094), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n11019) );
  MUX2_X1 U13613 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n9502), .S(n14231), .Z(
        n14234) );
  MUX2_X1 U13614 ( .A(n9477), .B(P2_REG1_REG_1__SCAN_IN), .S(n14220), .Z(
        n14227) );
  AND2_X1 U13615 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n14226) );
  NAND2_X1 U13616 ( .A1(n14227), .A2(n14226), .ZN(n14225) );
  NAND2_X1 U13617 ( .A1(n11007), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n11008) );
  NAND2_X1 U13618 ( .A1(n14225), .A2(n11008), .ZN(n14233) );
  NAND2_X1 U13619 ( .A1(n14234), .A2(n14233), .ZN(n14232) );
  NAND2_X1 U13620 ( .A1(n14231), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n11009) );
  NAND2_X1 U13621 ( .A1(n14232), .A2(n11009), .ZN(n15853) );
  MUX2_X1 U13622 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9518), .S(n15855), .Z(
        n15854) );
  NAND2_X1 U13623 ( .A1(n15853), .A2(n15854), .ZN(n15852) );
  NAND2_X1 U13624 ( .A1(n15855), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n11010) );
  NAND2_X1 U13625 ( .A1(n15852), .A2(n11010), .ZN(n14244) );
  MUX2_X1 U13626 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9529), .S(n14246), .Z(
        n14245) );
  NAND2_X1 U13627 ( .A1(n14244), .A2(n14245), .ZN(n14243) );
  NAND2_X1 U13628 ( .A1(n14246), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n11011) );
  NAND2_X1 U13629 ( .A1(n14243), .A2(n11011), .ZN(n15867) );
  MUX2_X1 U13630 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n9541), .S(n15869), .Z(
        n15868) );
  NAND2_X1 U13631 ( .A1(n15867), .A2(n15868), .ZN(n15866) );
  NAND2_X1 U13632 ( .A1(n15869), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n11012) );
  NAND2_X1 U13633 ( .A1(n15866), .A2(n11012), .ZN(n14258) );
  INV_X1 U13634 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n15942) );
  MUX2_X1 U13635 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n15942), .S(n14260), .Z(
        n14259) );
  NAND2_X1 U13636 ( .A1(n14258), .A2(n14259), .ZN(n14257) );
  NAND2_X1 U13637 ( .A1(n14260), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n11013) );
  NAND2_X1 U13638 ( .A1(n14257), .A2(n11013), .ZN(n14270) );
  XNOR2_X1 U13639 ( .A(n14272), .B(n11014), .ZN(n14271) );
  NAND2_X1 U13640 ( .A1(n14270), .A2(n14271), .ZN(n14269) );
  NAND2_X1 U13641 ( .A1(n14272), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n11015) );
  NAND2_X1 U13642 ( .A1(n14269), .A2(n11015), .ZN(n11063) );
  XNOR2_X1 U13643 ( .A(n11059), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n11064) );
  NAND2_X1 U13644 ( .A1(n11063), .A2(n11064), .ZN(n11062) );
  NAND2_X1 U13645 ( .A1(n11042), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n11016) );
  NAND2_X1 U13646 ( .A1(n11062), .A2(n11016), .ZN(n11018) );
  INV_X1 U13647 ( .A(n11096), .ZN(n11017) );
  AOI21_X1 U13648 ( .B1(n11019), .B2(n11018), .A(n11017), .ZN(n11053) );
  INV_X1 U13649 ( .A(n11020), .ZN(n11023) );
  OR2_X1 U13650 ( .A1(n11021), .A2(n11023), .ZN(n11025) );
  OAI21_X1 U13651 ( .B1(n11023), .B2(n11022), .A(n9507), .ZN(n11024) );
  NAND2_X1 U13652 ( .A1(n11025), .A2(n11024), .ZN(n11047) );
  NOR2_X1 U13653 ( .A1(n9478), .A2(P2_U3088), .ZN(n14829) );
  NAND2_X1 U13654 ( .A1(n11047), .A2(n6776), .ZN(n15873) );
  AND2_X1 U13655 ( .A1(n14829), .A2(n11026), .ZN(n11027) );
  NAND2_X1 U13656 ( .A1(n11047), .A2(n11027), .ZN(n14330) );
  MUX2_X1 U13657 ( .A(n11029), .B(P2_REG2_REG_1__SCAN_IN), .S(n14220), .Z(
        n11031) );
  AND2_X1 U13658 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n11030) );
  NAND2_X1 U13659 ( .A1(n11031), .A2(n11030), .ZN(n14224) );
  OAI21_X1 U13660 ( .B1(n11029), .B2(n14220), .A(n14224), .ZN(n14236) );
  NAND2_X1 U13661 ( .A1(n14231), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n11032) );
  MUX2_X1 U13662 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11033), .S(n15855), .Z(
        n15863) );
  NAND2_X1 U13663 ( .A1(n15862), .A2(n15863), .ZN(n15861) );
  NAND2_X1 U13664 ( .A1(n15855), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n14248) );
  NAND2_X1 U13665 ( .A1(n15861), .A2(n14248), .ZN(n11035) );
  INV_X1 U13666 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11995) );
  MUX2_X1 U13667 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n11995), .S(n14246), .Z(
        n11034) );
  NAND2_X1 U13668 ( .A1(n11035), .A2(n11034), .ZN(n14250) );
  NAND2_X1 U13669 ( .A1(n14246), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n11036) );
  NAND2_X1 U13670 ( .A1(n14250), .A2(n11036), .ZN(n15876) );
  MUX2_X1 U13671 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n12185), .S(n15869), .Z(
        n15877) );
  NAND2_X1 U13672 ( .A1(n15876), .A2(n15877), .ZN(n15875) );
  NAND2_X1 U13673 ( .A1(n15869), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n14262) );
  NAND2_X1 U13674 ( .A1(n15875), .A2(n14262), .ZN(n11038) );
  INV_X1 U13675 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11976) );
  MUX2_X1 U13676 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11976), .S(n14260), .Z(
        n11037) );
  NAND2_X1 U13677 ( .A1(n11038), .A2(n11037), .ZN(n14275) );
  NAND2_X1 U13678 ( .A1(n14260), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n14274) );
  NAND2_X1 U13679 ( .A1(n14275), .A2(n14274), .ZN(n11040) );
  INV_X1 U13680 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n12129) );
  MUX2_X1 U13681 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n12129), .S(n14272), .Z(
        n11039) );
  NAND2_X1 U13682 ( .A1(n11040), .A2(n11039), .ZN(n14277) );
  NAND2_X1 U13683 ( .A1(n14272), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n11056) );
  MUX2_X1 U13684 ( .A(n11054), .B(P2_REG2_REG_8__SCAN_IN), .S(n11059), .Z(
        n11041) );
  INV_X1 U13685 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11043) );
  MUX2_X1 U13686 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n11043), .S(n11094), .Z(
        n11045) );
  MUX2_X1 U13687 ( .A(n11043), .B(P2_REG2_REG_9__SCAN_IN), .S(n11094), .Z(
        n11044) );
  OAI21_X1 U13688 ( .B1(n6769), .B2(n11045), .A(n11086), .ZN(n11051) );
  AND2_X1 U13689 ( .A1(n9478), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11046) );
  NAND2_X1 U13690 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n12463) );
  NOR2_X2 U13691 ( .A1(n11047), .A2(P2_U3088), .ZN(n15851) );
  NAND2_X1 U13692 ( .A1(n15851), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n11048) );
  OAI211_X1 U13693 ( .C1(n14306), .C2(n11049), .A(n12463), .B(n11048), .ZN(
        n11050) );
  AOI21_X1 U13694 ( .B1(n15892), .B2(n11051), .A(n11050), .ZN(n11052) );
  OAI21_X1 U13695 ( .B1(n11053), .B2(n15873), .A(n11052), .ZN(P2_U3223) );
  INV_X1 U13696 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11054) );
  MUX2_X1 U13697 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n11054), .S(n11059), .Z(
        n11055) );
  NAND3_X1 U13698 ( .A1(n14277), .A2(n11056), .A3(n11055), .ZN(n11057) );
  AND3_X1 U13699 ( .A1(n15892), .A2(n11058), .A3(n11057), .ZN(n11061) );
  NAND2_X1 U13700 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n12552) );
  OAI21_X1 U13701 ( .B1(n14306), .B2(n11059), .A(n12552), .ZN(n11060) );
  AOI211_X1 U13702 ( .C1(n15851), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n11061), .B(
        n11060), .ZN(n11066) );
  OAI211_X1 U13703 ( .C1(n11064), .C2(n11063), .A(n15896), .B(n11062), .ZN(
        n11065) );
  NAND2_X1 U13704 ( .A1(n11066), .A2(n11065), .ZN(P2_U3222) );
  XNOR2_X1 U13705 ( .A(n11771), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n11072) );
  INV_X1 U13706 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n11070) );
  MUX2_X1 U13707 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n11070), .S(n15054), .Z(
        n15049) );
  AOI21_X1 U13708 ( .B1(n11072), .B2(n11071), .A(n11765), .ZN(n11084) );
  NOR2_X1 U13709 ( .A1(n11073), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14958) );
  NOR2_X1 U13710 ( .A1(n15699), .A2(n11767), .ZN(n11074) );
  AOI211_X1 U13711 ( .C1(n15680), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n14958), 
        .B(n11074), .ZN(n11083) );
  NOR2_X1 U13712 ( .A1(n11075), .A2(n12017), .ZN(n15055) );
  INV_X1 U13713 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n12028) );
  MUX2_X1 U13714 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n12028), .S(n15054), .Z(
        n11076) );
  OAI21_X1 U13715 ( .B1(n15060), .B2(n15055), .A(n11076), .ZN(n15058) );
  NAND2_X1 U13716 ( .A1(n15054), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n11079) );
  INV_X1 U13717 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11077) );
  MUX2_X1 U13718 ( .A(n11077), .B(P1_REG2_REG_11__SCAN_IN), .S(n11771), .Z(
        n11078) );
  AOI21_X1 U13719 ( .B1(n15058), .B2(n11079), .A(n11078), .ZN(n11770) );
  INV_X1 U13720 ( .A(n11770), .ZN(n11081) );
  NAND3_X1 U13721 ( .A1(n15058), .A2(n11079), .A3(n11078), .ZN(n11080) );
  NAND3_X1 U13722 ( .A1(n11081), .A2(n15724), .A3(n11080), .ZN(n11082) );
  OAI211_X1 U13723 ( .C1(n11084), .C2(n15102), .A(n11083), .B(n11082), .ZN(
        P1_U3254) );
  OR2_X1 U13724 ( .A1(n11094), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n11085) );
  NAND2_X1 U13725 ( .A1(n11086), .A2(n11085), .ZN(n11119) );
  INV_X1 U13726 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11087) );
  MUX2_X1 U13727 ( .A(n11087), .B(P2_REG2_REG_10__SCAN_IN), .S(n11114), .Z(
        n11118) );
  NAND2_X1 U13728 ( .A1(n11114), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n11088) );
  INV_X1 U13729 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n12508) );
  MUX2_X1 U13730 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n12508), .S(n11601), .Z(
        n11090) );
  INV_X1 U13731 ( .A(n15889), .ZN(n11089) );
  AOI21_X1 U13732 ( .B1(n11091), .B2(n11090), .A(n11089), .ZN(n11102) );
  AND2_X1 U13733 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n11093) );
  NOR2_X1 U13734 ( .A1(n14306), .A2(n11601), .ZN(n11092) );
  AOI211_X1 U13735 ( .C1(n15851), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n11093), 
        .B(n11092), .ZN(n11101) );
  XNOR2_X1 U13736 ( .A(n11601), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n11099) );
  OR2_X1 U13737 ( .A1(n11094), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n11095) );
  NAND2_X1 U13738 ( .A1(n11096), .A2(n11095), .ZN(n11112) );
  XNOR2_X1 U13739 ( .A(n11114), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n11113) );
  NAND2_X1 U13740 ( .A1(n11114), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n11097) );
  NAND2_X1 U13741 ( .A1(n11110), .A2(n11097), .ZN(n11098) );
  NAND2_X1 U13742 ( .A1(n11098), .A2(n11099), .ZN(n15882) );
  OAI211_X1 U13743 ( .C1(n11099), .C2(n11098), .A(n15882), .B(n15896), .ZN(
        n11100) );
  OAI211_X1 U13744 ( .C1(n11102), .C2(n14330), .A(n11101), .B(n11100), .ZN(
        P2_U3225) );
  AOI21_X1 U13745 ( .B1(n11105), .B2(n11104), .A(n11103), .ZN(n11109) );
  INV_X1 U13746 ( .A(n13428), .ZN(n13439) );
  AOI22_X1 U13747 ( .A1(n13400), .A2(n16006), .B1(n13439), .B2(n10901), .ZN(
        n11106) );
  NAND2_X1 U13748 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n11284) );
  OAI211_X1 U13749 ( .C1(n11664), .C2(n13441), .A(n11106), .B(n11284), .ZN(
        n11107) );
  AOI21_X1 U13750 ( .B1(n11460), .B2(n13443), .A(n11107), .ZN(n11108) );
  OAI21_X1 U13751 ( .B1(n11109), .B2(n13413), .A(n11108), .ZN(P3_U3170) );
  INV_X1 U13752 ( .A(n11110), .ZN(n11111) );
  AOI211_X1 U13753 ( .C1(n11113), .C2(n11112), .A(n15873), .B(n11111), .ZN(
        n11122) );
  INV_X1 U13754 ( .A(n15851), .ZN(n15900) );
  INV_X1 U13755 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n11616) );
  NAND2_X1 U13756 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n12661)
         );
  NAND2_X1 U13757 ( .A1(n15894), .A2(n11114), .ZN(n11115) );
  OAI211_X1 U13758 ( .C1(n15900), .C2(n11616), .A(n12661), .B(n11115), .ZN(
        n11121) );
  INV_X1 U13759 ( .A(n11116), .ZN(n11117) );
  AOI211_X1 U13760 ( .C1(n11119), .C2(n11118), .A(n14330), .B(n11117), .ZN(
        n11120) );
  OR3_X1 U13761 ( .A1(n11122), .A2(n11121), .A3(n11120), .ZN(P2_U3224) );
  INV_X1 U13762 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n11123) );
  MUX2_X1 U13763 ( .A(n11149), .B(n11123), .S(n13576), .Z(n11124) );
  AND2_X1 U13764 ( .A1(n11124), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11170) );
  NAND2_X1 U13765 ( .A1(n11171), .A2(n11170), .ZN(n11275) );
  INV_X1 U13766 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n11143) );
  MUX2_X1 U13767 ( .A(n15979), .B(n11143), .S(n13576), .Z(n11126) );
  INV_X1 U13768 ( .A(n11280), .ZN(n11125) );
  NAND2_X1 U13769 ( .A1(n11126), .A2(n11125), .ZN(n11129) );
  INV_X1 U13770 ( .A(n11126), .ZN(n11127) );
  NAND2_X1 U13771 ( .A1(n11127), .A2(n11280), .ZN(n11128) );
  NAND2_X1 U13772 ( .A1(n11129), .A2(n11128), .ZN(n11274) );
  AOI21_X1 U13773 ( .B1(n11275), .B2(n7334), .A(n11274), .ZN(n11277) );
  INV_X1 U13774 ( .A(n11129), .ZN(n11135) );
  INV_X1 U13775 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n11146) );
  MUX2_X1 U13776 ( .A(n11130), .B(n11146), .S(n13576), .Z(n11131) );
  NAND2_X1 U13777 ( .A1(n11131), .A2(n7100), .ZN(n11296) );
  INV_X1 U13778 ( .A(n11131), .ZN(n11132) );
  NAND2_X1 U13779 ( .A1(n11132), .A2(n11185), .ZN(n11133) );
  AND2_X1 U13780 ( .A1(n11296), .A2(n11133), .ZN(n11134) );
  OAI21_X1 U13781 ( .B1(n11277), .B2(n11135), .A(n11134), .ZN(n11297) );
  NOR3_X1 U13782 ( .A1(n11277), .A2(n11135), .A3(n11134), .ZN(n11136) );
  NAND2_X1 U13783 ( .A1(n13461), .A2(n12879), .ZN(n13622) );
  INV_X1 U13784 ( .A(n13622), .ZN(n13503) );
  OAI21_X1 U13785 ( .B1(n7360), .B2(n11136), .A(n13503), .ZN(n11163) );
  INV_X1 U13786 ( .A(n11139), .ZN(n11137) );
  OR2_X1 U13787 ( .A1(n13124), .A2(n11137), .ZN(n11138) );
  NAND2_X1 U13788 ( .A1(n11138), .A2(n8136), .ZN(n11157) );
  NOR2_X1 U13789 ( .A1(n11139), .A2(P3_U3151), .ZN(n13140) );
  INV_X1 U13790 ( .A(n13140), .ZN(n13145) );
  NAND2_X1 U13791 ( .A1(n13145), .A2(n11140), .ZN(n11156) );
  INV_X1 U13792 ( .A(n11156), .ZN(n11141) );
  INV_X1 U13793 ( .A(n11148), .ZN(n11142) );
  MUX2_X1 U13794 ( .A(P3_U3897), .B(n11142), .S(n12879), .Z(n13615) );
  NAND2_X1 U13795 ( .A1(n11142), .A2(n13576), .ZN(n13612) );
  MUX2_X1 U13796 ( .A(P3_REG1_REG_2__SCAN_IN), .B(n11143), .S(n11280), .Z(
        n11264) );
  NAND2_X1 U13797 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n11165), .ZN(n11144) );
  NAND2_X1 U13798 ( .A1(n11175), .A2(n6615), .ZN(n11263) );
  NAND2_X1 U13799 ( .A1(n11264), .A2(n11263), .ZN(n11262) );
  NAND2_X1 U13800 ( .A1(n11280), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n11145) );
  XNOR2_X1 U13801 ( .A(n11184), .B(n11146), .ZN(n11160) );
  NOR2_X2 U13802 ( .A1(n11148), .A2(n11147), .ZN(n13621) );
  NAND2_X1 U13803 ( .A1(n11177), .A2(n11151), .ZN(n11268) );
  XNOR2_X1 U13804 ( .A(n11280), .B(n15979), .ZN(n11269) );
  NAND2_X1 U13805 ( .A1(n11268), .A2(n11269), .ZN(n11267) );
  NAND2_X1 U13806 ( .A1(n11280), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n11152) );
  NAND2_X1 U13807 ( .A1(n11267), .A2(n11152), .ZN(n11153) );
  OAI21_X1 U13808 ( .B1(P3_REG2_REG_3__SCAN_IN), .B2(n11154), .A(n11289), .ZN(
        n11155) );
  NAND2_X1 U13809 ( .A1(n13621), .A2(n11155), .ZN(n11159) );
  AOI22_X1 U13810 ( .A1(n15945), .A2(P3_ADDR_REG_3__SCAN_IN), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(P3_U3151), .ZN(n11158) );
  OAI211_X1 U13811 ( .C1(n13612), .C2(n11160), .A(n11159), .B(n11158), .ZN(
        n11161) );
  AOI21_X1 U13812 ( .B1(n7100), .B2(n13615), .A(n11161), .ZN(n11162) );
  NAND2_X1 U13813 ( .A1(n11163), .A2(n11162), .ZN(P3_U3185) );
  INV_X1 U13814 ( .A(n13612), .ZN(n13589) );
  NOR3_X1 U13815 ( .A1(n13589), .A2(n13621), .A3(n13503), .ZN(n11169) );
  MUX2_X1 U13816 ( .A(P3_REG2_REG_0__SCAN_IN), .B(P3_REG1_REG_0__SCAN_IN), .S(
        n13576), .Z(n11164) );
  AOI21_X1 U13817 ( .B1(n11165), .B2(n11164), .A(n11170), .ZN(n11168) );
  AOI22_X1 U13818 ( .A1(n15945), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n11167) );
  NAND2_X1 U13819 ( .A1(n13615), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11166) );
  OAI211_X1 U13820 ( .C1(n11169), .C2(n11168), .A(n11167), .B(n11166), .ZN(
        P3_U3182) );
  OAI21_X1 U13821 ( .B1(n11171), .B2(n11170), .A(n11275), .ZN(n11174) );
  INV_X1 U13822 ( .A(n15945), .ZN(n13606) );
  INV_X1 U13823 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n11172) );
  OAI22_X1 U13824 ( .A1(n13606), .A2(n11172), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10057), .ZN(n11173) );
  AOI21_X1 U13825 ( .B1(n13503), .B2(n11174), .A(n11173), .ZN(n11182) );
  OAI21_X1 U13826 ( .B1(P3_REG1_REG_1__SCAN_IN), .B2(n11176), .A(n11175), .ZN(
        n11180) );
  OAI21_X1 U13827 ( .B1(P3_REG2_REG_1__SCAN_IN), .B2(n11178), .A(n11177), .ZN(
        n11179) );
  AOI22_X1 U13828 ( .A1(n13589), .A2(n11180), .B1(n13621), .B2(n11179), .ZN(
        n11181) );
  OAI211_X1 U13829 ( .C1(n11183), .C2(n13586), .A(n11182), .B(n11181), .ZN(
        P3_U3183) );
  INV_X1 U13830 ( .A(n11302), .ZN(n11195) );
  INV_X1 U13831 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n16021) );
  NAND2_X1 U13832 ( .A1(n11184), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n11188) );
  NAND2_X1 U13833 ( .A1(n11186), .A2(n11185), .ZN(n11187) );
  NAND2_X1 U13834 ( .A1(n11188), .A2(n11187), .ZN(n11282) );
  MUX2_X1 U13835 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n16021), .S(n11302), .Z(
        n11283) );
  NAND2_X1 U13836 ( .A1(n11282), .A2(n11283), .ZN(n11281) );
  INV_X1 U13837 ( .A(n11217), .ZN(n11201) );
  INV_X1 U13838 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n11200) );
  XNOR2_X1 U13839 ( .A(n11218), .B(n11200), .ZN(n11212) );
  XNOR2_X1 U13840 ( .A(n11302), .B(n11459), .ZN(n11286) );
  NAND2_X1 U13841 ( .A1(n11189), .A2(n11286), .ZN(n11291) );
  NAND2_X1 U13842 ( .A1(n11302), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n11190) );
  NAND2_X1 U13843 ( .A1(n11291), .A2(n11190), .ZN(n11191) );
  NAND2_X1 U13844 ( .A1(n11191), .A2(n11217), .ZN(n11252) );
  OAI21_X1 U13845 ( .B1(P3_REG2_REG_5__SCAN_IN), .B2(n6778), .A(n11253), .ZN(
        n11210) );
  NAND2_X1 U13846 ( .A1(n13615), .A2(n11201), .ZN(n11193) );
  NAND2_X1 U13847 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n11366) );
  OAI211_X1 U13848 ( .C1(n13606), .C2(n11194), .A(n11193), .B(n11366), .ZN(
        n11209) );
  MUX2_X1 U13849 ( .A(n11459), .B(n16021), .S(n13576), .Z(n11196) );
  NAND2_X1 U13850 ( .A1(n11196), .A2(n11195), .ZN(n11199) );
  INV_X1 U13851 ( .A(n11196), .ZN(n11197) );
  NAND2_X1 U13852 ( .A1(n11197), .A2(n11302), .ZN(n11198) );
  NAND2_X1 U13853 ( .A1(n11199), .A2(n11198), .ZN(n11295) );
  INV_X1 U13854 ( .A(n11199), .ZN(n11206) );
  MUX2_X1 U13855 ( .A(n7583), .B(n11200), .S(n13576), .Z(n11202) );
  NAND2_X1 U13856 ( .A1(n11202), .A2(n11201), .ZN(n11247) );
  INV_X1 U13857 ( .A(n11202), .ZN(n11203) );
  NAND2_X1 U13858 ( .A1(n11203), .A2(n11217), .ZN(n11204) );
  AND2_X1 U13859 ( .A1(n11247), .A2(n11204), .ZN(n11205) );
  OR3_X1 U13860 ( .A1(n11299), .A2(n11206), .A3(n11205), .ZN(n11207) );
  AOI21_X1 U13861 ( .B1(n11248), .B2(n11207), .A(n13622), .ZN(n11208) );
  AOI211_X1 U13862 ( .C1(n13621), .C2(n11210), .A(n11209), .B(n11208), .ZN(
        n11211) );
  OAI21_X1 U13863 ( .B1(n11212), .B2(n13612), .A(n11211), .ZN(P3_U3187) );
  INV_X1 U13864 ( .A(n11213), .ZN(n11215) );
  OAI22_X1 U13865 ( .A1(n6543), .A2(P3_U3151), .B1(SI_22_), .B2(n14006), .ZN(
        n11214) );
  AOI21_X1 U13866 ( .B1(n11215), .B2(n13999), .A(n11214), .ZN(P3_U3273) );
  INV_X1 U13867 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n11219) );
  MUX2_X1 U13868 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n11219), .S(n11258), .Z(
        n11245) );
  INV_X1 U13869 ( .A(n11327), .ZN(n11225) );
  INV_X1 U13870 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11642) );
  XNOR2_X1 U13871 ( .A(n11328), .B(n11642), .ZN(n11241) );
  MUX2_X1 U13872 ( .A(n15962), .B(n11219), .S(n13576), .Z(n11220) );
  NAND2_X1 U13873 ( .A1(n11220), .A2(n11258), .ZN(n11224) );
  INV_X1 U13874 ( .A(n11220), .ZN(n11222) );
  NAND2_X1 U13875 ( .A1(n11222), .A2(n11221), .ZN(n11223) );
  NAND2_X1 U13876 ( .A1(n11224), .A2(n11223), .ZN(n11246) );
  INV_X1 U13877 ( .A(n11224), .ZN(n11230) );
  MUX2_X1 U13878 ( .A(n7586), .B(n11642), .S(n13576), .Z(n11226) );
  NAND2_X1 U13879 ( .A1(n11226), .A2(n11225), .ZN(n11333) );
  INV_X1 U13880 ( .A(n11226), .ZN(n11227) );
  NAND2_X1 U13881 ( .A1(n11227), .A2(n11327), .ZN(n11228) );
  AND2_X1 U13882 ( .A1(n11333), .A2(n11228), .ZN(n11229) );
  INV_X1 U13883 ( .A(n11334), .ZN(n11232) );
  NOR3_X1 U13884 ( .A1(n11250), .A2(n11230), .A3(n11229), .ZN(n11231) );
  OAI21_X1 U13885 ( .B1(n11232), .B2(n11231), .A(n13503), .ZN(n11240) );
  OR2_X1 U13886 ( .A1(n11258), .A2(n15962), .ZN(n11233) );
  OAI21_X1 U13887 ( .B1(P3_REG2_REG_7__SCAN_IN), .B2(n6767), .A(n11338), .ZN(
        n11238) );
  AND2_X1 U13888 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n12058) );
  AOI21_X1 U13889 ( .B1(n15945), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n12058), .ZN(
        n11236) );
  OAI21_X1 U13890 ( .B1(n13586), .B2(n11327), .A(n11236), .ZN(n11237) );
  AOI21_X1 U13891 ( .B1(n11238), .B2(n13621), .A(n11237), .ZN(n11239) );
  OAI211_X1 U13892 ( .C1(n11241), .C2(n13612), .A(n11240), .B(n11239), .ZN(
        P3_U3189) );
  INV_X1 U13893 ( .A(n11242), .ZN(n11243) );
  AOI21_X1 U13894 ( .B1(n11245), .B2(n11244), .A(n11243), .ZN(n11261) );
  AND3_X1 U13895 ( .A1(n11248), .A2(n11247), .A3(n11246), .ZN(n11249) );
  OAI21_X1 U13896 ( .B1(n11250), .B2(n11249), .A(n13503), .ZN(n11260) );
  AND2_X1 U13897 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n11663) );
  INV_X1 U13898 ( .A(n11663), .ZN(n11251) );
  OAI21_X1 U13899 ( .B1(n13606), .B2(n10822), .A(n11251), .ZN(n11257) );
  NAND3_X1 U13900 ( .A1(n11253), .A2(n6781), .A3(n11252), .ZN(n11254) );
  INV_X1 U13901 ( .A(n13621), .ZN(n12143) );
  AOI21_X1 U13902 ( .B1(n11255), .B2(n11254), .A(n12143), .ZN(n11256) );
  AOI211_X1 U13903 ( .C1(n13615), .C2(n11258), .A(n11257), .B(n11256), .ZN(
        n11259) );
  OAI211_X1 U13904 ( .C1(n11261), .C2(n13612), .A(n11260), .B(n11259), .ZN(
        P3_U3188) );
  OAI21_X1 U13905 ( .B1(n11264), .B2(n11263), .A(n11262), .ZN(n11273) );
  NAND2_X1 U13906 ( .A1(n15945), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n11265) );
  OAI21_X1 U13907 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n11266), .A(n11265), .ZN(
        n11272) );
  OAI21_X1 U13908 ( .B1(n11269), .B2(n11268), .A(n11267), .ZN(n11270) );
  AND2_X1 U13909 ( .A1(n13621), .A2(n11270), .ZN(n11271) );
  AOI211_X1 U13910 ( .C1(n13589), .C2(n11273), .A(n11272), .B(n11271), .ZN(
        n11279) );
  AND3_X1 U13911 ( .A1(n11275), .A2(n7334), .A3(n11274), .ZN(n11276) );
  OAI21_X1 U13912 ( .B1(n11277), .B2(n11276), .A(n13503), .ZN(n11278) );
  OAI211_X1 U13913 ( .C1(n13586), .C2(n11280), .A(n11279), .B(n11278), .ZN(
        P3_U3184) );
  OAI21_X1 U13914 ( .B1(n11283), .B2(n11282), .A(n11281), .ZN(n11294) );
  OAI21_X1 U13915 ( .B1(n13606), .B2(n11285), .A(n11284), .ZN(n11293) );
  INV_X1 U13916 ( .A(n11286), .ZN(n11288) );
  NAND3_X1 U13917 ( .A1(n11289), .A2(n11288), .A3(n11287), .ZN(n11290) );
  AOI21_X1 U13918 ( .B1(n11291), .B2(n11290), .A(n12143), .ZN(n11292) );
  AOI211_X1 U13919 ( .C1(n13589), .C2(n11294), .A(n11293), .B(n11292), .ZN(
        n11301) );
  AND3_X1 U13920 ( .A1(n11297), .A2(n11296), .A3(n11295), .ZN(n11298) );
  OAI21_X1 U13921 ( .B1(n11299), .B2(n11298), .A(n13503), .ZN(n11300) );
  OAI211_X1 U13922 ( .C1(n13586), .C2(n11302), .A(n11301), .B(n11300), .ZN(
        P3_U3186) );
  XOR2_X1 U13923 ( .A(n11303), .B(n11304), .Z(n11310) );
  INV_X1 U13924 ( .A(n14971), .ZN(n14978) );
  AOI22_X1 U13925 ( .A1(n14978), .A2(n15751), .B1(n14983), .B2(n15425), .ZN(
        n11305) );
  OAI21_X1 U13926 ( .B1(n11307), .B2(n11306), .A(n11305), .ZN(n11308) );
  AOI21_X1 U13927 ( .B1(n14992), .B2(n15439), .A(n11308), .ZN(n11309) );
  OAI21_X1 U13928 ( .B1(n11310), .B2(n14994), .A(n11309), .ZN(P1_U3237) );
  OAI222_X1 U13929 ( .A1(n14826), .A2(n11311), .B1(P2_U3088), .B2(n9853), .C1(
        n14832), .C2(n12824), .ZN(P2_U3307) );
  NAND2_X1 U13930 ( .A1(n11315), .A2(n11312), .ZN(n11313) );
  INV_X1 U13931 ( .A(n11315), .ZN(n11316) );
  NAND2_X1 U13932 ( .A1(n11316), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n11317) );
  NAND2_X1 U13933 ( .A1(n11320), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n11321) );
  INV_X1 U13934 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n11562) );
  XNOR2_X1 U13935 ( .A(n11562), .B(P1_ADDR_REG_10__SCAN_IN), .ZN(n11619) );
  INV_X1 U13936 ( .A(n11619), .ZN(n11322) );
  NAND2_X1 U13937 ( .A1(n11618), .A2(n11617), .ZN(n11325) );
  XNOR2_X1 U13938 ( .A(n11325), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  XNOR2_X1 U13939 ( .A(n11464), .B(n11740), .ZN(n11465) );
  XOR2_X1 U13940 ( .A(n11466), .B(n11465), .Z(n11345) );
  INV_X1 U13941 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11729) );
  MUX2_X1 U13942 ( .A(n11729), .B(n11740), .S(n13576), .Z(n11329) );
  NAND2_X1 U13943 ( .A1(n11329), .A2(n11464), .ZN(n11471) );
  INV_X1 U13944 ( .A(n11329), .ZN(n11330) );
  NAND2_X1 U13945 ( .A1(n11330), .A2(n11467), .ZN(n11331) );
  NAND2_X1 U13946 ( .A1(n11471), .A2(n11331), .ZN(n11332) );
  AOI21_X1 U13947 ( .B1(n11334), .B2(n11333), .A(n11332), .ZN(n11477) );
  INV_X1 U13948 ( .A(n11477), .ZN(n11336) );
  NAND3_X1 U13949 ( .A1(n11334), .A2(n11333), .A3(n11332), .ZN(n11335) );
  AOI21_X1 U13950 ( .B1(n11336), .B2(n11335), .A(n13622), .ZN(n11343) );
  NAND3_X1 U13951 ( .A1(n11338), .A2(n6779), .A3(n11337), .ZN(n11339) );
  AOI21_X1 U13952 ( .B1(n11469), .B2(n11339), .A(n12143), .ZN(n11342) );
  AND2_X1 U13953 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n11847) );
  AOI21_X1 U13954 ( .B1(n15945), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11847), .ZN(
        n11340) );
  OAI21_X1 U13955 ( .B1(n13586), .B2(n11467), .A(n11340), .ZN(n11341) );
  NOR3_X1 U13956 ( .A1(n11343), .A2(n11342), .A3(n11341), .ZN(n11344) );
  OAI21_X1 U13957 ( .B1(n11345), .B2(n13612), .A(n11344), .ZN(P3_U3190) );
  INV_X1 U13958 ( .A(n11346), .ZN(n11400) );
  OAI222_X1 U13959 ( .A1(n15597), .A2(n11347), .B1(n15595), .B2(n11400), .C1(
        n6539), .C2(P1_U3086), .ZN(P1_U3336) );
  NAND2_X1 U13960 ( .A1(n11349), .A2(n11348), .ZN(n11350) );
  OAI22_X1 U13961 ( .A1(n11521), .A2(n13195), .B1(n11524), .B2(n13224), .ZN(
        n11352) );
  XNOR2_X1 U13962 ( .A(n11352), .B(n11908), .ZN(n11645) );
  NAND2_X1 U13963 ( .A1(n13235), .A2(n15018), .ZN(n11353) );
  OAI21_X1 U13964 ( .B1(n11521), .B2(n13224), .A(n11353), .ZN(n11646) );
  XNOR2_X1 U13965 ( .A(n11645), .B(n11646), .ZN(n11354) );
  XNOR2_X1 U13966 ( .A(n11644), .B(n11354), .ZN(n11361) );
  NAND2_X1 U13967 ( .A1(n11525), .A2(n15813), .ZN(n15795) );
  INV_X1 U13968 ( .A(n14989), .ZN(n14960) );
  NAND2_X1 U13969 ( .A1(n15746), .A2(n15017), .ZN(n11356) );
  NAND2_X1 U13970 ( .A1(n15426), .A2(n15425), .ZN(n11355) );
  NAND2_X1 U13971 ( .A1(n11356), .A2(n11355), .ZN(n11510) );
  AOI22_X1 U13972 ( .A1(n14960), .A2(n11510), .B1(P1_REG3_REG_4__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11359) );
  INV_X1 U13973 ( .A(n11357), .ZN(n11515) );
  NAND2_X1 U13974 ( .A1(n14928), .A2(n11515), .ZN(n11358) );
  OAI211_X1 U13975 ( .C1(n14980), .C2(n15795), .A(n11359), .B(n11358), .ZN(
        n11360) );
  AOI21_X1 U13976 ( .B1(n11361), .B2(n14969), .A(n11360), .ZN(n11362) );
  INV_X1 U13977 ( .A(n11362), .ZN(P1_U3230) );
  AOI21_X1 U13978 ( .B1(n11365), .B2(n11364), .A(n11363), .ZN(n11370) );
  AOI22_X1 U13979 ( .A1(n13400), .A2(n16012), .B1(n13439), .B2(n13460), .ZN(
        n11367) );
  OAI211_X1 U13980 ( .C1(n12059), .C2(n13441), .A(n11367), .B(n11366), .ZN(
        n11368) );
  AOI21_X1 U13981 ( .B1(n11416), .B2(n13443), .A(n11368), .ZN(n11369) );
  OAI21_X1 U13982 ( .B1(n11370), .B2(n13413), .A(n11369), .ZN(P3_U3167) );
  AND2_X1 U13983 ( .A1(n13124), .A2(n11371), .ZN(n11378) );
  INV_X1 U13984 ( .A(n11387), .ZN(n11392) );
  MUX2_X1 U13985 ( .A(n7391), .B(n11371), .S(n13124), .Z(n11388) );
  NAND2_X1 U13986 ( .A1(n11388), .A2(n11392), .ZN(n11377) );
  XNOR2_X1 U13987 ( .A(n11372), .B(n11387), .ZN(n11376) );
  AND2_X1 U13988 ( .A1(n11374), .A2(n11373), .ZN(n11375) );
  OAI211_X1 U13989 ( .C1(n11378), .C2(n11392), .A(n11377), .B(n11395), .ZN(
        n11381) );
  AND2_X2 U13990 ( .A1(n11381), .A2(n15985), .ZN(n15997) );
  AND2_X1 U13991 ( .A1(n15983), .A2(n8546), .ZN(n11403) );
  OR2_X1 U13992 ( .A1(n15969), .A2(n11403), .ZN(n15994) );
  INV_X1 U13993 ( .A(n15994), .ZN(n15956) );
  INV_X1 U13994 ( .A(n15981), .ZN(n16011) );
  INV_X1 U13995 ( .A(n15983), .ZN(n11379) );
  NAND2_X1 U13996 ( .A1(n16011), .A2(n11379), .ZN(n11380) );
  NOR2_X2 U13997 ( .A1(n11381), .A2(n11380), .ZN(n15958) );
  OAI22_X1 U13998 ( .A1(n13825), .A2(n11553), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n15985), .ZN(n11384) );
  MUX2_X1 U13999 ( .A(n11382), .B(P3_REG2_REG_3__SCAN_IN), .S(n15997), .Z(
        n11383) );
  AOI211_X1 U14000 ( .C1(n13837), .C2(n11385), .A(n11384), .B(n11383), .ZN(
        n11386) );
  INV_X1 U14001 ( .A(n11386), .ZN(P3_U3230) );
  NAND2_X1 U14002 ( .A1(n11388), .A2(n11387), .ZN(n11396) );
  OAI211_X1 U14003 ( .C1(n11390), .C2(n6543), .A(n11389), .B(n7391), .ZN(
        n11391) );
  NAND2_X1 U14004 ( .A1(n11391), .A2(n13124), .ZN(n11393) );
  NAND2_X1 U14005 ( .A1(n11393), .A2(n11392), .ZN(n11394) );
  INV_X2 U14006 ( .A(n16023), .ZN(n13911) );
  NOR2_X1 U14007 ( .A1(n13911), .A2(n11123), .ZN(n11397) );
  AOI21_X1 U14008 ( .B1(n13911), .B2(n12676), .A(n11397), .ZN(n11398) );
  OAI21_X1 U14009 ( .B1(n11399), .B2(n13905), .A(n11398), .ZN(P3_U3459) );
  INV_X1 U14010 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11401) );
  OAI222_X1 U14011 ( .A1(n14826), .A2(n11401), .B1(P2_U3088), .B2(n14332), 
        .C1(n14832), .C2(n11400), .ZN(P2_U3308) );
  NAND2_X1 U14012 ( .A1(n11408), .A2(n16006), .ZN(n13022) );
  NAND2_X1 U14013 ( .A1(n13460), .A2(n11407), .ZN(n13023) );
  AND2_X2 U14014 ( .A1(n13022), .A2(n13023), .ZN(n13019) );
  NAND2_X1 U14015 ( .A1(n11453), .A2(n13019), .ZN(n11452) );
  NAND2_X1 U14016 ( .A1(n11664), .A2(n16012), .ZN(n13028) );
  INV_X1 U14017 ( .A(n11664), .ZN(n13459) );
  INV_X1 U14018 ( .A(n16012), .ZN(n11425) );
  NAND2_X1 U14019 ( .A1(n13459), .A2(n11425), .ZN(n13027) );
  XNOR2_X1 U14020 ( .A(n11421), .B(n13025), .ZN(n16014) );
  INV_X1 U14021 ( .A(n16014), .ZN(n11420) );
  INV_X1 U14022 ( .A(n11403), .ZN(n15974) );
  NOR2_X1 U14023 ( .A1(n15997), .A2(n15974), .ZN(n13714) );
  INV_X1 U14024 ( .A(n13714), .ZN(n11419) );
  NAND2_X1 U14025 ( .A1(n16014), .A2(n15969), .ZN(n11415) );
  OAI22_X1 U14026 ( .A1(n11408), .A2(n15990), .B1(n12059), .B2(n15992), .ZN(
        n11404) );
  INV_X1 U14027 ( .A(n11404), .ZN(n11414) );
  INV_X1 U14028 ( .A(n13019), .ZN(n11405) );
  NAND3_X1 U14029 ( .A1(n11406), .A2(n11405), .A3(n12976), .ZN(n11411) );
  OR2_X1 U14030 ( .A1(n15967), .A2(n11553), .ZN(n11454) );
  OAI22_X1 U14031 ( .A1(n13019), .A2(n11454), .B1(n11408), .B2(n11407), .ZN(
        n11409) );
  INV_X1 U14032 ( .A(n11409), .ZN(n11410) );
  NAND2_X1 U14033 ( .A1(n11411), .A2(n11410), .ZN(n11426) );
  NOR2_X1 U14034 ( .A1(n11426), .A2(n13025), .ZN(n11586) );
  AND2_X1 U14035 ( .A1(n11426), .A2(n13025), .ZN(n11412) );
  OAI21_X1 U14036 ( .B1(n11586), .B2(n11412), .A(n13833), .ZN(n11413) );
  AND3_X1 U14037 ( .A1(n11415), .A2(n11414), .A3(n11413), .ZN(n16016) );
  INV_X2 U14038 ( .A(n15997), .ZN(n15995) );
  MUX2_X1 U14039 ( .A(n7583), .B(n16016), .S(n15995), .Z(n11418) );
  AOI22_X1 U14040 ( .A1(n15958), .A2(n16012), .B1(n15977), .B2(n11416), .ZN(
        n11417) );
  OAI211_X1 U14041 ( .C1(n11420), .C2(n11419), .A(n11418), .B(n11417), .ZN(
        P3_U3228) );
  NAND2_X1 U14042 ( .A1(n11421), .A2(n13025), .ZN(n11422) );
  NAND2_X1 U14043 ( .A1(n12059), .A2(n15959), .ZN(n13034) );
  INV_X1 U14044 ( .A(n12059), .ZN(n13458) );
  NAND2_X1 U14045 ( .A1(n11631), .A2(n13034), .ZN(n11424) );
  NAND2_X1 U14046 ( .A1(n11851), .A2(n15950), .ZN(n13039) );
  INV_X1 U14047 ( .A(n15950), .ZN(n12062) );
  NAND2_X1 U14048 ( .A1(n13457), .A2(n12062), .ZN(n13038) );
  NAND2_X1 U14049 ( .A1(n11424), .A2(n13037), .ZN(n11423) );
  OAI21_X1 U14050 ( .B1(n11424), .B2(n13037), .A(n11423), .ZN(n15947) );
  AND2_X1 U14051 ( .A1(n11664), .A2(n11425), .ZN(n11585) );
  NAND2_X1 U14052 ( .A1(n11426), .A2(n11427), .ZN(n11428) );
  OAI211_X1 U14053 ( .C1(n11430), .C2(n11429), .A(n11634), .B(n13833), .ZN(
        n11432) );
  AOI22_X1 U14054 ( .A1(n13458), .A2(n13828), .B1(n13830), .B2(n13456), .ZN(
        n11431) );
  NAND2_X1 U14055 ( .A1(n11432), .A2(n11431), .ZN(n15946) );
  AOI21_X1 U14056 ( .B1(n15947), .B2(n16007), .A(n15946), .ZN(n11641) );
  AOI22_X1 U14057 ( .A1(n13981), .A2(n15950), .B1(P3_REG0_REG_7__SCAN_IN), 
        .B2(n16018), .ZN(n11433) );
  OAI21_X1 U14058 ( .B1(n11641), .B2(n16018), .A(n11433), .ZN(P3_U3411) );
  INV_X1 U14059 ( .A(n11434), .ZN(n11442) );
  NAND4_X1 U14060 ( .A1(n11438), .A2(n11437), .A3(n11436), .A4(n11435), .ZN(
        n15180) );
  AND2_X2 U14061 ( .A1(n15180), .A2(n15393), .ZN(n15764) );
  NOR2_X1 U14062 ( .A1(n11441), .A2(n15598), .ZN(n15743) );
  AOI21_X1 U14063 ( .B1(n11442), .B2(n6544), .A(n15730), .ZN(n11451) );
  OAI22_X1 U14064 ( .A1(n6544), .A2(n8838), .B1(n11443), .B2(n15393), .ZN(
        n11444) );
  AOI21_X1 U14065 ( .B1(n11445), .B2(n6544), .A(n11444), .ZN(n11450) );
  NAND2_X1 U14066 ( .A1(n6544), .A2(n15754), .ZN(n15333) );
  INV_X1 U14067 ( .A(n15333), .ZN(n15313) );
  INV_X1 U14068 ( .A(n11447), .ZN(n11448) );
  OAI21_X1 U14069 ( .B1(n15313), .B2(n15383), .A(n11448), .ZN(n11449) );
  OAI211_X1 U14070 ( .C1(n11451), .C2(n11502), .A(n11450), .B(n11449), .ZN(
        P1_U3293) );
  OAI21_X1 U14071 ( .B1(n11453), .B2(n13019), .A(n11452), .ZN(n16008) );
  INV_X1 U14072 ( .A(n16008), .ZN(n11463) );
  NAND2_X1 U14073 ( .A1(n11455), .A2(n11454), .ZN(n11456) );
  XNOR2_X1 U14074 ( .A(n11456), .B(n13019), .ZN(n11458) );
  OAI22_X1 U14075 ( .A1(n15967), .A2(n15990), .B1(n11664), .B2(n15992), .ZN(
        n11457) );
  AOI21_X1 U14076 ( .B1(n11458), .B2(n13833), .A(n11457), .ZN(n16010) );
  MUX2_X1 U14077 ( .A(n11459), .B(n16010), .S(n15995), .Z(n11462) );
  AOI22_X1 U14078 ( .A1(n15958), .A2(n16006), .B1(n15977), .B2(n11460), .ZN(
        n11461) );
  OAI211_X1 U14079 ( .C1(n11463), .C2(n13807), .A(n11462), .B(n11461), .ZN(
        P3_U3229) );
  XNOR2_X1 U14080 ( .A(n11561), .B(P3_REG1_REG_9__SCAN_IN), .ZN(n11487) );
  NAND2_X1 U14081 ( .A1(n11467), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n11468) );
  NAND2_X1 U14082 ( .A1(n11469), .A2(n11468), .ZN(n11470) );
  INV_X1 U14083 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11840) );
  OAI21_X1 U14084 ( .B1(n6768), .B2(P3_REG2_REG_9__SCAN_IN), .A(n11576), .ZN(
        n11485) );
  INV_X1 U14085 ( .A(n11471), .ZN(n11476) );
  INV_X1 U14086 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11560) );
  MUX2_X1 U14087 ( .A(n11840), .B(n11560), .S(n13576), .Z(n11472) );
  INV_X1 U14088 ( .A(n11483), .ZN(n11559) );
  NAND2_X1 U14089 ( .A1(n11472), .A2(n11559), .ZN(n11567) );
  INV_X1 U14090 ( .A(n11472), .ZN(n11473) );
  NAND2_X1 U14091 ( .A1(n11473), .A2(n11483), .ZN(n11474) );
  AND2_X1 U14092 ( .A1(n11567), .A2(n11474), .ZN(n11475) );
  OAI21_X1 U14093 ( .B1(n11477), .B2(n11476), .A(n11475), .ZN(n11568) );
  INV_X1 U14094 ( .A(n11568), .ZN(n11479) );
  NOR3_X1 U14095 ( .A1(n11477), .A2(n11476), .A3(n11475), .ZN(n11478) );
  OAI21_X1 U14096 ( .B1(n11479), .B2(n11478), .A(n13503), .ZN(n11482) );
  NOR2_X1 U14097 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11480), .ZN(n12196) );
  AOI21_X1 U14098 ( .B1(n15945), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n12196), .ZN(
        n11481) );
  OAI211_X1 U14099 ( .C1(n13586), .C2(n11483), .A(n11482), .B(n11481), .ZN(
        n11484) );
  AOI21_X1 U14100 ( .B1(n13621), .B2(n11485), .A(n11484), .ZN(n11486) );
  OAI21_X1 U14101 ( .B1(n11487), .B2(n13612), .A(n11486), .ZN(P3_U3191) );
  INV_X1 U14102 ( .A(n11488), .ZN(n11489) );
  OAI222_X1 U14103 ( .A1(n11492), .A2(P3_U3151), .B1(n14006), .B2(n11490), 
        .C1(n13257), .C2(n11489), .ZN(P3_U3275) );
  NAND2_X1 U14104 ( .A1(n15750), .A2(n15738), .ZN(n11494) );
  OR2_X1 U14105 ( .A1(n15751), .A2(n15744), .ZN(n11493) );
  NAND2_X1 U14106 ( .A1(n11494), .A2(n11493), .ZN(n15424) );
  NAND2_X1 U14107 ( .A1(n15424), .A2(n11495), .ZN(n11497) );
  NAND2_X1 U14108 ( .A1(n11497), .A2(n11496), .ZN(n11538) );
  INV_X1 U14109 ( .A(n11539), .ZN(n11545) );
  NAND2_X1 U14110 ( .A1(n11538), .A2(n11545), .ZN(n11500) );
  NAND2_X1 U14111 ( .A1(n11541), .A2(n11498), .ZN(n11499) );
  NAND2_X2 U14112 ( .A1(n11500), .A2(n11499), .ZN(n11519) );
  XOR2_X1 U14113 ( .A(n11509), .B(n11519), .Z(n15797) );
  NAND2_X1 U14114 ( .A1(n15739), .A2(n15780), .ZN(n15435) );
  INV_X1 U14115 ( .A(n11533), .ZN(n11503) );
  AOI211_X1 U14116 ( .C1(n11525), .C2(n6906), .A(n15742), .B(n11503), .ZN(
        n15794) );
  NAND2_X1 U14117 ( .A1(n15427), .A2(n11506), .ZN(n11544) );
  NAND2_X1 U14118 ( .A1(n11544), .A2(n11539), .ZN(n11508) );
  NAND2_X1 U14119 ( .A1(n11508), .A2(n11507), .ZN(n11523) );
  XNOR2_X1 U14120 ( .A(n11523), .B(n11509), .ZN(n11512) );
  INV_X1 U14121 ( .A(n11510), .ZN(n11511) );
  OAI21_X1 U14122 ( .B1(n11512), .B2(n15829), .A(n11511), .ZN(n15798) );
  AOI21_X1 U14123 ( .B1(n15794), .B2(n6539), .A(n15798), .ZN(n11513) );
  MUX2_X1 U14124 ( .A(n11514), .B(n11513), .S(n6544), .Z(n11517) );
  INV_X1 U14125 ( .A(n15393), .ZN(n15760) );
  AOI22_X1 U14126 ( .A1(n15730), .A2(n11525), .B1(n15760), .B2(n11515), .ZN(
        n11516) );
  OAI211_X1 U14127 ( .C1(n15423), .C2(n15797), .A(n11517), .B(n11516), .ZN(
        P1_U3289) );
  NOR2_X1 U14128 ( .A1(n11525), .A2(n15018), .ZN(n11518) );
  NOR2_X1 U14129 ( .A1(n11748), .A2(n11709), .ZN(n11707) );
  AOI21_X1 U14130 ( .B1(n11709), .B2(n11748), .A(n11707), .ZN(n15802) );
  NAND2_X1 U14131 ( .A1(n11521), .A2(n15018), .ZN(n11522) );
  NAND2_X1 U14132 ( .A1(n11523), .A2(n11522), .ZN(n11527) );
  NAND2_X1 U14133 ( .A1(n11525), .A2(n11524), .ZN(n11526) );
  XOR2_X1 U14134 ( .A(n11710), .B(n11709), .Z(n11528) );
  NOR2_X1 U14135 ( .A1(n11528), .A2(n15829), .ZN(n15808) );
  NAND2_X1 U14136 ( .A1(n15016), .A2(n15746), .ZN(n11530) );
  NAND2_X1 U14137 ( .A1(n15426), .A2(n15018), .ZN(n11529) );
  NAND2_X1 U14138 ( .A1(n11530), .A2(n11529), .ZN(n15803) );
  NOR2_X1 U14139 ( .A1(n15808), .A2(n15803), .ZN(n11531) );
  MUX2_X1 U14140 ( .A(n10689), .B(n11531), .S(n6544), .Z(n11537) );
  AOI211_X1 U14141 ( .C1(n11742), .C2(n11533), .A(n15742), .B(n11532), .ZN(
        n15807) );
  NOR2_X2 U14142 ( .A1(n15180), .A2(n15748), .ZN(n15732) );
  OAI22_X1 U14143 ( .A1(n15418), .A2(n11534), .B1(n15393), .B2(n11653), .ZN(
        n11535) );
  AOI21_X1 U14144 ( .B1(n15807), .B2(n15732), .A(n11535), .ZN(n11536) );
  OAI211_X1 U14145 ( .C1(n15423), .C2(n15802), .A(n11537), .B(n11536), .ZN(
        P1_U3288) );
  XNOR2_X1 U14146 ( .A(n11538), .B(n11539), .ZN(n15788) );
  AOI211_X1 U14147 ( .C1(n15786), .C2(n15435), .A(n15742), .B(n11540), .ZN(
        n15785) );
  NOR2_X1 U14148 ( .A1(n15418), .A2(n11541), .ZN(n11543) );
  OAI22_X1 U14149 ( .A1(n6544), .A2(n7249), .B1(n15393), .B2(
        P1_REG3_REG_3__SCAN_IN), .ZN(n11542) );
  AOI211_X1 U14150 ( .C1(n15785), .C2(n15732), .A(n11543), .B(n11542), .ZN(
        n11549) );
  XNOR2_X1 U14151 ( .A(n11544), .B(n11545), .ZN(n11547) );
  OAI21_X1 U14152 ( .B1(n11547), .B2(n15829), .A(n11546), .ZN(n15790) );
  NAND2_X1 U14153 ( .A1(n15790), .A2(n6544), .ZN(n11548) );
  OAI211_X1 U14154 ( .C1(n15423), .C2(n15788), .A(n11549), .B(n11548), .ZN(
        P1_U3290) );
  INV_X1 U14155 ( .A(n11550), .ZN(n12748) );
  OAI222_X1 U14156 ( .A1(n14826), .A2(n11552), .B1(n12909), .B2(n12748), .C1(
        n11551), .C2(P2_U3088), .ZN(P2_U3306) );
  OAI22_X1 U14157 ( .A1(n13905), .A2(n11553), .B1(n13911), .B2(n11146), .ZN(
        n11554) );
  INV_X1 U14158 ( .A(n11554), .ZN(n11555) );
  OAI21_X1 U14159 ( .B1(n11556), .B2(n16023), .A(n11555), .ZN(P3_U3462) );
  INV_X1 U14160 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11815) );
  XNOR2_X1 U14161 ( .A(n11885), .B(n11815), .ZN(n11886) );
  INV_X1 U14162 ( .A(n11557), .ZN(n11558) );
  XOR2_X1 U14163 ( .A(n11887), .B(n11886), .Z(n11583) );
  INV_X1 U14164 ( .A(n11885), .ZN(n11573) );
  NAND2_X1 U14165 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n13301)
         );
  OAI21_X1 U14166 ( .B1(n13606), .B2(n11562), .A(n13301), .ZN(n11572) );
  INV_X1 U14167 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11574) );
  MUX2_X1 U14168 ( .A(n11574), .B(n11815), .S(n13576), .Z(n11563) );
  NAND2_X1 U14169 ( .A1(n11563), .A2(n11573), .ZN(n11876) );
  INV_X1 U14170 ( .A(n11563), .ZN(n11564) );
  NAND2_X1 U14171 ( .A1(n11564), .A2(n11885), .ZN(n11565) );
  NAND2_X1 U14172 ( .A1(n11876), .A2(n11565), .ZN(n11566) );
  AOI21_X1 U14173 ( .B1(n11568), .B2(n11567), .A(n11566), .ZN(n11878) );
  INV_X1 U14174 ( .A(n11878), .ZN(n11570) );
  NAND3_X1 U14175 ( .A1(n11568), .A2(n11567), .A3(n11566), .ZN(n11569) );
  AOI21_X1 U14176 ( .B1(n11570), .B2(n11569), .A(n13622), .ZN(n11571) );
  AOI211_X1 U14177 ( .C1(n13615), .C2(n11573), .A(n11572), .B(n11571), .ZN(
        n11582) );
  INV_X1 U14178 ( .A(n11576), .ZN(n11575) );
  XNOR2_X1 U14179 ( .A(n11885), .B(n11574), .ZN(n11577) );
  NOR3_X1 U14180 ( .A1(n11575), .A2(n7097), .A3(n11577), .ZN(n11580) );
  NAND2_X1 U14181 ( .A1(n11578), .A2(n11577), .ZN(n11871) );
  INV_X1 U14182 ( .A(n11871), .ZN(n11579) );
  OAI21_X1 U14183 ( .B1(n11580), .B2(n11579), .A(n13621), .ZN(n11581) );
  OAI211_X1 U14184 ( .C1(n11583), .C2(n13612), .A(n11582), .B(n11581), .ZN(
        P3_U3192) );
  OAI21_X1 U14185 ( .B1(n11584), .B2(n12973), .A(n11631), .ZN(n15953) );
  NOR2_X1 U14186 ( .A1(n11586), .A2(n11585), .ZN(n11587) );
  XNOR2_X1 U14187 ( .A(n11587), .B(n12973), .ZN(n11589) );
  OAI22_X1 U14188 ( .A1(n11851), .A2(n15992), .B1(n11664), .B2(n15990), .ZN(
        n11588) );
  AOI21_X1 U14189 ( .B1(n11589), .B2(n13833), .A(n11588), .ZN(n15954) );
  INV_X1 U14190 ( .A(n15954), .ZN(n11590) );
  AOI21_X1 U14191 ( .B1(n16007), .B2(n15953), .A(n11590), .ZN(n11593) );
  AOI22_X1 U14192 ( .A1(n13893), .A2(n15959), .B1(n16023), .B2(
        P3_REG1_REG_6__SCAN_IN), .ZN(n11591) );
  OAI21_X1 U14193 ( .B1(n11593), .B2(n16023), .A(n11591), .ZN(P3_U3465) );
  AOI22_X1 U14194 ( .A1(n13981), .A2(n15959), .B1(n16018), .B2(
        P3_REG0_REG_6__SCAN_IN), .ZN(n11592) );
  OAI21_X1 U14195 ( .B1(n11593), .B2(n16018), .A(n11592), .ZN(P3_U3408) );
  XNOR2_X1 U14196 ( .A(n11698), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n11600) );
  NAND2_X1 U14197 ( .A1(n11594), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n15881) );
  XNOR2_X1 U14198 ( .A(n15895), .B(n11595), .ZN(n15884) );
  AND2_X1 U14199 ( .A1(n15881), .A2(n15884), .ZN(n11596) );
  NAND2_X1 U14200 ( .A1(n15882), .A2(n11596), .ZN(n15883) );
  OR2_X1 U14201 ( .A1(n15895), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n11597) );
  NAND2_X1 U14202 ( .A1(n15883), .A2(n11597), .ZN(n11599) );
  INV_X1 U14203 ( .A(n11700), .ZN(n11598) );
  AOI211_X1 U14204 ( .C1(n11600), .C2(n11599), .A(n15873), .B(n11598), .ZN(
        n11612) );
  NAND2_X1 U14205 ( .A1(n11601), .A2(n12508), .ZN(n15887) );
  MUX2_X1 U14206 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n9639), .S(n15895), .Z(
        n15886) );
  NAND2_X1 U14207 ( .A1(n11602), .A2(n15886), .ZN(n15891) );
  OR2_X1 U14208 ( .A1(n15895), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n11603) );
  NAND2_X1 U14209 ( .A1(n15891), .A2(n11603), .ZN(n11606) );
  MUX2_X1 U14210 ( .A(n14644), .B(P2_REG2_REG_13__SCAN_IN), .S(n11698), .Z(
        n11605) );
  INV_X1 U14211 ( .A(n11693), .ZN(n11604) );
  AOI211_X1 U14212 ( .C1(n11606), .C2(n11605), .A(n14330), .B(n11604), .ZN(
        n11611) );
  NOR2_X1 U14213 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11607), .ZN(n11608) );
  AOI21_X1 U14214 ( .B1(n15894), .B2(n11698), .A(n11608), .ZN(n11609) );
  OAI21_X1 U14215 ( .B1(n15900), .B2(n7048), .A(n11609), .ZN(n11610) );
  OR3_X1 U14216 ( .A1(n11612), .A2(n11611), .A3(n11610), .ZN(P2_U3227) );
  NAND2_X1 U14217 ( .A1(n11613), .A2(n13999), .ZN(n11614) );
  OAI211_X1 U14218 ( .C1(n11615), .C2(n14006), .A(n11614), .B(n13145), .ZN(
        P3_U3272) );
  OR2_X1 U14219 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n15052), .ZN(n11621) );
  NAND2_X1 U14220 ( .A1(n11622), .A2(n11621), .ZN(n11829) );
  INV_X1 U14221 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n11827) );
  XNOR2_X1 U14222 ( .A(n11827), .B(P1_ADDR_REG_11__SCAN_IN), .ZN(n11828) );
  INV_X1 U14223 ( .A(n11828), .ZN(n11623) );
  XNOR2_X1 U14224 ( .A(n11829), .B(n11623), .ZN(n11624) );
  NAND2_X1 U14225 ( .A1(n11824), .A2(n11825), .ZN(n11626) );
  XNOR2_X1 U14226 ( .A(n11626), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  INV_X1 U14227 ( .A(n11627), .ZN(n11628) );
  OAI222_X1 U14228 ( .A1(n11630), .A2(P3_U3151), .B1(n14006), .B2(n11629), 
        .C1(n13257), .C2(n11628), .ZN(P3_U3274) );
  NAND2_X1 U14229 ( .A1(n11800), .A2(n13456), .ZN(n13043) );
  NAND2_X1 U14230 ( .A1(n11853), .A2(n12198), .ZN(n13042) );
  OAI21_X1 U14231 ( .B1(n11632), .B2(n13041), .A(n11798), .ZN(n11727) );
  NAND2_X1 U14232 ( .A1(n13457), .A2(n15950), .ZN(n11633) );
  NAND2_X1 U14233 ( .A1(n11635), .A2(n13041), .ZN(n11636) );
  NAND2_X1 U14234 ( .A1(n11802), .A2(n11636), .ZN(n11637) );
  NAND2_X1 U14235 ( .A1(n11637), .A2(n13833), .ZN(n11639) );
  AOI22_X1 U14236 ( .A1(n13457), .A2(n13828), .B1(n13830), .B2(n11848), .ZN(
        n11638) );
  NAND2_X1 U14237 ( .A1(n11639), .A2(n11638), .ZN(n11728) );
  AOI21_X1 U14238 ( .B1(n11727), .B2(n16007), .A(n11728), .ZN(n11739) );
  AOI22_X1 U14239 ( .A1(n13981), .A2(n11853), .B1(n16018), .B2(
        P3_REG0_REG_8__SCAN_IN), .ZN(n11640) );
  OAI21_X1 U14240 ( .B1(n11739), .B2(n16018), .A(n11640), .ZN(P3_U3414) );
  MUX2_X1 U14241 ( .A(n11642), .B(n11641), .S(n13911), .Z(n11643) );
  OAI21_X1 U14242 ( .B1(n13905), .B2(n12062), .A(n11643), .ZN(P3_U3466) );
  NAND2_X1 U14243 ( .A1(n11742), .A2(n10876), .ZN(n11648) );
  NAND2_X1 U14244 ( .A1(n13189), .A2(n15017), .ZN(n11647) );
  NAND2_X1 U14245 ( .A1(n11648), .A2(n11647), .ZN(n11649) );
  XNOR2_X1 U14246 ( .A(n11649), .B(n13233), .ZN(n11895) );
  NAND2_X1 U14247 ( .A1(n11742), .A2(n13189), .ZN(n11651) );
  NAND2_X1 U14248 ( .A1(n13235), .A2(n15017), .ZN(n11650) );
  XNOR2_X1 U14249 ( .A(n11895), .B(n11894), .ZN(n11652) );
  XNOR2_X1 U14250 ( .A(n11893), .B(n11652), .ZN(n11658) );
  NAND2_X1 U14251 ( .A1(n11742), .A2(n15813), .ZN(n15804) );
  AOI22_X1 U14252 ( .A1(n14960), .A2(n15803), .B1(P1_REG3_REG_5__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11656) );
  INV_X1 U14253 ( .A(n11653), .ZN(n11654) );
  NAND2_X1 U14254 ( .A1(n14928), .A2(n11654), .ZN(n11655) );
  OAI211_X1 U14255 ( .C1(n14980), .C2(n15804), .A(n11656), .B(n11655), .ZN(
        n11657) );
  AOI21_X1 U14256 ( .B1(n11658), .B2(n14969), .A(n11657), .ZN(n11659) );
  INV_X1 U14257 ( .A(n11659), .ZN(P1_U3227) );
  INV_X1 U14258 ( .A(n15957), .ZN(n11671) );
  INV_X1 U14259 ( .A(n13443), .ZN(n13323) );
  OAI211_X1 U14260 ( .C1(n11662), .C2(n11661), .A(n11660), .B(n13437), .ZN(
        n11670) );
  AOI21_X1 U14261 ( .B1(n13430), .B2(n13457), .A(n11663), .ZN(n11666) );
  OR2_X1 U14262 ( .A1(n13428), .A2(n11664), .ZN(n11665) );
  OAI211_X1 U14263 ( .C1(n13446), .C2(n11667), .A(n11666), .B(n11665), .ZN(
        n11668) );
  INV_X1 U14264 ( .A(n11668), .ZN(n11669) );
  OAI211_X1 U14265 ( .C1(n11671), .C2(n13323), .A(n11670), .B(n11669), .ZN(
        P3_U3179) );
  NAND2_X1 U14266 ( .A1(n14654), .A2(n14213), .ZN(n11673) );
  NAND2_X1 U14267 ( .A1(n14652), .A2(n14215), .ZN(n11672) );
  AND2_X1 U14268 ( .A1(n11673), .A2(n11672), .ZN(n12301) );
  OAI22_X1 U14269 ( .A1(n14147), .A2(n12301), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15856), .ZN(n11674) );
  AOI21_X1 U14270 ( .B1(n11676), .B2(n11675), .A(n14154), .ZN(n11677) );
  NAND2_X1 U14271 ( .A1(n11677), .A2(n14109), .ZN(n11678) );
  OAI211_X1 U14272 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n14186), .A(n11679), .B(
        n11678), .ZN(P2_U3190) );
  XOR2_X1 U14273 ( .A(n11681), .B(n11680), .Z(n11686) );
  INV_X1 U14274 ( .A(n14184), .ZN(n14160) );
  INV_X1 U14275 ( .A(n14185), .ZN(n14113) );
  AOI22_X1 U14276 ( .A1(n14160), .A2(n14215), .B1(n14113), .B2(n10168), .ZN(
        n11685) );
  NAND2_X1 U14277 ( .A1(n11683), .A2(n11682), .ZN(n13270) );
  AOI22_X1 U14278 ( .A1(n14189), .A2(n12099), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n13270), .ZN(n11684) );
  OAI211_X1 U14279 ( .C1(n11686), .C2(n14154), .A(n11685), .B(n11684), .ZN(
        P2_U3194) );
  XOR2_X1 U14280 ( .A(n11688), .B(n11687), .Z(n11691) );
  AOI22_X1 U14281 ( .A1(n14160), .A2(n14214), .B1(n14113), .B2(n14216), .ZN(
        n11690) );
  AOI22_X1 U14282 ( .A1(n14189), .A2(n12114), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n13270), .ZN(n11689) );
  OAI211_X1 U14283 ( .C1(n11691), .C2(n14154), .A(n11690), .B(n11689), .ZN(
        P2_U3209) );
  NAND2_X1 U14284 ( .A1(n11698), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11692) );
  NAND2_X1 U14285 ( .A1(n11693), .A2(n11692), .ZN(n11935) );
  XNOR2_X1 U14286 ( .A(n11935), .B(n11695), .ZN(n11934) );
  XNOR2_X1 U14287 ( .A(n11934), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n11706) );
  NOR2_X1 U14288 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11694), .ZN(n11697) );
  NOR2_X1 U14289 ( .A1(n14306), .A2(n11695), .ZN(n11696) );
  AOI211_X1 U14290 ( .C1(P2_ADDR_REG_14__SCAN_IN), .C2(n15851), .A(n11697), 
        .B(n11696), .ZN(n11705) );
  NAND2_X1 U14291 ( .A1(n11698), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11699) );
  NAND2_X1 U14292 ( .A1(n11700), .A2(n11699), .ZN(n11703) );
  XNOR2_X1 U14293 ( .A(n11940), .B(n11701), .ZN(n11702) );
  NAND2_X1 U14294 ( .A1(n11703), .A2(n11702), .ZN(n11942) );
  OAI211_X1 U14295 ( .C1(n11703), .C2(n11702), .A(n11942), .B(n15896), .ZN(
        n11704) );
  OAI211_X1 U14296 ( .C1(n11706), .C2(n14330), .A(n11705), .B(n11704), .ZN(
        P2_U3228) );
  NOR2_X1 U14297 ( .A1(n11742), .A2(n15017), .ZN(n11746) );
  NOR2_X1 U14298 ( .A1(n11707), .A2(n11746), .ZN(n11708) );
  XNOR2_X1 U14299 ( .A(n11708), .B(n11713), .ZN(n15734) );
  INV_X1 U14300 ( .A(n15734), .ZN(n11719) );
  INV_X1 U14301 ( .A(n15433), .ZN(n15792) );
  NAND2_X1 U14302 ( .A1(n11742), .A2(n11711), .ZN(n11712) );
  XOR2_X1 U14303 ( .A(n11754), .B(n11713), .Z(n11714) );
  AOI22_X1 U14304 ( .A1(n15015), .A2(n15746), .B1(n15426), .B2(n15017), .ZN(
        n11793) );
  OAI21_X1 U14305 ( .B1(n11714), .B2(n15829), .A(n11793), .ZN(n11715) );
  AOI21_X1 U14306 ( .B1(n15792), .B2(n15734), .A(n11715), .ZN(n15737) );
  INV_X1 U14307 ( .A(n11760), .ZN(n11716) );
  AOI211_X1 U14308 ( .C1(n15731), .C2(n11717), .A(n15742), .B(n11716), .ZN(
        n15733) );
  AOI21_X1 U14309 ( .B1(n15813), .B2(n15731), .A(n15733), .ZN(n11718) );
  OAI211_X1 U14310 ( .C1(n15815), .C2(n11719), .A(n15737), .B(n11718), .ZN(
        n11721) );
  NAND2_X1 U14311 ( .A1(n11721), .A2(n15838), .ZN(n11720) );
  OAI21_X1 U14312 ( .B1(n15838), .B2(n8796), .A(n11720), .ZN(P1_U3477) );
  INV_X2 U14313 ( .A(n15848), .ZN(n15850) );
  NAND2_X1 U14314 ( .A1(n11721), .A2(n15850), .ZN(n11722) );
  OAI21_X1 U14315 ( .B1(n15850), .B2(n11723), .A(n11722), .ZN(P1_U3534) );
  INV_X1 U14316 ( .A(n11724), .ZN(n11725) );
  OAI222_X1 U14317 ( .A1(n14826), .A2(n11726), .B1(P2_U3088), .B2(n9433), .C1(
        n14832), .C2(n11725), .ZN(P2_U3305) );
  INV_X1 U14318 ( .A(n11727), .ZN(n11733) );
  AOI22_X1 U14319 ( .A1(n15958), .A2(n11853), .B1(n15977), .B2(n11846), .ZN(
        n11732) );
  INV_X1 U14320 ( .A(n11728), .ZN(n11730) );
  MUX2_X1 U14321 ( .A(n11730), .B(n11729), .S(n15997), .Z(n11731) );
  OAI211_X1 U14322 ( .C1(n11733), .C2(n13807), .A(n11732), .B(n11731), .ZN(
        P3_U3225) );
  INV_X1 U14323 ( .A(n11734), .ZN(n11738) );
  AOI21_X1 U14324 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n14830), .A(n6782), 
        .ZN(n11735) );
  OAI21_X1 U14325 ( .B1(n11738), .B2(n14832), .A(n11735), .ZN(P2_U3304) );
  AOI21_X1 U14326 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n15588), .A(n11736), 
        .ZN(n11737) );
  OAI21_X1 U14327 ( .B1(n11738), .B2(n15595), .A(n11737), .ZN(P1_U3332) );
  MUX2_X1 U14328 ( .A(n11740), .B(n11739), .S(n13911), .Z(n11741) );
  OAI21_X1 U14329 ( .B1(n11800), .B2(n13905), .A(n11741), .ZN(P3_U3467) );
  NAND2_X1 U14330 ( .A1(n15731), .A2(n15016), .ZN(n11745) );
  NAND2_X1 U14331 ( .A1(n11742), .A2(n15017), .ZN(n11743) );
  NOR2_X1 U14332 ( .A1(n15731), .A2(n15016), .ZN(n11744) );
  AOI21_X1 U14333 ( .B1(n11746), .B2(n11745), .A(n11744), .ZN(n11747) );
  OR2_X1 U14334 ( .A1(n11749), .A2(n11755), .ZN(n11750) );
  AND2_X1 U14335 ( .A1(n12005), .A2(n11750), .ZN(n15816) );
  INV_X1 U14336 ( .A(n11751), .ZN(n11752) );
  NAND2_X1 U14337 ( .A1(n6544), .A2(n11752), .ZN(n15438) );
  NAND2_X1 U14338 ( .A1(n11797), .A2(n15016), .ZN(n11753) );
  XNOR2_X1 U14339 ( .A(n11954), .B(n11755), .ZN(n11756) );
  NAND2_X1 U14340 ( .A1(n11756), .A2(n15754), .ZN(n11758) );
  AOI22_X1 U14341 ( .A1(n15016), .A2(n15426), .B1(n15746), .B2(n15014), .ZN(
        n11757) );
  OAI211_X1 U14342 ( .C1(n15816), .C2(n15433), .A(n11758), .B(n11757), .ZN(
        n15818) );
  MUX2_X1 U14343 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n15818), .S(n6544), .Z(
        n11759) );
  INV_X1 U14344 ( .A(n11759), .ZN(n11764) );
  AOI211_X1 U14345 ( .C1(n15812), .C2(n11760), .A(n15742), .B(n11950), .ZN(
        n15811) );
  OAI22_X1 U14346 ( .A1(n15418), .A2(n11761), .B1(n15393), .B2(n14843), .ZN(
        n11762) );
  AOI21_X1 U14347 ( .B1(n15811), .B2(n15732), .A(n11762), .ZN(n11763) );
  OAI211_X1 U14348 ( .C1(n15816), .C2(n15438), .A(n11764), .B(n11763), .ZN(
        P1_U3286) );
  XNOR2_X1 U14349 ( .A(n15066), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n11769) );
  XNOR2_X1 U14350 ( .A(n15710), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n15708) );
  AOI211_X1 U14351 ( .C1(n11769), .C2(n11768), .A(n15102), .B(n15065), .ZN(
        n11780) );
  MUX2_X1 U14352 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n12386), .S(n15710), .Z(
        n15707) );
  INV_X1 U14353 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11772) );
  MUX2_X1 U14354 ( .A(n11772), .B(P1_REG2_REG_13__SCAN_IN), .S(n15066), .Z(
        n11773) );
  AOI211_X1 U14355 ( .C1(n11774), .C2(n11773), .A(n15142), .B(n15075), .ZN(
        n11779) );
  NOR2_X1 U14356 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11775), .ZN(n11776) );
  AOI21_X1 U14357 ( .B1(n15680), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n11776), 
        .ZN(n11777) );
  OAI21_X1 U14358 ( .B1(n15072), .B2(n15699), .A(n11777), .ZN(n11778) );
  OR3_X1 U14359 ( .A1(n11780), .A2(n11779), .A3(n11778), .ZN(P1_U3256) );
  INV_X1 U14360 ( .A(n11893), .ZN(n11782) );
  INV_X1 U14361 ( .A(n11894), .ZN(n11899) );
  INV_X1 U14362 ( .A(n11895), .ZN(n11900) );
  OAI21_X1 U14363 ( .B1(n11893), .B2(n11899), .A(n11900), .ZN(n11781) );
  OAI21_X1 U14364 ( .B1(n11782), .B2(n11894), .A(n11781), .ZN(n11789) );
  NAND2_X1 U14365 ( .A1(n15731), .A2(n10876), .ZN(n11784) );
  NAND2_X1 U14366 ( .A1(n15016), .A2(n13189), .ZN(n11783) );
  NAND2_X1 U14367 ( .A1(n11784), .A2(n11783), .ZN(n11785) );
  XNOR2_X1 U14368 ( .A(n11785), .B(n13233), .ZN(n11896) );
  NAND2_X1 U14369 ( .A1(n15731), .A2(n13189), .ZN(n11787) );
  OR2_X1 U14370 ( .A1(n13223), .A2(n14839), .ZN(n11786) );
  XNOR2_X1 U14371 ( .A(n11896), .B(n11897), .ZN(n11788) );
  XNOR2_X1 U14372 ( .A(n11789), .B(n11788), .ZN(n11790) );
  NAND2_X1 U14373 ( .A1(n11790), .A2(n14969), .ZN(n11796) );
  INV_X1 U14374 ( .A(n11791), .ZN(n15729) );
  OAI21_X1 U14375 ( .B1(n14989), .B2(n11793), .A(n11792), .ZN(n11794) );
  AOI21_X1 U14376 ( .B1(n15729), .B2(n14928), .A(n11794), .ZN(n11795) );
  OAI211_X1 U14377 ( .C1(n11797), .C2(n14963), .A(n11796), .B(n11795), .ZN(
        P1_U3239) );
  NAND2_X1 U14378 ( .A1(n12203), .A2(n11848), .ZN(n13047) );
  OR2_X1 U14379 ( .A1(n12203), .A2(n11848), .ZN(n13048) );
  XNOR2_X1 U14380 ( .A(n13308), .B(n13455), .ZN(n11804) );
  OAI21_X1 U14381 ( .B1(n7979), .B2(n7944), .A(n12527), .ZN(n11822) );
  INV_X1 U14382 ( .A(n16007), .ZN(n13909) );
  NOR2_X1 U14383 ( .A1(n16018), .A2(n13909), .ZN(n13992) );
  INV_X1 U14384 ( .A(n13992), .ZN(n13988) );
  INV_X1 U14385 ( .A(n13308), .ZN(n11799) );
  AOI22_X1 U14386 ( .A1(n13981), .A2(n11799), .B1(P3_REG0_REG_10__SCAN_IN), 
        .B2(n16018), .ZN(n11810) );
  NAND2_X1 U14387 ( .A1(n11800), .A2(n12198), .ZN(n11801) );
  NAND2_X1 U14388 ( .A1(n13048), .A2(n13047), .ZN(n12979) );
  OR2_X1 U14389 ( .A1(n12203), .A2(n13303), .ZN(n11805) );
  NAND3_X1 U14390 ( .A1(n11837), .A2(n7944), .A3(n11805), .ZN(n11806) );
  NAND3_X1 U14391 ( .A1(n12070), .A2(n13833), .A3(n11806), .ZN(n11808) );
  AOI22_X1 U14392 ( .A1(n13828), .A2(n11848), .B1(n13454), .B2(n13830), .ZN(
        n11807) );
  NAND2_X1 U14393 ( .A1(n11808), .A2(n11807), .ZN(n11820) );
  NAND2_X1 U14394 ( .A1(n11820), .A2(n16017), .ZN(n11809) );
  OAI211_X1 U14395 ( .C1(n11822), .C2(n13988), .A(n11810), .B(n11809), .ZN(
        P3_U3420) );
  INV_X1 U14396 ( .A(n11811), .ZN(n11813) );
  OAI222_X1 U14397 ( .A1(P3_U3151), .A2(n11814), .B1(n13257), .B2(n11813), 
        .C1(n11812), .C2(n14006), .ZN(P3_U3271) );
  INV_X1 U14398 ( .A(n13902), .ZN(n13900) );
  OAI22_X1 U14399 ( .A1(n13905), .A2(n13308), .B1(n13911), .B2(n11815), .ZN(
        n11816) );
  AOI21_X1 U14400 ( .B1(n11820), .B2(n13911), .A(n11816), .ZN(n11817) );
  OAI21_X1 U14401 ( .B1(n11822), .B2(n13900), .A(n11817), .ZN(P3_U3469) );
  AOI22_X1 U14402 ( .A1(n15997), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n15977), 
        .B2(n13305), .ZN(n11818) );
  OAI21_X1 U14403 ( .B1(n13825), .B2(n13308), .A(n11818), .ZN(n11819) );
  AOI21_X1 U14404 ( .B1(n11820), .B2(n15995), .A(n11819), .ZN(n11821) );
  OAI21_X1 U14405 ( .B1(n11822), .B2(n13807), .A(n11821), .ZN(P3_U3223) );
  INV_X1 U14406 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n11823) );
  NAND2_X1 U14407 ( .A1(n11824), .A2(n11823), .ZN(n11826) );
  OAI22_X1 U14408 ( .A1(n11829), .A2(n11828), .B1(P1_ADDR_REG_11__SCAN_IN), 
        .B2(n11827), .ZN(n12292) );
  XNOR2_X1 U14409 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n12291) );
  INV_X1 U14410 ( .A(n12291), .ZN(n11830) );
  XNOR2_X1 U14411 ( .A(n12292), .B(n11830), .ZN(n11831) );
  NAND2_X1 U14412 ( .A1(n12289), .A2(n12290), .ZN(n11833) );
  XNOR2_X1 U14413 ( .A(n11833), .B(P2_ADDR_REG_12__SCAN_IN), .ZN(SUB_1596_U68)
         );
  XNOR2_X1 U14414 ( .A(n11834), .B(n12979), .ZN(n13910) );
  NAND2_X1 U14415 ( .A1(n11835), .A2(n13045), .ZN(n11836) );
  NAND3_X1 U14416 ( .A1(n11837), .A2(n13833), .A3(n11836), .ZN(n11839) );
  AOI22_X1 U14417 ( .A1(n13828), .A2(n13456), .B1(n13455), .B2(n13830), .ZN(
        n11838) );
  NAND2_X1 U14418 ( .A1(n11839), .A2(n11838), .ZN(n13906) );
  INV_X1 U14419 ( .A(n13906), .ZN(n11841) );
  MUX2_X1 U14420 ( .A(n11841), .B(n11840), .S(n15997), .Z(n11843) );
  INV_X1 U14421 ( .A(n12203), .ZN(n13907) );
  AOI22_X1 U14422 ( .A1(n15958), .A2(n13907), .B1(n15977), .B2(n12200), .ZN(
        n11842) );
  OAI211_X1 U14423 ( .C1(n13807), .C2(n13910), .A(n11843), .B(n11842), .ZN(
        P3_U3224) );
  XNOR2_X1 U14424 ( .A(n11845), .B(n11844), .ZN(n11855) );
  NAND2_X1 U14425 ( .A1(n13443), .A2(n11846), .ZN(n11850) );
  AOI21_X1 U14426 ( .B1(n13430), .B2(n11848), .A(n11847), .ZN(n11849) );
  OAI211_X1 U14427 ( .C1(n11851), .C2(n13428), .A(n11850), .B(n11849), .ZN(
        n11852) );
  AOI21_X1 U14428 ( .B1(n11853), .B2(n13400), .A(n11852), .ZN(n11854) );
  OAI21_X1 U14429 ( .B1(n11855), .B2(n13413), .A(n11854), .ZN(P3_U3161) );
  INV_X1 U14430 ( .A(n15913), .ZN(n11856) );
  NAND2_X1 U14431 ( .A1(n15910), .A2(n11856), .ZN(n11857) );
  AND2_X1 U14432 ( .A1(n11861), .A2(n11860), .ZN(n11862) );
  NAND2_X1 U14433 ( .A1(n14645), .A2(n11862), .ZN(n14554) );
  INV_X1 U14434 ( .A(n14554), .ZN(n12112) );
  INV_X1 U14435 ( .A(n14784), .ZN(n11863) );
  NAND2_X1 U14436 ( .A1(n12112), .A2(n11863), .ZN(n11869) );
  NAND2_X1 U14437 ( .A1(n11864), .A2(n13267), .ZN(n14782) );
  AOI21_X1 U14438 ( .B1(n14634), .B2(n11968), .A(n14784), .ZN(n11865) );
  AOI21_X1 U14439 ( .B1(n14654), .B2(n14216), .A(n11865), .ZN(n14783) );
  OAI21_X1 U14440 ( .B1(n11866), .B2(n14782), .A(n14783), .ZN(n11867) );
  INV_X1 U14441 ( .A(n14642), .ZN(n14661) );
  AOI22_X1 U14442 ( .A1(n14645), .A2(n11867), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n14661), .ZN(n11868) );
  OAI211_X1 U14443 ( .C1(n12668), .C2(n14645), .A(n11869), .B(n11868), .ZN(
        P2_U3265) );
  NAND2_X1 U14444 ( .A1(n11885), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n11870) );
  OR2_X1 U14445 ( .A1(n11872), .A2(n12145), .ZN(n11873) );
  OAI21_X1 U14446 ( .B1(P3_REG2_REG_11__SCAN_IN), .B2(n11874), .A(n12142), 
        .ZN(n11884) );
  NAND2_X1 U14447 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n13405)
         );
  NAND2_X1 U14448 ( .A1(n15945), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n11875) );
  OAI211_X1 U14449 ( .C1(n13586), .C2(n12145), .A(n13405), .B(n11875), .ZN(
        n11883) );
  INV_X1 U14450 ( .A(n11876), .ZN(n11877) );
  NOR2_X1 U14451 ( .A1(n11878), .A2(n11877), .ZN(n11880) );
  MUX2_X1 U14452 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13576), .Z(n12146) );
  XNOR2_X1 U14453 ( .A(n12146), .B(n12145), .ZN(n11879) );
  NOR2_X1 U14454 ( .A1(n11880), .A2(n11879), .ZN(n12149) );
  AOI21_X1 U14455 ( .B1(n11880), .B2(n11879), .A(n12149), .ZN(n11881) );
  NOR2_X1 U14456 ( .A1(n11881), .A2(n13622), .ZN(n11882) );
  AOI211_X1 U14457 ( .C1(n13621), .C2(n11884), .A(n11883), .B(n11882), .ZN(
        n11891) );
  NAND2_X1 U14458 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n11888), .ZN(n12137) );
  OAI21_X1 U14459 ( .B1(n11888), .B2(P3_REG1_REG_11__SCAN_IN), .A(n12137), 
        .ZN(n11889) );
  NAND2_X1 U14460 ( .A1(n11889), .A2(n13589), .ZN(n11890) );
  NAND2_X1 U14461 ( .A1(n11891), .A2(n11890), .ZN(P3_U3193) );
  AOI22_X1 U14462 ( .A1(n11895), .A2(n11894), .B1(n11896), .B2(n11897), .ZN(
        n11892) );
  OAI21_X1 U14463 ( .B1(n11895), .B2(n11894), .A(n11897), .ZN(n11903) );
  INV_X1 U14464 ( .A(n11896), .ZN(n11902) );
  INV_X1 U14465 ( .A(n11897), .ZN(n11898) );
  AND2_X1 U14466 ( .A1(n11899), .A2(n11898), .ZN(n11901) );
  AOI22_X1 U14467 ( .A1(n11903), .A2(n11902), .B1(n11901), .B2(n11900), .ZN(
        n11904) );
  NAND2_X1 U14468 ( .A1(n11905), .A2(n11904), .ZN(n14836) );
  NAND2_X1 U14469 ( .A1(n15812), .A2(n10876), .ZN(n11907) );
  NAND2_X1 U14470 ( .A1(n15015), .A2(n13189), .ZN(n11906) );
  NAND2_X1 U14471 ( .A1(n11907), .A2(n11906), .ZN(n11909) );
  XNOR2_X1 U14472 ( .A(n11909), .B(n11908), .ZN(n11911) );
  NOR2_X1 U14473 ( .A1(n13223), .A2(n11955), .ZN(n11910) );
  AOI21_X1 U14474 ( .B1(n15812), .B2(n13189), .A(n11910), .ZN(n11912) );
  XNOR2_X1 U14475 ( .A(n11911), .B(n11912), .ZN(n14837) );
  INV_X1 U14476 ( .A(n11911), .ZN(n11913) );
  OR2_X1 U14477 ( .A1(n11913), .A2(n11912), .ZN(n11914) );
  NAND2_X1 U14478 ( .A1(n12001), .A2(n10876), .ZN(n11917) );
  NAND2_X1 U14479 ( .A1(n13189), .A2(n15014), .ZN(n11916) );
  NAND2_X1 U14480 ( .A1(n11917), .A2(n11916), .ZN(n11918) );
  XNOR2_X1 U14481 ( .A(n11918), .B(n13233), .ZN(n11920) );
  INV_X1 U14482 ( .A(n15014), .ZN(n14840) );
  NOR2_X1 U14483 ( .A1(n13223), .A2(n14840), .ZN(n11919) );
  AOI21_X1 U14484 ( .B1(n12001), .B2(n13189), .A(n11919), .ZN(n11921) );
  NAND2_X1 U14485 ( .A1(n11920), .A2(n11921), .ZN(n12416) );
  INV_X1 U14486 ( .A(n11920), .ZN(n11923) );
  INV_X1 U14487 ( .A(n11921), .ZN(n11922) );
  NAND2_X1 U14488 ( .A1(n11923), .A2(n11922), .ZN(n11924) );
  NAND2_X1 U14489 ( .A1(n12416), .A2(n11924), .ZN(n11928) );
  INV_X1 U14490 ( .A(n11928), .ZN(n11926) );
  INV_X1 U14491 ( .A(n12417), .ZN(n11927) );
  AOI21_X1 U14492 ( .B1(n11925), .B2(n11928), .A(n11927), .ZN(n11933) );
  OAI21_X1 U14493 ( .B1(n14971), .B2(n11955), .A(n11929), .ZN(n11931) );
  INV_X1 U14494 ( .A(n14928), .ZN(n14988) );
  OAI22_X1 U14495 ( .A1(n14963), .A2(n15821), .B1(n14988), .B2(n11951), .ZN(
        n11930) );
  AOI211_X1 U14496 ( .C1(n14983), .C2(n15013), .A(n11931), .B(n11930), .ZN(
        n11932) );
  OAI21_X1 U14497 ( .B1(n11933), .B2(n14994), .A(n11932), .ZN(P1_U3221) );
  NAND2_X1 U14498 ( .A1(n11934), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n11937) );
  NAND2_X1 U14499 ( .A1(n11935), .A2(n11940), .ZN(n11936) );
  NAND2_X1 U14500 ( .A1(n11937), .A2(n11936), .ZN(n12205) );
  XNOR2_X1 U14501 ( .A(n12205), .B(n11943), .ZN(n12204) );
  XNOR2_X1 U14502 ( .A(n12204), .B(P2_REG2_REG_15__SCAN_IN), .ZN(n11947) );
  NOR2_X1 U14503 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14183), .ZN(n11939) );
  NOR2_X1 U14504 ( .A1(n14306), .A2(n11943), .ZN(n11938) );
  AOI211_X1 U14505 ( .C1(n15851), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n11939), 
        .B(n11938), .ZN(n11946) );
  NAND2_X1 U14506 ( .A1(n11940), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n11941) );
  NAND2_X1 U14507 ( .A1(n11942), .A2(n11941), .ZN(n12211) );
  XNOR2_X1 U14508 ( .A(n12211), .B(n11943), .ZN(n11944) );
  NAND2_X1 U14509 ( .A1(n11944), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n12213) );
  OAI211_X1 U14510 ( .C1(n11944), .C2(P2_REG1_REG_15__SCAN_IN), .A(n12213), 
        .B(n15896), .ZN(n11945) );
  OAI211_X1 U14511 ( .C1(n11947), .C2(n14330), .A(n11946), .B(n11945), .ZN(
        P2_U3229) );
  OR2_X1 U14512 ( .A1(n15812), .A2(n15015), .ZN(n12003) );
  NAND2_X1 U14513 ( .A1(n12005), .A2(n12003), .ZN(n11949) );
  INV_X1 U14514 ( .A(n11959), .ZN(n11948) );
  NAND2_X1 U14515 ( .A1(n11949), .A2(n11948), .ZN(n12002) );
  OAI21_X1 U14516 ( .B1(n11949), .B2(n11948), .A(n12002), .ZN(n15824) );
  OAI211_X1 U14517 ( .C1(n11950), .C2(n15821), .A(n12029), .B(n10870), .ZN(
        n15820) );
  INV_X1 U14518 ( .A(n15732), .ZN(n15304) );
  INV_X1 U14519 ( .A(n11951), .ZN(n11952) );
  AOI22_X1 U14520 ( .A1(n15730), .A2(n12001), .B1(n15760), .B2(n11952), .ZN(
        n11953) );
  OAI21_X1 U14521 ( .B1(n15820), .B2(n15304), .A(n11953), .ZN(n11964) );
  NAND2_X1 U14522 ( .A1(n15812), .A2(n11955), .ZN(n11956) );
  AND2_X1 U14523 ( .A1(n11958), .A2(n11956), .ZN(n11960) );
  AND2_X1 U14524 ( .A1(n11959), .A2(n11956), .ZN(n11957) );
  OAI211_X1 U14525 ( .C1(n11960), .C2(n11959), .A(n12010), .B(n15754), .ZN(
        n11962) );
  AOI22_X1 U14526 ( .A1(n15426), .A2(n15015), .B1(n15013), .B2(n15746), .ZN(
        n11961) );
  NAND2_X1 U14527 ( .A1(n11962), .A2(n11961), .ZN(n15822) );
  MUX2_X1 U14528 ( .A(n15822), .B(P1_REG2_REG_8__SCAN_IN), .S(n15764), .Z(
        n11963) );
  AOI211_X1 U14529 ( .C1(n15383), .C2(n15824), .A(n11964), .B(n11963), .ZN(
        n11965) );
  INV_X1 U14530 ( .A(n11965), .ZN(P1_U3285) );
  OAI21_X1 U14531 ( .B1(n11967), .B2(n11971), .A(n11966), .ZN(n15936) );
  INV_X1 U14532 ( .A(n15936), .ZN(n11982) );
  INV_X1 U14533 ( .A(n11968), .ZN(n14547) );
  OAI22_X1 U14534 ( .A1(n12548), .A2(n14638), .B1(n14636), .B2(n14104), .ZN(
        n11975) );
  NAND3_X1 U14535 ( .A1(n11969), .A2(n11971), .A3(n11970), .ZN(n11972) );
  AOI21_X1 U14536 ( .B1(n11973), .B2(n11972), .A(n14634), .ZN(n11974) );
  AOI211_X1 U14537 ( .C1(n14547), .C2(n15936), .A(n11975), .B(n11974), .ZN(
        n15933) );
  MUX2_X1 U14538 ( .A(n11976), .B(n15933), .S(n14645), .Z(n11981) );
  NAND2_X1 U14539 ( .A1(n14645), .A2(n14332), .ZN(n14360) );
  AOI21_X1 U14540 ( .B1(n12186), .B2(n12350), .A(n14658), .ZN(n11978) );
  NAND2_X1 U14541 ( .A1(n11978), .A2(n12130), .ZN(n15930) );
  OAI22_X1 U14542 ( .A1(n14360), .A2(n15930), .B1(n12352), .B2(n14642), .ZN(
        n11979) );
  AOI21_X1 U14543 ( .B1(n14433), .B2(n12350), .A(n11979), .ZN(n11980) );
  OAI211_X1 U14544 ( .C1(n11982), .C2(n14554), .A(n11981), .B(n11980), .ZN(
        P2_U3259) );
  INV_X1 U14545 ( .A(n11983), .ZN(n11984) );
  OAI222_X1 U14546 ( .A1(n14006), .A2(n11985), .B1(n13257), .B2(n11984), .C1(
        n8091), .C2(P3_U3151), .ZN(P3_U3270) );
  NAND2_X1 U14547 ( .A1(n14645), .A2(n14547), .ZN(n11986) );
  OAI21_X1 U14548 ( .B1(n11988), .B2(n11992), .A(n11987), .ZN(n15928) );
  INV_X1 U14549 ( .A(n15928), .ZN(n12000) );
  NAND3_X1 U14550 ( .A1(n11990), .A2(n11992), .A3(n11991), .ZN(n11993) );
  NAND2_X1 U14551 ( .A1(n11989), .A2(n11993), .ZN(n11994) );
  AOI222_X1 U14552 ( .A1(n14657), .A2(n11994), .B1(n14212), .B2(n14654), .C1(
        n14214), .C2(n14652), .ZN(n15925) );
  MUX2_X1 U14553 ( .A(n11995), .B(n15925), .S(n14645), .Z(n11999) );
  OAI211_X1 U14554 ( .C1(n11996), .C2(n15924), .A(n12187), .B(n10450), .ZN(
        n15923) );
  OAI22_X1 U14555 ( .A1(n14360), .A2(n15923), .B1(n14105), .B2(n14642), .ZN(
        n11997) );
  AOI21_X1 U14556 ( .B1(n14433), .B2(n14107), .A(n11997), .ZN(n11998) );
  OAI211_X1 U14557 ( .C1(n14669), .C2(n12000), .A(n11999), .B(n11998), .ZN(
        P2_U3261) );
  OR2_X1 U14558 ( .A1(n12001), .A2(n15014), .ZN(n12004) );
  NAND2_X1 U14559 ( .A1(n12002), .A2(n12004), .ZN(n12008) );
  OAI21_X1 U14560 ( .B1(n12008), .B2(n12011), .A(n12023), .ZN(n12016) );
  INV_X1 U14561 ( .A(n12016), .ZN(n12042) );
  OAI22_X1 U14562 ( .A1(n14840), .A2(n15758), .B1(n15411), .B2(n12170), .ZN(
        n12015) );
  NAND2_X1 U14563 ( .A1(n15821), .A2(n15014), .ZN(n12009) );
  NAND2_X1 U14564 ( .A1(n12012), .A2(n12011), .ZN(n12013) );
  AOI21_X1 U14565 ( .B1(n7655), .B2(n12013), .A(n15829), .ZN(n12014) );
  AOI211_X1 U14566 ( .C1(n15792), .C2(n12016), .A(n12015), .B(n12014), .ZN(
        n12041) );
  MUX2_X1 U14567 ( .A(n12017), .B(n12041), .S(n6544), .Z(n12022) );
  XNOR2_X1 U14568 ( .A(n12029), .B(n12655), .ZN(n12018) );
  NOR2_X1 U14569 ( .A1(n12018), .A2(n15742), .ZN(n12039) );
  INV_X1 U14570 ( .A(n12655), .ZN(n12019) );
  OAI22_X1 U14571 ( .A1(n12019), .A2(n15418), .B1(n12643), .B2(n15393), .ZN(
        n12020) );
  AOI21_X1 U14572 ( .B1(n12039), .B2(n15732), .A(n12020), .ZN(n12021) );
  OAI211_X1 U14573 ( .C1(n12042), .C2(n15438), .A(n12022), .B(n12021), .ZN(
        P1_U3284) );
  INV_X1 U14574 ( .A(n12026), .ZN(n12024) );
  NAND2_X1 U14575 ( .A1(n12025), .A2(n12024), .ZN(n12172) );
  OAI21_X1 U14576 ( .B1(n12025), .B2(n12024), .A(n12172), .ZN(n15834) );
  INV_X1 U14577 ( .A(n15834), .ZN(n12038) );
  INV_X1 U14578 ( .A(n12158), .ZN(n15830) );
  NOR2_X1 U14579 ( .A1(n12027), .A2(n12026), .ZN(n15831) );
  OR3_X1 U14580 ( .A1(n15830), .A2(n15831), .A3(n15333), .ZN(n12037) );
  OAI22_X1 U14581 ( .A1(n6544), .A2(n12028), .B1(n12576), .B2(n15393), .ZN(
        n12035) );
  NAND2_X1 U14582 ( .A1(n12031), .A2(n12426), .ZN(n12030) );
  NAND2_X1 U14583 ( .A1(n12030), .A2(n10870), .ZN(n12032) );
  OR2_X1 U14584 ( .A1(n12032), .A2(n12165), .ZN(n12033) );
  AOI22_X1 U14585 ( .A1(n15013), .A2(n15426), .B1(n15746), .B2(n15011), .ZN(
        n12577) );
  AND2_X1 U14586 ( .A1(n12033), .A2(n12577), .ZN(n15826) );
  NOR3_X1 U14587 ( .A1(n15826), .A2(n15748), .A3(n15764), .ZN(n12034) );
  AOI211_X1 U14588 ( .C1(n15730), .C2(n12426), .A(n12035), .B(n12034), .ZN(
        n12036) );
  OAI211_X1 U14589 ( .C1(n12038), .C2(n15423), .A(n12037), .B(n12036), .ZN(
        P1_U3283) );
  INV_X1 U14590 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n12044) );
  AOI21_X1 U14591 ( .B1(n15813), .B2(n12655), .A(n12039), .ZN(n12040) );
  OAI211_X1 U14592 ( .C1(n12042), .C2(n15815), .A(n12041), .B(n12040), .ZN(
        n12045) );
  NAND2_X1 U14593 ( .A1(n12045), .A2(n15838), .ZN(n12043) );
  OAI21_X1 U14594 ( .B1(n15838), .B2(n12044), .A(n12043), .ZN(P1_U3486) );
  NAND2_X1 U14595 ( .A1(n12045), .A2(n15850), .ZN(n12046) );
  OAI21_X1 U14596 ( .B1(n15850), .B2(n11068), .A(n12046), .ZN(P1_U3537) );
  NAND2_X1 U14597 ( .A1(n14180), .A2(n14658), .ZN(n14164) );
  INV_X1 U14598 ( .A(n14164), .ZN(n14179) );
  INV_X1 U14599 ( .A(n12047), .ZN(n12048) );
  AOI22_X1 U14600 ( .A1(n14179), .A2(n14213), .B1(n14180), .B2(n12048), .ZN(
        n12050) );
  NOR2_X1 U14601 ( .A1(n12050), .A2(n12049), .ZN(n12055) );
  OAI22_X1 U14602 ( .A1(n12179), .A2(n14185), .B1(n14184), .B2(n12336), .ZN(
        n12054) );
  NAND2_X1 U14603 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n15870) );
  INV_X1 U14604 ( .A(n12188), .ZN(n12051) );
  NAND2_X1 U14605 ( .A1(n14168), .A2(n12051), .ZN(n12052) );
  OAI211_X1 U14606 ( .C1(n14173), .C2(n12412), .A(n15870), .B(n12052), .ZN(
        n12053) );
  AOI211_X1 U14607 ( .C1(n12055), .C2(n14108), .A(n12054), .B(n12053), .ZN(
        n12056) );
  OAI21_X1 U14608 ( .B1(n12057), .B2(n14154), .A(n12056), .ZN(P2_U3199) );
  AOI21_X1 U14609 ( .B1(n13430), .B2(n13456), .A(n12058), .ZN(n12061) );
  OR2_X1 U14610 ( .A1(n13428), .A2(n12059), .ZN(n12060) );
  OAI211_X1 U14611 ( .C1(n13446), .C2(n12062), .A(n12061), .B(n12060), .ZN(
        n12066) );
  XNOR2_X1 U14612 ( .A(n6757), .B(n12063), .ZN(n12064) );
  NOR2_X1 U14613 ( .A1(n12064), .A2(n13413), .ZN(n12065) );
  AOI211_X1 U14614 ( .C1(n15949), .C2(n13443), .A(n12066), .B(n12065), .ZN(
        n12067) );
  INV_X1 U14615 ( .A(n12067), .ZN(P3_U3153) );
  INV_X1 U14616 ( .A(n13408), .ZN(n12490) );
  INV_X1 U14617 ( .A(n13454), .ZN(n13342) );
  AND2_X1 U14618 ( .A1(n12490), .A2(n13342), .ZN(n12529) );
  INV_X1 U14619 ( .A(n12529), .ZN(n13056) );
  NAND2_X1 U14620 ( .A1(n13408), .A2(n13454), .ZN(n13060) );
  NAND2_X1 U14621 ( .A1(n13056), .A2(n13060), .ZN(n13055) );
  NAND2_X1 U14622 ( .A1(n13308), .A2(n13455), .ZN(n12526) );
  NAND2_X1 U14623 ( .A1(n12527), .A2(n12526), .ZN(n12068) );
  NOR2_X1 U14624 ( .A1(n12068), .A2(n13055), .ZN(n12488) );
  AOI21_X1 U14625 ( .B1(n13055), .B2(n12068), .A(n12488), .ZN(n12083) );
  OR2_X1 U14626 ( .A1(n13308), .A2(n13407), .ZN(n12069) );
  INV_X1 U14627 ( .A(n13055), .ZN(n12071) );
  XNOR2_X1 U14628 ( .A(n12492), .B(n12071), .ZN(n12072) );
  NAND2_X1 U14629 ( .A1(n12072), .A2(n13833), .ZN(n12074) );
  AOI22_X1 U14630 ( .A1(n13453), .A2(n13830), .B1(n13828), .B2(n13455), .ZN(
        n12073) );
  NAND2_X1 U14631 ( .A1(n12074), .A2(n12073), .ZN(n12080) );
  AOI22_X1 U14632 ( .A1(n15997), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n15977), 
        .B2(n13411), .ZN(n12075) );
  OAI21_X1 U14633 ( .B1(n13825), .B2(n13408), .A(n12075), .ZN(n12076) );
  AOI21_X1 U14634 ( .B1(n12080), .B2(n15995), .A(n12076), .ZN(n12077) );
  OAI21_X1 U14635 ( .B1(n12083), .B2(n13807), .A(n12077), .ZN(P3_U3222) );
  AOI22_X1 U14636 ( .A1(n12490), .A2(n13893), .B1(P3_REG1_REG_11__SCAN_IN), 
        .B2(n16023), .ZN(n12079) );
  NAND2_X1 U14637 ( .A1(n12080), .A2(n13911), .ZN(n12078) );
  OAI211_X1 U14638 ( .C1(n12083), .C2(n13900), .A(n12079), .B(n12078), .ZN(
        P3_U3470) );
  AOI22_X1 U14639 ( .A1(n13981), .A2(n12490), .B1(P3_REG0_REG_11__SCAN_IN), 
        .B2(n16018), .ZN(n12082) );
  NAND2_X1 U14640 ( .A1(n12080), .A2(n16017), .ZN(n12081) );
  OAI211_X1 U14641 ( .C1(n12083), .C2(n13988), .A(n12082), .B(n12081), .ZN(
        P3_U3423) );
  INV_X2 U14642 ( .A(n10450), .ZN(n14658) );
  AOI211_X1 U14643 ( .C1(n13267), .C2(n12099), .A(n12113), .B(n14658), .ZN(
        n12682) );
  INV_X2 U14644 ( .A(n14360), .ZN(n14672) );
  NOR2_X1 U14645 ( .A1(n14645), .A2(n11029), .ZN(n12098) );
  OAI21_X1 U14646 ( .B1(n12084), .B2(n12091), .A(n12107), .ZN(n12088) );
  OAI22_X1 U14647 ( .A1(n12086), .A2(n14636), .B1(n14638), .B2(n12085), .ZN(
        n12087) );
  AOI21_X1 U14648 ( .B1(n12088), .B2(n14657), .A(n12087), .ZN(n12095) );
  INV_X1 U14649 ( .A(n12089), .ZN(n12090) );
  NAND2_X1 U14650 ( .A1(n12091), .A2(n12090), .ZN(n12092) );
  NAND2_X1 U14651 ( .A1(n12093), .A2(n12092), .ZN(n12684) );
  NAND2_X1 U14652 ( .A1(n12684), .A2(n14547), .ZN(n12094) );
  NAND2_X1 U14653 ( .A1(n12095), .A2(n12094), .ZN(n12683) );
  NAND2_X1 U14654 ( .A1(n14645), .A2(n12683), .ZN(n12096) );
  OAI21_X1 U14655 ( .B1(n7530), .B2(n14642), .A(n12096), .ZN(n12097) );
  AOI211_X1 U14656 ( .C1(n12682), .C2(n14672), .A(n12098), .B(n12097), .ZN(
        n12101) );
  AOI22_X1 U14657 ( .A1(n12112), .A2(n12684), .B1(n14433), .B2(n12099), .ZN(
        n12100) );
  NAND2_X1 U14658 ( .A1(n12101), .A2(n12100), .ZN(P2_U3264) );
  INV_X2 U14659 ( .A(n14645), .ZN(n14674) );
  INV_X1 U14660 ( .A(n12102), .ZN(n12106) );
  NAND2_X1 U14661 ( .A1(n12103), .A2(n12106), .ZN(n12249) );
  OAI21_X1 U14662 ( .B1(n12103), .B2(n12106), .A(n12249), .ZN(n15921) );
  OAI22_X1 U14663 ( .A1(n12104), .A2(n14638), .B1(n14636), .B2(n13274), .ZN(
        n12111) );
  NAND3_X1 U14664 ( .A1(n12107), .A2(n12106), .A3(n12105), .ZN(n12108) );
  AOI21_X1 U14665 ( .B1(n12109), .B2(n12108), .A(n14634), .ZN(n12110) );
  AOI211_X1 U14666 ( .C1(n14547), .C2(n15921), .A(n12111), .B(n12110), .ZN(
        n15918) );
  AOI22_X1 U14667 ( .A1(n12112), .A2(n15921), .B1(n14433), .B2(n12114), .ZN(
        n12120) );
  INV_X1 U14668 ( .A(n12113), .ZN(n12115) );
  NAND2_X1 U14669 ( .A1(n12115), .A2(n12114), .ZN(n12116) );
  AND3_X1 U14670 ( .A1(n10450), .A2(n12251), .A3(n12116), .ZN(n15915) );
  OAI22_X1 U14671 ( .A1(n14645), .A2(n11028), .B1(n12117), .B2(n14642), .ZN(
        n12118) );
  AOI21_X1 U14672 ( .B1(n14672), .B2(n15915), .A(n12118), .ZN(n12119) );
  OAI211_X1 U14673 ( .C1(n14674), .C2(n15918), .A(n12120), .B(n12119), .ZN(
        P2_U3263) );
  INV_X1 U14674 ( .A(n12125), .ZN(n12124) );
  INV_X1 U14675 ( .A(n12123), .ZN(n12121) );
  NOR2_X1 U14676 ( .A1(n12121), .A2(n12125), .ZN(n12318) );
  INV_X1 U14677 ( .A(n12318), .ZN(n12122) );
  OAI21_X1 U14678 ( .B1(n12124), .B2(n12123), .A(n12122), .ZN(n12309) );
  INV_X1 U14679 ( .A(n12309), .ZN(n12134) );
  XOR2_X1 U14680 ( .A(n12126), .B(n12125), .Z(n12127) );
  AOI22_X1 U14681 ( .A1(n14654), .A2(n14209), .B1(n14652), .B2(n14211), .ZN(
        n12340) );
  OAI21_X1 U14682 ( .B1(n12127), .B2(n14634), .A(n12340), .ZN(n12307) );
  INV_X1 U14683 ( .A(n12307), .ZN(n12128) );
  MUX2_X1 U14684 ( .A(n12129), .B(n12128), .S(n14645), .Z(n12133) );
  AOI211_X1 U14685 ( .C1(n12342), .C2(n12130), .A(n14658), .B(n12321), .ZN(
        n12308) );
  OAI22_X1 U14686 ( .A1(n14664), .A2(n12398), .B1(n14642), .B2(n12345), .ZN(
        n12131) );
  AOI21_X1 U14687 ( .B1(n14672), .B2(n12308), .A(n12131), .ZN(n12132) );
  OAI211_X1 U14688 ( .C1(n14669), .C2(n12134), .A(n12133), .B(n12132), .ZN(
        P2_U3258) );
  INV_X1 U14689 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n13466) );
  AOI22_X1 U14690 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n13467), .B1(n13475), 
        .B2(n13466), .ZN(n12140) );
  INV_X1 U14691 ( .A(n12135), .ZN(n12136) );
  NAND2_X1 U14692 ( .A1(n12136), .A2(n12145), .ZN(n12138) );
  NAND2_X1 U14693 ( .A1(n12138), .A2(n12137), .ZN(n12139) );
  OAI21_X1 U14694 ( .B1(n12140), .B2(n12139), .A(n13465), .ZN(n12155) );
  NAND3_X1 U14695 ( .A1(n12142), .A2(n6780), .A3(n12141), .ZN(n12144) );
  AOI21_X1 U14696 ( .B1(n13469), .B2(n12144), .A(n12143), .ZN(n12154) );
  NOR2_X1 U14697 ( .A1(n12146), .A2(n12145), .ZN(n12148) );
  MUX2_X1 U14698 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n13576), .Z(n13474) );
  XNOR2_X1 U14699 ( .A(n13474), .B(n13467), .ZN(n12147) );
  OAI21_X1 U14700 ( .B1(n12149), .B2(n12148), .A(n12147), .ZN(n12150) );
  NAND3_X1 U14701 ( .A1(n7352), .A2(n13503), .A3(n12150), .ZN(n12152) );
  AND2_X1 U14702 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n13339) );
  AOI21_X1 U14703 ( .B1(n15945), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n13339), 
        .ZN(n12151) );
  OAI211_X1 U14704 ( .C1(n13586), .C2(n13467), .A(n12152), .B(n12151), .ZN(
        n12153) );
  AOI211_X1 U14705 ( .C1(n12155), .C2(n13589), .A(n12154), .B(n12153), .ZN(
        n12156) );
  INV_X1 U14706 ( .A(n12156), .ZN(P3_U3194) );
  NAND2_X1 U14707 ( .A1(n15828), .A2(n15012), .ZN(n12157) );
  NAND2_X1 U14708 ( .A1(n12158), .A2(n12157), .ZN(n12161) );
  INV_X1 U14709 ( .A(n12161), .ZN(n12159) );
  AOI21_X1 U14710 ( .B1(n12159), .B2(n12173), .A(n15829), .ZN(n12164) );
  NAND2_X1 U14711 ( .A1(n12161), .A2(n12160), .ZN(n12381) );
  NAND2_X1 U14712 ( .A1(n15746), .A2(n15010), .ZN(n12163) );
  NAND2_X1 U14713 ( .A1(n15426), .A2(n15012), .ZN(n12162) );
  NAND2_X1 U14714 ( .A1(n12163), .A2(n12162), .ZN(n14959) );
  AOI21_X1 U14715 ( .B1(n12164), .B2(n12381), .A(n14959), .ZN(n15561) );
  INV_X1 U14716 ( .A(n12165), .ZN(n12167) );
  INV_X1 U14717 ( .A(n15559), .ZN(n14964) );
  INV_X1 U14718 ( .A(n12387), .ZN(n12166) );
  AOI211_X1 U14719 ( .C1(n15559), .C2(n12167), .A(n15742), .B(n12166), .ZN(
        n15558) );
  NOR2_X1 U14720 ( .A1(n14964), .A2(n15418), .ZN(n12169) );
  OAI22_X1 U14721 ( .A1(n6544), .A2(n11077), .B1(n14956), .B2(n15393), .ZN(
        n12168) );
  AOI211_X1 U14722 ( .C1(n15558), .C2(n15732), .A(n12169), .B(n12168), .ZN(
        n12176) );
  NAND2_X1 U14723 ( .A1(n15828), .A2(n12170), .ZN(n12171) );
  NAND2_X1 U14724 ( .A1(n12172), .A2(n12171), .ZN(n12174) );
  NAND2_X1 U14725 ( .A1(n12174), .A2(n12173), .ZN(n12376) );
  OAI21_X1 U14726 ( .B1(n12174), .B2(n12173), .A(n12376), .ZN(n15557) );
  NAND2_X1 U14727 ( .A1(n15557), .A2(n15383), .ZN(n12175) );
  OAI211_X1 U14728 ( .C1(n15561), .C2(n15764), .A(n12176), .B(n12175), .ZN(
        P1_U3282) );
  OAI21_X1 U14729 ( .B1(n12178), .B2(n12181), .A(n12177), .ZN(n12314) );
  INV_X1 U14730 ( .A(n12314), .ZN(n12192) );
  OAI22_X1 U14731 ( .A1(n12179), .A2(n14636), .B1(n14638), .B2(n12336), .ZN(
        n12184) );
  NAND3_X1 U14732 ( .A1(n11989), .A2(n12181), .A3(n12180), .ZN(n12182) );
  AOI21_X1 U14733 ( .B1(n11969), .B2(n12182), .A(n14634), .ZN(n12183) );
  AOI211_X1 U14734 ( .C1(n14547), .C2(n12314), .A(n12184), .B(n12183), .ZN(
        n12311) );
  MUX2_X1 U14735 ( .A(n12185), .B(n12311), .S(n14645), .Z(n12191) );
  AOI211_X1 U14736 ( .C1(n12315), .C2(n12187), .A(n14658), .B(n7615), .ZN(
        n12313) );
  OAI22_X1 U14737 ( .A1(n14664), .A2(n12412), .B1(n14642), .B2(n12188), .ZN(
        n12189) );
  AOI21_X1 U14738 ( .B1(n14672), .B2(n12313), .A(n12189), .ZN(n12190) );
  OAI211_X1 U14739 ( .C1(n12192), .C2(n14554), .A(n12191), .B(n12190), .ZN(
        P2_U3260) );
  OAI21_X1 U14740 ( .B1(n12194), .B2(n12193), .A(n13297), .ZN(n12195) );
  NAND2_X1 U14741 ( .A1(n12195), .A2(n13437), .ZN(n12202) );
  AOI21_X1 U14742 ( .B1(n13455), .B2(n13430), .A(n12196), .ZN(n12197) );
  OAI21_X1 U14743 ( .B1(n12198), .B2(n13428), .A(n12197), .ZN(n12199) );
  AOI21_X1 U14744 ( .B1(n12200), .B2(n13443), .A(n12199), .ZN(n12201) );
  OAI211_X1 U14745 ( .C1(n13446), .C2(n12203), .A(n12202), .B(n12201), .ZN(
        P3_U3171) );
  NAND2_X1 U14746 ( .A1(n12204), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n12207) );
  NAND2_X1 U14747 ( .A1(n12205), .A2(n12210), .ZN(n12206) );
  NAND2_X1 U14748 ( .A1(n12207), .A2(n12206), .ZN(n14283) );
  XNOR2_X1 U14749 ( .A(n14291), .B(n14583), .ZN(n14282) );
  XNOR2_X1 U14750 ( .A(n14283), .B(n14282), .ZN(n12219) );
  NAND2_X1 U14751 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n14088)
         );
  OAI21_X1 U14752 ( .B1(n14306), .B2(n12208), .A(n14088), .ZN(n12209) );
  AOI21_X1 U14753 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(n15851), .A(n12209), 
        .ZN(n12218) );
  NAND2_X1 U14754 ( .A1(n12211), .A2(n12210), .ZN(n12212) );
  NAND2_X1 U14755 ( .A1(n12213), .A2(n12212), .ZN(n12216) );
  INV_X1 U14756 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n12214) );
  XNOR2_X1 U14757 ( .A(n14291), .B(n12214), .ZN(n12215) );
  NAND2_X1 U14758 ( .A1(n12216), .A2(n12215), .ZN(n14293) );
  OAI211_X1 U14759 ( .C1(n12216), .C2(n12215), .A(n14293), .B(n15896), .ZN(
        n12217) );
  OAI211_X1 U14760 ( .C1(n12219), .C2(n14330), .A(n12218), .B(n12217), .ZN(
        P2_U3230) );
  INV_X1 U14761 ( .A(n12220), .ZN(n12224) );
  OAI222_X1 U14762 ( .A1(P1_U3086), .A2(n12222), .B1(n15595), .B2(n12224), 
        .C1(n12221), .C2(n15597), .ZN(P1_U3331) );
  OAI222_X1 U14763 ( .A1(P2_U3088), .A2(n12225), .B1(n12909), .B2(n12224), 
        .C1(n12223), .C2(n14826), .ZN(P2_U3303) );
  NAND2_X1 U14764 ( .A1(n12939), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n12228) );
  NAND2_X1 U14765 ( .A1(n12938), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n12227) );
  OAI211_X1 U14766 ( .C1(n6545), .C2(n12883), .A(n12228), .B(n12227), .ZN(
        n12229) );
  INV_X1 U14767 ( .A(n12229), .ZN(n12230) );
  NAND2_X1 U14768 ( .A1(n13463), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n12231) );
  OAI21_X1 U14769 ( .B1(n13640), .B2(n13463), .A(n12231), .ZN(P3_U3520) );
  NOR2_X1 U14770 ( .A1(n12232), .A2(n12236), .ZN(n12499) );
  AOI21_X1 U14771 ( .B1(n12232), .B2(n12236), .A(n12499), .ZN(n12513) );
  NAND2_X1 U14772 ( .A1(n12233), .A2(n12275), .ZN(n12269) );
  NAND2_X1 U14773 ( .A1(n12269), .A2(n12234), .ZN(n12237) );
  OAI211_X1 U14774 ( .C1(n12237), .C2(n12236), .A(n12235), .B(n14657), .ZN(
        n12240) );
  NAND2_X1 U14775 ( .A1(n14652), .A2(n14208), .ZN(n12239) );
  NAND2_X1 U14776 ( .A1(n14654), .A2(n14653), .ZN(n12238) );
  AND2_X1 U14777 ( .A1(n12239), .A2(n12238), .ZN(n12662) );
  NAND2_X1 U14778 ( .A1(n12240), .A2(n12662), .ZN(n12514) );
  NAND2_X1 U14779 ( .A1(n12514), .A2(n14645), .ZN(n12247) );
  INV_X1 U14780 ( .A(n12241), .ZN(n12278) );
  AOI211_X1 U14781 ( .C1(n12242), .C2(n12278), .A(n14658), .B(n12506), .ZN(
        n12515) );
  INV_X1 U14782 ( .A(n12243), .ZN(n12664) );
  AOI22_X1 U14783 ( .A1(n14674), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n12664), 
        .B2(n14661), .ZN(n12244) );
  OAI21_X1 U14784 ( .B1(n9865), .B2(n14664), .A(n12244), .ZN(n12245) );
  AOI21_X1 U14785 ( .B1(n12515), .B2(n14672), .A(n12245), .ZN(n12246) );
  OAI211_X1 U14786 ( .C1(n14669), .C2(n12513), .A(n12247), .B(n12246), .ZN(
        P2_U3255) );
  NAND2_X1 U14787 ( .A1(n12249), .A2(n12248), .ZN(n12250) );
  NAND2_X1 U14788 ( .A1(n10450), .A2(n12252), .ZN(n12253) );
  NOR2_X1 U14789 ( .A1(n11996), .A2(n12253), .ZN(n12303) );
  NAND2_X1 U14790 ( .A1(n11990), .A2(n12255), .ZN(n12256) );
  NAND2_X1 U14791 ( .A1(n12256), .A2(n14657), .ZN(n12300) );
  OAI211_X1 U14792 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n14642), .A(n12300), .B(
        n12301), .ZN(n12257) );
  MUX2_X1 U14793 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n12257), .S(n14645), .Z(
        n12258) );
  INV_X1 U14794 ( .A(n12258), .ZN(n12259) );
  OAI211_X1 U14795 ( .C1(n14669), .C2(n12299), .A(n12260), .B(n12259), .ZN(
        P2_U3262) );
  INV_X1 U14796 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n12265) );
  NAND2_X1 U14797 ( .A1(n12939), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n12263) );
  NAND2_X1 U14798 ( .A1(n12261), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n12262) );
  OAI211_X1 U14799 ( .C1(n12265), .C2(n12264), .A(n12263), .B(n12262), .ZN(
        n12266) );
  INV_X1 U14800 ( .A(n12266), .ZN(n12267) );
  NAND2_X1 U14801 ( .A1(n13463), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n12268) );
  OAI21_X1 U14802 ( .B1(n12958), .B2(n13463), .A(n12268), .ZN(P3_U3521) );
  OAI211_X1 U14803 ( .C1(n12233), .C2(n12275), .A(n12269), .B(n14657), .ZN(
        n12272) );
  NAND2_X1 U14804 ( .A1(n14654), .A2(n14207), .ZN(n12271) );
  NAND2_X1 U14805 ( .A1(n14652), .A2(n14209), .ZN(n12270) );
  AND2_X1 U14806 ( .A1(n12271), .A2(n12270), .ZN(n12464) );
  NAND2_X1 U14807 ( .A1(n12272), .A2(n12464), .ZN(n12367) );
  INV_X1 U14808 ( .A(n12367), .ZN(n12284) );
  NAND2_X1 U14809 ( .A1(n12274), .A2(n12273), .ZN(n12276) );
  XNOR2_X1 U14810 ( .A(n12276), .B(n12275), .ZN(n12369) );
  INV_X1 U14811 ( .A(n14669), .ZN(n14588) );
  AOI21_X1 U14812 ( .B1(n12277), .B2(n12468), .A(n14658), .ZN(n12279) );
  NAND2_X1 U14813 ( .A1(n12279), .A2(n12278), .ZN(n12365) );
  OAI22_X1 U14814 ( .A1(n14645), .A2(n11043), .B1(n12465), .B2(n14642), .ZN(
        n12280) );
  AOI21_X1 U14815 ( .B1(n14433), .B2(n12468), .A(n12280), .ZN(n12281) );
  OAI21_X1 U14816 ( .B1(n14360), .B2(n12365), .A(n12281), .ZN(n12282) );
  AOI21_X1 U14817 ( .B1(n12369), .B2(n14588), .A(n12282), .ZN(n12283) );
  OAI21_X1 U14818 ( .B1(n12284), .B2(n14674), .A(n12283), .ZN(P2_U3256) );
  INV_X1 U14819 ( .A(n12285), .ZN(n12287) );
  OAI222_X1 U14820 ( .A1(P3_U3151), .A2(n12288), .B1(n13257), .B2(n12287), 
        .C1(n14006), .C2(n12286), .ZN(P3_U3269) );
  INV_X1 U14821 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15901) );
  NAND2_X1 U14822 ( .A1(n12292), .A2(n12291), .ZN(n12294) );
  NAND2_X1 U14823 ( .A1(n15715), .A2(P3_ADDR_REG_12__SCAN_IN), .ZN(n12293) );
  NAND2_X1 U14824 ( .A1(n12294), .A2(n12293), .ZN(n12585) );
  XNOR2_X1 U14825 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n12584) );
  INV_X1 U14826 ( .A(n12584), .ZN(n12295) );
  XNOR2_X1 U14827 ( .A(n12585), .B(n12295), .ZN(n12296) );
  NAND2_X1 U14828 ( .A1(n12297), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n12298) );
  NAND2_X1 U14829 ( .A1(n12583), .A2(n12298), .ZN(SUB_1596_U67) );
  NOR2_X1 U14830 ( .A1(n12299), .A2(n14774), .ZN(n12305) );
  INV_X1 U14831 ( .A(n12300), .ZN(n12304) );
  INV_X1 U14832 ( .A(n12301), .ZN(n12302) );
  NOR4_X1 U14833 ( .A1(n12305), .A2(n12304), .A3(n12303), .A4(n12302), .ZN(
        n12410) );
  OAI21_X1 U14834 ( .B1(n12410), .B2(n15941), .A(n12306), .ZN(P2_U3502) );
  AOI211_X1 U14835 ( .C1(n15929), .C2(n12309), .A(n12308), .B(n12307), .ZN(
        n12401) );
  AOI22_X1 U14836 ( .A1(n14682), .A2(n12342), .B1(n15941), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n12310) );
  OAI21_X1 U14837 ( .B1(n12401), .B2(n15941), .A(n12310), .ZN(P2_U3506) );
  INV_X1 U14838 ( .A(n10166), .ZN(n15937) );
  INV_X1 U14839 ( .A(n12311), .ZN(n12312) );
  AOI211_X1 U14840 ( .C1(n15937), .C2(n12314), .A(n12313), .B(n12312), .ZN(
        n12415) );
  AOI22_X1 U14841 ( .A1(n14682), .A2(n12315), .B1(n15941), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n12316) );
  OAI21_X1 U14842 ( .B1(n12415), .B2(n15941), .A(n12316), .ZN(P2_U3504) );
  NOR2_X1 U14843 ( .A1(n12318), .A2(n12317), .ZN(n12320) );
  XNOR2_X1 U14844 ( .A(n12320), .B(n12319), .ZN(n12362) );
  INV_X1 U14845 ( .A(n12321), .ZN(n12323) );
  INV_X1 U14846 ( .A(n12277), .ZN(n12322) );
  AOI211_X1 U14847 ( .C1(n12331), .C2(n12323), .A(n14658), .B(n12322), .ZN(
        n12357) );
  INV_X1 U14848 ( .A(n12324), .ZN(n12325) );
  AOI211_X1 U14849 ( .C1(n12327), .C2(n12326), .A(n14634), .B(n12325), .ZN(
        n12330) );
  NAND2_X1 U14850 ( .A1(n14652), .A2(n14210), .ZN(n12328) );
  OAI21_X1 U14851 ( .B1(n12329), .B2(n14638), .A(n12328), .ZN(n12551) );
  OR2_X1 U14852 ( .A1(n12330), .A2(n12551), .ZN(n12356) );
  AOI211_X1 U14853 ( .C1(n12362), .C2(n15929), .A(n12357), .B(n12356), .ZN(
        n12405) );
  AOI22_X1 U14854 ( .A1(n14682), .A2(n12331), .B1(n15941), .B2(
        P2_REG1_REG_8__SCAN_IN), .ZN(n12332) );
  OAI21_X1 U14855 ( .B1(n12405), .B2(n15941), .A(n12332), .ZN(P2_U3507) );
  INV_X1 U14856 ( .A(n12333), .ZN(n12334) );
  AOI21_X1 U14857 ( .B1(n12346), .B2(n12334), .A(n14154), .ZN(n12338) );
  NOR3_X1 U14858 ( .A1(n14164), .A2(n12336), .A3(n12335), .ZN(n12337) );
  OAI21_X1 U14859 ( .B1(n12338), .B2(n12337), .A(n12546), .ZN(n12344) );
  OAI22_X1 U14860 ( .A1(n14147), .A2(n12340), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12339), .ZN(n12341) );
  AOI21_X1 U14861 ( .B1(n14189), .B2(n12342), .A(n12341), .ZN(n12343) );
  OAI211_X1 U14862 ( .C1(n14186), .C2(n12345), .A(n12344), .B(n12343), .ZN(
        P2_U3185) );
  INV_X1 U14863 ( .A(n12346), .ZN(n12347) );
  AOI211_X1 U14864 ( .C1(n12349), .C2(n12348), .A(n14154), .B(n12347), .ZN(
        n12355) );
  OAI22_X1 U14865 ( .A1(n12548), .A2(n14184), .B1(n14185), .B2(n14104), .ZN(
        n12354) );
  NAND2_X1 U14866 ( .A1(n14189), .A2(n12350), .ZN(n12351) );
  NAND2_X1 U14867 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n14255) );
  OAI211_X1 U14868 ( .C1(n14186), .C2(n12352), .A(n12351), .B(n14255), .ZN(
        n12353) );
  OR3_X1 U14869 ( .A1(n12355), .A2(n12354), .A3(n12353), .ZN(P2_U3211) );
  INV_X1 U14870 ( .A(n12356), .ZN(n12364) );
  NAND2_X1 U14871 ( .A1(n12357), .A2(n14672), .ZN(n12360) );
  INV_X1 U14872 ( .A(n12358), .ZN(n12558) );
  AOI22_X1 U14873 ( .A1(n14674), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n12558), 
        .B2(n14661), .ZN(n12359) );
  OAI211_X1 U14874 ( .C1(n12554), .C2(n14664), .A(n12360), .B(n12359), .ZN(
        n12361) );
  AOI21_X1 U14875 ( .B1(n12362), .B2(n14588), .A(n12361), .ZN(n12363) );
  OAI21_X1 U14876 ( .B1(n12364), .B2(n14674), .A(n12363), .ZN(P2_U3257) );
  OAI21_X1 U14877 ( .B1(n12366), .B2(n15931), .A(n12365), .ZN(n12368) );
  AOI211_X1 U14878 ( .C1(n15929), .C2(n12369), .A(n12368), .B(n12367), .ZN(
        n12374) );
  NAND2_X1 U14879 ( .A1(n15941), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n12370) );
  OAI21_X1 U14880 ( .B1(n12374), .B2(n15941), .A(n12370), .ZN(P2_U3508) );
  NOR2_X4 U14881 ( .A1(n12372), .A2(n12371), .ZN(n14818) );
  NAND2_X1 U14882 ( .A1(n15938), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n12373) );
  OAI21_X1 U14883 ( .B1(n12374), .B2(n15938), .A(n12373), .ZN(P2_U3457) );
  OR2_X1 U14884 ( .A1(n15559), .A2(n15011), .ZN(n12375) );
  NAND2_X1 U14885 ( .A1(n12376), .A2(n12375), .ZN(n12378) );
  NAND2_X1 U14886 ( .A1(n12378), .A2(n12377), .ZN(n12601) );
  OR2_X1 U14887 ( .A1(n12378), .A2(n12377), .ZN(n12379) );
  NAND2_X1 U14888 ( .A1(n12601), .A2(n12379), .ZN(n12536) );
  INV_X1 U14889 ( .A(n12536), .ZN(n12393) );
  INV_X1 U14890 ( .A(n15011), .ZN(n14892) );
  OR2_X1 U14891 ( .A1(n15559), .A2(n14892), .ZN(n12380) );
  NAND2_X1 U14892 ( .A1(n12381), .A2(n12380), .ZN(n12383) );
  NAND2_X1 U14893 ( .A1(n12383), .A2(n12382), .ZN(n12607) );
  OAI211_X1 U14894 ( .C1(n12383), .C2(n12382), .A(n12607), .B(n15754), .ZN(
        n12385) );
  AOI22_X1 U14895 ( .A1(n15426), .A2(n15011), .B1(n15746), .B2(n15009), .ZN(
        n12384) );
  NAND2_X1 U14896 ( .A1(n12385), .A2(n12384), .ZN(n12540) );
  NAND2_X1 U14897 ( .A1(n12540), .A2(n6544), .ZN(n12392) );
  OAI22_X1 U14898 ( .A1(n6544), .A2(n12386), .B1(n14893), .B2(n15393), .ZN(
        n12390) );
  AOI21_X1 U14899 ( .B1(n12387), .B2(n12605), .A(n15742), .ZN(n12388) );
  NAND2_X1 U14900 ( .A1(n12388), .A2(n12617), .ZN(n12537) );
  NOR2_X1 U14901 ( .A1(n12537), .A2(n15304), .ZN(n12389) );
  AOI211_X1 U14902 ( .C1(n15730), .C2(n12605), .A(n12390), .B(n12389), .ZN(
        n12391) );
  OAI211_X1 U14903 ( .C1(n15423), .C2(n12393), .A(n12392), .B(n12391), .ZN(
        P1_U3281) );
  INV_X1 U14904 ( .A(n12394), .ZN(n12396) );
  OAI222_X1 U14905 ( .A1(n13576), .A2(P3_U3151), .B1(n13257), .B2(n12396), 
        .C1(n12395), .C2(n14006), .ZN(P3_U3268) );
  OAI22_X1 U14906 ( .A1(n14822), .A2(n12398), .B1(n14818), .B2(n12397), .ZN(
        n12399) );
  INV_X1 U14907 ( .A(n12399), .ZN(n12400) );
  OAI21_X1 U14908 ( .B1(n12401), .B2(n15938), .A(n12400), .ZN(P2_U3451) );
  OAI22_X1 U14909 ( .A1(n14822), .A2(n12554), .B1(n14818), .B2(n12402), .ZN(
        n12403) );
  INV_X1 U14910 ( .A(n12403), .ZN(n12404) );
  OAI21_X1 U14911 ( .B1(n12405), .B2(n15938), .A(n12404), .ZN(P2_U3454) );
  INV_X1 U14912 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n12406) );
  OAI22_X1 U14913 ( .A1(n14822), .A2(n12407), .B1(n14818), .B2(n12406), .ZN(
        n12408) );
  INV_X1 U14914 ( .A(n12408), .ZN(n12409) );
  OAI21_X1 U14915 ( .B1(n12410), .B2(n15938), .A(n12409), .ZN(P2_U3439) );
  INV_X1 U14916 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n12411) );
  OAI22_X1 U14917 ( .A1(n14822), .A2(n12412), .B1(n14818), .B2(n12411), .ZN(
        n12413) );
  INV_X1 U14918 ( .A(n12413), .ZN(n12414) );
  OAI21_X1 U14919 ( .B1(n12415), .B2(n15938), .A(n12414), .ZN(P2_U3445) );
  NAND2_X1 U14920 ( .A1(n15559), .A2(n10876), .ZN(n12419) );
  NAND2_X1 U14921 ( .A1(n13189), .A2(n15011), .ZN(n12418) );
  NAND2_X1 U14922 ( .A1(n12419), .A2(n12418), .ZN(n12420) );
  XNOR2_X1 U14923 ( .A(n12420), .B(n11908), .ZN(n14884) );
  NAND2_X1 U14924 ( .A1(n15559), .A2(n13189), .ZN(n12422) );
  NAND2_X1 U14925 ( .A1(n13235), .A2(n15011), .ZN(n12421) );
  NAND2_X1 U14926 ( .A1(n12422), .A2(n12421), .ZN(n14883) );
  NAND2_X1 U14927 ( .A1(n14884), .A2(n14883), .ZN(n12436) );
  NAND2_X1 U14928 ( .A1(n12426), .A2(n10876), .ZN(n12424) );
  NAND2_X1 U14929 ( .A1(n13189), .A2(n15012), .ZN(n12423) );
  NAND2_X1 U14930 ( .A1(n12424), .A2(n12423), .ZN(n12425) );
  XNOR2_X1 U14931 ( .A(n12425), .B(n11908), .ZN(n12572) );
  NAND2_X1 U14932 ( .A1(n12426), .A2(n13189), .ZN(n12428) );
  NAND2_X1 U14933 ( .A1(n13235), .A2(n15012), .ZN(n12427) );
  NAND2_X1 U14934 ( .A1(n12428), .A2(n12427), .ZN(n12571) );
  NAND2_X1 U14935 ( .A1(n12572), .A2(n12571), .ZN(n14952) );
  NAND2_X1 U14936 ( .A1(n12655), .A2(n10876), .ZN(n12430) );
  NAND2_X1 U14937 ( .A1(n15013), .A2(n13189), .ZN(n12429) );
  NAND2_X1 U14938 ( .A1(n12430), .A2(n12429), .ZN(n12431) );
  XNOR2_X1 U14939 ( .A(n12431), .B(n11908), .ZN(n12650) );
  NAND2_X1 U14940 ( .A1(n12655), .A2(n13189), .ZN(n12434) );
  OR2_X1 U14941 ( .A1(n13223), .A2(n12432), .ZN(n12433) );
  NAND2_X1 U14942 ( .A1(n12434), .A2(n12433), .ZN(n12569) );
  NAND2_X1 U14943 ( .A1(n12650), .A2(n12569), .ZN(n12435) );
  INV_X1 U14944 ( .A(n12569), .ZN(n12567) );
  INV_X1 U14945 ( .A(n12571), .ZN(n12439) );
  INV_X1 U14946 ( .A(n12437), .ZN(n12438) );
  NAND2_X1 U14947 ( .A1(n12439), .A2(n12438), .ZN(n12440) );
  NAND2_X1 U14948 ( .A1(n12441), .A2(n12440), .ZN(n12442) );
  INV_X1 U14949 ( .A(n14883), .ZN(n14887) );
  INV_X1 U14950 ( .A(n14884), .ZN(n14888) );
  NAND2_X1 U14951 ( .A1(n12605), .A2(n10876), .ZN(n12444) );
  NAND2_X1 U14952 ( .A1(n13189), .A2(n15010), .ZN(n12443) );
  NAND2_X1 U14953 ( .A1(n12444), .A2(n12443), .ZN(n12445) );
  XNOR2_X1 U14954 ( .A(n12445), .B(n11908), .ZN(n12451) );
  INV_X1 U14955 ( .A(n15010), .ZN(n12604) );
  NOR2_X1 U14956 ( .A1(n13223), .A2(n12604), .ZN(n12446) );
  AOI21_X1 U14957 ( .B1(n12605), .B2(n13189), .A(n12446), .ZN(n12449) );
  XNOR2_X1 U14958 ( .A(n12451), .B(n12449), .ZN(n14890) );
  INV_X1 U14959 ( .A(n12449), .ZN(n12450) );
  NAND2_X1 U14960 ( .A1(n12451), .A2(n12450), .ZN(n12452) );
  NAND2_X1 U14961 ( .A1(n15553), .A2(n10876), .ZN(n12454) );
  NAND2_X1 U14962 ( .A1(n13189), .A2(n15009), .ZN(n12453) );
  NAND2_X1 U14963 ( .A1(n12454), .A2(n12453), .ZN(n12455) );
  XNOR2_X1 U14964 ( .A(n12455), .B(n11908), .ZN(n12633) );
  NOR2_X1 U14965 ( .A1(n13223), .A2(n15410), .ZN(n12456) );
  AOI21_X1 U14966 ( .B1(n15553), .B2(n13189), .A(n12456), .ZN(n12631) );
  XNOR2_X1 U14967 ( .A(n12633), .B(n12631), .ZN(n12629) );
  XNOR2_X1 U14968 ( .A(n12630), .B(n12629), .ZN(n12462) );
  NAND2_X1 U14969 ( .A1(n15426), .A2(n15010), .ZN(n12458) );
  NAND2_X1 U14970 ( .A1(n15746), .A2(n15008), .ZN(n12457) );
  NAND2_X1 U14971 ( .A1(n12458), .A2(n12457), .ZN(n12612) );
  AOI22_X1 U14972 ( .A1(n14960), .A2(n12612), .B1(P1_REG3_REG_13__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12459) );
  OAI21_X1 U14973 ( .B1(n14988), .B2(n12614), .A(n12459), .ZN(n12460) );
  AOI21_X1 U14974 ( .B1(n15553), .B2(n14992), .A(n12460), .ZN(n12461) );
  OAI21_X1 U14975 ( .B1(n12462), .B2(n14994), .A(n12461), .ZN(P1_U3234) );
  OAI21_X1 U14976 ( .B1(n14147), .B2(n12464), .A(n12463), .ZN(n12467) );
  NOR2_X1 U14977 ( .A1(n14186), .A2(n12465), .ZN(n12466) );
  AOI211_X1 U14978 ( .C1(n12468), .C2(n14189), .A(n12467), .B(n12466), .ZN(
        n12475) );
  INV_X1 U14979 ( .A(n12469), .ZN(n12473) );
  OAI22_X1 U14980 ( .A1(n14164), .A2(n12471), .B1(n12470), .B2(n14154), .ZN(
        n12472) );
  NAND3_X1 U14981 ( .A1(n12555), .A2(n12473), .A3(n12472), .ZN(n12474) );
  OAI211_X1 U14982 ( .C1(n12476), .C2(n14154), .A(n12475), .B(n12474), .ZN(
        P2_U3203) );
  INV_X1 U14983 ( .A(n12477), .ZN(n12481) );
  OAI222_X1 U14984 ( .A1(n14826), .A2(n12479), .B1(n12909), .B2(n12481), .C1(
        P2_U3088), .C2(n12478), .ZN(P2_U3302) );
  OAI222_X1 U14985 ( .A1(n15597), .A2(n12482), .B1(n15595), .B2(n12481), .C1(
        P1_U3086), .C2(n12480), .ZN(P1_U3330) );
  OAI222_X1 U14986 ( .A1(P2_U3088), .A2(n12484), .B1(n12909), .B2(n12486), 
        .C1(n12483), .C2(n14826), .ZN(P2_U3301) );
  OAI222_X1 U14987 ( .A1(P1_U3086), .A2(n12487), .B1(n15595), .B2(n12486), 
        .C1(n12485), .C2(n15597), .ZN(P1_U3329) );
  NOR2_X1 U14988 ( .A1(n12488), .A2(n12529), .ZN(n12489) );
  NAND2_X1 U14989 ( .A1(n13344), .A2(n13388), .ZN(n13067) );
  XNOR2_X1 U14990 ( .A(n12489), .B(n12983), .ZN(n12599) );
  NAND2_X1 U14991 ( .A1(n13408), .A2(n13342), .ZN(n12491) );
  XNOR2_X1 U14992 ( .A(n12523), .B(n12983), .ZN(n12493) );
  INV_X1 U14993 ( .A(n13833), .ZN(n15988) );
  OAI222_X1 U14994 ( .A1(n15992), .A2(n13284), .B1(n15990), .B2(n13342), .C1(
        n12493), .C2(n15988), .ZN(n12596) );
  INV_X1 U14995 ( .A(n12596), .ZN(n12494) );
  MUX2_X1 U14996 ( .A(n12495), .B(n12494), .S(n15995), .Z(n12497) );
  AOI22_X1 U14997 ( .A1(n13344), .A2(n15958), .B1(n15977), .B2(n13338), .ZN(
        n12496) );
  OAI211_X1 U14998 ( .C1(n12599), .C2(n13807), .A(n12497), .B(n12496), .ZN(
        P3_U3221) );
  NOR2_X1 U14999 ( .A1(n12499), .A2(n12498), .ZN(n12500) );
  NAND2_X1 U15000 ( .A1(n12500), .A2(n12504), .ZN(n14666) );
  OAI21_X1 U15001 ( .B1(n12500), .B2(n12504), .A(n14666), .ZN(n14775) );
  INV_X1 U15002 ( .A(n12502), .ZN(n12503) );
  AOI21_X1 U15003 ( .B1(n12504), .B2(n12501), .A(n12503), .ZN(n12505) );
  AOI22_X1 U15004 ( .A1(n14654), .A2(n14206), .B1(n14652), .B2(n14207), .ZN(
        n14146) );
  OAI21_X1 U15005 ( .B1(n12505), .B2(n14634), .A(n14146), .ZN(n14776) );
  NAND2_X1 U15006 ( .A1(n14776), .A2(n14645), .ZN(n12512) );
  INV_X1 U15007 ( .A(n14659), .ZN(n12507) );
  AOI211_X1 U15008 ( .C1(n14151), .C2(n9866), .A(n14658), .B(n12507), .ZN(
        n14777) );
  NOR2_X1 U15009 ( .A1(n14664), .A2(n14823), .ZN(n12510) );
  OAI22_X1 U15010 ( .A1(n14645), .A2(n12508), .B1(n14148), .B2(n14642), .ZN(
        n12509) );
  AOI211_X1 U15011 ( .C1(n14777), .C2(n14672), .A(n12510), .B(n12509), .ZN(
        n12511) );
  OAI211_X1 U15012 ( .C1(n14669), .C2(n14775), .A(n12512), .B(n12511), .ZN(
        P2_U3254) );
  INV_X1 U15013 ( .A(n12513), .ZN(n12516) );
  AOI211_X1 U15014 ( .C1(n15929), .C2(n12516), .A(n12515), .B(n12514), .ZN(
        n12519) );
  MUX2_X1 U15015 ( .A(n12517), .B(n12519), .S(n14818), .Z(n12518) );
  OAI21_X1 U15016 ( .B1(n9865), .B2(n14822), .A(n12518), .ZN(P2_U3460) );
  MUX2_X1 U15017 ( .A(n12520), .B(n12519), .S(n15944), .Z(n12521) );
  OAI21_X1 U15018 ( .B1(n9865), .B2(n14781), .A(n12521), .ZN(P2_U3509) );
  INV_X1 U15019 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n12525) );
  INV_X1 U15020 ( .A(n13344), .ZN(n12522) );
  XNOR2_X1 U15021 ( .A(n13389), .B(n13829), .ZN(n12985) );
  INV_X1 U15022 ( .A(n12985), .ZN(n13065) );
  XNOR2_X1 U15023 ( .A(n12851), .B(n13065), .ZN(n12524) );
  AOI222_X1 U15024 ( .A1(n13833), .A2(n12524), .B1(n13452), .B2(n13830), .C1(
        n13453), .C2(n13828), .ZN(n12563) );
  MUX2_X1 U15025 ( .A(n12525), .B(n12563), .S(n13911), .Z(n12532) );
  INV_X1 U15026 ( .A(n13067), .ZN(n12528) );
  AOI21_X1 U15027 ( .B1(n12983), .B2(n12529), .A(n12528), .ZN(n12530) );
  XNOR2_X1 U15028 ( .A(n12885), .B(n13065), .ZN(n12562) );
  INV_X1 U15029 ( .A(n13389), .ZN(n12850) );
  AOI22_X1 U15030 ( .A1(n12562), .A2(n13902), .B1(n12850), .B2(n13893), .ZN(
        n12531) );
  NAND2_X1 U15031 ( .A1(n12532), .A2(n12531), .ZN(P3_U3472) );
  MUX2_X1 U15032 ( .A(n12533), .B(n12563), .S(n16017), .Z(n12535) );
  AOI22_X1 U15033 ( .A1(n12562), .A2(n13992), .B1(n12850), .B2(n13981), .ZN(
        n12534) );
  NAND2_X1 U15034 ( .A1(n12535), .A2(n12534), .ZN(P3_U3429) );
  INV_X1 U15035 ( .A(n15813), .ZN(n15827) );
  NAND2_X1 U15036 ( .A1(n12536), .A2(n15835), .ZN(n12538) );
  OAI211_X1 U15037 ( .C1(n7830), .C2(n15827), .A(n12538), .B(n12537), .ZN(
        n12539) );
  NOR2_X1 U15038 ( .A1(n12540), .A2(n12539), .ZN(n12543) );
  MUX2_X1 U15039 ( .A(n12541), .B(n12543), .S(n15850), .Z(n12542) );
  INV_X1 U15040 ( .A(n12542), .ZN(P1_U3540) );
  INV_X1 U15041 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n12544) );
  MUX2_X1 U15042 ( .A(n12544), .B(n12543), .S(n15838), .Z(n12545) );
  INV_X1 U15043 ( .A(n12545), .ZN(P1_U3495) );
  INV_X1 U15044 ( .A(n12546), .ZN(n12550) );
  NOR3_X1 U15045 ( .A1(n14164), .A2(n12548), .A3(n12547), .ZN(n12549) );
  AOI21_X1 U15046 ( .B1(n12550), .B2(n14180), .A(n12549), .ZN(n12561) );
  INV_X1 U15047 ( .A(n14147), .ZN(n14170) );
  NAND2_X1 U15048 ( .A1(n14170), .A2(n12551), .ZN(n12553) );
  OAI211_X1 U15049 ( .C1(n14173), .C2(n12554), .A(n12553), .B(n12552), .ZN(
        n12557) );
  NOR2_X1 U15050 ( .A1(n12555), .A2(n14154), .ZN(n12556) );
  AOI211_X1 U15051 ( .C1(n14168), .C2(n12558), .A(n12557), .B(n12556), .ZN(
        n12559) );
  OAI21_X1 U15052 ( .B1(n12561), .B2(n12560), .A(n12559), .ZN(P2_U3193) );
  INV_X1 U15053 ( .A(n12562), .ZN(n12566) );
  MUX2_X1 U15054 ( .A(n7581), .B(n12563), .S(n15995), .Z(n12565) );
  AOI22_X1 U15055 ( .A1(n12850), .A2(n15958), .B1(n15977), .B2(n13392), .ZN(
        n12564) );
  OAI211_X1 U15056 ( .C1(n12566), .C2(n13807), .A(n12565), .B(n12564), .ZN(
        P3_U3220) );
  XNOR2_X1 U15057 ( .A(n12568), .B(n12567), .ZN(n12651) );
  NOR2_X1 U15058 ( .A1(n12651), .A2(n12650), .ZN(n12649) );
  NOR2_X1 U15059 ( .A1(n12570), .A2(n12569), .ZN(n12574) );
  XNOR2_X1 U15060 ( .A(n12572), .B(n12571), .ZN(n12573) );
  NOR3_X1 U15061 ( .A1(n12649), .A2(n12574), .A3(n12573), .ZN(n14886) );
  INV_X1 U15062 ( .A(n14886), .ZN(n14953) );
  OAI21_X1 U15063 ( .B1(n12649), .B2(n12574), .A(n12573), .ZN(n12575) );
  NAND3_X1 U15064 ( .A1(n14953), .A2(n14969), .A3(n12575), .ZN(n12581) );
  INV_X1 U15065 ( .A(n12576), .ZN(n12579) );
  NAND2_X1 U15066 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n15051)
         );
  OAI21_X1 U15067 ( .B1(n14989), .B2(n12577), .A(n15051), .ZN(n12578) );
  AOI21_X1 U15068 ( .B1(n12579), .B2(n14928), .A(n12578), .ZN(n12580) );
  OAI211_X1 U15069 ( .C1(n15828), .C2(n14963), .A(n12581), .B(n12580), .ZN(
        P1_U3217) );
  NAND2_X1 U15070 ( .A1(n12583), .A2(n12582), .ZN(n12591) );
  NAND2_X1 U15071 ( .A1(n12585), .A2(n12584), .ZN(n12588) );
  INV_X1 U15072 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n12586) );
  NAND2_X1 U15073 ( .A1(n12586), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n12587) );
  NAND2_X1 U15074 ( .A1(n12588), .A2(n12587), .ZN(n15613) );
  XNOR2_X1 U15075 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n15612) );
  INV_X1 U15076 ( .A(n15612), .ZN(n12589) );
  XNOR2_X1 U15077 ( .A(n15613), .B(n12589), .ZN(n12590) );
  NAND2_X1 U15078 ( .A1(n12592), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n12593) );
  NAND2_X1 U15079 ( .A1(n15611), .A2(n12593), .ZN(SUB_1596_U66) );
  MUX2_X1 U15080 ( .A(P3_REG1_REG_12__SCAN_IN), .B(n12596), .S(n13911), .Z(
        n12594) );
  AOI21_X1 U15081 ( .B1(n13893), .B2(n13344), .A(n12594), .ZN(n12595) );
  OAI21_X1 U15082 ( .B1(n13900), .B2(n12599), .A(n12595), .ZN(P3_U3471) );
  MUX2_X1 U15083 ( .A(P3_REG0_REG_12__SCAN_IN), .B(n12596), .S(n16017), .Z(
        n12597) );
  AOI21_X1 U15084 ( .B1(n13981), .B2(n13344), .A(n12597), .ZN(n12598) );
  OAI21_X1 U15085 ( .B1(n13988), .B2(n12599), .A(n12598), .ZN(P3_U3426) );
  OR2_X1 U15086 ( .A1(n12605), .A2(n15010), .ZN(n12600) );
  NAND2_X1 U15087 ( .A1(n12601), .A2(n12600), .ZN(n12602) );
  INV_X1 U15088 ( .A(n12610), .ZN(n12608) );
  OAI21_X1 U15089 ( .B1(n12602), .B2(n12608), .A(n12690), .ZN(n12603) );
  INV_X1 U15090 ( .A(n12603), .ZN(n15556) );
  NAND2_X1 U15091 ( .A1(n12607), .A2(n12606), .ZN(n12611) );
  INV_X1 U15092 ( .A(n12611), .ZN(n12609) );
  AOI21_X1 U15093 ( .B1(n12609), .B2(n12608), .A(n15829), .ZN(n12613) );
  AOI21_X1 U15094 ( .B1(n12613), .B2(n12712), .A(n12612), .ZN(n15555) );
  OAI21_X1 U15095 ( .B1(n12614), .B2(n15393), .A(n15555), .ZN(n12615) );
  NAND2_X1 U15096 ( .A1(n12615), .A2(n6544), .ZN(n12620) );
  INV_X1 U15097 ( .A(n15415), .ZN(n12616) );
  AOI211_X1 U15098 ( .C1(n15553), .C2(n12617), .A(n15742), .B(n12616), .ZN(
        n15552) );
  OAI22_X1 U15099 ( .A1(n7829), .A2(n15418), .B1(n11772), .B2(n6544), .ZN(
        n12618) );
  AOI21_X1 U15100 ( .B1(n15552), .B2(n15732), .A(n12618), .ZN(n12619) );
  OAI211_X1 U15101 ( .C1(n15556), .C2(n15423), .A(n12620), .B(n12619), .ZN(
        P1_U3280) );
  OAI22_X1 U15102 ( .A1(n15419), .A2(n13195), .B1(n12622), .B2(n13224), .ZN(
        n12621) );
  XNOR2_X1 U15103 ( .A(n12621), .B(n13233), .ZN(n12624) );
  NOR2_X1 U15104 ( .A1(n13223), .A2(n12622), .ZN(n12623) );
  AOI21_X1 U15105 ( .B1(n15548), .B2(n13189), .A(n12623), .ZN(n12625) );
  NAND2_X1 U15106 ( .A1(n12624), .A2(n12625), .ZN(n13164) );
  INV_X1 U15107 ( .A(n12624), .ZN(n12627) );
  INV_X1 U15108 ( .A(n12625), .ZN(n12626) );
  NAND2_X1 U15109 ( .A1(n12627), .A2(n12626), .ZN(n12628) );
  NAND2_X1 U15110 ( .A1(n13164), .A2(n12628), .ZN(n12637) );
  NAND2_X1 U15111 ( .A1(n12630), .A2(n12629), .ZN(n12635) );
  INV_X1 U15112 ( .A(n12631), .ZN(n12632) );
  NAND2_X1 U15113 ( .A1(n12633), .A2(n12632), .ZN(n12634) );
  AOI21_X1 U15114 ( .B1(n12637), .B2(n12636), .A(n13165), .ZN(n12642) );
  INV_X1 U15115 ( .A(n15412), .ZN(n15007) );
  NAND2_X1 U15116 ( .A1(n14983), .A2(n15007), .ZN(n12638) );
  NAND2_X1 U15117 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n15070)
         );
  OAI211_X1 U15118 ( .C1(n15410), .C2(n14971), .A(n12638), .B(n15070), .ZN(
        n12640) );
  NOR2_X1 U15119 ( .A1(n15419), .A2(n14963), .ZN(n12639) );
  AOI211_X1 U15120 ( .C1(n14928), .C2(n15416), .A(n12640), .B(n12639), .ZN(
        n12641) );
  OAI21_X1 U15121 ( .B1(n12642), .B2(n14994), .A(n12641), .ZN(P1_U3215) );
  NAND2_X1 U15122 ( .A1(n14983), .A2(n15012), .ZN(n12648) );
  NAND2_X1 U15123 ( .A1(n14978), .A2(n15014), .ZN(n12647) );
  INV_X1 U15124 ( .A(n12643), .ZN(n12644) );
  NAND2_X1 U15125 ( .A1(n14928), .A2(n12644), .ZN(n12646) );
  NAND4_X1 U15126 ( .A1(n12648), .A2(n12647), .A3(n12646), .A4(n12645), .ZN(
        n12654) );
  AOI21_X1 U15127 ( .B1(n12651), .B2(n12650), .A(n12649), .ZN(n12652) );
  NOR2_X1 U15128 ( .A1(n12652), .A2(n14994), .ZN(n12653) );
  AOI211_X1 U15129 ( .C1(n14992), .C2(n12655), .A(n12654), .B(n12653), .ZN(
        n12656) );
  INV_X1 U15130 ( .A(n12656), .ZN(P1_U3231) );
  AOI21_X1 U15131 ( .B1(n12658), .B2(n12657), .A(n14154), .ZN(n12660) );
  NAND2_X1 U15132 ( .A1(n12660), .A2(n12659), .ZN(n12666) );
  OAI21_X1 U15133 ( .B1(n14147), .B2(n12662), .A(n12661), .ZN(n12663) );
  AOI21_X1 U15134 ( .B1(n12664), .B2(n14168), .A(n12663), .ZN(n12665) );
  OAI211_X1 U15135 ( .C1(n9865), .C2(n14173), .A(n12666), .B(n12665), .ZN(
        P2_U3189) );
  NAND2_X1 U15136 ( .A1(n15892), .A2(n12668), .ZN(n12667) );
  OAI211_X1 U15137 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n15873), .A(n12667), .B(
        n14306), .ZN(n12671) );
  OAI22_X1 U15138 ( .A1(n12669), .A2(n15873), .B1(n14330), .B2(n12668), .ZN(
        n12670) );
  MUX2_X1 U15139 ( .A(n12671), .B(n12670), .S(n14222), .Z(n12675) );
  NAND2_X1 U15140 ( .A1(n15851), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n12672) );
  OAI21_X1 U15141 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n12673), .A(n12672), .ZN(
        n12674) );
  OR2_X1 U15142 ( .A1(n12675), .A2(n12674), .ZN(P2_U3214) );
  MUX2_X1 U15143 ( .A(n12676), .B(P3_REG2_REG_0__SCAN_IN), .S(n15997), .Z(
        n12681) );
  INV_X1 U15144 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n12679) );
  NAND2_X1 U15145 ( .A1(n15958), .A2(n12677), .ZN(n12678) );
  OAI21_X1 U15146 ( .B1(n12679), .B2(n15985), .A(n12678), .ZN(n12680) );
  OR2_X1 U15147 ( .A1(n12681), .A2(n12680), .ZN(P3_U3233) );
  AOI211_X1 U15148 ( .C1(n15937), .C2(n12684), .A(n12683), .B(n12682), .ZN(
        n12686) );
  MUX2_X1 U15149 ( .A(n9476), .B(n12686), .S(n14818), .Z(n12685) );
  OAI21_X1 U15150 ( .B1(n12688), .B2(n14822), .A(n12685), .ZN(P2_U3433) );
  MUX2_X1 U15151 ( .A(n9477), .B(n12686), .S(n15944), .Z(n12687) );
  OAI21_X1 U15152 ( .B1(n12688), .B2(n14781), .A(n12687), .ZN(P2_U3500) );
  OR2_X1 U15153 ( .A1(n15553), .A2(n15009), .ZN(n12689) );
  NAND2_X1 U15154 ( .A1(n15548), .A2(n15008), .ZN(n12691) );
  INV_X1 U15155 ( .A(n12691), .ZN(n15395) );
  NOR2_X1 U15156 ( .A1(n15405), .A2(n15395), .ZN(n12693) );
  NOR2_X1 U15157 ( .A1(n15543), .A2(n15007), .ZN(n12692) );
  AOI21_X1 U15158 ( .B1(n12694), .B2(n12693), .A(n12692), .ZN(n12695) );
  OR2_X1 U15159 ( .A1(n15537), .A2(n15006), .ZN(n12696) );
  NAND2_X1 U15160 ( .A1(n14965), .A2(n15359), .ZN(n12698) );
  INV_X1 U15161 ( .A(n15341), .ZN(n15004) );
  OR2_X1 U15162 ( .A1(n15519), .A2(n15004), .ZN(n12700) );
  NAND2_X1 U15163 ( .A1(n15305), .A2(n15003), .ZN(n12701) );
  OR2_X1 U15164 ( .A1(n15507), .A2(n15002), .ZN(n12702) );
  INV_X1 U15165 ( .A(n12729), .ZN(n15280) );
  NAND2_X1 U15166 ( .A1(n15281), .A2(n15280), .ZN(n15279) );
  NAND2_X1 U15167 ( .A1(n15277), .A2(n13194), .ZN(n12703) );
  NAND2_X2 U15168 ( .A1(n15279), .A2(n12703), .ZN(n15258) );
  NAND2_X1 U15169 ( .A1(n15265), .A2(n15000), .ZN(n12704) );
  OR2_X1 U15170 ( .A1(n15265), .A2(n15000), .ZN(n12705) );
  INV_X1 U15171 ( .A(n15244), .ZN(n12706) );
  NAND2_X1 U15172 ( .A1(n15222), .A2(n14998), .ZN(n12708) );
  NAND3_X1 U15173 ( .A1(n12715), .A2(n12714), .A3(n15370), .ZN(n15355) );
  NOR2_X1 U15174 ( .A1(n15531), .A2(n15340), .ZN(n12719) );
  AND2_X1 U15175 ( .A1(n12717), .A2(n12716), .ZN(n15353) );
  INV_X1 U15176 ( .A(n15006), .ZN(n15361) );
  NAND2_X1 U15177 ( .A1(n15537), .A2(n15361), .ZN(n15354) );
  NAND2_X1 U15178 ( .A1(n15531), .A2(n15340), .ZN(n12718) );
  OAI211_X1 U15179 ( .C1(n15355), .C2(n15353), .A(n15354), .B(n12718), .ZN(
        n15337) );
  INV_X1 U15180 ( .A(n12719), .ZN(n15336) );
  INV_X1 U15181 ( .A(n12722), .ZN(n12723) );
  INV_X1 U15182 ( .A(n15507), .ZN(n15288) );
  INV_X1 U15183 ( .A(n12730), .ZN(n15245) );
  INV_X1 U15184 ( .A(n15488), .ZN(n15255) );
  INV_X1 U15185 ( .A(n14999), .ZN(n12731) );
  INV_X1 U15186 ( .A(n15212), .ZN(n12733) );
  NAND2_X1 U15187 ( .A1(n15482), .A2(n12733), .ZN(n15210) );
  INV_X1 U15188 ( .A(n14998), .ZN(n14852) );
  NAND2_X1 U15189 ( .A1(n15222), .A2(n14852), .ZN(n12738) );
  AOI22_X1 U15190 ( .A1(n15181), .A2(n15746), .B1(n15426), .B2(n14998), .ZN(
        n12740) );
  NAND2_X1 U15191 ( .A1(n15468), .A2(n6544), .ZN(n12747) );
  NOR2_X2 U15192 ( .A1(n15415), .A2(n15548), .ZN(n15414) );
  INV_X1 U15193 ( .A(n15543), .ZN(n12742) );
  OAI211_X1 U15194 ( .C1(n15161), .C2(n15216), .A(n10870), .B(n15195), .ZN(
        n15470) );
  INV_X1 U15195 ( .A(n15470), .ZN(n12745) );
  AOI22_X1 U15196 ( .A1(n14854), .A2(n15760), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n15764), .ZN(n12743) );
  OAI21_X1 U15197 ( .B1(n15161), .B2(n15418), .A(n12743), .ZN(n12744) );
  AOI21_X1 U15198 ( .B1(n12745), .B2(n15732), .A(n12744), .ZN(n12746) );
  OAI211_X1 U15199 ( .C1(n15472), .C2(n15438), .A(n12747), .B(n12746), .ZN(
        P1_U3266) );
  OAI222_X1 U15200 ( .A1(n15597), .A2(n12749), .B1(n15595), .B2(n12748), .C1(
        P1_U3086), .C2(n10808), .ZN(P1_U3334) );
  NAND2_X1 U15201 ( .A1(n14485), .A2(n14658), .ZN(n14132) );
  INV_X1 U15202 ( .A(n14132), .ZN(n12794) );
  XNOR2_X1 U15203 ( .A(n12750), .B(n12751), .ZN(n14130) );
  INV_X1 U15204 ( .A(n14130), .ZN(n12793) );
  XNOR2_X1 U15205 ( .A(n14620), .B(n10413), .ZN(n12835) );
  NOR2_X1 U15206 ( .A1(n10450), .A2(n14637), .ZN(n12756) );
  INV_X1 U15207 ( .A(n12756), .ZN(n12834) );
  OAI21_X1 U15208 ( .B1(n12835), .B2(n12834), .A(n12832), .ZN(n12759) );
  XNOR2_X1 U15209 ( .A(n14605), .B(n10413), .ZN(n12839) );
  OR2_X1 U15210 ( .A1(n10450), .A2(n14089), .ZN(n12761) );
  NAND2_X1 U15211 ( .A1(n12755), .A2(n12756), .ZN(n12752) );
  NAND2_X1 U15212 ( .A1(n12835), .A2(n12752), .ZN(n12754) );
  XNOR2_X1 U15213 ( .A(n14580), .B(n12750), .ZN(n12841) );
  OR2_X1 U15214 ( .A1(n14594), .A2(n10450), .ZN(n12840) );
  NAND2_X1 U15215 ( .A1(n12841), .A2(n12840), .ZN(n12753) );
  OAI211_X1 U15216 ( .C1(n12756), .C2(n12755), .A(n12754), .B(n12753), .ZN(
        n12757) );
  AOI21_X1 U15217 ( .B1(n12839), .B2(n12761), .A(n12757), .ZN(n12758) );
  INV_X1 U15218 ( .A(n12839), .ZN(n12762) );
  INV_X1 U15219 ( .A(n12761), .ZN(n12837) );
  NAND2_X1 U15220 ( .A1(n12762), .A2(n12837), .ZN(n12763) );
  XNOR2_X1 U15221 ( .A(n14566), .B(n10413), .ZN(n12768) );
  OR2_X1 U15222 ( .A1(n14538), .A2(n10450), .ZN(n12769) );
  XNOR2_X1 U15223 ( .A(n12768), .B(n12769), .ZN(n12843) );
  OAI21_X1 U15224 ( .B1(n12763), .B2(n12840), .A(n12843), .ZN(n12765) );
  AOI21_X1 U15225 ( .B1(n12763), .B2(n12840), .A(n12841), .ZN(n12764) );
  NOR2_X1 U15226 ( .A1(n12765), .A2(n12764), .ZN(n12766) );
  INV_X1 U15227 ( .A(n12768), .ZN(n12770) );
  NAND2_X1 U15228 ( .A1(n12770), .A2(n12769), .ZN(n12771) );
  XNOR2_X1 U15229 ( .A(n14552), .B(n10413), .ZN(n12773) );
  NAND2_X1 U15230 ( .A1(n14202), .A2(n14658), .ZN(n12774) );
  XNOR2_X1 U15231 ( .A(n12773), .B(n12774), .ZN(n14155) );
  INV_X1 U15232 ( .A(n14155), .ZN(n12772) );
  INV_X1 U15233 ( .A(n12773), .ZN(n12776) );
  INV_X1 U15234 ( .A(n12774), .ZN(n12775) );
  NAND2_X1 U15235 ( .A1(n12776), .A2(n12775), .ZN(n12777) );
  XNOR2_X1 U15236 ( .A(n14732), .B(n12750), .ZN(n12778) );
  NAND2_X1 U15237 ( .A1(n14201), .A2(n14658), .ZN(n12779) );
  NAND2_X1 U15238 ( .A1(n12778), .A2(n12779), .ZN(n14031) );
  INV_X1 U15239 ( .A(n12778), .ZN(n12781) );
  INV_X1 U15240 ( .A(n12779), .ZN(n12780) );
  NAND2_X1 U15241 ( .A1(n12781), .A2(n12780), .ZN(n14030) );
  XNOR2_X1 U15242 ( .A(n14515), .B(n12750), .ZN(n12783) );
  NAND2_X1 U15243 ( .A1(n14484), .A2(n14658), .ZN(n12784) );
  NAND2_X1 U15244 ( .A1(n12783), .A2(n12784), .ZN(n14118) );
  INV_X1 U15245 ( .A(n12783), .ZN(n12786) );
  INV_X1 U15246 ( .A(n12784), .ZN(n12785) );
  NAND2_X1 U15247 ( .A1(n12786), .A2(n12785), .ZN(n14119) );
  XNOR2_X1 U15248 ( .A(n14491), .B(n10413), .ZN(n12789) );
  NAND2_X1 U15249 ( .A1(n14200), .A2(n14658), .ZN(n12787) );
  XNOR2_X1 U15250 ( .A(n12789), .B(n12787), .ZN(n14055) );
  INV_X1 U15251 ( .A(n12787), .ZN(n12788) );
  NAND2_X1 U15252 ( .A1(n12789), .A2(n12788), .ZN(n14128) );
  INV_X1 U15253 ( .A(n14128), .ZN(n12791) );
  NOR2_X1 U15254 ( .A1(n12795), .A2(n10450), .ZN(n14022) );
  XNOR2_X1 U15255 ( .A(n14710), .B(n10413), .ZN(n14071) );
  XNOR2_X1 U15256 ( .A(n14705), .B(n10413), .ZN(n12797) );
  AND2_X1 U15257 ( .A1(n14198), .A2(n14658), .ZN(n12798) );
  NOR2_X1 U15258 ( .A1(n12797), .A2(n12798), .ZN(n14075) );
  INV_X1 U15259 ( .A(n14075), .ZN(n12796) );
  OAI21_X1 U15260 ( .B1(n14022), .B2(n14071), .A(n12796), .ZN(n12802) );
  NAND3_X1 U15261 ( .A1(n12796), .A2(n14022), .A3(n14071), .ZN(n12801) );
  INV_X1 U15262 ( .A(n12797), .ZN(n14078) );
  INV_X1 U15263 ( .A(n12798), .ZN(n12799) );
  NOR2_X1 U15264 ( .A1(n14078), .A2(n12799), .ZN(n14074) );
  INV_X1 U15265 ( .A(n14074), .ZN(n12800) );
  XNOR2_X1 U15266 ( .A(n14700), .B(n10413), .ZN(n12803) );
  AND2_X1 U15267 ( .A1(n14197), .A2(n14658), .ZN(n12804) );
  NAND2_X1 U15268 ( .A1(n12803), .A2(n12804), .ZN(n12807) );
  INV_X1 U15269 ( .A(n12803), .ZN(n14165) );
  INV_X1 U15270 ( .A(n12804), .ZN(n12805) );
  NAND2_X1 U15271 ( .A1(n14165), .A2(n12805), .ZN(n12806) );
  NAND2_X1 U15272 ( .A1(n12807), .A2(n12806), .ZN(n14076) );
  XNOR2_X1 U15273 ( .A(n14695), .B(n10413), .ZN(n12809) );
  NAND2_X1 U15274 ( .A1(n14196), .A2(n14658), .ZN(n12810) );
  XNOR2_X1 U15275 ( .A(n12809), .B(n12810), .ZN(n14177) );
  INV_X1 U15276 ( .A(n12809), .ZN(n12811) );
  XNOR2_X1 U15277 ( .A(n14690), .B(n10413), .ZN(n12813) );
  INV_X1 U15278 ( .A(n12813), .ZN(n12815) );
  AND2_X1 U15279 ( .A1(n14195), .A2(n14658), .ZN(n12812) );
  INV_X1 U15280 ( .A(n12812), .ZN(n12814) );
  NAND2_X1 U15281 ( .A1(n12817), .A2(n12816), .ZN(n14052) );
  INV_X1 U15282 ( .A(n14355), .ZN(n12819) );
  OAI22_X1 U15283 ( .A1(n12819), .A2(n14638), .B1(n12818), .B2(n14636), .ZN(
        n14378) );
  INV_X1 U15284 ( .A(n14378), .ZN(n12821) );
  OAI22_X1 U15285 ( .A1(n12821), .A2(n14147), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12820), .ZN(n12822) );
  AOI21_X1 U15286 ( .B1(n14385), .B2(n14168), .A(n12822), .ZN(n12823) );
  OAI222_X1 U15287 ( .A1(n15597), .A2(n12825), .B1(n15595), .B2(n12824), .C1(
        n8722), .C2(P1_U3086), .ZN(P1_U3335) );
  NOR2_X1 U15288 ( .A1(n15596), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12826) );
  NAND2_X1 U15289 ( .A1(n15596), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12828) );
  INV_X1 U15290 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n12871) );
  XNOR2_X1 U15291 ( .A(n12871), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n12830) );
  XNOR2_X1 U15292 ( .A(n12870), .B(n12830), .ZN(n12864) );
  INV_X1 U15293 ( .A(n12864), .ZN(n12831) );
  OAI222_X1 U15294 ( .A1(n13257), .A2(n12831), .B1(P3_U3151), .B2(n12879), 
        .C1(n12865), .C2(n14006), .ZN(P3_U3267) );
  INV_X1 U15295 ( .A(n12832), .ZN(n12833) );
  XNOR2_X1 U15296 ( .A(n12835), .B(n12834), .ZN(n14013) );
  NOR3_X1 U15297 ( .A1(n14012), .A2(n12833), .A3(n14013), .ZN(n14018) );
  AOI21_X1 U15298 ( .B1(n12835), .B2(n12834), .A(n14018), .ZN(n12836) );
  INV_X1 U15299 ( .A(n12836), .ZN(n12838) );
  XNOR2_X1 U15300 ( .A(n12836), .B(n12839), .ZN(n14181) );
  NAND2_X1 U15301 ( .A1(n14181), .A2(n12837), .ZN(n14182) );
  OAI21_X1 U15302 ( .B1(n12839), .B2(n12838), .A(n14182), .ZN(n14086) );
  XNOR2_X1 U15303 ( .A(n12841), .B(n12840), .ZN(n14087) );
  NOR2_X1 U15304 ( .A1(n14086), .A2(n14087), .ZN(n14085) );
  INV_X1 U15305 ( .A(n12841), .ZN(n12842) );
  AOI22_X1 U15306 ( .A1(n12842), .A2(n14180), .B1(n14179), .B2(n14203), .ZN(
        n12844) );
  OR3_X1 U15307 ( .A1(n14085), .A2(n12844), .A3(n12843), .ZN(n12848) );
  NAND2_X1 U15308 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n14288)
         );
  OAI21_X1 U15309 ( .B1(n14184), .B2(n14563), .A(n14288), .ZN(n12846) );
  OAI22_X1 U15310 ( .A1(n14567), .A2(n14186), .B1(n14185), .B2(n14594), .ZN(
        n12845) );
  AOI211_X1 U15311 ( .C1(n14566), .C2(n14189), .A(n12846), .B(n12845), .ZN(
        n12847) );
  OAI211_X1 U15312 ( .C1(n14154), .C2(n12849), .A(n12848), .B(n12847), .ZN(
        P2_U3200) );
  NAND2_X1 U15313 ( .A1(n13817), .A2(n13831), .ZN(n13075) );
  INV_X1 U15314 ( .A(n13817), .ZN(n13897) );
  OR2_X1 U15315 ( .A1(n13980), .A2(n13812), .ZN(n13078) );
  NAND2_X1 U15316 ( .A1(n13980), .A2(n13812), .ZN(n13079) );
  INV_X1 U15317 ( .A(n13980), .ZN(n13361) );
  INV_X1 U15318 ( .A(n13751), .ZN(n13084) );
  INV_X1 U15319 ( .A(n13974), .ZN(n13371) );
  INV_X1 U15320 ( .A(n12890), .ZN(n12852) );
  NAND2_X1 U15321 ( .A1(n13084), .A2(n12852), .ZN(n13750) );
  OR2_X1 U15322 ( .A1(n13782), .A2(n13759), .ZN(n13752) );
  NAND2_X1 U15323 ( .A1(n13964), .A2(n13743), .ZN(n13741) );
  NAND2_X1 U15324 ( .A1(n13964), .A2(n13772), .ZN(n13091) );
  NOR2_X1 U15325 ( .A1(n13782), .A2(n13789), .ZN(n13756) );
  NOR2_X1 U15326 ( .A1(n13755), .A2(n13756), .ZN(n13740) );
  INV_X1 U15327 ( .A(n13740), .ZN(n12854) );
  NAND2_X1 U15328 ( .A1(n12854), .A2(n13741), .ZN(n12855) );
  AND2_X1 U15329 ( .A1(n7852), .A2(n12855), .ZN(n12856) );
  INV_X1 U15330 ( .A(n13958), .ZN(n12857) );
  INV_X1 U15331 ( .A(n13874), .ZN(n13327) );
  INV_X1 U15332 ( .A(n13948), .ZN(n12859) );
  INV_X1 U15333 ( .A(n13702), .ZN(n12989) );
  INV_X1 U15334 ( .A(n13683), .ZN(n13678) );
  NAND2_X1 U15335 ( .A1(n13664), .A2(n7984), .ZN(n12863) );
  NAND2_X1 U15336 ( .A1(n13667), .A2(n13422), .ZN(n12862) );
  NAND2_X1 U15337 ( .A1(n12864), .A2(n12935), .ZN(n12867) );
  OR2_X1 U15338 ( .A1(n7252), .A2(n12865), .ZN(n12866) );
  NOR2_X1 U15339 ( .A1(n13927), .A2(n13666), .ZN(n13636) );
  AND2_X1 U15340 ( .A1(n13259), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12869) );
  NAND2_X1 U15341 ( .A1(n12871), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12872) );
  NAND2_X1 U15342 ( .A1(n15593), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12928) );
  NAND2_X1 U15343 ( .A1(n14827), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12873) );
  NAND2_X1 U15344 ( .A1(n12928), .A2(n12873), .ZN(n12874) );
  NAND2_X1 U15345 ( .A1(n12875), .A2(n12874), .ZN(n12876) );
  NAND2_X1 U15346 ( .A1(n12929), .A2(n12876), .ZN(n14009) );
  OR2_X1 U15347 ( .A1(n7252), .A2(n14007), .ZN(n12877) );
  NAND2_X1 U15348 ( .A1(n13844), .A2(n13640), .ZN(n12954) );
  NOR2_X1 U15349 ( .A1(n12879), .A2(n8086), .ZN(n12880) );
  OR2_X1 U15350 ( .A1(n15992), .A2(n12880), .ZN(n13623) );
  OAI22_X1 U15351 ( .A1(n13655), .A2(n15990), .B1(n12958), .B2(n13623), .ZN(
        n12881) );
  AOI21_X1 U15352 ( .B1(n12882), .B2(n13833), .A(n12881), .ZN(n13842) );
  MUX2_X1 U15353 ( .A(n12883), .B(n13842), .S(n16017), .Z(n12900) );
  NOR2_X1 U15354 ( .A1(n13389), .A2(n13829), .ZN(n12884) );
  NAND2_X1 U15355 ( .A1(n13389), .A2(n13829), .ZN(n12886) );
  AND2_X1 U15356 ( .A1(n13996), .A2(n13452), .ZN(n12888) );
  NAND2_X1 U15357 ( .A1(n13798), .A2(n13797), .ZN(n13796) );
  NAND2_X1 U15358 ( .A1(n13083), .A2(n12890), .ZN(n12891) );
  AND2_X1 U15359 ( .A1(n12891), .A2(n13752), .ZN(n12892) );
  OR2_X1 U15360 ( .A1(n13958), .A2(n13760), .ZN(n13096) );
  NAND2_X1 U15361 ( .A1(n13874), .A2(n13398), .ZN(n12896) );
  AND2_X1 U15362 ( .A1(n13948), .A2(n13731), .ZN(n12971) );
  XNOR2_X1 U15363 ( .A(n12898), .B(n13704), .ZN(n13118) );
  NAND2_X1 U15364 ( .A1(n12898), .A2(n13704), .ZN(n13113) );
  INV_X1 U15365 ( .A(n13665), .ZN(n13692) );
  NAND2_X1 U15366 ( .A1(n13119), .A2(n13692), .ZN(n13121) );
  NAND2_X1 U15367 ( .A1(n12899), .A2(n13120), .ZN(n13648) );
  INV_X1 U15368 ( .A(n13666), .ZN(n13639) );
  NAND2_X1 U15369 ( .A1(n13927), .A2(n13639), .ZN(n13127) );
  NAND2_X1 U15370 ( .A1(n13921), .A2(n13655), .ZN(n13133) );
  INV_X1 U15371 ( .A(n14822), .ZN(n12906) );
  NAND2_X1 U15372 ( .A1(n14681), .A2(n14358), .ZN(n12901) );
  INV_X1 U15373 ( .A(n14352), .ZN(n12903) );
  NAND2_X1 U15374 ( .A1(n14193), .A2(n12903), .ZN(n12904) );
  NOR2_X1 U15375 ( .A1(n14638), .A2(n12904), .ZN(n14675) );
  INV_X1 U15376 ( .A(n14675), .ZN(n14337) );
  MUX2_X1 U15377 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n14679), .S(n14818), .Z(
        n12905) );
  INV_X1 U15378 ( .A(n12907), .ZN(P2_U3497) );
  INV_X1 U15379 ( .A(n12908), .ZN(n15594) );
  XNOR2_X1 U15380 ( .A(n13448), .B(n12911), .ZN(n12912) );
  XNOR2_X1 U15381 ( .A(n13921), .B(n12912), .ZN(n12919) );
  INV_X1 U15382 ( .A(n12919), .ZN(n12913) );
  NAND2_X1 U15383 ( .A1(n12913), .A2(n13437), .ZN(n12925) );
  INV_X1 U15384 ( .A(n12914), .ZN(n12915) );
  NAND4_X1 U15385 ( .A1(n12924), .A2(n13437), .A3(n12919), .A4(n12915), .ZN(
        n12923) );
  AOI22_X1 U15386 ( .A1(n13645), .A2(n13443), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12917) );
  NAND2_X1 U15387 ( .A1(n13666), .A2(n13439), .ZN(n12916) );
  OAI211_X1 U15388 ( .C1(n13640), .C2(n13441), .A(n12917), .B(n12916), .ZN(
        n12921) );
  NOR4_X1 U15389 ( .A1(n12919), .A2(n12918), .A3(n13666), .A4(n13413), .ZN(
        n12920) );
  AOI211_X1 U15390 ( .C1(n13921), .C2(n13400), .A(n12921), .B(n12920), .ZN(
        n12922) );
  OAI211_X1 U15391 ( .C1(n12925), .C2(n12924), .A(n12923), .B(n12922), .ZN(
        P3_U3160) );
  NAND2_X1 U15392 ( .A1(n13277), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12931) );
  NAND2_X1 U15393 ( .A1(n13280), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12930) );
  AND2_X1 U15394 ( .A1(n12931), .A2(n12930), .ZN(n12946) );
  NAND2_X1 U15395 ( .A1(n12949), .A2(n12931), .ZN(n12934) );
  INV_X1 U15396 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n12932) );
  XNOR2_X1 U15397 ( .A(n12932), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n12933) );
  XNOR2_X1 U15398 ( .A(n12934), .B(n12933), .ZN(n14000) );
  NAND2_X1 U15399 ( .A1(n14000), .A2(n12935), .ZN(n12937) );
  INV_X1 U15400 ( .A(SI_31_), .ZN(n14005) );
  OR2_X1 U15401 ( .A1(n7252), .A2(n14005), .ZN(n12936) );
  NAND2_X1 U15402 ( .A1(n12938), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12941) );
  NAND2_X1 U15403 ( .A1(n12939), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12940) );
  OAI211_X1 U15404 ( .C1(n12942), .C2(n6545), .A(n12941), .B(n12940), .ZN(
        n12943) );
  INV_X1 U15405 ( .A(n12943), .ZN(n12944) );
  NAND2_X1 U15406 ( .A1(n12949), .A2(n12948), .ZN(n13256) );
  INV_X1 U15407 ( .A(SI_30_), .ZN(n13254) );
  OR2_X1 U15408 ( .A1(n7252), .A2(n13254), .ZN(n12952) );
  INV_X1 U15409 ( .A(n12954), .ZN(n12955) );
  AOI21_X1 U15410 ( .B1(n13915), .B2(n12958), .A(n12955), .ZN(n12956) );
  INV_X1 U15411 ( .A(n12993), .ZN(n13137) );
  NAND2_X1 U15412 ( .A1(n13915), .A2(n13624), .ZN(n12962) );
  INV_X1 U15413 ( .A(n12962), .ZN(n12957) );
  NOR2_X1 U15414 ( .A1(n13137), .A2(n12957), .ZN(n12961) );
  INV_X1 U15415 ( .A(n13624), .ZN(n13447) );
  NAND2_X1 U15416 ( .A1(n12969), .A2(n12959), .ZN(n12965) );
  NAND2_X1 U15417 ( .A1(n12965), .A2(n13616), .ZN(n12960) );
  AOI21_X1 U15418 ( .B1(n12964), .B2(n12961), .A(n12960), .ZN(n12999) );
  NAND2_X1 U15419 ( .A1(n12968), .A2(n12967), .ZN(n12998) );
  INV_X1 U15420 ( .A(n12969), .ZN(n13135) );
  INV_X1 U15421 ( .A(n12970), .ZN(n13132) );
  INV_X1 U15422 ( .A(n13649), .ZN(n13652) );
  INV_X1 U15423 ( .A(n12971), .ZN(n13107) );
  NAND2_X1 U15424 ( .A1(n13106), .A2(n13107), .ZN(n13100) );
  INV_X1 U15425 ( .A(n13025), .ZN(n12977) );
  NAND4_X1 U15426 ( .A1(n15965), .A2(n10905), .A3(n13019), .A4(n12972), .ZN(
        n12975) );
  INV_X1 U15427 ( .A(n12973), .ZN(n12974) );
  NOR4_X1 U15428 ( .A1(n12977), .A2(n12976), .A3(n12975), .A4(n12974), .ZN(
        n12978) );
  NAND2_X1 U15429 ( .A1(n12978), .A2(n13037), .ZN(n12981) );
  INV_X1 U15430 ( .A(n13041), .ZN(n12980) );
  NOR4_X1 U15431 ( .A1(n12981), .A2(n12980), .A3(n12979), .A4(n13055), .ZN(
        n12982) );
  NAND4_X1 U15432 ( .A1(n12984), .A2(n7944), .A3(n12983), .A4(n12982), .ZN(
        n12986) );
  INV_X1 U15433 ( .A(n13797), .ZN(n13799) );
  NOR4_X1 U15434 ( .A1(n13750), .A2(n12986), .A3(n13799), .A4(n12985), .ZN(
        n12987) );
  NAND4_X1 U15435 ( .A1(n13755), .A2(n13777), .A3(n13826), .A4(n12987), .ZN(
        n12988) );
  NOR4_X1 U15436 ( .A1(n12989), .A2(n7852), .A3(n13100), .A4(n12988), .ZN(
        n12990) );
  INV_X1 U15437 ( .A(n13118), .ZN(n13695) );
  XNOR2_X1 U15438 ( .A(n13874), .B(n13744), .ZN(n13728) );
  NAND4_X1 U15439 ( .A1(n13683), .A2(n12990), .A3(n13695), .A4(n13728), .ZN(
        n12991) );
  NOR4_X1 U15440 ( .A1(n13132), .A2(n13652), .A3(n13663), .A4(n12991), .ZN(
        n12992) );
  NAND4_X1 U15441 ( .A1(n12993), .A2(n13135), .A3(n12992), .A4(n13635), .ZN(
        n12994) );
  XNOR2_X1 U15442 ( .A(n12994), .B(n13599), .ZN(n12996) );
  OR2_X2 U15443 ( .A1(n12996), .A2(n12995), .ZN(n12997) );
  OAI21_X1 U15444 ( .B1(n12999), .B2(n12998), .A(n12997), .ZN(n13141) );
  NAND2_X1 U15445 ( .A1(n13000), .A2(n6543), .ZN(n13003) );
  NAND2_X1 U15446 ( .A1(n13000), .A2(n8546), .ZN(n13001) );
  NAND3_X1 U15447 ( .A1(n13007), .A2(n13001), .A3(n13124), .ZN(n13002) );
  OAI21_X1 U15448 ( .B1(n13004), .B2(n13003), .A(n13002), .ZN(n13005) );
  MUX2_X1 U15449 ( .A(n13008), .B(n13007), .S(n13101), .Z(n13009) );
  NAND2_X1 U15450 ( .A1(n13010), .A2(n13124), .ZN(n13012) );
  INV_X1 U15451 ( .A(n13015), .ZN(n13011) );
  AOI21_X1 U15452 ( .B1(n13013), .B2(n13012), .A(n13011), .ZN(n13021) );
  AOI21_X1 U15453 ( .B1(n13015), .B2(n13014), .A(n13124), .ZN(n13020) );
  INV_X1 U15454 ( .A(n13016), .ZN(n13017) );
  NAND2_X1 U15455 ( .A1(n13017), .A2(n13101), .ZN(n13018) );
  MUX2_X1 U15456 ( .A(n13023), .B(n13022), .S(n13124), .Z(n13024) );
  NAND3_X1 U15457 ( .A1(n13026), .A2(n13025), .A3(n13024), .ZN(n13033) );
  NAND2_X1 U15458 ( .A1(n13035), .A2(n13027), .ZN(n13030) );
  NAND2_X1 U15459 ( .A1(n13034), .A2(n13028), .ZN(n13029) );
  MUX2_X1 U15460 ( .A(n13030), .B(n13029), .S(n13101), .Z(n13031) );
  INV_X1 U15461 ( .A(n13031), .ZN(n13032) );
  MUX2_X1 U15462 ( .A(n13035), .B(n13034), .S(n13124), .Z(n13036) );
  MUX2_X1 U15463 ( .A(n13039), .B(n13038), .S(n13124), .Z(n13040) );
  MUX2_X1 U15464 ( .A(n13043), .B(n13042), .S(n13124), .Z(n13044) );
  NAND3_X1 U15465 ( .A1(n13046), .A2(n13045), .A3(n13044), .ZN(n13050) );
  MUX2_X1 U15466 ( .A(n13048), .B(n13047), .S(n13124), .Z(n13049) );
  NAND2_X1 U15467 ( .A1(n13050), .A2(n13049), .ZN(n13051) );
  NAND2_X1 U15468 ( .A1(n13051), .A2(n7944), .ZN(n13059) );
  NOR2_X1 U15469 ( .A1(n13308), .A2(n13124), .ZN(n13053) );
  AND2_X1 U15470 ( .A1(n13308), .A2(n13124), .ZN(n13052) );
  MUX2_X1 U15471 ( .A(n13053), .B(n13052), .S(n13455), .Z(n13054) );
  NOR2_X1 U15472 ( .A1(n13055), .A2(n13054), .ZN(n13058) );
  AOI21_X1 U15473 ( .B1(n13067), .B2(n13056), .A(n13101), .ZN(n13057) );
  AOI21_X1 U15474 ( .B1(n13059), .B2(n13058), .A(n13057), .ZN(n13064) );
  INV_X1 U15475 ( .A(n13061), .ZN(n13063) );
  AND2_X1 U15476 ( .A1(n13061), .A2(n13060), .ZN(n13062) );
  OAI22_X1 U15477 ( .A1(n13064), .A2(n13063), .B1(n13062), .B2(n13124), .ZN(
        n13066) );
  MUX2_X1 U15478 ( .A(n13284), .B(n13101), .S(n13389), .Z(n13068) );
  OAI21_X1 U15479 ( .B1(n13829), .B2(n13124), .A(n13068), .ZN(n13069) );
  NAND2_X1 U15480 ( .A1(n13996), .A2(n13124), .ZN(n13071) );
  OR2_X1 U15481 ( .A1(n13996), .A2(n13124), .ZN(n13070) );
  MUX2_X1 U15482 ( .A(n13071), .B(n13070), .S(n13811), .Z(n13072) );
  AOI21_X1 U15483 ( .B1(n13073), .B2(n13072), .A(n13814), .ZN(n13082) );
  NAND2_X1 U15484 ( .A1(n13079), .A2(n13074), .ZN(n13077) );
  NAND2_X1 U15485 ( .A1(n13078), .A2(n13075), .ZN(n13076) );
  MUX2_X1 U15486 ( .A(n13077), .B(n13076), .S(n13124), .Z(n13081) );
  MUX2_X1 U15487 ( .A(n13079), .B(n13078), .S(n13101), .Z(n13080) );
  OAI21_X1 U15488 ( .B1(n13082), .B2(n13081), .A(n13080), .ZN(n13090) );
  NOR2_X1 U15489 ( .A1(n13739), .A2(n13750), .ZN(n13089) );
  OAI211_X1 U15490 ( .C1(n13739), .C2(n13084), .A(n13083), .B(n13091), .ZN(
        n13087) );
  INV_X1 U15491 ( .A(n13085), .ZN(n13086) );
  MUX2_X1 U15492 ( .A(n13087), .B(n13086), .S(n13101), .Z(n13088) );
  AOI21_X1 U15493 ( .B1(n13090), .B2(n13089), .A(n13088), .ZN(n13095) );
  INV_X1 U15494 ( .A(n13092), .ZN(n13093) );
  MUX2_X1 U15495 ( .A(n12893), .B(n13093), .S(n13124), .Z(n13094) );
  OAI21_X1 U15496 ( .B1(n13095), .B2(n13094), .A(n12895), .ZN(n13099) );
  NAND2_X1 U15497 ( .A1(n13958), .A2(n13760), .ZN(n13097) );
  MUX2_X1 U15498 ( .A(n13097), .B(n13096), .S(n13124), .Z(n13098) );
  INV_X1 U15499 ( .A(n13100), .ZN(n13718) );
  NAND2_X1 U15500 ( .A1(n13744), .A2(n13101), .ZN(n13103) );
  OR2_X1 U15501 ( .A1(n13744), .A2(n13101), .ZN(n13102) );
  MUX2_X1 U15502 ( .A(n13103), .B(n13102), .S(n13874), .Z(n13104) );
  NAND3_X1 U15503 ( .A1(n13105), .A2(n13718), .A3(n13104), .ZN(n13109) );
  MUX2_X1 U15504 ( .A(n13107), .B(n13106), .S(n13124), .Z(n13108) );
  NAND2_X1 U15505 ( .A1(n13109), .A2(n13108), .ZN(n13111) );
  NOR2_X1 U15506 ( .A1(n13720), .A2(n13124), .ZN(n13110) );
  AOI22_X1 U15507 ( .A1(n13111), .A2(n13702), .B1(n13110), .B2(n13710), .ZN(
        n13117) );
  NAND2_X1 U15508 ( .A1(n13695), .A2(n13112), .ZN(n13115) );
  XNOR2_X1 U15509 ( .A(n13113), .B(n13124), .ZN(n13114) );
  NAND2_X1 U15510 ( .A1(n13115), .A2(n13114), .ZN(n13116) );
  INV_X1 U15511 ( .A(n13119), .ZN(n13937) );
  NAND3_X1 U15512 ( .A1(n13120), .A2(n13937), .A3(n13665), .ZN(n13122) );
  MUX2_X1 U15513 ( .A(n13122), .B(n13121), .S(n8579), .Z(n13126) );
  INV_X1 U15514 ( .A(n13123), .ZN(n13125) );
  NOR2_X1 U15515 ( .A1(n13128), .A2(n6930), .ZN(n13131) );
  INV_X1 U15516 ( .A(n13128), .ZN(n13129) );
  INV_X1 U15517 ( .A(n13134), .ZN(n13136) );
  NAND2_X1 U15518 ( .A1(n13143), .A2(n13142), .ZN(n13144) );
  OAI211_X1 U15519 ( .C1(n6543), .C2(n13145), .A(n13144), .B(P3_B_REG_SCAN_IN), 
        .ZN(n13147) );
  NAND2_X1 U15520 ( .A1(n13148), .A2(n13147), .ZN(P3_U3296) );
  NAND2_X1 U15521 ( .A1(n15462), .A2(n10876), .ZN(n13150) );
  NAND2_X1 U15522 ( .A1(n15181), .A2(n13189), .ZN(n13149) );
  NAND2_X1 U15523 ( .A1(n13150), .A2(n13149), .ZN(n13151) );
  XNOR2_X1 U15524 ( .A(n13151), .B(n13233), .ZN(n13153) );
  AOI22_X1 U15525 ( .A1(n15462), .A2(n13189), .B1(n13235), .B2(n15181), .ZN(
        n13152) );
  XNOR2_X1 U15526 ( .A(n13153), .B(n13152), .ZN(n13247) );
  INV_X1 U15527 ( .A(n13247), .ZN(n13154) );
  NAND2_X1 U15528 ( .A1(n13154), .A2(n14969), .ZN(n13253) );
  AND2_X1 U15529 ( .A1(n15003), .A2(n13235), .ZN(n13155) );
  AOI21_X1 U15530 ( .B1(n15305), .B2(n13189), .A(n13155), .ZN(n13186) );
  INV_X1 U15531 ( .A(n13186), .ZN(n13188) );
  OAI22_X1 U15532 ( .A1(n15512), .A2(n13195), .B1(n15322), .B2(n13224), .ZN(
        n13156) );
  XNOR2_X1 U15533 ( .A(n13156), .B(n11908), .ZN(n13187) );
  OAI22_X1 U15534 ( .A1(n15345), .A2(n13224), .B1(n15321), .B2(n13223), .ZN(
        n13182) );
  NAND2_X1 U15535 ( .A1(n14965), .A2(n10876), .ZN(n13158) );
  NAND2_X1 U15536 ( .A1(n15359), .A2(n13189), .ZN(n13157) );
  NAND2_X1 U15537 ( .A1(n13158), .A2(n13157), .ZN(n13159) );
  XNOR2_X1 U15538 ( .A(n13159), .B(n11908), .ZN(n13181) );
  NAND2_X1 U15539 ( .A1(n15537), .A2(n10876), .ZN(n13161) );
  NAND2_X1 U15540 ( .A1(n15006), .A2(n13189), .ZN(n13160) );
  NAND2_X1 U15541 ( .A1(n13161), .A2(n13160), .ZN(n13162) );
  XNOR2_X1 U15542 ( .A(n13162), .B(n11908), .ZN(n13170) );
  INV_X1 U15543 ( .A(n13170), .ZN(n13174) );
  AND2_X1 U15544 ( .A1(n13235), .A2(n15006), .ZN(n13163) );
  AOI21_X1 U15545 ( .B1(n15537), .B2(n13189), .A(n13163), .ZN(n13173) );
  NAND2_X1 U15546 ( .A1(n15543), .A2(n10876), .ZN(n13167) );
  NAND2_X1 U15547 ( .A1(n15007), .A2(n13189), .ZN(n13166) );
  NAND2_X1 U15548 ( .A1(n13167), .A2(n13166), .ZN(n13168) );
  XNOR2_X1 U15549 ( .A(n13168), .B(n13233), .ZN(n14905) );
  NOR2_X1 U15550 ( .A1(n15412), .A2(n13223), .ZN(n13169) );
  AOI21_X1 U15551 ( .B1(n15543), .B2(n13189), .A(n13169), .ZN(n14906) );
  NAND2_X1 U15552 ( .A1(n14905), .A2(n14906), .ZN(n13172) );
  XNOR2_X1 U15553 ( .A(n13170), .B(n13173), .ZN(n14909) );
  OAI21_X1 U15554 ( .B1(n14905), .B2(n14906), .A(n14909), .ZN(n13171) );
  NAND2_X1 U15555 ( .A1(n15531), .A2(n10876), .ZN(n13176) );
  OR2_X1 U15556 ( .A1(n15340), .A2(n13224), .ZN(n13175) );
  NAND2_X1 U15557 ( .A1(n13176), .A2(n13175), .ZN(n13177) );
  XNOR2_X1 U15558 ( .A(n13177), .B(n13233), .ZN(n13180) );
  NOR2_X1 U15559 ( .A1(n15340), .A2(n13223), .ZN(n13178) );
  AOI21_X1 U15560 ( .B1(n15531), .B2(n13189), .A(n13178), .ZN(n13179) );
  NOR2_X1 U15561 ( .A1(n13180), .A2(n13179), .ZN(n14918) );
  NAND2_X1 U15562 ( .A1(n13180), .A2(n13179), .ZN(n14916) );
  XOR2_X1 U15563 ( .A(n13182), .B(n13181), .Z(n14968) );
  NAND2_X1 U15564 ( .A1(n14967), .A2(n14968), .ZN(n14966) );
  OAI22_X1 U15565 ( .A1(n15327), .A2(n13195), .B1(n15341), .B2(n13224), .ZN(
        n13183) );
  XNOR2_X1 U15566 ( .A(n13183), .B(n11908), .ZN(n13185) );
  OAI22_X1 U15567 ( .A1(n15327), .A2(n13224), .B1(n15341), .B2(n13223), .ZN(
        n13184) );
  XNOR2_X1 U15568 ( .A(n13185), .B(n13184), .ZN(n14869) );
  XOR2_X1 U15569 ( .A(n13186), .B(n13187), .Z(n14937) );
  AOI22_X1 U15570 ( .A1(n15507), .A2(n13189), .B1(n13235), .B2(n15002), .ZN(
        n13192) );
  AOI22_X1 U15571 ( .A1(n15507), .A2(n10876), .B1(n13189), .B2(n15002), .ZN(
        n13190) );
  XNOR2_X1 U15572 ( .A(n13190), .B(n11908), .ZN(n13191) );
  XOR2_X1 U15573 ( .A(n13192), .B(n13191), .Z(n14877) );
  NAND2_X1 U15574 ( .A1(n13191), .A2(n13192), .ZN(n13193) );
  OAI22_X1 U15575 ( .A1(n15277), .A2(n13224), .B1(n13194), .B2(n13223), .ZN(
        n13198) );
  OAI22_X1 U15576 ( .A1(n15277), .A2(n13195), .B1(n13194), .B2(n13224), .ZN(
        n13196) );
  XNOR2_X1 U15577 ( .A(n13196), .B(n11908), .ZN(n13197) );
  XOR2_X1 U15578 ( .A(n13198), .B(n13197), .Z(n14943) );
  INV_X1 U15579 ( .A(n13197), .ZN(n13200) );
  OAI22_X1 U15580 ( .A1(n15493), .A2(n13224), .B1(n15274), .B2(n13223), .ZN(
        n13205) );
  NAND2_X1 U15581 ( .A1(n15265), .A2(n10876), .ZN(n13203) );
  NAND2_X1 U15582 ( .A1(n15000), .A2(n13189), .ZN(n13202) );
  NAND2_X1 U15583 ( .A1(n13203), .A2(n13202), .ZN(n13204) );
  XNOR2_X1 U15584 ( .A(n13204), .B(n11908), .ZN(n13206) );
  XOR2_X1 U15585 ( .A(n13205), .B(n13206), .Z(n14861) );
  NAND2_X1 U15586 ( .A1(n14860), .A2(n14861), .ZN(n13208) );
  NAND2_X1 U15587 ( .A1(n15488), .A2(n10876), .ZN(n13210) );
  NAND2_X1 U15588 ( .A1(n14999), .A2(n13189), .ZN(n13209) );
  NAND2_X1 U15589 ( .A1(n13210), .A2(n13209), .ZN(n13211) );
  XNOR2_X1 U15590 ( .A(n13211), .B(n11908), .ZN(n13212) );
  AOI22_X1 U15591 ( .A1(n15488), .A2(n13189), .B1(n13235), .B2(n14999), .ZN(
        n13214) );
  XNOR2_X1 U15592 ( .A(n13212), .B(n13214), .ZN(n14927) );
  INV_X1 U15593 ( .A(n13212), .ZN(n13213) );
  AOI22_X1 U15594 ( .A1(n15482), .A2(n13189), .B1(n13235), .B2(n15212), .ZN(
        n13219) );
  NAND2_X1 U15595 ( .A1(n15482), .A2(n10876), .ZN(n13216) );
  NAND2_X1 U15596 ( .A1(n15212), .A2(n13189), .ZN(n13215) );
  NAND2_X1 U15597 ( .A1(n13216), .A2(n13215), .ZN(n13218) );
  XOR2_X1 U15598 ( .A(n13219), .B(n13221), .Z(n14898) );
  INV_X1 U15599 ( .A(n13219), .ZN(n13220) );
  NAND2_X1 U15600 ( .A1(n15222), .A2(n10876), .ZN(n13227) );
  NAND2_X1 U15601 ( .A1(n14998), .A2(n13189), .ZN(n13226) );
  NAND2_X1 U15602 ( .A1(n13227), .A2(n13226), .ZN(n13228) );
  NAND2_X1 U15603 ( .A1(n15469), .A2(n10876), .ZN(n13232) );
  NAND2_X1 U15604 ( .A1(n15213), .A2(n13189), .ZN(n13231) );
  NAND2_X1 U15605 ( .A1(n13232), .A2(n13231), .ZN(n13234) );
  XNOR2_X1 U15606 ( .A(n13234), .B(n13233), .ZN(n13239) );
  AND2_X1 U15607 ( .A1(n15213), .A2(n13235), .ZN(n13236) );
  AOI21_X1 U15608 ( .B1(n15469), .B2(n13189), .A(n13236), .ZN(n13238) );
  XNOR2_X1 U15609 ( .A(n13239), .B(n13238), .ZN(n14849) );
  INV_X1 U15610 ( .A(n14849), .ZN(n13237) );
  NAND2_X1 U15611 ( .A1(n14850), .A2(n13237), .ZN(n13252) );
  NAND2_X1 U15612 ( .A1(n13239), .A2(n13238), .ZN(n13246) );
  INV_X1 U15613 ( .A(n13246), .ZN(n13240) );
  AND2_X1 U15614 ( .A1(n13247), .A2(n13241), .ZN(n13242) );
  NAND2_X1 U15615 ( .A1(n13252), .A2(n13242), .ZN(n13251) );
  NAND2_X1 U15616 ( .A1(n15213), .A2(n15426), .ZN(n13244) );
  NAND2_X1 U15617 ( .A1(n14997), .A2(n15746), .ZN(n13243) );
  NAND2_X1 U15618 ( .A1(n13244), .A2(n13243), .ZN(n15461) );
  INV_X1 U15619 ( .A(n15461), .ZN(n15194) );
  AOI22_X1 U15620 ( .A1(n15192), .A2(n14928), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13245) );
  OAI21_X1 U15621 ( .B1(n15194), .B2(n14989), .A(n13245), .ZN(n13249) );
  NOR3_X1 U15622 ( .A1(n13247), .A2(n14994), .A3(n13246), .ZN(n13248) );
  AOI211_X1 U15623 ( .C1(n14992), .C2(n15462), .A(n13249), .B(n13248), .ZN(
        n13250) );
  OAI211_X1 U15624 ( .C1(n13253), .C2(n13252), .A(n13251), .B(n13250), .ZN(
        P1_U3220) );
  OAI222_X1 U15625 ( .A1(n13257), .A2(n13256), .B1(n13255), .B2(P3_U3151), 
        .C1(n13254), .C2(n14006), .ZN(P3_U3265) );
  INV_X1 U15626 ( .A(n13258), .ZN(n14833) );
  OAI222_X1 U15627 ( .A1(n15597), .A2(n13259), .B1(n15595), .B2(n14833), .C1(
        P1_U3086), .C2(n8855), .ZN(P1_U3327) );
  NAND3_X1 U15628 ( .A1(n13260), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n13264) );
  NAND2_X1 U15629 ( .A1(n15583), .A2(n13261), .ZN(n13263) );
  NAND2_X1 U15630 ( .A1(n14830), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n13262) );
  OAI211_X1 U15631 ( .C1(n13265), .C2(n13264), .A(n13263), .B(n13262), .ZN(
        P2_U3296) );
  INV_X1 U15632 ( .A(n13266), .ZN(n13268) );
  AOI22_X1 U15633 ( .A1(n14179), .A2(n13268), .B1(n14189), .B2(n13267), .ZN(
        n13273) );
  INV_X1 U15634 ( .A(n13269), .ZN(n13271) );
  AOI22_X1 U15635 ( .A1(n14180), .A2(n13271), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n13270), .ZN(n13272) );
  OAI211_X1 U15636 ( .C1(n13274), .C2(n14184), .A(n13273), .B(n13272), .ZN(
        P2_U3204) );
  INV_X1 U15637 ( .A(n13275), .ZN(n13278) );
  OAI222_X1 U15638 ( .A1(n14826), .A2(n13280), .B1(P2_U3088), .B2(n13279), 
        .C1(n14832), .C2(n13278), .ZN(P2_U3297) );
  NOR2_X1 U15639 ( .A1(n6760), .A2(n13281), .ZN(n13282) );
  OAI21_X1 U15640 ( .B1(n13282), .B2(n13435), .A(n13437), .ZN(n13287) );
  AND2_X1 U15641 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n13505) );
  AOI21_X1 U15642 ( .B1(n13831), .B2(n13430), .A(n13505), .ZN(n13283) );
  OAI21_X1 U15643 ( .B1(n13284), .B2(n13428), .A(n13283), .ZN(n13285) );
  AOI21_X1 U15644 ( .B1(n13823), .B2(n13443), .A(n13285), .ZN(n13286) );
  OAI211_X1 U15645 ( .C1(n13446), .C2(n13996), .A(n13287), .B(n13286), .ZN(
        P3_U3155) );
  NAND2_X1 U15646 ( .A1(n13288), .A2(n13720), .ZN(n13289) );
  AND2_X1 U15647 ( .A1(n13290), .A2(n13289), .ZN(n13295) );
  AOI22_X1 U15648 ( .A1(n13711), .A2(n13443), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13292) );
  NAND2_X1 U15649 ( .A1(n13450), .A2(n13439), .ZN(n13291) );
  OAI211_X1 U15650 ( .C1(n13704), .C2(n13441), .A(n13292), .B(n13291), .ZN(
        n13293) );
  AOI21_X1 U15651 ( .B1(n13710), .B2(n13400), .A(n13293), .ZN(n13294) );
  OAI21_X1 U15652 ( .B1(n13295), .B2(n13413), .A(n13294), .ZN(P3_U3156) );
  AND2_X1 U15653 ( .A1(n13297), .A2(n13296), .ZN(n13300) );
  OAI211_X1 U15654 ( .C1(n13300), .C2(n13299), .A(n13437), .B(n13298), .ZN(
        n13307) );
  NAND2_X1 U15655 ( .A1(n13430), .A2(n13454), .ZN(n13302) );
  OAI211_X1 U15656 ( .C1(n13428), .C2(n13303), .A(n13302), .B(n13301), .ZN(
        n13304) );
  AOI21_X1 U15657 ( .B1(n13305), .B2(n13443), .A(n13304), .ZN(n13306) );
  OAI211_X1 U15658 ( .C1(n13446), .C2(n13308), .A(n13307), .B(n13306), .ZN(
        P3_U3157) );
  INV_X1 U15659 ( .A(n13964), .ZN(n13316) );
  OAI211_X1 U15660 ( .C1(n13311), .C2(n13310), .A(n13309), .B(n13437), .ZN(
        n13315) );
  NAND2_X1 U15661 ( .A1(n13789), .A2(n13439), .ZN(n13312) );
  NAND2_X1 U15662 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13605)
         );
  OAI211_X1 U15663 ( .C1(n13760), .C2(n13441), .A(n13312), .B(n13605), .ZN(
        n13313) );
  AOI21_X1 U15664 ( .B1(n13764), .B2(n13443), .A(n13313), .ZN(n13314) );
  OAI211_X1 U15665 ( .C1(n13316), .C2(n13446), .A(n13315), .B(n13314), .ZN(
        P3_U3159) );
  OAI21_X1 U15666 ( .B1(n13319), .B2(n13318), .A(n13317), .ZN(n13320) );
  NAND2_X1 U15667 ( .A1(n13320), .A2(n13437), .ZN(n13326) );
  INV_X1 U15668 ( .A(n13321), .ZN(n13733) );
  INV_X1 U15669 ( .A(n13760), .ZN(n13451) );
  AOI22_X1 U15670 ( .A1(n13451), .A2(n13439), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13322) );
  OAI21_X1 U15671 ( .B1(n13733), .B2(n13323), .A(n13322), .ZN(n13324) );
  AOI21_X1 U15672 ( .B1(n13430), .B2(n13450), .A(n13324), .ZN(n13325) );
  OAI211_X1 U15673 ( .C1(n13327), .C2(n13446), .A(n13326), .B(n13325), .ZN(
        P3_U3163) );
  NAND2_X1 U15674 ( .A1(n13329), .A2(n13328), .ZN(n13337) );
  INV_X1 U15675 ( .A(n13331), .ZN(n13333) );
  INV_X1 U15676 ( .A(n13330), .ZN(n13332) );
  OR2_X1 U15677 ( .A1(n13331), .A2(n13330), .ZN(n13334) );
  OAI21_X1 U15678 ( .B1(n13333), .B2(n13332), .A(n13334), .ZN(n13404) );
  NOR2_X1 U15679 ( .A1(n13404), .A2(n13454), .ZN(n13403) );
  INV_X1 U15680 ( .A(n13334), .ZN(n13335) );
  NOR2_X1 U15681 ( .A1(n13403), .A2(n13335), .ZN(n13336) );
  XOR2_X1 U15682 ( .A(n13337), .B(n13336), .Z(n13346) );
  NAND2_X1 U15683 ( .A1(n13443), .A2(n13338), .ZN(n13341) );
  AOI21_X1 U15684 ( .B1(n13430), .B2(n13829), .A(n13339), .ZN(n13340) );
  OAI211_X1 U15685 ( .C1(n13342), .C2(n13428), .A(n13341), .B(n13340), .ZN(
        n13343) );
  AOI21_X1 U15686 ( .B1(n13344), .B2(n13400), .A(n13343), .ZN(n13345) );
  OAI21_X1 U15687 ( .B1(n13346), .B2(n13413), .A(n13345), .ZN(P3_U3164) );
  INV_X1 U15688 ( .A(n13348), .ZN(n13350) );
  NOR3_X1 U15689 ( .A1(n7921), .A2(n13350), .A3(n13349), .ZN(n13353) );
  INV_X1 U15690 ( .A(n13351), .ZN(n13352) );
  OAI21_X1 U15691 ( .B1(n13353), .B2(n13352), .A(n13437), .ZN(n13357) );
  AOI22_X1 U15692 ( .A1(n13685), .A2(n13443), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13354) );
  OAI21_X1 U15693 ( .B1(n13704), .B2(n13428), .A(n13354), .ZN(n13355) );
  AOI21_X1 U15694 ( .B1(n6960), .B2(n13430), .A(n13355), .ZN(n13356) );
  OAI211_X1 U15695 ( .C1(n13937), .C2(n13446), .A(n13357), .B(n13356), .ZN(
        P3_U3165) );
  XNOR2_X1 U15696 ( .A(n13358), .B(n13359), .ZN(n13365) );
  NAND2_X1 U15697 ( .A1(n13439), .A2(n13831), .ZN(n13360) );
  NAND2_X1 U15698 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n13544)
         );
  OAI211_X1 U15699 ( .C1(n13773), .C2(n13441), .A(n13360), .B(n13544), .ZN(
        n13363) );
  NOR2_X1 U15700 ( .A1(n13361), .A2(n13446), .ZN(n13362) );
  AOI211_X1 U15701 ( .C1(n13804), .C2(n13443), .A(n13363), .B(n13362), .ZN(
        n13364) );
  OAI21_X1 U15702 ( .B1(n13365), .B2(n13413), .A(n13364), .ZN(P3_U3166) );
  NAND2_X1 U15703 ( .A1(n13367), .A2(n13366), .ZN(n13369) );
  XOR2_X1 U15704 ( .A(n13369), .B(n13368), .Z(n13375) );
  NAND2_X1 U15705 ( .A1(n13788), .A2(n13439), .ZN(n13370) );
  NAND2_X1 U15706 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13560)
         );
  OAI211_X1 U15707 ( .C1(n13759), .C2(n13441), .A(n13370), .B(n13560), .ZN(
        n13373) );
  NOR2_X1 U15708 ( .A1(n13371), .A2(n13446), .ZN(n13372) );
  AOI211_X1 U15709 ( .C1(n13792), .C2(n13443), .A(n13373), .B(n13372), .ZN(
        n13374) );
  OAI21_X1 U15710 ( .B1(n13375), .B2(n13413), .A(n13374), .ZN(P3_U3168) );
  NOR2_X1 U15711 ( .A1(n13377), .A2(n6748), .ZN(n13378) );
  XNOR2_X1 U15712 ( .A(n13376), .B(n13378), .ZN(n13383) );
  AOI22_X1 U15713 ( .A1(n13743), .A2(n13439), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13380) );
  NAND2_X1 U15714 ( .A1(n13747), .A2(n13443), .ZN(n13379) );
  OAI211_X1 U15715 ( .C1(n13398), .C2(n13441), .A(n13380), .B(n13379), .ZN(
        n13381) );
  AOI21_X1 U15716 ( .B1(n13958), .B2(n13400), .A(n13381), .ZN(n13382) );
  OAI21_X1 U15717 ( .B1(n13383), .B2(n13413), .A(n13382), .ZN(P3_U3173) );
  XNOR2_X1 U15718 ( .A(n13384), .B(n13829), .ZN(n13385) );
  XNOR2_X1 U15719 ( .A(n13386), .B(n13385), .ZN(n13394) );
  NAND2_X1 U15720 ( .A1(n13430), .A2(n13452), .ZN(n13387) );
  NAND2_X1 U15721 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n13473)
         );
  OAI211_X1 U15722 ( .C1(n13428), .C2(n13388), .A(n13387), .B(n13473), .ZN(
        n13391) );
  NOR2_X1 U15723 ( .A1(n13389), .A2(n13446), .ZN(n13390) );
  AOI211_X1 U15724 ( .C1(n13392), .C2(n13443), .A(n13391), .B(n13390), .ZN(
        n13393) );
  OAI21_X1 U15725 ( .B1(n13394), .B2(n13413), .A(n13393), .ZN(P3_U3174) );
  AOI21_X1 U15726 ( .B1(n13450), .B2(n13395), .A(n6673), .ZN(n13402) );
  NAND2_X1 U15727 ( .A1(n13720), .A2(n13430), .ZN(n13397) );
  AOI22_X1 U15728 ( .A1(n13723), .A2(n13443), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13396) );
  OAI211_X1 U15729 ( .C1(n13398), .C2(n13428), .A(n13397), .B(n13396), .ZN(
        n13399) );
  AOI21_X1 U15730 ( .B1(n13948), .B2(n13400), .A(n13399), .ZN(n13401) );
  OAI21_X1 U15731 ( .B1(n13402), .B2(n13413), .A(n13401), .ZN(P3_U3175) );
  AOI21_X1 U15732 ( .B1(n13454), .B2(n13404), .A(n13403), .ZN(n13414) );
  NAND2_X1 U15733 ( .A1(n13430), .A2(n13453), .ZN(n13406) );
  OAI211_X1 U15734 ( .C1(n13428), .C2(n13407), .A(n13406), .B(n13405), .ZN(
        n13410) );
  NOR2_X1 U15735 ( .A1(n13408), .A2(n13446), .ZN(n13409) );
  AOI211_X1 U15736 ( .C1(n13411), .C2(n13443), .A(n13410), .B(n13409), .ZN(
        n13412) );
  OAI21_X1 U15737 ( .B1(n13414), .B2(n13413), .A(n13412), .ZN(P3_U3176) );
  INV_X1 U15738 ( .A(n13782), .ZN(n13971) );
  OAI211_X1 U15739 ( .C1(n13417), .C2(n13416), .A(n13415), .B(n13437), .ZN(
        n13421) );
  NAND2_X1 U15740 ( .A1(n13801), .A2(n13439), .ZN(n13418) );
  NAND2_X1 U15741 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13584)
         );
  OAI211_X1 U15742 ( .C1(n13772), .C2(n13441), .A(n13418), .B(n13584), .ZN(
        n13419) );
  AOI21_X1 U15743 ( .B1(n13774), .B2(n13443), .A(n13419), .ZN(n13420) );
  OAI211_X1 U15744 ( .C1(n13971), .C2(n13446), .A(n13421), .B(n13420), .ZN(
        P3_U3178) );
  OAI21_X1 U15745 ( .B1(n13425), .B2(n13424), .A(n13423), .ZN(n13426) );
  NAND2_X1 U15746 ( .A1(n13426), .A2(n13437), .ZN(n13432) );
  AOI22_X1 U15747 ( .A1(n13672), .A2(n13443), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13427) );
  OAI21_X1 U15748 ( .B1(n13692), .B2(n13428), .A(n13427), .ZN(n13429) );
  AOI21_X1 U15749 ( .B1(n13430), .B2(n13666), .A(n13429), .ZN(n13431) );
  OAI211_X1 U15750 ( .C1(n6961), .C2(n13446), .A(n13432), .B(n13431), .ZN(
        P3_U3180) );
  OAI21_X1 U15751 ( .B1(n13435), .B2(n13434), .A(n13433), .ZN(n13438) );
  NAND3_X1 U15752 ( .A1(n13438), .A2(n13437), .A3(n13436), .ZN(n13445) );
  NAND2_X1 U15753 ( .A1(n13439), .A2(n13452), .ZN(n13440) );
  NAND2_X1 U15754 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n13521)
         );
  OAI211_X1 U15755 ( .C1(n13812), .C2(n13441), .A(n13440), .B(n13521), .ZN(
        n13442) );
  AOI21_X1 U15756 ( .B1(n13815), .B2(n13443), .A(n13442), .ZN(n13444) );
  OAI211_X1 U15757 ( .C1(n13446), .C2(n13817), .A(n13445), .B(n13444), .ZN(
        P3_U3181) );
  MUX2_X1 U15758 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n13447), .S(n13461), .Z(
        P3_U3522) );
  MUX2_X1 U15759 ( .A(n13448), .B(P3_DATAO_REG_28__SCAN_IN), .S(n13463), .Z(
        P3_U3519) );
  MUX2_X1 U15760 ( .A(n13666), .B(P3_DATAO_REG_27__SCAN_IN), .S(n13463), .Z(
        P3_U3518) );
  MUX2_X1 U15761 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n6960), .S(n13461), .Z(
        P3_U3517) );
  MUX2_X1 U15762 ( .A(n13665), .B(P3_DATAO_REG_25__SCAN_IN), .S(n13463), .Z(
        P3_U3516) );
  MUX2_X1 U15763 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n13449), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U15764 ( .A(n13720), .B(P3_DATAO_REG_23__SCAN_IN), .S(n13463), .Z(
        P3_U3514) );
  MUX2_X1 U15765 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n13450), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15766 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n13744), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U15767 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13451), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15768 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n13743), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U15769 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13789), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15770 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13801), .S(n13461), .Z(
        P3_U3508) );
  MUX2_X1 U15771 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n13788), .S(n13461), .Z(
        P3_U3507) );
  MUX2_X1 U15772 ( .A(n13831), .B(P3_DATAO_REG_15__SCAN_IN), .S(n13463), .Z(
        P3_U3506) );
  MUX2_X1 U15773 ( .A(n13452), .B(P3_DATAO_REG_14__SCAN_IN), .S(n13463), .Z(
        P3_U3505) );
  MUX2_X1 U15774 ( .A(n13829), .B(P3_DATAO_REG_13__SCAN_IN), .S(n13463), .Z(
        P3_U3504) );
  MUX2_X1 U15775 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n13453), .S(n13461), .Z(
        P3_U3503) );
  MUX2_X1 U15776 ( .A(n13454), .B(P3_DATAO_REG_11__SCAN_IN), .S(n13463), .Z(
        P3_U3502) );
  MUX2_X1 U15777 ( .A(n13455), .B(P3_DATAO_REG_10__SCAN_IN), .S(n13463), .Z(
        P3_U3501) );
  MUX2_X1 U15778 ( .A(n13456), .B(P3_DATAO_REG_8__SCAN_IN), .S(n13463), .Z(
        P3_U3499) );
  MUX2_X1 U15779 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n13457), .S(n13461), .Z(
        P3_U3498) );
  MUX2_X1 U15780 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n13458), .S(n13461), .Z(
        P3_U3497) );
  MUX2_X1 U15781 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n13459), .S(n13461), .Z(
        P3_U3496) );
  MUX2_X1 U15782 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n13460), .S(n13461), .Z(
        P3_U3495) );
  MUX2_X1 U15783 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n10901), .S(n13461), .Z(
        P3_U3494) );
  MUX2_X1 U15784 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n13462), .S(n13461), .Z(
        P3_U3493) );
  MUX2_X1 U15785 ( .A(n8170), .B(P3_DATAO_REG_1__SCAN_IN), .S(n13463), .Z(
        P3_U3492) );
  MUX2_X1 U15786 ( .A(n13464), .B(P3_DATAO_REG_0__SCAN_IN), .S(n13463), .Z(
        P3_U3491) );
  INV_X1 U15787 ( .A(n13486), .ZN(n13496) );
  XOR2_X1 U15788 ( .A(P3_REG1_REG_13__SCAN_IN), .B(n13487), .Z(n13485) );
  NAND2_X1 U15789 ( .A1(n13467), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n13468) );
  NAND2_X1 U15790 ( .A1(n13469), .A2(n13468), .ZN(n13470) );
  OAI21_X1 U15791 ( .B1(P3_REG2_REG_13__SCAN_IN), .B2(n13471), .A(n13493), 
        .ZN(n13483) );
  NAND2_X1 U15792 ( .A1(n15945), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n13472) );
  OAI211_X1 U15793 ( .C1(n13586), .C2(n13486), .A(n13473), .B(n13472), .ZN(
        n13482) );
  INV_X1 U15794 ( .A(n13474), .ZN(n13476) );
  NOR2_X1 U15795 ( .A1(n13476), .A2(n13475), .ZN(n13478) );
  MUX2_X1 U15796 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13576), .Z(n13495) );
  XNOR2_X1 U15797 ( .A(n13495), .B(n13486), .ZN(n13477) );
  OAI21_X1 U15798 ( .B1(n13479), .B2(n13478), .A(n13477), .ZN(n13480) );
  AOI21_X1 U15799 ( .B1(n7350), .B2(n13480), .A(n13622), .ZN(n13481) );
  AOI211_X1 U15800 ( .C1(n13621), .C2(n13483), .A(n13482), .B(n13481), .ZN(
        n13484) );
  OAI21_X1 U15801 ( .B1(n13485), .B2(n13612), .A(n13484), .ZN(P3_U3195) );
  NAND2_X1 U15802 ( .A1(n13508), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n13517) );
  OAI21_X1 U15803 ( .B1(n13508), .B2(P3_REG1_REG_14__SCAN_IN), .A(n13517), 
        .ZN(n13498) );
  INV_X1 U15804 ( .A(n13518), .ZN(n13490) );
  AOI21_X1 U15805 ( .B1(n13491), .B2(n13498), .A(n13490), .ZN(n13512) );
  NAND2_X1 U15806 ( .A1(n13508), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n13525) );
  OAI21_X1 U15807 ( .B1(n13508), .B2(P3_REG2_REG_14__SCAN_IN), .A(n13525), 
        .ZN(n13499) );
  NAND3_X1 U15808 ( .A1(n13493), .A2(n13499), .A3(n13492), .ZN(n13494) );
  NAND2_X1 U15809 ( .A1(n13526), .A2(n13494), .ZN(n13510) );
  INV_X1 U15810 ( .A(n13495), .ZN(n13497) );
  AND2_X1 U15811 ( .A1(n13497), .A2(n13496), .ZN(n13501) );
  MUX2_X1 U15812 ( .A(n13499), .B(n13498), .S(n13576), .Z(n13500) );
  OAI21_X1 U15813 ( .B1(n13502), .B2(n13501), .A(n13500), .ZN(n13504) );
  NAND3_X1 U15814 ( .A1(n13504), .A2(n13503), .A3(n13514), .ZN(n13507) );
  AOI21_X1 U15815 ( .B1(n15945), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n13505), 
        .ZN(n13506) );
  OAI211_X1 U15816 ( .C1(n13586), .C2(n13508), .A(n13507), .B(n13506), .ZN(
        n13509) );
  AOI21_X1 U15817 ( .B1(n13621), .B2(n13510), .A(n13509), .ZN(n13511) );
  OAI21_X1 U15818 ( .B1(n13512), .B2(n13612), .A(n13511), .ZN(P3_U3196) );
  MUX2_X1 U15819 ( .A(n13525), .B(n13517), .S(n13576), .Z(n13513) );
  XNOR2_X1 U15820 ( .A(n13539), .B(n13534), .ZN(n13516) );
  MUX2_X1 U15821 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n13576), .Z(n13515) );
  NOR2_X1 U15822 ( .A1(n13516), .A2(n13515), .ZN(n13540) );
  AOI21_X1 U15823 ( .B1(n13516), .B2(n13515), .A(n13540), .ZN(n13532) );
  INV_X1 U15824 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n13523) );
  OAI21_X1 U15825 ( .B1(n13519), .B2(P3_REG1_REG_15__SCAN_IN), .A(n13535), 
        .ZN(n13520) );
  NAND2_X1 U15826 ( .A1(n13589), .A2(n13520), .ZN(n13522) );
  OAI211_X1 U15827 ( .C1(n13606), .C2(n13523), .A(n13522), .B(n13521), .ZN(
        n13524) );
  AOI21_X1 U15828 ( .B1(n7708), .B2(n13615), .A(n13524), .ZN(n13531) );
  OAI21_X1 U15829 ( .B1(P3_REG2_REG_15__SCAN_IN), .B2(n13528), .A(n13548), 
        .ZN(n13529) );
  NAND2_X1 U15830 ( .A1(n13529), .A2(n13621), .ZN(n13530) );
  OAI211_X1 U15831 ( .C1(n13532), .C2(n13622), .A(n13531), .B(n13530), .ZN(
        P3_U3197) );
  NAND2_X1 U15832 ( .A1(n13534), .A2(n13533), .ZN(n13536) );
  XNOR2_X1 U15833 ( .A(n13556), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n13537) );
  OAI21_X1 U15834 ( .B1(n13538), .B2(n13537), .A(n13557), .ZN(n13554) );
  INV_X1 U15835 ( .A(n13539), .ZN(n13541) );
  INV_X1 U15836 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13803) );
  INV_X1 U15837 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13892) );
  MUX2_X1 U15838 ( .A(n13803), .B(n13892), .S(n13576), .Z(n13542) );
  NOR2_X1 U15839 ( .A1(n13556), .A2(n13542), .ZN(n13561) );
  NOR2_X1 U15840 ( .A1(n13561), .A2(n6765), .ZN(n13543) );
  XNOR2_X1 U15841 ( .A(n13562), .B(n13543), .ZN(n13552) );
  INV_X1 U15842 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n15636) );
  OAI21_X1 U15843 ( .B1(n13606), .B2(n15636), .A(n13544), .ZN(n13545) );
  AOI21_X1 U15844 ( .B1(n13556), .B2(n13615), .A(n13545), .ZN(n13551) );
  XNOR2_X1 U15845 ( .A(n13556), .B(n13803), .ZN(n13547) );
  AND3_X1 U15846 ( .A1(n13548), .A2(n13547), .A3(n13546), .ZN(n13549) );
  OAI21_X1 U15847 ( .B1(n13568), .B2(n13549), .A(n13621), .ZN(n13550) );
  OAI211_X1 U15848 ( .C1(n13552), .C2(n13622), .A(n13551), .B(n13550), .ZN(
        n13553) );
  AOI21_X1 U15849 ( .B1(n13589), .B2(n13554), .A(n13553), .ZN(n13555) );
  INV_X1 U15850 ( .A(n13555), .ZN(P3_U3198) );
  OR2_X1 U15851 ( .A1(n13556), .A2(n13892), .ZN(n13558) );
  XNOR2_X1 U15852 ( .A(n13582), .B(P3_REG1_REG_17__SCAN_IN), .ZN(n13567) );
  NAND2_X1 U15853 ( .A1(n15945), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n13559) );
  OAI211_X1 U15854 ( .C1(n13586), .C2(n13581), .A(n13560), .B(n13559), .ZN(
        n13566) );
  MUX2_X1 U15855 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13576), .Z(n13577) );
  XNOR2_X1 U15856 ( .A(n13581), .B(n13577), .ZN(n13564) );
  AOI211_X1 U15857 ( .C1(n13564), .C2(n13563), .A(n13622), .B(n6669), .ZN(
        n13565) );
  AOI211_X1 U15858 ( .C1(n13589), .C2(n13567), .A(n13566), .B(n13565), .ZN(
        n13575) );
  INV_X1 U15859 ( .A(n13581), .ZN(n13570) );
  AOI21_X1 U15860 ( .B1(n13571), .B2(n13570), .A(n13590), .ZN(n13572) );
  NAND2_X1 U15861 ( .A1(n13572), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n13594) );
  OAI21_X1 U15862 ( .B1(P3_REG2_REG_17__SCAN_IN), .B2(n13572), .A(n13594), 
        .ZN(n13573) );
  NAND2_X1 U15863 ( .A1(n13573), .A2(n13621), .ZN(n13574) );
  NAND2_X1 U15864 ( .A1(n13575), .A2(n13574), .ZN(P3_U3199) );
  MUX2_X1 U15865 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n13576), .Z(n13579) );
  XNOR2_X1 U15866 ( .A(n13602), .B(n13607), .ZN(n13578) );
  NOR2_X1 U15867 ( .A1(n13578), .A2(n13579), .ZN(n13601) );
  AOI21_X1 U15868 ( .B1(n13579), .B2(n13578), .A(n13601), .ZN(n13598) );
  XOR2_X1 U15869 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n13607), .Z(n13608) );
  XNOR2_X1 U15870 ( .A(n13609), .B(n13608), .ZN(n13588) );
  NAND2_X1 U15871 ( .A1(n15945), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n13583) );
  OAI211_X1 U15872 ( .C1(n13586), .C2(n13585), .A(n13584), .B(n13583), .ZN(
        n13587) );
  AOI21_X1 U15873 ( .B1(n13589), .B2(n13588), .A(n13587), .ZN(n13597) );
  INV_X1 U15874 ( .A(n13590), .ZN(n13593) );
  INV_X1 U15875 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13776) );
  OR2_X1 U15876 ( .A1(n13607), .A2(n13776), .ZN(n13617) );
  NAND2_X1 U15877 ( .A1(n13607), .A2(n13776), .ZN(n13591) );
  NAND2_X1 U15878 ( .A1(n13617), .A2(n13591), .ZN(n13592) );
  AND3_X1 U15879 ( .A1(n13594), .A2(n13593), .A3(n13592), .ZN(n13595) );
  OAI21_X1 U15880 ( .B1(n13619), .B2(n13595), .A(n13621), .ZN(n13596) );
  OAI211_X1 U15881 ( .C1(n13598), .C2(n13622), .A(n13597), .B(n13596), .ZN(
        P3_U3200) );
  XNOR2_X1 U15882 ( .A(n13599), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13610) );
  XNOR2_X1 U15883 ( .A(n13599), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n13620) );
  MUX2_X1 U15884 ( .A(n13610), .B(n13620), .S(n13600), .Z(n13604) );
  AOI21_X1 U15885 ( .B1(n13602), .B2(n13607), .A(n13601), .ZN(n13603) );
  OAI21_X1 U15886 ( .B1(n13606), .B2(n15661), .A(n13605), .ZN(n13614) );
  XNOR2_X1 U15887 ( .A(n13611), .B(n13610), .ZN(n13613) );
  INV_X1 U15888 ( .A(n13617), .ZN(n13618) );
  NOR2_X1 U15889 ( .A1(n13625), .A2(n15985), .ZN(n13630) );
  AOI21_X1 U15890 ( .B1(n13912), .B2(n15995), .A(n13630), .ZN(n13628) );
  NAND2_X1 U15891 ( .A1(n15997), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n13626) );
  OAI211_X1 U15892 ( .C1(n13914), .C2(n13825), .A(n13628), .B(n13626), .ZN(
        P3_U3202) );
  INV_X1 U15893 ( .A(n13915), .ZN(n13629) );
  NAND2_X1 U15894 ( .A1(n15997), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n13627) );
  OAI211_X1 U15895 ( .C1(n13629), .C2(n13825), .A(n13628), .B(n13627), .ZN(
        P3_U3203) );
  AOI21_X1 U15896 ( .B1(n13844), .B2(n15958), .A(n13630), .ZN(n13632) );
  NAND2_X1 U15897 ( .A1(n13845), .A2(n13837), .ZN(n13631) );
  NAND3_X1 U15898 ( .A1(n13633), .A2(n13632), .A3(n13631), .ZN(P3_U3204) );
  INV_X1 U15899 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n13644) );
  INV_X1 U15900 ( .A(n13651), .ZN(n13637) );
  OAI22_X1 U15901 ( .A1(n13640), .A2(n15992), .B1(n13639), .B2(n15990), .ZN(
        n13641) );
  AOI21_X1 U15902 ( .B1(n13643), .B2(n13642), .A(n13641), .ZN(n13919) );
  AOI22_X1 U15903 ( .A1(n13921), .A2(n15958), .B1(n15977), .B2(n13645), .ZN(
        n13646) );
  INV_X1 U15904 ( .A(n13928), .ZN(n13662) );
  INV_X1 U15905 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n13658) );
  INV_X1 U15906 ( .A(n13650), .ZN(n13653) );
  OAI22_X1 U15907 ( .A1(n13655), .A2(n15992), .B1(n13654), .B2(n15990), .ZN(
        n13656) );
  MUX2_X1 U15908 ( .A(n13658), .B(n13925), .S(n15995), .Z(n13661) );
  AOI22_X1 U15909 ( .A1(n13927), .A2(n15958), .B1(n15977), .B2(n13659), .ZN(
        n13660) );
  OAI211_X1 U15910 ( .C1(n13662), .C2(n13807), .A(n13661), .B(n13660), .ZN(
        P3_U3206) );
  XNOR2_X1 U15911 ( .A(n13664), .B(n13663), .ZN(n13671) );
  AOI22_X1 U15912 ( .A1(n13666), .A2(n13830), .B1(n13828), .B2(n13665), .ZN(
        n13670) );
  NAND2_X1 U15913 ( .A1(n13855), .A2(n15969), .ZN(n13669) );
  INV_X1 U15914 ( .A(n13854), .ZN(n13676) );
  AOI22_X1 U15915 ( .A1(n13672), .A2(n15977), .B1(n15997), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n13673) );
  OAI21_X1 U15916 ( .B1(n6961), .B2(n13825), .A(n13673), .ZN(n13674) );
  AOI21_X1 U15917 ( .B1(n13855), .B2(n13714), .A(n13674), .ZN(n13675) );
  OAI21_X1 U15918 ( .B1(n13676), .B2(n15997), .A(n13675), .ZN(P3_U3207) );
  OAI211_X1 U15919 ( .C1(n13679), .C2(n13678), .A(n13677), .B(n13833), .ZN(
        n13681) );
  NAND2_X1 U15920 ( .A1(n6960), .A2(n13830), .ZN(n13680) );
  OAI211_X1 U15921 ( .C1(n13704), .C2(n15990), .A(n13681), .B(n13680), .ZN(
        n13858) );
  INV_X1 U15922 ( .A(n13858), .ZN(n13689) );
  OAI21_X1 U15923 ( .B1(n13684), .B2(n13683), .A(n13682), .ZN(n13859) );
  AOI22_X1 U15924 ( .A1(n13685), .A2(n15977), .B1(n15997), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n13686) );
  OAI21_X1 U15925 ( .B1(n13937), .B2(n13825), .A(n13686), .ZN(n13687) );
  AOI21_X1 U15926 ( .B1(n13859), .B2(n13837), .A(n13687), .ZN(n13688) );
  OAI21_X1 U15927 ( .B1(n13689), .B2(n15997), .A(n13688), .ZN(P3_U3208) );
  XNOR2_X1 U15928 ( .A(n13690), .B(n13695), .ZN(n13691) );
  OAI222_X1 U15929 ( .A1(n15990), .A2(n13693), .B1(n15992), .B2(n13692), .C1(
        n15988), .C2(n13691), .ZN(n13862) );
  INV_X1 U15930 ( .A(n13862), .ZN(n13700) );
  OAI21_X1 U15931 ( .B1(n6647), .B2(n13695), .A(n13694), .ZN(n13863) );
  AOI22_X1 U15932 ( .A1(n13696), .A2(n15977), .B1(n15997), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n13697) );
  OAI21_X1 U15933 ( .B1(n13941), .B2(n13825), .A(n13697), .ZN(n13698) );
  AOI21_X1 U15934 ( .B1(n13863), .B2(n13837), .A(n13698), .ZN(n13699) );
  OAI21_X1 U15935 ( .B1(n13700), .B2(n15997), .A(n13699), .ZN(P3_U3209) );
  INV_X1 U15936 ( .A(n15969), .ZN(n13708) );
  XNOR2_X1 U15937 ( .A(n13701), .B(n13702), .ZN(n13709) );
  XNOR2_X1 U15938 ( .A(n16036), .B(n13702), .ZN(n13706) );
  OAI22_X1 U15939 ( .A1(n13704), .A2(n15992), .B1(n13731), .B2(n15990), .ZN(
        n13705) );
  AOI21_X1 U15940 ( .B1(n13706), .B2(n13833), .A(n13705), .ZN(n13707) );
  OAI21_X1 U15941 ( .B1(n13708), .B2(n13709), .A(n13707), .ZN(n13866) );
  INV_X1 U15942 ( .A(n13866), .ZN(n13716) );
  INV_X1 U15943 ( .A(n13709), .ZN(n13867) );
  INV_X1 U15944 ( .A(n13710), .ZN(n13945) );
  AOI22_X1 U15945 ( .A1(n13711), .A2(n15977), .B1(n15997), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n13712) );
  OAI21_X1 U15946 ( .B1(n13945), .B2(n13825), .A(n13712), .ZN(n13713) );
  AOI21_X1 U15947 ( .B1(n13867), .B2(n13714), .A(n13713), .ZN(n13715) );
  OAI21_X1 U15948 ( .B1(n13716), .B2(n15997), .A(n13715), .ZN(P3_U3210) );
  XNOR2_X1 U15949 ( .A(n13717), .B(n13718), .ZN(n13949) );
  INV_X1 U15950 ( .A(n13949), .ZN(n13726) );
  XNOR2_X1 U15951 ( .A(n13719), .B(n13718), .ZN(n13721) );
  AOI222_X1 U15952 ( .A1(n13833), .A2(n13721), .B1(n13720), .B2(n13830), .C1(
        n13744), .C2(n13828), .ZN(n13946) );
  MUX2_X1 U15953 ( .A(n13722), .B(n13946), .S(n15995), .Z(n13725) );
  AOI22_X1 U15954 ( .A1(n13948), .A2(n15958), .B1(n15977), .B2(n13723), .ZN(
        n13724) );
  OAI211_X1 U15955 ( .C1(n13726), .C2(n13807), .A(n13725), .B(n13724), .ZN(
        P3_U3211) );
  XNOR2_X1 U15956 ( .A(n13727), .B(n13728), .ZN(n13955) );
  XOR2_X1 U15957 ( .A(n13729), .B(n13728), .Z(n13730) );
  OAI222_X1 U15958 ( .A1(n15990), .A2(n13760), .B1(n15992), .B2(n13731), .C1(
        n15988), .C2(n13730), .ZN(n13873) );
  NAND2_X1 U15959 ( .A1(n13873), .A2(n15995), .ZN(n13736) );
  OAI22_X1 U15960 ( .A1(n13733), .A2(n15985), .B1(n15995), .B2(n13732), .ZN(
        n13734) );
  AOI21_X1 U15961 ( .B1(n13874), .B2(n15958), .A(n13734), .ZN(n13735) );
  OAI211_X1 U15962 ( .C1(n13955), .C2(n13807), .A(n13736), .B(n13735), .ZN(
        P3_U3212) );
  OAI21_X1 U15963 ( .B1(n13738), .B2(n12895), .A(n13737), .ZN(n13961) );
  INV_X1 U15964 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n13746) );
  NAND2_X1 U15965 ( .A1(n13768), .A2(n13739), .ZN(n13754) );
  NAND2_X1 U15966 ( .A1(n13754), .A2(n13740), .ZN(n13757) );
  NAND2_X1 U15967 ( .A1(n13757), .A2(n13741), .ZN(n13742) );
  XNOR2_X1 U15968 ( .A(n13742), .B(n12895), .ZN(n13745) );
  AOI222_X1 U15969 ( .A1(n13833), .A2(n13745), .B1(n13744), .B2(n13830), .C1(
        n13743), .C2(n13828), .ZN(n13956) );
  MUX2_X1 U15970 ( .A(n13746), .B(n13956), .S(n15995), .Z(n13749) );
  AOI22_X1 U15971 ( .A1(n13958), .A2(n15958), .B1(n15977), .B2(n13747), .ZN(
        n13748) );
  OAI211_X1 U15972 ( .C1(n13961), .C2(n13807), .A(n13749), .B(n13748), .ZN(
        P3_U3213) );
  INV_X1 U15973 ( .A(n13750), .ZN(n13786) );
  AOI21_X1 U15974 ( .B1(n13785), .B2(n13786), .A(n13751), .ZN(n13778) );
  NAND2_X1 U15975 ( .A1(n13778), .A2(n13777), .ZN(n13885) );
  NAND2_X1 U15976 ( .A1(n13885), .A2(n13752), .ZN(n13753) );
  XOR2_X1 U15977 ( .A(n13755), .B(n13753), .Z(n13965) );
  INV_X1 U15978 ( .A(n13965), .ZN(n13767) );
  INV_X1 U15979 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13763) );
  INV_X1 U15980 ( .A(n13754), .ZN(n13769) );
  OAI21_X1 U15981 ( .B1(n13769), .B2(n13756), .A(n13755), .ZN(n13758) );
  AND3_X1 U15982 ( .A1(n13758), .A2(n13833), .A3(n13757), .ZN(n13762) );
  OAI22_X1 U15983 ( .A1(n13760), .A2(n15992), .B1(n13759), .B2(n15990), .ZN(
        n13761) );
  NOR2_X1 U15984 ( .A1(n13762), .A2(n13761), .ZN(n13962) );
  MUX2_X1 U15985 ( .A(n13763), .B(n13962), .S(n15995), .Z(n13766) );
  AOI22_X1 U15986 ( .A1(n13964), .A2(n15958), .B1(n15977), .B2(n13764), .ZN(
        n13765) );
  OAI211_X1 U15987 ( .C1(n13767), .C2(n13807), .A(n13766), .B(n13765), .ZN(
        P3_U3214) );
  INV_X1 U15988 ( .A(n13768), .ZN(n13770) );
  AOI21_X1 U15989 ( .B1(n13777), .B2(n13770), .A(n13769), .ZN(n13771) );
  OAI222_X1 U15990 ( .A1(n15990), .A2(n13773), .B1(n15992), .B2(n13772), .C1(
        n15988), .C2(n13771), .ZN(n13884) );
  INV_X1 U15991 ( .A(n13884), .ZN(n13784) );
  INV_X1 U15992 ( .A(n13774), .ZN(n13775) );
  OAI22_X1 U15993 ( .A1(n15995), .A2(n13776), .B1(n13775), .B2(n15985), .ZN(
        n13781) );
  NOR2_X1 U15994 ( .A1(n13778), .A2(n13777), .ZN(n13883) );
  INV_X1 U15995 ( .A(n13885), .ZN(n13779) );
  NOR3_X1 U15996 ( .A1(n13883), .A2(n13779), .A3(n13807), .ZN(n13780) );
  AOI211_X1 U15997 ( .C1(n15958), .C2(n13782), .A(n13781), .B(n13780), .ZN(
        n13783) );
  OAI21_X1 U15998 ( .B1(n13784), .B2(n15997), .A(n13783), .ZN(P3_U3215) );
  XNOR2_X1 U15999 ( .A(n13785), .B(n13786), .ZN(n13975) );
  INV_X1 U16000 ( .A(n13975), .ZN(n13795) );
  INV_X1 U16001 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13791) );
  XNOR2_X1 U16002 ( .A(n13787), .B(n13786), .ZN(n13790) );
  AOI222_X1 U16003 ( .A1(n13833), .A2(n13790), .B1(n13789), .B2(n13830), .C1(
        n13788), .C2(n13828), .ZN(n13972) );
  MUX2_X1 U16004 ( .A(n13791), .B(n13972), .S(n15995), .Z(n13794) );
  AOI22_X1 U16005 ( .A1(n13974), .A2(n15958), .B1(n15977), .B2(n13792), .ZN(
        n13793) );
  OAI211_X1 U16006 ( .C1(n13795), .C2(n13807), .A(n13794), .B(n13793), .ZN(
        P3_U3216) );
  OAI21_X1 U16007 ( .B1(n13798), .B2(n13797), .A(n13796), .ZN(n13982) );
  INV_X1 U16008 ( .A(n13982), .ZN(n13808) );
  XNOR2_X1 U16009 ( .A(n13800), .B(n13799), .ZN(n13802) );
  AOI222_X1 U16010 ( .A1(n13833), .A2(n13802), .B1(n13801), .B2(n13830), .C1(
        n13831), .C2(n13828), .ZN(n13978) );
  MUX2_X1 U16011 ( .A(n13803), .B(n13978), .S(n15995), .Z(n13806) );
  AOI22_X1 U16012 ( .A1(n13980), .A2(n15958), .B1(n15977), .B2(n13804), .ZN(
        n13805) );
  OAI211_X1 U16013 ( .C1(n13808), .C2(n13807), .A(n13806), .B(n13805), .ZN(
        P3_U3217) );
  XNOR2_X1 U16014 ( .A(n13809), .B(n13814), .ZN(n13810) );
  OAI222_X1 U16015 ( .A1(n15992), .A2(n13812), .B1(n15990), .B2(n13811), .C1(
        n13810), .C2(n15988), .ZN(n13896) );
  INV_X1 U16016 ( .A(n13896), .ZN(n13821) );
  XNOR2_X1 U16017 ( .A(n13813), .B(n13814), .ZN(n13989) );
  INV_X1 U16018 ( .A(n13989), .ZN(n13819) );
  AOI22_X1 U16019 ( .A1(n15997), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15977), 
        .B2(n13815), .ZN(n13816) );
  OAI21_X1 U16020 ( .B1(n13817), .B2(n13825), .A(n13816), .ZN(n13818) );
  AOI21_X1 U16021 ( .B1(n13819), .B2(n13837), .A(n13818), .ZN(n13820) );
  OAI21_X1 U16022 ( .B1(n13821), .B2(n15997), .A(n13820), .ZN(P3_U3218) );
  XOR2_X1 U16023 ( .A(n13826), .B(n13822), .Z(n13993) );
  INV_X1 U16024 ( .A(n13823), .ZN(n13824) );
  OAI22_X1 U16025 ( .A1(n13996), .A2(n13825), .B1(n13824), .B2(n15985), .ZN(
        n13836) );
  XOR2_X1 U16026 ( .A(n13827), .B(n13826), .Z(n13832) );
  AOI222_X1 U16027 ( .A1(n13833), .A2(n13832), .B1(n13831), .B2(n13830), .C1(
        n13829), .C2(n13828), .ZN(n13990) );
  INV_X1 U16028 ( .A(n13990), .ZN(n13834) );
  MUX2_X1 U16029 ( .A(P3_REG2_REG_14__SCAN_IN), .B(n13834), .S(n15995), .Z(
        n13835) );
  AOI211_X1 U16030 ( .C1(n13837), .C2(n13993), .A(n13836), .B(n13835), .ZN(
        n13838) );
  INV_X1 U16031 ( .A(n13838), .ZN(P3_U3219) );
  NAND2_X1 U16032 ( .A1(n13912), .A2(n13911), .ZN(n13840) );
  NAND2_X1 U16033 ( .A1(n16023), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n13839) );
  OAI211_X1 U16034 ( .C1(n13914), .C2(n13905), .A(n13840), .B(n13839), .ZN(
        P3_U3490) );
  NAND2_X1 U16035 ( .A1(n13915), .A2(n13893), .ZN(n13841) );
  OAI211_X1 U16036 ( .C1(n13911), .C2(n12265), .A(n13841), .B(n13840), .ZN(
        P3_U3489) );
  INV_X1 U16037 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n13843) );
  MUX2_X1 U16038 ( .A(n13843), .B(n13842), .S(n13911), .Z(n13847) );
  MUX2_X1 U16039 ( .A(n13848), .B(n13919), .S(n13911), .Z(n13850) );
  NAND2_X1 U16040 ( .A1(n13850), .A2(n13849), .ZN(P3_U3487) );
  MUX2_X1 U16041 ( .A(n13851), .B(n13925), .S(n13911), .Z(n13853) );
  AOI22_X1 U16042 ( .A1(n13928), .A2(n13902), .B1(n13893), .B2(n13927), .ZN(
        n13852) );
  NAND2_X1 U16043 ( .A1(n13853), .A2(n13852), .ZN(P3_U3486) );
  MUX2_X1 U16044 ( .A(n13856), .B(n13931), .S(n13911), .Z(n13857) );
  OAI21_X1 U16045 ( .B1(n6961), .B2(n13905), .A(n13857), .ZN(P3_U3485) );
  AOI21_X1 U16046 ( .B1(n16007), .B2(n13859), .A(n13858), .ZN(n13934) );
  MUX2_X1 U16047 ( .A(n13860), .B(n13934), .S(n13911), .Z(n13861) );
  OAI21_X1 U16048 ( .B1(n13937), .B2(n13905), .A(n13861), .ZN(P3_U3484) );
  AOI21_X1 U16049 ( .B1(n16007), .B2(n13863), .A(n13862), .ZN(n13938) );
  MUX2_X1 U16050 ( .A(n13864), .B(n13938), .S(n13911), .Z(n13865) );
  OAI21_X1 U16051 ( .B1(n13941), .B2(n13905), .A(n13865), .ZN(P3_U3483) );
  AOI21_X1 U16052 ( .B1(n16013), .B2(n13867), .A(n13866), .ZN(n13942) );
  MUX2_X1 U16053 ( .A(n13868), .B(n13942), .S(n13911), .Z(n13869) );
  OAI21_X1 U16054 ( .B1(n13945), .B2(n13905), .A(n13869), .ZN(P3_U3482) );
  INV_X1 U16055 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13870) );
  MUX2_X1 U16056 ( .A(n13870), .B(n13946), .S(n13911), .Z(n13872) );
  AOI22_X1 U16057 ( .A1(n13949), .A2(n13902), .B1(n13893), .B2(n13948), .ZN(
        n13871) );
  NAND2_X1 U16058 ( .A1(n13872), .A2(n13871), .ZN(P3_U3481) );
  INV_X1 U16059 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13875) );
  AOI21_X1 U16060 ( .B1(n16011), .B2(n13874), .A(n13873), .ZN(n13952) );
  MUX2_X1 U16061 ( .A(n13875), .B(n13952), .S(n13911), .Z(n13876) );
  OAI21_X1 U16062 ( .B1(n13900), .B2(n13955), .A(n13876), .ZN(P3_U3480) );
  MUX2_X1 U16063 ( .A(n13877), .B(n13956), .S(n13911), .Z(n13879) );
  NAND2_X1 U16064 ( .A1(n13958), .A2(n13893), .ZN(n13878) );
  OAI211_X1 U16065 ( .C1(n13900), .C2(n13961), .A(n13879), .B(n13878), .ZN(
        P3_U3479) );
  MUX2_X1 U16066 ( .A(n13880), .B(n13962), .S(n13911), .Z(n13882) );
  AOI22_X1 U16067 ( .A1(n13965), .A2(n13902), .B1(n13893), .B2(n13964), .ZN(
        n13881) );
  NAND2_X1 U16068 ( .A1(n13882), .A2(n13881), .ZN(P3_U3478) );
  NOR2_X1 U16069 ( .A1(n13883), .A2(n13909), .ZN(n13886) );
  AOI21_X1 U16070 ( .B1(n13886), .B2(n13885), .A(n13884), .ZN(n13968) );
  MUX2_X1 U16071 ( .A(n13887), .B(n13968), .S(n13911), .Z(n13888) );
  OAI21_X1 U16072 ( .B1(n13971), .B2(n13905), .A(n13888), .ZN(P3_U3477) );
  MUX2_X1 U16073 ( .A(n13889), .B(n13972), .S(n13911), .Z(n13891) );
  AOI22_X1 U16074 ( .A1(n13975), .A2(n13902), .B1(n13974), .B2(n13893), .ZN(
        n13890) );
  NAND2_X1 U16075 ( .A1(n13891), .A2(n13890), .ZN(P3_U3476) );
  MUX2_X1 U16076 ( .A(n13892), .B(n13978), .S(n13911), .Z(n13895) );
  AOI22_X1 U16077 ( .A1(n13982), .A2(n13902), .B1(n13893), .B2(n13980), .ZN(
        n13894) );
  NAND2_X1 U16078 ( .A1(n13895), .A2(n13894), .ZN(P3_U3475) );
  AOI21_X1 U16079 ( .B1(n13897), .B2(n16011), .A(n13896), .ZN(n13985) );
  MUX2_X1 U16080 ( .A(n13898), .B(n13985), .S(n13911), .Z(n13899) );
  OAI21_X1 U16081 ( .B1(n13900), .B2(n13989), .A(n13899), .ZN(P3_U3474) );
  MUX2_X1 U16082 ( .A(n13901), .B(n13990), .S(n13911), .Z(n13904) );
  NAND2_X1 U16083 ( .A1(n13993), .A2(n13902), .ZN(n13903) );
  OAI211_X1 U16084 ( .C1(n13905), .C2(n13996), .A(n13904), .B(n13903), .ZN(
        P3_U3473) );
  AOI21_X1 U16085 ( .B1(n13907), .B2(n16011), .A(n13906), .ZN(n13908) );
  OAI21_X1 U16086 ( .B1(n13910), .B2(n13909), .A(n13908), .ZN(n13998) );
  MUX2_X1 U16087 ( .A(P3_REG1_REG_9__SCAN_IN), .B(n13998), .S(n13911), .Z(
        P3_U3468) );
  NAND2_X1 U16088 ( .A1(n16018), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n13913) );
  NAND2_X1 U16089 ( .A1(n13912), .A2(n16017), .ZN(n13916) );
  OAI211_X1 U16090 ( .C1(n13914), .C2(n13997), .A(n13913), .B(n13916), .ZN(
        P3_U3458) );
  INV_X1 U16091 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n13918) );
  NAND2_X1 U16092 ( .A1(n13915), .A2(n13981), .ZN(n13917) );
  OAI211_X1 U16093 ( .C1(n13918), .C2(n16017), .A(n13917), .B(n13916), .ZN(
        P3_U3457) );
  INV_X1 U16094 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13920) );
  MUX2_X1 U16095 ( .A(n13920), .B(n13919), .S(n16017), .Z(n13924) );
  NAND2_X1 U16096 ( .A1(n13924), .A2(n13923), .ZN(P3_U3455) );
  INV_X1 U16097 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13926) );
  MUX2_X1 U16098 ( .A(n13926), .B(n13925), .S(n16017), .Z(n13930) );
  AOI22_X1 U16099 ( .A1(n13928), .A2(n13992), .B1(n13981), .B2(n13927), .ZN(
        n13929) );
  NAND2_X1 U16100 ( .A1(n13930), .A2(n13929), .ZN(P3_U3454) );
  INV_X1 U16101 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13932) );
  MUX2_X1 U16102 ( .A(n13932), .B(n13931), .S(n16017), .Z(n13933) );
  OAI21_X1 U16103 ( .B1(n6961), .B2(n13997), .A(n13933), .ZN(P3_U3453) );
  INV_X1 U16104 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13935) );
  MUX2_X1 U16105 ( .A(n13935), .B(n13934), .S(n16017), .Z(n13936) );
  OAI21_X1 U16106 ( .B1(n13937), .B2(n13997), .A(n13936), .ZN(P3_U3452) );
  INV_X1 U16107 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13939) );
  MUX2_X1 U16108 ( .A(n13939), .B(n13938), .S(n16017), .Z(n13940) );
  OAI21_X1 U16109 ( .B1(n13941), .B2(n13997), .A(n13940), .ZN(P3_U3451) );
  INV_X1 U16110 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13943) );
  MUX2_X1 U16111 ( .A(n13943), .B(n13942), .S(n16017), .Z(n13944) );
  OAI21_X1 U16112 ( .B1(n13945), .B2(n13997), .A(n13944), .ZN(P3_U3450) );
  INV_X1 U16113 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13947) );
  MUX2_X1 U16114 ( .A(n13947), .B(n13946), .S(n16017), .Z(n13951) );
  AOI22_X1 U16115 ( .A1(n13949), .A2(n13992), .B1(n13981), .B2(n13948), .ZN(
        n13950) );
  NAND2_X1 U16116 ( .A1(n13951), .A2(n13950), .ZN(P3_U3449) );
  INV_X1 U16117 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13953) );
  MUX2_X1 U16118 ( .A(n13953), .B(n13952), .S(n16017), .Z(n13954) );
  OAI21_X1 U16119 ( .B1(n13955), .B2(n13988), .A(n13954), .ZN(P3_U3448) );
  INV_X1 U16120 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13957) );
  MUX2_X1 U16121 ( .A(n13957), .B(n13956), .S(n16017), .Z(n13960) );
  NAND2_X1 U16122 ( .A1(n13958), .A2(n13981), .ZN(n13959) );
  OAI211_X1 U16123 ( .C1(n13961), .C2(n13988), .A(n13960), .B(n13959), .ZN(
        P3_U3447) );
  INV_X1 U16124 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13963) );
  MUX2_X1 U16125 ( .A(n13963), .B(n13962), .S(n16017), .Z(n13967) );
  AOI22_X1 U16126 ( .A1(n13965), .A2(n13992), .B1(n13981), .B2(n13964), .ZN(
        n13966) );
  NAND2_X1 U16127 ( .A1(n13967), .A2(n13966), .ZN(P3_U3446) );
  INV_X1 U16128 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13969) );
  MUX2_X1 U16129 ( .A(n13969), .B(n13968), .S(n16017), .Z(n13970) );
  OAI21_X1 U16130 ( .B1(n13971), .B2(n13997), .A(n13970), .ZN(P3_U3444) );
  INV_X1 U16131 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13973) );
  MUX2_X1 U16132 ( .A(n13973), .B(n13972), .S(n16017), .Z(n13977) );
  AOI22_X1 U16133 ( .A1(n13975), .A2(n13992), .B1(n13974), .B2(n13981), .ZN(
        n13976) );
  NAND2_X1 U16134 ( .A1(n13977), .A2(n13976), .ZN(P3_U3441) );
  INV_X1 U16135 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13979) );
  MUX2_X1 U16136 ( .A(n13979), .B(n13978), .S(n16017), .Z(n13984) );
  AOI22_X1 U16137 ( .A1(n13982), .A2(n13992), .B1(n13981), .B2(n13980), .ZN(
        n13983) );
  NAND2_X1 U16138 ( .A1(n13984), .A2(n13983), .ZN(P3_U3438) );
  INV_X1 U16139 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13986) );
  MUX2_X1 U16140 ( .A(n13986), .B(n13985), .S(n16017), .Z(n13987) );
  OAI21_X1 U16141 ( .B1(n13989), .B2(n13988), .A(n13987), .ZN(P3_U3435) );
  MUX2_X1 U16142 ( .A(n13991), .B(n13990), .S(n16017), .Z(n13995) );
  NAND2_X1 U16143 ( .A1(n13993), .A2(n13992), .ZN(n13994) );
  OAI211_X1 U16144 ( .C1(n13997), .C2(n13996), .A(n13995), .B(n13994), .ZN(
        P3_U3432) );
  MUX2_X1 U16145 ( .A(P3_REG0_REG_9__SCAN_IN), .B(n13998), .S(n16017), .Z(
        P3_U3417) );
  NAND2_X1 U16146 ( .A1(n14000), .A2(n13999), .ZN(n14004) );
  NAND4_X1 U16147 ( .A1(n8125), .A2(P3_STATE_REG_SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .A4(n14002), .ZN(n14003) );
  OAI211_X1 U16148 ( .C1(n14005), .C2(n14006), .A(n14004), .B(n14003), .ZN(
        P3_U3264) );
  OAI222_X1 U16149 ( .A1(n13257), .A2(n14009), .B1(n14008), .B2(P3_U3151), 
        .C1(n14007), .C2(n14006), .ZN(P3_U3266) );
  NOR3_X1 U16150 ( .A1(n14010), .A2(n14164), .A3(n14205), .ZN(n14011) );
  AOI21_X1 U16151 ( .B1(n14012), .B2(n14180), .A(n14011), .ZN(n14021) );
  INV_X1 U16152 ( .A(n14013), .ZN(n14020) );
  NAND2_X1 U16153 ( .A1(n14759), .A2(n14189), .ZN(n14016) );
  NAND2_X1 U16154 ( .A1(n14654), .A2(n14576), .ZN(n14014) );
  OAI21_X1 U16155 ( .B1(n14205), .B2(n14636), .A(n14014), .ZN(n14614) );
  AOI22_X1 U16156 ( .A1(n14170), .A2(n14614), .B1(P2_REG3_REG_14__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14015) );
  OAI211_X1 U16157 ( .C1(n14186), .C2(n14617), .A(n14016), .B(n14015), .ZN(
        n14017) );
  AOI21_X1 U16158 ( .B1(n14018), .B2(n14180), .A(n14017), .ZN(n14019) );
  OAI21_X1 U16159 ( .B1(n14021), .B2(n14020), .A(n14019), .ZN(P2_U3187) );
  AOI22_X1 U16160 ( .A1(n14023), .A2(n14180), .B1(n14179), .B2(n14199), .ZN(
        n14029) );
  INV_X1 U16161 ( .A(n14072), .ZN(n14028) );
  NOR2_X1 U16162 ( .A1(n14186), .A2(n14454), .ZN(n14026) );
  AOI22_X1 U16163 ( .A1(n14198), .A2(n14654), .B1(n14652), .B2(n14485), .ZN(
        n14448) );
  OAI22_X1 U16164 ( .A1(n14448), .A2(n14147), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14024), .ZN(n14025) );
  AOI211_X1 U16165 ( .C1(n14710), .C2(n14189), .A(n14026), .B(n14025), .ZN(
        n14027) );
  OAI21_X1 U16166 ( .B1(n14029), .B2(n14028), .A(n14027), .ZN(P2_U3188) );
  NAND2_X1 U16167 ( .A1(n14031), .A2(n14030), .ZN(n14033) );
  XOR2_X1 U16168 ( .A(n14033), .B(n14032), .Z(n14039) );
  INV_X1 U16169 ( .A(n14528), .ZN(n14036) );
  OAI22_X1 U16170 ( .A1(n14057), .A2(n14638), .B1(n14563), .B2(n14636), .ZN(
        n14524) );
  NOR2_X1 U16171 ( .A1(n14034), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14334) );
  AOI21_X1 U16172 ( .B1(n14170), .B2(n14524), .A(n14334), .ZN(n14035) );
  OAI21_X1 U16173 ( .B1(n14036), .B2(n14186), .A(n14035), .ZN(n14037) );
  AOI21_X1 U16174 ( .B1(n14732), .B2(n14189), .A(n14037), .ZN(n14038) );
  OAI21_X1 U16175 ( .B1(n14039), .B2(n14154), .A(n14038), .ZN(P2_U3191) );
  NAND2_X1 U16176 ( .A1(n14355), .A2(n14658), .ZN(n14040) );
  XNOR2_X1 U16177 ( .A(n14040), .B(n6546), .ZN(n14041) );
  XNOR2_X1 U16178 ( .A(n14369), .B(n14041), .ZN(n14043) );
  INV_X1 U16179 ( .A(n14043), .ZN(n14042) );
  INV_X1 U16180 ( .A(n14050), .ZN(n14053) );
  INV_X1 U16181 ( .A(n14049), .ZN(n14044) );
  INV_X1 U16182 ( .A(n14369), .ZN(n14346) );
  AOI22_X1 U16183 ( .A1(n14366), .A2(n14168), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14047) );
  NAND2_X1 U16184 ( .A1(n14045), .A2(n14170), .ZN(n14046) );
  OAI211_X1 U16185 ( .C1(n14346), .C2(n14173), .A(n14047), .B(n14046), .ZN(
        n14048) );
  AOI21_X1 U16186 ( .B1(n14050), .B2(n14049), .A(n14048), .ZN(n14051) );
  OAI211_X1 U16187 ( .C1(n14055), .C2(n14054), .A(n14129), .B(n14180), .ZN(
        n14061) );
  NOR2_X1 U16188 ( .A1(n14184), .A2(n14056), .ZN(n14059) );
  OAI22_X1 U16189 ( .A1(n14186), .A2(n14492), .B1(n14185), .B2(n14057), .ZN(
        n14058) );
  AOI211_X1 U16190 ( .C1(P2_REG3_REG_21__SCAN_IN), .C2(P2_U3088), .A(n14059), 
        .B(n14058), .ZN(n14060) );
  OAI211_X1 U16191 ( .C1(n14799), .C2(n14173), .A(n14061), .B(n14060), .ZN(
        P2_U3195) );
  NAND2_X1 U16192 ( .A1(n14063), .A2(n14062), .ZN(n14065) );
  XOR2_X1 U16193 ( .A(n14065), .B(n14064), .Z(n14070) );
  NAND2_X1 U16194 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n15898)
         );
  OAI21_X1 U16195 ( .B1(n14185), .B2(n14066), .A(n15898), .ZN(n14068) );
  OAI22_X1 U16196 ( .A1(n14186), .A2(n14660), .B1(n14184), .B2(n14205), .ZN(
        n14067) );
  AOI211_X1 U16197 ( .C1(n14769), .C2(n14189), .A(n14068), .B(n14067), .ZN(
        n14069) );
  OAI21_X1 U16198 ( .B1(n14070), .B2(n14154), .A(n14069), .ZN(P2_U3196) );
  NOR2_X1 U16199 ( .A1(n14075), .A2(n14074), .ZN(n14095) );
  NAND2_X1 U16200 ( .A1(n14096), .A2(n14095), .ZN(n14094) );
  AOI21_X1 U16201 ( .B1(n14094), .B2(n14076), .A(n14154), .ZN(n14080) );
  NOR3_X1 U16202 ( .A1(n14078), .A2(n14077), .A3(n14164), .ZN(n14079) );
  OAI21_X1 U16203 ( .B1(n14080), .B2(n14079), .A(n14163), .ZN(n14084) );
  AOI22_X1 U16204 ( .A1(n14196), .A2(n14654), .B1(n14652), .B2(n14198), .ZN(
        n14409) );
  OAI22_X1 U16205 ( .A1(n14409), .A2(n14147), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14081), .ZN(n14082) );
  AOI21_X1 U16206 ( .B1(n14413), .B2(n14168), .A(n14082), .ZN(n14083) );
  OAI211_X1 U16207 ( .C1(n14415), .C2(n14173), .A(n14084), .B(n14083), .ZN(
        P2_U3197) );
  AOI21_X1 U16208 ( .B1(n14087), .B2(n14086), .A(n14085), .ZN(n14093) );
  OAI21_X1 U16209 ( .B1(n14184), .B2(n14538), .A(n14088), .ZN(n14091) );
  OAI22_X1 U16210 ( .A1(n14572), .A2(n14186), .B1(n14185), .B2(n14089), .ZN(
        n14090) );
  AOI211_X1 U16211 ( .C1(n14580), .C2(n14189), .A(n14091), .B(n14090), .ZN(
        n14092) );
  OAI21_X1 U16212 ( .B1(n14093), .B2(n14154), .A(n14092), .ZN(P2_U3198) );
  OAI211_X1 U16213 ( .C1(n14096), .C2(n14095), .A(n14094), .B(n14180), .ZN(
        n14102) );
  INV_X1 U16214 ( .A(n14430), .ZN(n14100) );
  AND2_X1 U16215 ( .A1(n14199), .A2(n14652), .ZN(n14097) );
  AOI21_X1 U16216 ( .B1(n14197), .B2(n14654), .A(n14097), .ZN(n14424) );
  OAI22_X1 U16217 ( .A1(n14424), .A2(n14147), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14098), .ZN(n14099) );
  AOI21_X1 U16218 ( .B1(n14100), .B2(n14168), .A(n14099), .ZN(n14101) );
  OAI211_X1 U16219 ( .C1(n14103), .C2(n14173), .A(n14102), .B(n14101), .ZN(
        P2_U3201) );
  AND2_X1 U16220 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n14242) );
  OAI22_X1 U16221 ( .A1(n14186), .A2(n14105), .B1(n14184), .B2(n14104), .ZN(
        n14106) );
  AOI211_X1 U16222 ( .C1(n14107), .C2(n14189), .A(n14242), .B(n14106), .ZN(
        n14117) );
  OAI21_X1 U16223 ( .B1(n14111), .B2(n14109), .A(n14108), .ZN(n14110) );
  NAND2_X1 U16224 ( .A1(n14110), .A2(n14180), .ZN(n14116) );
  NOR3_X1 U16225 ( .A1(n14164), .A2(n14112), .A3(n14111), .ZN(n14114) );
  OAI21_X1 U16226 ( .B1(n14114), .B2(n14113), .A(n14214), .ZN(n14115) );
  NAND3_X1 U16227 ( .A1(n14117), .A2(n14116), .A3(n14115), .ZN(P2_U3202) );
  NAND2_X1 U16228 ( .A1(n14119), .A2(n14118), .ZN(n14121) );
  XOR2_X1 U16229 ( .A(n14121), .B(n14120), .Z(n14127) );
  OAI22_X1 U16230 ( .A1(n14185), .A2(n14539), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14122), .ZN(n14125) );
  INV_X1 U16231 ( .A(n14516), .ZN(n14123) );
  INV_X1 U16232 ( .A(n14200), .ZN(n14511) );
  OAI22_X1 U16233 ( .A1(n14123), .A2(n14186), .B1(n14184), .B2(n14511), .ZN(
        n14124) );
  AOI211_X1 U16234 ( .C1(n14515), .C2(n14189), .A(n14125), .B(n14124), .ZN(
        n14126) );
  OAI21_X1 U16235 ( .B1(n14127), .B2(n14154), .A(n14126), .ZN(P2_U3205) );
  NAND2_X1 U16236 ( .A1(n14129), .A2(n14128), .ZN(n14131) );
  XNOR2_X1 U16237 ( .A(n14131), .B(n14130), .ZN(n14133) );
  NAND3_X1 U16238 ( .A1(n14133), .A2(n14180), .A3(n14132), .ZN(n14140) );
  INV_X1 U16239 ( .A(n14133), .ZN(n14134) );
  NAND3_X1 U16240 ( .A1(n14134), .A2(n14179), .A3(n14485), .ZN(n14139) );
  AOI22_X1 U16241 ( .A1(n14199), .A2(n14654), .B1(n14652), .B2(n14200), .ZN(
        n14473) );
  OAI22_X1 U16242 ( .A1(n14147), .A2(n14473), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14135), .ZN(n14137) );
  NOR2_X1 U16243 ( .A1(n14716), .A2(n14173), .ZN(n14136) );
  AOI211_X1 U16244 ( .C1(n14168), .C2(n14475), .A(n14137), .B(n14136), .ZN(
        n14138) );
  NAND3_X1 U16245 ( .A1(n14140), .A2(n14139), .A3(n14138), .ZN(P2_U3207) );
  NAND2_X1 U16246 ( .A1(n14142), .A2(n14141), .ZN(n14144) );
  XOR2_X1 U16247 ( .A(n14144), .B(n14143), .Z(n14153) );
  OAI22_X1 U16248 ( .A1(n14147), .A2(n14146), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14145), .ZN(n14150) );
  NOR2_X1 U16249 ( .A1(n14186), .A2(n14148), .ZN(n14149) );
  AOI211_X1 U16250 ( .C1(n14151), .C2(n14189), .A(n14150), .B(n14149), .ZN(
        n14152) );
  OAI21_X1 U16251 ( .B1(n14153), .B2(n14154), .A(n14152), .ZN(P2_U3208) );
  AOI21_X1 U16252 ( .B1(n14156), .B2(n14155), .A(n14154), .ZN(n14158) );
  NAND2_X1 U16253 ( .A1(n14158), .A2(n14157), .ZN(n14162) );
  AND2_X1 U16254 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14308) );
  OAI22_X1 U16255 ( .A1(n14549), .A2(n14186), .B1(n14185), .B2(n14538), .ZN(
        n14159) );
  AOI211_X1 U16256 ( .C1(n14160), .C2(n14201), .A(n14308), .B(n14159), .ZN(
        n14161) );
  OAI211_X1 U16257 ( .C1(n14552), .C2(n14173), .A(n14162), .B(n14161), .ZN(
        P2_U3210) );
  NOR3_X1 U16258 ( .A1(n14165), .A2(n14169), .A3(n14164), .ZN(n14166) );
  AOI21_X1 U16259 ( .B1(n12808), .B2(n14180), .A(n14166), .ZN(n14178) );
  INV_X1 U16260 ( .A(n14167), .ZN(n14399) );
  AOI22_X1 U16261 ( .A1(n14168), .A2(n14399), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14172) );
  OAI22_X1 U16262 ( .A1(n7884), .A2(n14638), .B1(n14169), .B2(n14636), .ZN(
        n14393) );
  NAND2_X1 U16263 ( .A1(n14393), .A2(n14170), .ZN(n14171) );
  OAI211_X1 U16264 ( .C1(n14401), .C2(n14173), .A(n14172), .B(n14171), .ZN(
        n14174) );
  AOI21_X1 U16265 ( .B1(n14175), .B2(n14180), .A(n14174), .ZN(n14176) );
  OAI21_X1 U16266 ( .B1(n14178), .B2(n14177), .A(n14176), .ZN(P2_U3212) );
  AOI22_X1 U16267 ( .A1(n14181), .A2(n14180), .B1(n14179), .B2(n14576), .ZN(
        n14192) );
  INV_X1 U16268 ( .A(n14182), .ZN(n14191) );
  OAI22_X1 U16269 ( .A1(n14184), .A2(n14594), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14183), .ZN(n14188) );
  OAI22_X1 U16270 ( .A1(n14602), .A2(n14186), .B1(n14185), .B2(n14637), .ZN(
        n14187) );
  AOI211_X1 U16271 ( .C1(n14754), .C2(n14189), .A(n14188), .B(n14187), .ZN(
        n14190) );
  OAI21_X1 U16272 ( .B1(n14192), .B2(n14191), .A(n14190), .ZN(P2_U3213) );
  MUX2_X1 U16273 ( .A(n14193), .B(P2_DATAO_REG_31__SCAN_IN), .S(n14217), .Z(
        P2_U3562) );
  MUX2_X1 U16274 ( .A(n14351), .B(P2_DATAO_REG_30__SCAN_IN), .S(n14217), .Z(
        P2_U3561) );
  MUX2_X1 U16275 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n14194), .S(P2_U3947), .Z(
        P2_U3560) );
  MUX2_X1 U16276 ( .A(n14355), .B(P2_DATAO_REG_28__SCAN_IN), .S(n14217), .Z(
        P2_U3559) );
  MUX2_X1 U16277 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n14195), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U16278 ( .A(n14196), .B(P2_DATAO_REG_26__SCAN_IN), .S(n14217), .Z(
        P2_U3557) );
  MUX2_X1 U16279 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n14197), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U16280 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n14198), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U16281 ( .A(n14199), .B(P2_DATAO_REG_23__SCAN_IN), .S(n14217), .Z(
        P2_U3554) );
  MUX2_X1 U16282 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n14485), .S(P2_U3947), .Z(
        P2_U3553) );
  MUX2_X1 U16283 ( .A(n14200), .B(P2_DATAO_REG_21__SCAN_IN), .S(n14217), .Z(
        P2_U3552) );
  MUX2_X1 U16284 ( .A(n14484), .B(P2_DATAO_REG_20__SCAN_IN), .S(n14217), .Z(
        P2_U3551) );
  MUX2_X1 U16285 ( .A(n14201), .B(P2_DATAO_REG_19__SCAN_IN), .S(n14217), .Z(
        P2_U3550) );
  MUX2_X1 U16286 ( .A(n14202), .B(P2_DATAO_REG_18__SCAN_IN), .S(n14217), .Z(
        P2_U3549) );
  MUX2_X1 U16287 ( .A(n14575), .B(P2_DATAO_REG_17__SCAN_IN), .S(n14217), .Z(
        P2_U3548) );
  MUX2_X1 U16288 ( .A(n14203), .B(P2_DATAO_REG_16__SCAN_IN), .S(n14217), .Z(
        P2_U3547) );
  MUX2_X1 U16289 ( .A(n14576), .B(P2_DATAO_REG_15__SCAN_IN), .S(n14217), .Z(
        P2_U3546) );
  MUX2_X1 U16290 ( .A(n14204), .B(P2_DATAO_REG_14__SCAN_IN), .S(n14217), .Z(
        P2_U3545) );
  INV_X1 U16291 ( .A(n14205), .ZN(n14655) );
  MUX2_X1 U16292 ( .A(n14655), .B(P2_DATAO_REG_13__SCAN_IN), .S(n14217), .Z(
        P2_U3544) );
  MUX2_X1 U16293 ( .A(n14206), .B(P2_DATAO_REG_12__SCAN_IN), .S(n14217), .Z(
        P2_U3543) );
  MUX2_X1 U16294 ( .A(n14653), .B(P2_DATAO_REG_11__SCAN_IN), .S(n14217), .Z(
        P2_U3542) );
  MUX2_X1 U16295 ( .A(n14207), .B(P2_DATAO_REG_10__SCAN_IN), .S(n14217), .Z(
        P2_U3541) );
  MUX2_X1 U16296 ( .A(n14208), .B(P2_DATAO_REG_9__SCAN_IN), .S(n14217), .Z(
        P2_U3540) );
  MUX2_X1 U16297 ( .A(n14209), .B(P2_DATAO_REG_8__SCAN_IN), .S(n14217), .Z(
        P2_U3539) );
  MUX2_X1 U16298 ( .A(n14210), .B(P2_DATAO_REG_7__SCAN_IN), .S(n14217), .Z(
        P2_U3538) );
  MUX2_X1 U16299 ( .A(n14211), .B(P2_DATAO_REG_6__SCAN_IN), .S(n14217), .Z(
        P2_U3537) );
  MUX2_X1 U16300 ( .A(n14212), .B(P2_DATAO_REG_5__SCAN_IN), .S(n14217), .Z(
        P2_U3536) );
  MUX2_X1 U16301 ( .A(n14213), .B(P2_DATAO_REG_4__SCAN_IN), .S(n14217), .Z(
        P2_U3535) );
  MUX2_X1 U16302 ( .A(n14214), .B(P2_DATAO_REG_3__SCAN_IN), .S(n14217), .Z(
        P2_U3534) );
  MUX2_X1 U16303 ( .A(n14215), .B(P2_DATAO_REG_2__SCAN_IN), .S(n14217), .Z(
        P2_U3533) );
  MUX2_X1 U16304 ( .A(n14216), .B(P2_DATAO_REG_1__SCAN_IN), .S(n14217), .Z(
        P2_U3532) );
  MUX2_X1 U16305 ( .A(n10168), .B(P2_DATAO_REG_0__SCAN_IN), .S(n14217), .Z(
        P2_U3531) );
  NOR2_X1 U16306 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7530), .ZN(n14219) );
  NOR2_X1 U16307 ( .A1(n14306), .A2(n14220), .ZN(n14218) );
  AOI211_X1 U16308 ( .C1(n15851), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n14219), .B(
        n14218), .ZN(n14230) );
  MUX2_X1 U16309 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n11029), .S(n14220), .Z(
        n14221) );
  OAI21_X1 U16310 ( .B1(n12668), .B2(n14222), .A(n14221), .ZN(n14223) );
  NAND3_X1 U16311 ( .A1(n15892), .A2(n14224), .A3(n14223), .ZN(n14229) );
  OAI211_X1 U16312 ( .C1(n14227), .C2(n14226), .A(n15896), .B(n14225), .ZN(
        n14228) );
  NAND3_X1 U16313 ( .A1(n14230), .A2(n14229), .A3(n14228), .ZN(P2_U3215) );
  AOI22_X1 U16314 ( .A1(n15894), .A2(n14231), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(P2_U3088), .ZN(n14241) );
  NAND2_X1 U16315 ( .A1(n15851), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n14240) );
  OAI211_X1 U16316 ( .C1(n14234), .C2(n14233), .A(n15896), .B(n14232), .ZN(
        n14239) );
  OAI211_X1 U16317 ( .C1(n14237), .C2(n14236), .A(n15892), .B(n14235), .ZN(
        n14238) );
  NAND4_X1 U16318 ( .A1(n14241), .A2(n14240), .A3(n14239), .A4(n14238), .ZN(
        P2_U3216) );
  NAND2_X1 U16319 ( .A1(n15851), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n14254) );
  AOI21_X1 U16320 ( .B1(n15894), .B2(n14246), .A(n14242), .ZN(n14253) );
  OAI211_X1 U16321 ( .C1(n14245), .C2(n14244), .A(n15896), .B(n14243), .ZN(
        n14252) );
  MUX2_X1 U16322 ( .A(n11995), .B(P2_REG2_REG_4__SCAN_IN), .S(n14246), .Z(
        n14247) );
  NAND3_X1 U16323 ( .A1(n15861), .A2(n14248), .A3(n14247), .ZN(n14249) );
  NAND3_X1 U16324 ( .A1(n15892), .A2(n14250), .A3(n14249), .ZN(n14251) );
  NAND4_X1 U16325 ( .A1(n14254), .A2(n14253), .A3(n14252), .A4(n14251), .ZN(
        P2_U3218) );
  NAND2_X1 U16326 ( .A1(n15851), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14267) );
  INV_X1 U16327 ( .A(n14255), .ZN(n14256) );
  AOI21_X1 U16328 ( .B1(n15894), .B2(n14260), .A(n14256), .ZN(n14266) );
  OAI211_X1 U16329 ( .C1(n14259), .C2(n14258), .A(n15896), .B(n14257), .ZN(
        n14265) );
  MUX2_X1 U16330 ( .A(n11976), .B(P2_REG2_REG_6__SCAN_IN), .S(n14260), .Z(
        n14261) );
  NAND3_X1 U16331 ( .A1(n15875), .A2(n14262), .A3(n14261), .ZN(n14263) );
  NAND3_X1 U16332 ( .A1(n15892), .A2(n14275), .A3(n14263), .ZN(n14264) );
  NAND4_X1 U16333 ( .A1(n14267), .A2(n14266), .A3(n14265), .A4(n14264), .ZN(
        P2_U3220) );
  NAND2_X1 U16334 ( .A1(n15851), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n14281) );
  AND2_X1 U16335 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n14268) );
  AOI21_X1 U16336 ( .B1(n15894), .B2(n14272), .A(n14268), .ZN(n14280) );
  OAI211_X1 U16337 ( .C1(n14271), .C2(n14270), .A(n15896), .B(n14269), .ZN(
        n14279) );
  MUX2_X1 U16338 ( .A(n12129), .B(P2_REG2_REG_7__SCAN_IN), .S(n14272), .Z(
        n14273) );
  NAND3_X1 U16339 ( .A1(n14275), .A2(n14274), .A3(n14273), .ZN(n14276) );
  NAND3_X1 U16340 ( .A1(n15892), .A2(n14277), .A3(n14276), .ZN(n14278) );
  NAND4_X1 U16341 ( .A1(n14281), .A2(n14280), .A3(n14279), .A4(n14278), .ZN(
        P2_U3221) );
  NAND2_X1 U16342 ( .A1(n14283), .A2(n14282), .ZN(n14285) );
  NAND2_X1 U16343 ( .A1(n14291), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n14284) );
  NAND2_X1 U16344 ( .A1(n14285), .A2(n14284), .ZN(n14287) );
  MUX2_X1 U16345 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n9959), .S(n14309), .Z(
        n14286) );
  NAND2_X1 U16346 ( .A1(n14287), .A2(n14286), .ZN(n14300) );
  OAI211_X1 U16347 ( .C1(n14287), .C2(n14286), .A(n14300), .B(n15892), .ZN(
        n14298) );
  OAI21_X1 U16348 ( .B1(n14306), .B2(n14289), .A(n14288), .ZN(n14290) );
  AOI21_X1 U16349 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(n15851), .A(n14290), 
        .ZN(n14297) );
  NAND2_X1 U16350 ( .A1(n14291), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n14292) );
  NAND2_X1 U16351 ( .A1(n14293), .A2(n14292), .ZN(n14295) );
  INV_X1 U16352 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n14745) );
  XNOR2_X1 U16353 ( .A(n14309), .B(n14745), .ZN(n14294) );
  NAND2_X1 U16354 ( .A1(n14295), .A2(n14294), .ZN(n14311) );
  OAI211_X1 U16355 ( .C1(n14295), .C2(n14294), .A(n14311), .B(n15896), .ZN(
        n14296) );
  NAND3_X1 U16356 ( .A1(n14298), .A2(n14297), .A3(n14296), .ZN(P2_U3231) );
  NAND2_X1 U16357 ( .A1(n14309), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n14299) );
  NAND2_X1 U16358 ( .A1(n14300), .A2(n14299), .ZN(n14301) );
  NAND2_X1 U16359 ( .A1(n14301), .A2(n14312), .ZN(n14302) );
  INV_X1 U16360 ( .A(n14321), .ZN(n14303) );
  AOI21_X1 U16361 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n14304), .A(n14303), 
        .ZN(n14320) );
  NOR2_X1 U16362 ( .A1(n14306), .A2(n14305), .ZN(n14307) );
  AOI211_X1 U16363 ( .C1(n15851), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n14308), 
        .B(n14307), .ZN(n14319) );
  NAND2_X1 U16364 ( .A1(n14309), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n14310) );
  NAND2_X1 U16365 ( .A1(n14311), .A2(n14310), .ZN(n14313) );
  NAND2_X1 U16366 ( .A1(n14313), .A2(n14312), .ZN(n14324) );
  OR2_X1 U16367 ( .A1(n14313), .A2(n14312), .ZN(n14314) );
  NAND2_X1 U16368 ( .A1(n14324), .A2(n14314), .ZN(n14316) );
  INV_X1 U16369 ( .A(n14316), .ZN(n14317) );
  INV_X1 U16370 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n14315) );
  OR2_X1 U16371 ( .A1(n14316), .A2(n14315), .ZN(n14325) );
  OAI211_X1 U16372 ( .C1(n14317), .C2(P2_REG1_REG_18__SCAN_IN), .A(n15896), 
        .B(n14325), .ZN(n14318) );
  OAI211_X1 U16373 ( .C1(n14320), .C2(n14330), .A(n14319), .B(n14318), .ZN(
        P2_U3232) );
  INV_X1 U16374 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n14322) );
  XNOR2_X1 U16375 ( .A(n14323), .B(n14322), .ZN(n14331) );
  INV_X1 U16376 ( .A(n14331), .ZN(n14328) );
  NAND2_X1 U16377 ( .A1(n14325), .A2(n14324), .ZN(n14326) );
  XNOR2_X1 U16378 ( .A(n14326), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n14329) );
  AOI21_X1 U16379 ( .B1(n14329), .B2(n15896), .A(n15894), .ZN(n14327) );
  OAI21_X1 U16380 ( .B1(n14328), .B2(n14330), .A(n14327), .ZN(n14333) );
  XNOR2_X1 U16381 ( .A(n14335), .B(n14788), .ZN(n14336) );
  NAND2_X1 U16382 ( .A1(n14676), .A2(n14672), .ZN(n14339) );
  NOR2_X1 U16383 ( .A1(n14674), .A2(n14337), .ZN(n14340) );
  AOI21_X1 U16384 ( .B1(n14674), .B2(P2_REG2_REG_31__SCAN_IN), .A(n14340), 
        .ZN(n14338) );
  OAI211_X1 U16385 ( .C1(n14788), .C2(n14664), .A(n14339), .B(n14338), .ZN(
        P2_U3234) );
  AOI21_X1 U16386 ( .B1(n14674), .B2(P2_REG2_REG_30__SCAN_IN), .A(n14340), 
        .ZN(n14342) );
  NAND2_X1 U16387 ( .A1(n14681), .A2(n14433), .ZN(n14341) );
  OAI211_X1 U16388 ( .C1(n14343), .C2(n14360), .A(n14342), .B(n14341), .ZN(
        P2_U3235) );
  INV_X1 U16389 ( .A(n14351), .ZN(n14353) );
  NOR3_X1 U16390 ( .A1(n14638), .A2(n14353), .A3(n14352), .ZN(n14354) );
  AOI21_X1 U16391 ( .B1(n14355), .B2(n14652), .A(n14354), .ZN(n14356) );
  OAI211_X1 U16392 ( .C1(n14686), .C2(n14359), .A(n10450), .B(n14358), .ZN(
        n14685) );
  NOR2_X1 U16393 ( .A1(n14685), .A2(n14360), .ZN(n14364) );
  AOI22_X1 U16394 ( .A1(n14674), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n14361), 
        .B2(n14661), .ZN(n14362) );
  OAI21_X1 U16395 ( .B1(n14686), .B2(n14664), .A(n14362), .ZN(n14363) );
  AOI211_X1 U16396 ( .C1(n14688), .C2(n14645), .A(n14364), .B(n14363), .ZN(
        n14365) );
  OAI21_X1 U16397 ( .B1(n14684), .B2(n14669), .A(n14365), .ZN(P2_U3236) );
  INV_X1 U16398 ( .A(n14366), .ZN(n14368) );
  OAI21_X1 U16399 ( .B1(n14368), .B2(n14642), .A(n14367), .ZN(n14375) );
  AOI22_X1 U16400 ( .A1(n14369), .A2(n14433), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n14674), .ZN(n14372) );
  NAND2_X1 U16401 ( .A1(n14370), .A2(n14672), .ZN(n14371) );
  OAI211_X1 U16402 ( .C1(n14373), .C2(n14669), .A(n14372), .B(n14371), .ZN(
        n14374) );
  AOI21_X1 U16403 ( .B1(n14375), .B2(n14645), .A(n14374), .ZN(n14376) );
  INV_X1 U16404 ( .A(n14376), .ZN(P2_U3237) );
  XNOR2_X1 U16405 ( .A(n14377), .B(n14381), .ZN(n14379) );
  OAI21_X1 U16406 ( .B1(n14382), .B2(n14381), .A(n14380), .ZN(n14693) );
  INV_X1 U16407 ( .A(n14693), .ZN(n14389) );
  AOI21_X1 U16408 ( .B1(n14396), .B2(n14690), .A(n14658), .ZN(n14384) );
  NAND2_X1 U16409 ( .A1(n14689), .A2(n14672), .ZN(n14387) );
  AOI22_X1 U16410 ( .A1(n14674), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n14385), 
        .B2(n14661), .ZN(n14386) );
  OAI211_X1 U16411 ( .C1(n7622), .C2(n14664), .A(n14387), .B(n14386), .ZN(
        n14388) );
  AOI21_X1 U16412 ( .B1(n14389), .B2(n14588), .A(n14388), .ZN(n14390) );
  OAI21_X1 U16413 ( .B1(n14692), .B2(n14674), .A(n14390), .ZN(P2_U3238) );
  XNOR2_X1 U16414 ( .A(n14391), .B(n14392), .ZN(n14394) );
  INV_X1 U16415 ( .A(n14395), .ZN(n14398) );
  INV_X1 U16416 ( .A(n14396), .ZN(n14397) );
  AOI211_X1 U16417 ( .C1(n14695), .C2(n14398), .A(n14658), .B(n14397), .ZN(
        n14694) );
  AOI22_X1 U16418 ( .A1(n14674), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n14399), 
        .B2(n14661), .ZN(n14400) );
  OAI21_X1 U16419 ( .B1(n14401), .B2(n14664), .A(n14400), .ZN(n14406) );
  OAI21_X1 U16420 ( .B1(n14404), .B2(n14403), .A(n14402), .ZN(n14698) );
  NOR2_X1 U16421 ( .A1(n14698), .A2(n14669), .ZN(n14405) );
  AOI211_X1 U16422 ( .C1(n14694), .C2(n14672), .A(n14406), .B(n14405), .ZN(
        n14407) );
  OAI21_X1 U16423 ( .B1(n14674), .B2(n14697), .A(n14407), .ZN(P2_U3239) );
  XNOR2_X1 U16424 ( .A(n14408), .B(n14417), .ZN(n14411) );
  INV_X1 U16425 ( .A(n14409), .ZN(n14410) );
  AOI21_X1 U16426 ( .B1(n14411), .B2(n14657), .A(n14410), .ZN(n14702) );
  INV_X1 U16427 ( .A(n14436), .ZN(n14412) );
  AOI211_X1 U16428 ( .C1(n14700), .C2(n14412), .A(n14658), .B(n14395), .ZN(
        n14699) );
  AOI22_X1 U16429 ( .A1(n14674), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n14413), 
        .B2(n14661), .ZN(n14414) );
  OAI21_X1 U16430 ( .B1(n14415), .B2(n14664), .A(n14414), .ZN(n14420) );
  OAI21_X1 U16431 ( .B1(n14418), .B2(n14417), .A(n14416), .ZN(n14703) );
  NOR2_X1 U16432 ( .A1(n14703), .A2(n14669), .ZN(n14419) );
  AOI211_X1 U16433 ( .C1(n14699), .C2(n14672), .A(n14420), .B(n14419), .ZN(
        n14421) );
  OAI21_X1 U16434 ( .B1(n14674), .B2(n14702), .A(n14421), .ZN(P2_U3240) );
  XNOR2_X1 U16435 ( .A(n14422), .B(n14423), .ZN(n14426) );
  INV_X1 U16436 ( .A(n14424), .ZN(n14425) );
  AOI21_X1 U16437 ( .B1(n14426), .B2(n14657), .A(n14425), .ZN(n14707) );
  OAI21_X1 U16438 ( .B1(n14429), .B2(n14428), .A(n14427), .ZN(n14708) );
  OAI22_X1 U16439 ( .A1(n14645), .A2(n14431), .B1(n14430), .B2(n14642), .ZN(
        n14432) );
  AOI21_X1 U16440 ( .B1(n14705), .B2(n14433), .A(n14432), .ZN(n14438) );
  NAND2_X1 U16441 ( .A1(n14452), .A2(n14705), .ZN(n14434) );
  NAND2_X1 U16442 ( .A1(n14434), .A2(n10450), .ZN(n14435) );
  NOR2_X1 U16443 ( .A1(n14436), .A2(n14435), .ZN(n14704) );
  NAND2_X1 U16444 ( .A1(n14704), .A2(n14672), .ZN(n14437) );
  OAI211_X1 U16445 ( .C1(n14708), .C2(n14669), .A(n14438), .B(n14437), .ZN(
        n14439) );
  INV_X1 U16446 ( .A(n14439), .ZN(n14440) );
  OAI21_X1 U16447 ( .B1(n14707), .B2(n14674), .A(n14440), .ZN(P2_U3241) );
  OAI21_X1 U16448 ( .B1(n14441), .B2(n14443), .A(n14442), .ZN(n14445) );
  NAND2_X1 U16449 ( .A1(n14445), .A2(n9843), .ZN(n14447) );
  XNOR2_X1 U16450 ( .A(n14447), .B(n14446), .ZN(n14450) );
  INV_X1 U16451 ( .A(n14448), .ZN(n14449) );
  AOI21_X1 U16452 ( .B1(n14450), .B2(n14657), .A(n14449), .ZN(n14712) );
  INV_X1 U16453 ( .A(n14452), .ZN(n14453) );
  AOI211_X1 U16454 ( .C1(n14710), .C2(n14451), .A(n14658), .B(n14453), .ZN(
        n14709) );
  INV_X1 U16455 ( .A(n14454), .ZN(n14455) );
  AOI22_X1 U16456 ( .A1(n14674), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n14455), 
        .B2(n14661), .ZN(n14456) );
  OAI21_X1 U16457 ( .B1(n14457), .B2(n14664), .A(n14456), .ZN(n14462) );
  OAI21_X1 U16458 ( .B1(n14460), .B2(n14459), .A(n14458), .ZN(n14713) );
  NOR2_X1 U16459 ( .A1(n14713), .A2(n14669), .ZN(n14461) );
  AOI211_X1 U16460 ( .C1(n14709), .C2(n14672), .A(n14462), .B(n14461), .ZN(
        n14463) );
  OAI21_X1 U16461 ( .B1(n14674), .B2(n14712), .A(n14463), .ZN(P2_U3242) );
  NAND2_X1 U16462 ( .A1(n14465), .A2(n14464), .ZN(n14466) );
  NAND2_X1 U16463 ( .A1(n14467), .A2(n14466), .ZN(n14714) );
  INV_X1 U16464 ( .A(n14508), .ZN(n14498) );
  NAND2_X1 U16465 ( .A1(n14441), .A2(n14498), .ZN(n14509) );
  NAND2_X1 U16466 ( .A1(n14509), .A2(n14468), .ZN(n14481) );
  INV_X1 U16467 ( .A(n14488), .ZN(n14469) );
  OAI21_X1 U16468 ( .B1(n14511), .B2(n14491), .A(n14482), .ZN(n14471) );
  XNOR2_X1 U16469 ( .A(n14471), .B(n14470), .ZN(n14472) );
  NAND2_X1 U16470 ( .A1(n14472), .A2(n14657), .ZN(n14474) );
  NAND2_X1 U16471 ( .A1(n14474), .A2(n14473), .ZN(n14719) );
  NAND2_X1 U16472 ( .A1(n14719), .A2(n14645), .ZN(n14480) );
  OAI211_X1 U16473 ( .C1(n14490), .C2(n14716), .A(n10450), .B(n14451), .ZN(
        n14715) );
  INV_X1 U16474 ( .A(n14715), .ZN(n14478) );
  AOI22_X1 U16475 ( .A1(n14674), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n14475), 
        .B2(n14661), .ZN(n14476) );
  OAI21_X1 U16476 ( .B1(n14716), .B2(n14664), .A(n14476), .ZN(n14477) );
  AOI21_X1 U16477 ( .B1(n14478), .B2(n14672), .A(n14477), .ZN(n14479) );
  OAI211_X1 U16478 ( .C1(n14669), .C2(n14714), .A(n14480), .B(n14479), .ZN(
        P2_U3243) );
  INV_X1 U16479 ( .A(n14481), .ZN(n14483) );
  OAI211_X1 U16480 ( .C1(n14483), .C2(n14488), .A(n14657), .B(n14482), .ZN(
        n14487) );
  AOI22_X1 U16481 ( .A1(n14485), .A2(n14654), .B1(n14652), .B2(n14484), .ZN(
        n14486) );
  NAND2_X1 U16482 ( .A1(n14487), .A2(n14486), .ZN(n14720) );
  INV_X1 U16483 ( .A(n14720), .ZN(n14497) );
  NAND2_X1 U16484 ( .A1(n14501), .A2(n6750), .ZN(n14489) );
  XNOR2_X1 U16485 ( .A(n14489), .B(n14488), .ZN(n14722) );
  AOI211_X1 U16486 ( .C1(n14491), .C2(n14513), .A(n14658), .B(n14490), .ZN(
        n14721) );
  NAND2_X1 U16487 ( .A1(n14721), .A2(n14672), .ZN(n14494) );
  AOI22_X1 U16488 ( .A1(n14674), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n6858), 
        .B2(n14661), .ZN(n14493) );
  OAI211_X1 U16489 ( .C1(n14799), .C2(n14664), .A(n14494), .B(n14493), .ZN(
        n14495) );
  AOI21_X1 U16490 ( .B1(n14722), .B2(n14588), .A(n14495), .ZN(n14496) );
  OAI21_X1 U16491 ( .B1(n14497), .B2(n14674), .A(n14496), .ZN(P2_U3244) );
  NAND2_X1 U16492 ( .A1(n14499), .A2(n14498), .ZN(n14500) );
  NAND2_X1 U16493 ( .A1(n14501), .A2(n14500), .ZN(n14725) );
  INV_X1 U16494 ( .A(n14541), .ZN(n14504) );
  INV_X1 U16495 ( .A(n14505), .ZN(n14506) );
  OAI222_X1 U16496 ( .A1(n14636), .A2(n14539), .B1(n14638), .B2(n14511), .C1(
        n14634), .C2(n14510), .ZN(n14726) );
  NAND2_X1 U16497 ( .A1(n14726), .A2(n14645), .ZN(n14520) );
  INV_X1 U16498 ( .A(n14513), .ZN(n14514) );
  AOI211_X1 U16499 ( .C1(n14515), .C2(n14512), .A(n14658), .B(n14514), .ZN(
        n14727) );
  AOI22_X1 U16500 ( .A1(n14674), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14516), 
        .B2(n14661), .ZN(n14517) );
  OAI21_X1 U16501 ( .B1(n14803), .B2(n14664), .A(n14517), .ZN(n14518) );
  AOI21_X1 U16502 ( .B1(n14727), .B2(n14672), .A(n14518), .ZN(n14519) );
  OAI211_X1 U16503 ( .C1(n14669), .C2(n14725), .A(n14520), .B(n14519), .ZN(
        P2_U3245) );
  OAI21_X1 U16504 ( .B1(n14523), .B2(n14522), .A(n14521), .ZN(n14525) );
  AOI21_X1 U16505 ( .B1(n14525), .B2(n14657), .A(n14524), .ZN(n14734) );
  INV_X1 U16506 ( .A(n14548), .ZN(n14527) );
  INV_X1 U16507 ( .A(n14512), .ZN(n14526) );
  AOI211_X1 U16508 ( .C1(n14732), .C2(n14527), .A(n14658), .B(n14526), .ZN(
        n14731) );
  AOI22_X1 U16509 ( .A1(n14674), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n14528), 
        .B2(n14661), .ZN(n14529) );
  OAI21_X1 U16510 ( .B1(n14530), .B2(n14664), .A(n14529), .ZN(n14535) );
  OAI21_X1 U16511 ( .B1(n14533), .B2(n14532), .A(n14531), .ZN(n14735) );
  NOR2_X1 U16512 ( .A1(n14735), .A2(n14669), .ZN(n14534) );
  AOI211_X1 U16513 ( .C1(n14731), .C2(n14672), .A(n14535), .B(n14534), .ZN(
        n14536) );
  OAI21_X1 U16514 ( .B1(n14734), .B2(n14674), .A(n14536), .ZN(P2_U3246) );
  XNOR2_X1 U16515 ( .A(n14537), .B(n14540), .ZN(n14553) );
  OAI22_X1 U16516 ( .A1(n14539), .A2(n14638), .B1(n14538), .B2(n14636), .ZN(
        n14546) );
  INV_X1 U16517 ( .A(n14560), .ZN(n14542) );
  AOI21_X1 U16518 ( .B1(n14542), .B2(n14541), .A(n14540), .ZN(n14543) );
  NOR3_X1 U16519 ( .A1(n14544), .A2(n14543), .A3(n14634), .ZN(n14545) );
  AOI211_X1 U16520 ( .C1(n14547), .C2(n14553), .A(n14546), .B(n14545), .ZN(
        n14739) );
  AOI211_X1 U16521 ( .C1(n14737), .C2(n14564), .A(n14658), .B(n14548), .ZN(
        n14736) );
  INV_X1 U16522 ( .A(n14549), .ZN(n14550) );
  AOI22_X1 U16523 ( .A1(n14674), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n14550), 
        .B2(n14661), .ZN(n14551) );
  OAI21_X1 U16524 ( .B1(n14552), .B2(n14664), .A(n14551), .ZN(n14556) );
  INV_X1 U16525 ( .A(n14553), .ZN(n14740) );
  NOR2_X1 U16526 ( .A1(n14740), .A2(n14554), .ZN(n14555) );
  AOI211_X1 U16527 ( .C1(n14736), .C2(n14672), .A(n14556), .B(n14555), .ZN(
        n14557) );
  OAI21_X1 U16528 ( .B1(n14739), .B2(n14674), .A(n14557), .ZN(P2_U3247) );
  OAI21_X1 U16529 ( .B1(n14559), .B2(n14561), .A(n14558), .ZN(n14741) );
  OAI222_X1 U16530 ( .A1(n14638), .A2(n14563), .B1(n14636), .B2(n14594), .C1(
        n14634), .C2(n14562), .ZN(n14742) );
  NAND2_X1 U16531 ( .A1(n14742), .A2(n14645), .ZN(n14571) );
  INV_X1 U16532 ( .A(n14564), .ZN(n14565) );
  AOI211_X1 U16533 ( .C1(n14566), .C2(n14581), .A(n14658), .B(n14565), .ZN(
        n14743) );
  NOR2_X1 U16534 ( .A1(n14809), .A2(n14664), .ZN(n14569) );
  OAI22_X1 U16535 ( .A1(n14645), .A2(n9959), .B1(n14567), .B2(n14642), .ZN(
        n14568) );
  AOI211_X1 U16536 ( .C1(n14743), .C2(n14672), .A(n14569), .B(n14568), .ZN(
        n14570) );
  OAI211_X1 U16537 ( .C1(n14669), .C2(n14741), .A(n14571), .B(n14570), .ZN(
        P2_U3248) );
  INV_X1 U16538 ( .A(n14572), .ZN(n14579) );
  XNOR2_X1 U16539 ( .A(n14573), .B(n9705), .ZN(n14574) );
  NAND2_X1 U16540 ( .A1(n14574), .A2(n14657), .ZN(n14578) );
  AOI22_X1 U16541 ( .A1(n14652), .A2(n14576), .B1(n14654), .B2(n14575), .ZN(
        n14577) );
  NAND2_X1 U16542 ( .A1(n14578), .A2(n14577), .ZN(n14752) );
  AOI21_X1 U16543 ( .B1(n14579), .B2(n14661), .A(n14752), .ZN(n14591) );
  AOI21_X1 U16544 ( .B1(n14599), .B2(n14580), .A(n14658), .ZN(n14582) );
  NAND2_X1 U16545 ( .A1(n14582), .A2(n14581), .ZN(n14749) );
  INV_X1 U16546 ( .A(n14749), .ZN(n14585) );
  OAI22_X1 U16547 ( .A1(n7627), .A2(n14664), .B1(n14645), .B2(n14583), .ZN(
        n14584) );
  AOI21_X1 U16548 ( .B1(n14585), .B2(n14672), .A(n14584), .ZN(n14590) );
  NAND2_X1 U16549 ( .A1(n14587), .A2(n14586), .ZN(n14747) );
  NAND3_X1 U16550 ( .A1(n14748), .A2(n14747), .A3(n14588), .ZN(n14589) );
  OAI211_X1 U16551 ( .C1(n14591), .C2(n14674), .A(n14590), .B(n14589), .ZN(
        P2_U3249) );
  AOI21_X1 U16552 ( .B1(n14593), .B2(n14592), .A(n14634), .ZN(n14597) );
  OAI22_X1 U16553 ( .A1(n14637), .A2(n14636), .B1(n14638), .B2(n14594), .ZN(
        n14595) );
  AOI21_X1 U16554 ( .B1(n14597), .B2(n14596), .A(n14595), .ZN(n14756) );
  INV_X1 U16555 ( .A(n14598), .ZN(n14601) );
  INV_X1 U16556 ( .A(n14599), .ZN(n14600) );
  AOI211_X1 U16557 ( .C1(n14754), .C2(n14601), .A(n14658), .B(n14600), .ZN(
        n14753) );
  INV_X1 U16558 ( .A(n14602), .ZN(n14603) );
  AOI22_X1 U16559 ( .A1(n14674), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n14603), 
        .B2(n14661), .ZN(n14604) );
  OAI21_X1 U16560 ( .B1(n14605), .B2(n14664), .A(n14604), .ZN(n14611) );
  AND2_X1 U16561 ( .A1(n14607), .A2(n14606), .ZN(n14608) );
  XNOR2_X1 U16562 ( .A(n14609), .B(n14608), .ZN(n14757) );
  NOR2_X1 U16563 ( .A1(n14757), .A2(n14669), .ZN(n14610) );
  AOI211_X1 U16564 ( .C1(n14753), .C2(n14672), .A(n14611), .B(n14610), .ZN(
        n14612) );
  OAI21_X1 U16565 ( .B1(n14756), .B2(n14674), .A(n14612), .ZN(P2_U3250) );
  XOR2_X1 U16566 ( .A(n14613), .B(n14625), .Z(n14615) );
  AOI21_X1 U16567 ( .B1(n14615), .B2(n14657), .A(n14614), .ZN(n14761) );
  INV_X1 U16568 ( .A(n14640), .ZN(n14616) );
  AOI211_X1 U16569 ( .C1(n14759), .C2(n14616), .A(n14658), .B(n14598), .ZN(
        n14758) );
  INV_X1 U16570 ( .A(n14617), .ZN(n14618) );
  AOI22_X1 U16571 ( .A1(n14674), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n14618), 
        .B2(n14661), .ZN(n14619) );
  OAI21_X1 U16572 ( .B1(n14620), .B2(n14664), .A(n14619), .ZN(n14628) );
  NAND2_X1 U16573 ( .A1(n14622), .A2(n14621), .ZN(n14630) );
  NAND2_X1 U16574 ( .A1(n14630), .A2(n14632), .ZN(n14624) );
  NAND2_X1 U16575 ( .A1(n14624), .A2(n14623), .ZN(n14626) );
  XOR2_X1 U16576 ( .A(n14626), .B(n14625), .Z(n14762) );
  NOR2_X1 U16577 ( .A1(n14762), .A2(n14669), .ZN(n14627) );
  AOI211_X1 U16578 ( .C1(n14758), .C2(n14672), .A(n14628), .B(n14627), .ZN(
        n14629) );
  OAI21_X1 U16579 ( .B1(n14761), .B2(n14674), .A(n14629), .ZN(P2_U3251) );
  XNOR2_X1 U16580 ( .A(n14630), .B(n14632), .ZN(n14765) );
  INV_X1 U16581 ( .A(n14765), .ZN(n14650) );
  AOI21_X1 U16582 ( .B1(n14632), .B2(n14631), .A(n6666), .ZN(n14633) );
  OAI222_X1 U16583 ( .A1(n14638), .A2(n14637), .B1(n14636), .B2(n14635), .C1(
        n14634), .C2(n14633), .ZN(n14763) );
  NAND2_X1 U16584 ( .A1(n14763), .A2(n14645), .ZN(n14649) );
  AOI211_X1 U16585 ( .C1(n14641), .C2(n14639), .A(n14658), .B(n14640), .ZN(
        n14764) );
  NOR2_X1 U16586 ( .A1(n14664), .A2(n14816), .ZN(n14647) );
  OAI22_X1 U16587 ( .A1(n14645), .A2(n14644), .B1(n14643), .B2(n14642), .ZN(
        n14646) );
  AOI211_X1 U16588 ( .C1(n14764), .C2(n14672), .A(n14647), .B(n14646), .ZN(
        n14648) );
  OAI211_X1 U16589 ( .C1(n14669), .C2(n14650), .A(n14649), .B(n14648), .ZN(
        P2_U3252) );
  XNOR2_X1 U16590 ( .A(n14651), .B(n14668), .ZN(n14656) );
  AOI222_X1 U16591 ( .A1(n14657), .A2(n14656), .B1(n14655), .B2(n14654), .C1(
        n14653), .C2(n14652), .ZN(n14772) );
  AOI211_X1 U16592 ( .C1(n14769), .C2(n14659), .A(n14658), .B(n9867), .ZN(
        n14768) );
  INV_X1 U16593 ( .A(n14660), .ZN(n14662) );
  AOI22_X1 U16594 ( .A1(n14674), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n14662), 
        .B2(n14661), .ZN(n14663) );
  OAI21_X1 U16595 ( .B1(n7619), .B2(n14664), .A(n14663), .ZN(n14671) );
  NAND2_X1 U16596 ( .A1(n14666), .A2(n14665), .ZN(n14667) );
  XOR2_X1 U16597 ( .A(n14668), .B(n14667), .Z(n14773) );
  NOR2_X1 U16598 ( .A1(n14773), .A2(n14669), .ZN(n14670) );
  AOI211_X1 U16599 ( .C1(n14768), .C2(n14672), .A(n14671), .B(n14670), .ZN(
        n14673) );
  OAI21_X1 U16600 ( .B1(n14674), .B2(n14772), .A(n14673), .ZN(P2_U3253) );
  INV_X1 U16601 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n14677) );
  NOR2_X1 U16602 ( .A1(n14676), .A2(n14675), .ZN(n14785) );
  MUX2_X1 U16603 ( .A(n14677), .B(n14785), .S(n15944), .Z(n14678) );
  OAI21_X1 U16604 ( .B1(n14788), .B2(n14781), .A(n14678), .ZN(P2_U3530) );
  MUX2_X1 U16605 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n14679), .S(n15944), .Z(
        n14680) );
  INV_X1 U16606 ( .A(n14683), .ZN(P2_U3529) );
  OAI21_X1 U16607 ( .B1(n14686), .B2(n15931), .A(n14685), .ZN(n14687) );
  MUX2_X1 U16608 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n14789), .S(n15944), .Z(
        P2_U3528) );
  AOI21_X1 U16609 ( .B1(n14770), .B2(n14690), .A(n14689), .ZN(n14691) );
  OAI211_X1 U16610 ( .C1(n14774), .C2(n14693), .A(n14692), .B(n14691), .ZN(
        n14790) );
  MUX2_X1 U16611 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14790), .S(n15944), .Z(
        P2_U3526) );
  AOI21_X1 U16612 ( .B1(n14770), .B2(n14695), .A(n14694), .ZN(n14696) );
  OAI211_X1 U16613 ( .C1(n14774), .C2(n14698), .A(n14697), .B(n14696), .ZN(
        n14791) );
  MUX2_X1 U16614 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14791), .S(n15944), .Z(
        P2_U3525) );
  AOI21_X1 U16615 ( .B1(n14770), .B2(n14700), .A(n14699), .ZN(n14701) );
  OAI211_X1 U16616 ( .C1(n14774), .C2(n14703), .A(n14702), .B(n14701), .ZN(
        n14792) );
  MUX2_X1 U16617 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n14792), .S(n15944), .Z(
        P2_U3524) );
  AOI21_X1 U16618 ( .B1(n14770), .B2(n14705), .A(n14704), .ZN(n14706) );
  OAI211_X1 U16619 ( .C1(n14708), .C2(n14774), .A(n14707), .B(n14706), .ZN(
        n14793) );
  MUX2_X1 U16620 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14793), .S(n15944), .Z(
        P2_U3523) );
  AOI21_X1 U16621 ( .B1(n14770), .B2(n14710), .A(n14709), .ZN(n14711) );
  OAI211_X1 U16622 ( .C1(n14774), .C2(n14713), .A(n14712), .B(n14711), .ZN(
        n14794) );
  MUX2_X1 U16623 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14794), .S(n15944), .Z(
        P2_U3522) );
  NOR2_X1 U16624 ( .A1(n14714), .A2(n14774), .ZN(n14718) );
  OAI21_X1 U16625 ( .B1(n14716), .B2(n15931), .A(n14715), .ZN(n14717) );
  MUX2_X1 U16626 ( .A(n14795), .B(P2_REG1_REG_22__SCAN_IN), .S(n15941), .Z(
        P2_U3521) );
  AOI211_X1 U16627 ( .C1(n15929), .C2(n14722), .A(n14721), .B(n14720), .ZN(
        n14796) );
  MUX2_X1 U16628 ( .A(n14723), .B(n14796), .S(n15944), .Z(n14724) );
  OAI21_X1 U16629 ( .B1(n14799), .B2(n14781), .A(n14724), .ZN(P2_U3520) );
  INV_X1 U16630 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n14729) );
  INV_X1 U16631 ( .A(n14725), .ZN(n14728) );
  AOI211_X1 U16632 ( .C1(n14728), .C2(n15929), .A(n14727), .B(n14726), .ZN(
        n14800) );
  MUX2_X1 U16633 ( .A(n14729), .B(n14800), .S(n15944), .Z(n14730) );
  OAI21_X1 U16634 ( .B1(n14803), .B2(n14781), .A(n14730), .ZN(P2_U3519) );
  AOI21_X1 U16635 ( .B1(n14770), .B2(n14732), .A(n14731), .ZN(n14733) );
  OAI211_X1 U16636 ( .C1(n14774), .C2(n14735), .A(n14734), .B(n14733), .ZN(
        n14804) );
  MUX2_X1 U16637 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n14804), .S(n15944), .Z(
        P2_U3518) );
  AOI21_X1 U16638 ( .B1(n14770), .B2(n14737), .A(n14736), .ZN(n14738) );
  OAI211_X1 U16639 ( .C1(n10166), .C2(n14740), .A(n14739), .B(n14738), .ZN(
        n14805) );
  MUX2_X1 U16640 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14805), .S(n15944), .Z(
        P2_U3517) );
  INV_X1 U16641 ( .A(n14741), .ZN(n14744) );
  AOI211_X1 U16642 ( .C1(n14744), .C2(n15929), .A(n14743), .B(n14742), .ZN(
        n14806) );
  MUX2_X1 U16643 ( .A(n14745), .B(n14806), .S(n15944), .Z(n14746) );
  OAI21_X1 U16644 ( .B1(n14809), .B2(n14781), .A(n14746), .ZN(P2_U3516) );
  NAND3_X1 U16645 ( .A1(n14748), .A2(n14747), .A3(n15929), .ZN(n14750) );
  OAI211_X1 U16646 ( .C1(n7627), .C2(n15931), .A(n14750), .B(n14749), .ZN(
        n14751) );
  MUX2_X1 U16647 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14810), .S(n15944), .Z(
        P2_U3515) );
  AOI21_X1 U16648 ( .B1(n14770), .B2(n14754), .A(n14753), .ZN(n14755) );
  OAI211_X1 U16649 ( .C1(n14774), .C2(n14757), .A(n14756), .B(n14755), .ZN(
        n14811) );
  MUX2_X1 U16650 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n14811), .S(n15944), .Z(
        P2_U3514) );
  AOI21_X1 U16651 ( .B1(n14770), .B2(n14759), .A(n14758), .ZN(n14760) );
  OAI211_X1 U16652 ( .C1(n14774), .C2(n14762), .A(n14761), .B(n14760), .ZN(
        n14812) );
  MUX2_X1 U16653 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n14812), .S(n15944), .Z(
        P2_U3513) );
  AOI211_X1 U16654 ( .C1(n15929), .C2(n14765), .A(n14764), .B(n14763), .ZN(
        n14813) );
  MUX2_X1 U16655 ( .A(n14766), .B(n14813), .S(n15944), .Z(n14767) );
  OAI21_X1 U16656 ( .B1(n14816), .B2(n14781), .A(n14767), .ZN(P2_U3512) );
  AOI21_X1 U16657 ( .B1(n14770), .B2(n14769), .A(n14768), .ZN(n14771) );
  OAI211_X1 U16658 ( .C1(n14774), .C2(n14773), .A(n14772), .B(n14771), .ZN(
        n14817) );
  MUX2_X1 U16659 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n14817), .S(n15944), .Z(
        P2_U3511) );
  INV_X1 U16660 ( .A(n14775), .ZN(n14778) );
  AOI211_X1 U16661 ( .C1(n14778), .C2(n15929), .A(n14777), .B(n14776), .ZN(
        n14819) );
  MUX2_X1 U16662 ( .A(n14779), .B(n14819), .S(n15944), .Z(n14780) );
  OAI21_X1 U16663 ( .B1(n14823), .B2(n14781), .A(n14780), .ZN(P2_U3510) );
  OAI211_X1 U16664 ( .C1(n14784), .C2(n10166), .A(n14783), .B(n14782), .ZN(
        n14824) );
  MUX2_X1 U16665 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n14824), .S(n15944), .Z(
        P2_U3499) );
  INV_X1 U16666 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n14786) );
  MUX2_X1 U16667 ( .A(n14786), .B(n14785), .S(n14818), .Z(n14787) );
  OAI21_X1 U16668 ( .B1(n14788), .B2(n14822), .A(n14787), .ZN(P2_U3498) );
  MUX2_X1 U16669 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n14790), .S(n14818), .Z(
        P2_U3494) );
  MUX2_X1 U16670 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14791), .S(n14818), .Z(
        P2_U3493) );
  MUX2_X1 U16671 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n14792), .S(n14818), .Z(
        P2_U3492) );
  MUX2_X1 U16672 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14793), .S(n14818), .Z(
        P2_U3491) );
  MUX2_X1 U16673 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14794), .S(n14818), .Z(
        P2_U3490) );
  MUX2_X1 U16674 ( .A(n14795), .B(P2_REG0_REG_22__SCAN_IN), .S(n15938), .Z(
        P2_U3489) );
  INV_X1 U16675 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n14797) );
  MUX2_X1 U16676 ( .A(n14797), .B(n14796), .S(n14818), .Z(n14798) );
  OAI21_X1 U16677 ( .B1(n14799), .B2(n14822), .A(n14798), .ZN(P2_U3488) );
  MUX2_X1 U16678 ( .A(n14801), .B(n14800), .S(n14818), .Z(n14802) );
  OAI21_X1 U16679 ( .B1(n14803), .B2(n14822), .A(n14802), .ZN(P2_U3487) );
  MUX2_X1 U16680 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n14804), .S(n14818), .Z(
        P2_U3486) );
  MUX2_X1 U16681 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14805), .S(n14818), .Z(
        P2_U3484) );
  INV_X1 U16682 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n14807) );
  MUX2_X1 U16683 ( .A(n14807), .B(n14806), .S(n14818), .Z(n14808) );
  OAI21_X1 U16684 ( .B1(n14809), .B2(n14822), .A(n14808), .ZN(P2_U3481) );
  MUX2_X1 U16685 ( .A(n14810), .B(P2_REG0_REG_16__SCAN_IN), .S(n15938), .Z(
        P2_U3478) );
  MUX2_X1 U16686 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n14811), .S(n14818), .Z(
        P2_U3475) );
  MUX2_X1 U16687 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n14812), .S(n14818), .Z(
        P2_U3472) );
  INV_X1 U16688 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n14814) );
  MUX2_X1 U16689 ( .A(n14814), .B(n14813), .S(n14818), .Z(n14815) );
  OAI21_X1 U16690 ( .B1(n14816), .B2(n14822), .A(n14815), .ZN(P2_U3469) );
  MUX2_X1 U16691 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n14817), .S(n14818), .Z(
        P2_U3466) );
  MUX2_X1 U16692 ( .A(n14820), .B(n14819), .S(n14818), .Z(n14821) );
  OAI21_X1 U16693 ( .B1(n14823), .B2(n14822), .A(n14821), .ZN(P2_U3463) );
  MUX2_X1 U16694 ( .A(P2_REG0_REG_0__SCAN_IN), .B(n14824), .S(n14818), .Z(
        P2_U3430) );
  INV_X1 U16695 ( .A(n14825), .ZN(n15592) );
  OAI222_X1 U16696 ( .A1(P2_U3088), .A2(n14828), .B1(n14832), .B2(n15592), 
        .C1(n14827), .C2(n14826), .ZN(P2_U3298) );
  AOI21_X1 U16697 ( .B1(n14830), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n14829), 
        .ZN(n14831) );
  OAI21_X1 U16698 ( .B1(n14833), .B2(n14832), .A(n14831), .ZN(P2_U3299) );
  INV_X1 U16699 ( .A(n14834), .ZN(n14835) );
  MUX2_X1 U16700 ( .A(n14835), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XOR2_X1 U16701 ( .A(n14836), .B(n14837), .Z(n14838) );
  NAND2_X1 U16702 ( .A1(n14838), .A2(n14969), .ZN(n14848) );
  OAI22_X1 U16703 ( .A1(n14971), .A2(n14839), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8821), .ZN(n14842) );
  NOR2_X1 U16704 ( .A1(n14921), .A2(n14840), .ZN(n14841) );
  NOR2_X1 U16705 ( .A1(n14842), .A2(n14841), .ZN(n14847) );
  NAND2_X1 U16706 ( .A1(n14992), .A2(n15812), .ZN(n14846) );
  INV_X1 U16707 ( .A(n14843), .ZN(n14844) );
  NAND2_X1 U16708 ( .A1(n14928), .A2(n14844), .ZN(n14845) );
  NAND4_X1 U16709 ( .A1(n14848), .A2(n14847), .A3(n14846), .A4(n14845), .ZN(
        P1_U3213) );
  XNOR2_X1 U16710 ( .A(n14850), .B(n14849), .ZN(n14859) );
  INV_X1 U16711 ( .A(n15181), .ZN(n14856) );
  OAI22_X1 U16712 ( .A1(n14852), .A2(n14971), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14851), .ZN(n14853) );
  AOI21_X1 U16713 ( .B1(n14854), .B2(n14928), .A(n14853), .ZN(n14855) );
  OAI21_X1 U16714 ( .B1(n14856), .B2(n14921), .A(n14855), .ZN(n14857) );
  AOI21_X1 U16715 ( .B1(n15469), .B2(n14992), .A(n14857), .ZN(n14858) );
  OAI21_X1 U16716 ( .B1(n14859), .B2(n14994), .A(n14858), .ZN(P1_U3214) );
  XOR2_X1 U16717 ( .A(n14861), .B(n14860), .Z(n14866) );
  AOI22_X1 U16718 ( .A1(n14999), .A2(n15746), .B1(n15426), .B2(n15001), .ZN(
        n15491) );
  NOR2_X1 U16719 ( .A1(n15491), .A2(n14989), .ZN(n14864) );
  OAI22_X1 U16720 ( .A1(n15262), .A2(n14988), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14862), .ZN(n14863) );
  AOI211_X1 U16721 ( .C1(n15265), .C2(n14992), .A(n14864), .B(n14863), .ZN(
        n14865) );
  OAI21_X1 U16722 ( .B1(n14866), .B2(n14994), .A(n14865), .ZN(P1_U3216) );
  AOI211_X1 U16723 ( .C1(n14869), .C2(n14868), .A(n14994), .B(n14867), .ZN(
        n14870) );
  INV_X1 U16724 ( .A(n14870), .ZN(n14874) );
  NAND2_X1 U16725 ( .A1(n14983), .A2(n15003), .ZN(n14871) );
  NAND2_X1 U16726 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n15146)
         );
  OAI211_X1 U16727 ( .C1(n15321), .C2(n14971), .A(n14871), .B(n15146), .ZN(
        n14872) );
  AOI21_X1 U16728 ( .B1(n15323), .B2(n14928), .A(n14872), .ZN(n14873) );
  OAI211_X1 U16729 ( .C1(n15327), .C2(n14963), .A(n14874), .B(n14873), .ZN(
        P1_U3219) );
  OAI21_X1 U16730 ( .B1(n14877), .B2(n14876), .A(n14875), .ZN(n14878) );
  NAND2_X1 U16731 ( .A1(n14878), .A2(n14969), .ZN(n14882) );
  AOI22_X1 U16732 ( .A1(n15001), .A2(n15746), .B1(n15426), .B2(n15003), .ZN(
        n15291) );
  OAI22_X1 U16733 ( .A1(n15291), .A2(n14989), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14879), .ZN(n14880) );
  AOI21_X1 U16734 ( .B1(n15293), .B2(n14928), .A(n14880), .ZN(n14881) );
  OAI211_X1 U16735 ( .C1(n15288), .C2(n14963), .A(n14882), .B(n14881), .ZN(
        P1_U3223) );
  INV_X1 U16736 ( .A(n14952), .ZN(n14885) );
  XNOR2_X1 U16737 ( .A(n14884), .B(n14883), .ZN(n14950) );
  NOR3_X1 U16738 ( .A1(n14886), .A2(n14885), .A3(n14950), .ZN(n14955) );
  AOI21_X1 U16739 ( .B1(n14888), .B2(n14887), .A(n14955), .ZN(n14891) );
  OAI211_X1 U16740 ( .C1(n14891), .C2(n14890), .A(n14969), .B(n14889), .ZN(
        n14897) );
  NAND2_X1 U16741 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n15713)
         );
  OAI21_X1 U16742 ( .B1(n14971), .B2(n14892), .A(n15713), .ZN(n14895) );
  NOR2_X1 U16743 ( .A1(n14988), .A2(n14893), .ZN(n14894) );
  AOI211_X1 U16744 ( .C1(n14983), .C2(n15009), .A(n14895), .B(n14894), .ZN(
        n14896) );
  OAI211_X1 U16745 ( .C1(n7830), .C2(n14963), .A(n14897), .B(n14896), .ZN(
        P1_U3224) );
  AND2_X1 U16746 ( .A1(n14999), .A2(n15426), .ZN(n14899) );
  AOI21_X1 U16747 ( .B1(n14998), .B2(n15746), .A(n14899), .ZN(n15479) );
  INV_X1 U16748 ( .A(n14900), .ZN(n15232) );
  AOI22_X1 U16749 ( .A1(n15232), .A2(n14928), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14901) );
  OAI21_X1 U16750 ( .B1(n15479), .B2(n14989), .A(n14901), .ZN(n14902) );
  AOI21_X1 U16751 ( .B1(n15482), .B2(n14992), .A(n14902), .ZN(n14903) );
  OAI21_X1 U16752 ( .B1(n14904), .B2(n14994), .A(n14903), .ZN(P1_U3225) );
  NAND2_X1 U16753 ( .A1(n6602), .A2(n14905), .ZN(n14907) );
  OAI21_X1 U16754 ( .B1(n6602), .B2(n14905), .A(n14907), .ZN(n14986) );
  INV_X1 U16755 ( .A(n14906), .ZN(n14987) );
  NOR2_X1 U16756 ( .A1(n14986), .A2(n14987), .ZN(n14985) );
  INV_X1 U16757 ( .A(n14907), .ZN(n14908) );
  NOR3_X1 U16758 ( .A1(n14985), .A2(n14909), .A3(n14908), .ZN(n14911) );
  OAI21_X1 U16759 ( .B1(n14911), .B2(n14910), .A(n14969), .ZN(n14915) );
  OAI22_X1 U16760 ( .A1(n15340), .A2(n15411), .B1(n15412), .B2(n15758), .ZN(
        n15372) );
  INV_X1 U16761 ( .A(n15372), .ZN(n14912) );
  NAND2_X1 U16762 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n15096)
         );
  OAI21_X1 U16763 ( .B1(n14912), .B2(n14989), .A(n15096), .ZN(n14913) );
  AOI21_X1 U16764 ( .B1(n15379), .B2(n14928), .A(n14913), .ZN(n14914) );
  OAI211_X1 U16765 ( .C1(n7825), .C2(n14963), .A(n14915), .B(n14914), .ZN(
        P1_U3226) );
  INV_X1 U16766 ( .A(n14916), .ZN(n14917) );
  NOR2_X1 U16767 ( .A1(n14918), .A2(n14917), .ZN(n14919) );
  XNOR2_X1 U16768 ( .A(n6745), .B(n14919), .ZN(n14925) );
  NAND2_X1 U16769 ( .A1(n14978), .A2(n15006), .ZN(n14920) );
  NAND2_X1 U16770 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n15110)
         );
  OAI211_X1 U16771 ( .C1(n15321), .C2(n14921), .A(n14920), .B(n15110), .ZN(
        n14923) );
  NOR2_X1 U16772 ( .A1(n7824), .A2(n14963), .ZN(n14922) );
  AOI211_X1 U16773 ( .C1(n14928), .C2(n15364), .A(n14923), .B(n14922), .ZN(
        n14924) );
  OAI21_X1 U16774 ( .B1(n14925), .B2(n14994), .A(n14924), .ZN(P1_U3228) );
  XOR2_X1 U16775 ( .A(n14927), .B(n14926), .Z(n14932) );
  AOI22_X1 U16776 ( .A1(n15212), .A2(n15746), .B1(n15426), .B2(n15000), .ZN(
        n15248) );
  AOI22_X1 U16777 ( .A1(n15252), .A2(n14928), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14929) );
  OAI21_X1 U16778 ( .B1(n15248), .B2(n14989), .A(n14929), .ZN(n14930) );
  AOI21_X1 U16779 ( .B1(n15488), .B2(n14992), .A(n14930), .ZN(n14931) );
  OAI21_X1 U16780 ( .B1(n14932), .B2(n14994), .A(n14931), .ZN(P1_U3229) );
  NOR2_X1 U16781 ( .A1(n15341), .A2(n15758), .ZN(n14933) );
  AOI21_X1 U16782 ( .B1(n15002), .B2(n15746), .A(n14933), .ZN(n15510) );
  INV_X1 U16783 ( .A(n15510), .ZN(n14934) );
  AOI22_X1 U16784 ( .A1(n14934), .A2(n14960), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14935) );
  OAI21_X1 U16785 ( .B1(n15306), .B2(n14988), .A(n14935), .ZN(n14939) );
  AOI211_X1 U16786 ( .C1(n6559), .C2(n14937), .A(n14994), .B(n14936), .ZN(
        n14938) );
  AOI211_X1 U16787 ( .C1(n14992), .C2(n15305), .A(n14939), .B(n14938), .ZN(
        n14940) );
  INV_X1 U16788 ( .A(n14940), .ZN(P1_U3233) );
  OAI21_X1 U16789 ( .B1(n14943), .B2(n14942), .A(n14941), .ZN(n14944) );
  NAND2_X1 U16790 ( .A1(n14944), .A2(n14969), .ZN(n14949) );
  NOR2_X1 U16791 ( .A1(n14988), .A2(n15272), .ZN(n14947) );
  OAI22_X1 U16792 ( .A1(n12727), .A2(n14971), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14945), .ZN(n14946) );
  AOI211_X1 U16793 ( .C1(n15000), .C2(n14983), .A(n14947), .B(n14946), .ZN(
        n14948) );
  OAI211_X1 U16794 ( .C1(n14963), .C2(n15277), .A(n14949), .B(n14948), .ZN(
        P1_U3235) );
  INV_X1 U16795 ( .A(n14950), .ZN(n14951) );
  AOI21_X1 U16796 ( .B1(n14953), .B2(n14952), .A(n14951), .ZN(n14954) );
  OAI21_X1 U16797 ( .B1(n14955), .B2(n14954), .A(n14969), .ZN(n14962) );
  NOR2_X1 U16798 ( .A1(n14988), .A2(n14956), .ZN(n14957) );
  AOI211_X1 U16799 ( .C1(n14960), .C2(n14959), .A(n14958), .B(n14957), .ZN(
        n14961) );
  OAI211_X1 U16800 ( .C1(n14964), .C2(n14963), .A(n14962), .B(n14961), .ZN(
        P1_U3236) );
  AND2_X1 U16801 ( .A1(n14965), .A2(n15813), .ZN(n15525) );
  INV_X1 U16802 ( .A(n15525), .ZN(n14976) );
  OAI21_X1 U16803 ( .B1(n14968), .B2(n14967), .A(n14966), .ZN(n14970) );
  NAND2_X1 U16804 ( .A1(n14970), .A2(n14969), .ZN(n14975) );
  OAI22_X1 U16805 ( .A1(n14971), .A2(n15340), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15116), .ZN(n14973) );
  NOR2_X1 U16806 ( .A1(n14988), .A2(n15346), .ZN(n14972) );
  AOI211_X1 U16807 ( .C1(n14983), .C2(n15004), .A(n14973), .B(n14972), .ZN(
        n14974) );
  OAI211_X1 U16808 ( .C1(n14976), .C2(n14980), .A(n14975), .B(n14974), .ZN(
        P1_U3238) );
  AOI22_X1 U16809 ( .A1(n15212), .A2(n14978), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14979) );
  OAI21_X1 U16810 ( .B1(n15220), .B2(n14988), .A(n14979), .ZN(n14982) );
  NAND2_X1 U16811 ( .A1(n15222), .A2(n15813), .ZN(n15477) );
  NOR2_X1 U16812 ( .A1(n15477), .A2(n14980), .ZN(n14981) );
  AOI211_X1 U16813 ( .C1(n14983), .C2(n15213), .A(n14982), .B(n14981), .ZN(
        n14984) );
  AOI21_X1 U16814 ( .B1(n14987), .B2(n14986), .A(n14985), .ZN(n14995) );
  NOR2_X1 U16815 ( .A1(n14988), .A2(n15394), .ZN(n14991) );
  AOI22_X1 U16816 ( .A1(n15006), .A2(n15746), .B1(n15426), .B2(n15008), .ZN(
        n15390) );
  NAND2_X1 U16817 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n15726)
         );
  OAI21_X1 U16818 ( .B1(n14989), .B2(n15390), .A(n15726), .ZN(n14990) );
  AOI211_X1 U16819 ( .C1(n15543), .C2(n14992), .A(n14991), .B(n14990), .ZN(
        n14993) );
  OAI21_X1 U16820 ( .B1(n14995), .B2(n14994), .A(n14993), .ZN(P1_U3241) );
  INV_X1 U16821 ( .A(n14996), .ZN(n15151) );
  MUX2_X1 U16822 ( .A(n15151), .B(P1_DATAO_REG_31__SCAN_IN), .S(n15019), .Z(
        P1_U3591) );
  MUX2_X1 U16823 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n15177), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16824 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14997), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16825 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n15181), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16826 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n15213), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16827 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14998), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16828 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n15212), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16829 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14999), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16830 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n15000), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16831 ( .A(n15001), .B(P1_DATAO_REG_22__SCAN_IN), .S(n15019), .Z(
        P1_U3582) );
  MUX2_X1 U16832 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n15002), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16833 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n15003), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16834 ( .A(n15004), .B(P1_DATAO_REG_19__SCAN_IN), .S(n15019), .Z(
        P1_U3579) );
  MUX2_X1 U16835 ( .A(n15359), .B(P1_DATAO_REG_18__SCAN_IN), .S(n15019), .Z(
        P1_U3578) );
  MUX2_X1 U16836 ( .A(n15005), .B(P1_DATAO_REG_17__SCAN_IN), .S(n15019), .Z(
        P1_U3577) );
  MUX2_X1 U16837 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n15006), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16838 ( .A(n15007), .B(P1_DATAO_REG_15__SCAN_IN), .S(n15019), .Z(
        P1_U3575) );
  MUX2_X1 U16839 ( .A(n15008), .B(P1_DATAO_REG_14__SCAN_IN), .S(n15019), .Z(
        P1_U3574) );
  MUX2_X1 U16840 ( .A(n15009), .B(P1_DATAO_REG_13__SCAN_IN), .S(n15019), .Z(
        P1_U3573) );
  MUX2_X1 U16841 ( .A(n15010), .B(P1_DATAO_REG_12__SCAN_IN), .S(n15019), .Z(
        P1_U3572) );
  MUX2_X1 U16842 ( .A(n15011), .B(P1_DATAO_REG_11__SCAN_IN), .S(n15019), .Z(
        P1_U3571) );
  MUX2_X1 U16843 ( .A(n15012), .B(P1_DATAO_REG_10__SCAN_IN), .S(n15019), .Z(
        P1_U3570) );
  MUX2_X1 U16844 ( .A(n15013), .B(P1_DATAO_REG_9__SCAN_IN), .S(n15019), .Z(
        P1_U3569) );
  MUX2_X1 U16845 ( .A(n15014), .B(P1_DATAO_REG_8__SCAN_IN), .S(n15019), .Z(
        P1_U3568) );
  MUX2_X1 U16846 ( .A(n15015), .B(P1_DATAO_REG_7__SCAN_IN), .S(n15019), .Z(
        P1_U3567) );
  MUX2_X1 U16847 ( .A(n15016), .B(P1_DATAO_REG_6__SCAN_IN), .S(n15019), .Z(
        P1_U3566) );
  MUX2_X1 U16848 ( .A(n15017), .B(P1_DATAO_REG_5__SCAN_IN), .S(n15019), .Z(
        P1_U3565) );
  MUX2_X1 U16849 ( .A(n15018), .B(P1_DATAO_REG_4__SCAN_IN), .S(n15019), .Z(
        P1_U3564) );
  MUX2_X1 U16850 ( .A(n15425), .B(P1_DATAO_REG_3__SCAN_IN), .S(n15019), .Z(
        P1_U3563) );
  MUX2_X1 U16851 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n15745), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16852 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n15751), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16853 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n15753), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI22_X1 U16854 ( .A1(n15728), .A2(n15021), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15020), .ZN(n15022) );
  AOI21_X1 U16855 ( .B1(n15023), .B2(n15720), .A(n15022), .ZN(n15033) );
  OAI211_X1 U16856 ( .C1(n15026), .C2(n15025), .A(n15723), .B(n15024), .ZN(
        n15032) );
  INV_X1 U16857 ( .A(n15027), .ZN(n15030) );
  OAI211_X1 U16858 ( .C1(n15030), .C2(n15029), .A(n15724), .B(n15028), .ZN(
        n15031) );
  NAND3_X1 U16859 ( .A1(n15033), .A2(n15032), .A3(n15031), .ZN(P1_U3244) );
  NOR2_X1 U16860 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n15034), .ZN(n15037) );
  NOR2_X1 U16861 ( .A1(n15728), .A2(n15035), .ZN(n15036) );
  AOI211_X1 U16862 ( .C1(n15720), .C2(n15040), .A(n15037), .B(n15036), .ZN(
        n15047) );
  OAI211_X1 U16863 ( .C1(n15039), .C2(n15038), .A(n15723), .B(n15691), .ZN(
        n15046) );
  MUX2_X1 U16864 ( .A(n7249), .B(P1_REG2_REG_3__SCAN_IN), .S(n15040), .Z(
        n15043) );
  NAND3_X1 U16865 ( .A1(n15043), .A2(n15042), .A3(n15041), .ZN(n15044) );
  NAND3_X1 U16866 ( .A1(n15724), .A2(n15687), .A3(n15044), .ZN(n15045) );
  NAND3_X1 U16867 ( .A1(n15047), .A2(n15046), .A3(n15045), .ZN(P1_U3246) );
  OAI211_X1 U16868 ( .C1(n15050), .C2(n15049), .A(n15048), .B(n15723), .ZN(
        n15063) );
  OAI21_X1 U16869 ( .B1(n15728), .B2(n15052), .A(n15051), .ZN(n15053) );
  AOI21_X1 U16870 ( .B1(n15054), .B2(n15720), .A(n15053), .ZN(n15062) );
  MUX2_X1 U16871 ( .A(n12028), .B(P1_REG2_REG_10__SCAN_IN), .S(n15054), .Z(
        n15057) );
  INV_X1 U16872 ( .A(n15055), .ZN(n15056) );
  NAND2_X1 U16873 ( .A1(n15057), .A2(n15056), .ZN(n15059) );
  OAI211_X1 U16874 ( .C1(n15060), .C2(n15059), .A(n15058), .B(n15724), .ZN(
        n15061) );
  NAND3_X1 U16875 ( .A1(n15063), .A2(n15062), .A3(n15061), .ZN(P1_U3253) );
  XNOR2_X1 U16876 ( .A(n15081), .B(n15064), .ZN(n15068) );
  OAI21_X1 U16877 ( .B1(n15068), .B2(n15067), .A(n15080), .ZN(n15069) );
  NAND2_X1 U16878 ( .A1(n15069), .A2(n15723), .ZN(n15079) );
  OAI21_X1 U16879 ( .B1(n15728), .B2(n15614), .A(n15070), .ZN(n15071) );
  AOI21_X1 U16880 ( .B1(n15081), .B2(n15720), .A(n15071), .ZN(n15078) );
  NOR2_X1 U16881 ( .A1(n15072), .A2(n11772), .ZN(n15074) );
  INV_X1 U16882 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n15088) );
  MUX2_X1 U16883 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n15088), .S(n15081), .Z(
        n15073) );
  OAI21_X1 U16884 ( .B1(n15075), .B2(n15074), .A(n15073), .ZN(n15086) );
  OR3_X1 U16885 ( .A1(n15075), .A2(n15074), .A3(n15073), .ZN(n15076) );
  NAND3_X1 U16886 ( .A1(n15086), .A2(n15724), .A3(n15076), .ZN(n15077) );
  NAND3_X1 U16887 ( .A1(n15079), .A2(n15078), .A3(n15077), .ZN(P1_U3257) );
  XNOR2_X1 U16888 ( .A(n15101), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n15085) );
  INV_X1 U16889 ( .A(n15082), .ZN(n15083) );
  AOI211_X1 U16890 ( .C1(n15085), .C2(n15084), .A(n15102), .B(n6759), .ZN(
        n15100) );
  OAI21_X1 U16891 ( .B1(n15088), .B2(n15087), .A(n15086), .ZN(n15089) );
  NOR2_X1 U16892 ( .A1(n15089), .A2(n15721), .ZN(n15090) );
  AOI21_X1 U16893 ( .B1(n15721), .B2(n15089), .A(n15090), .ZN(n15718) );
  INV_X1 U16894 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n15717) );
  INV_X1 U16895 ( .A(n15090), .ZN(n15091) );
  INV_X1 U16896 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n15092) );
  MUX2_X1 U16897 ( .A(n15092), .B(P1_REG2_REG_16__SCAN_IN), .S(n15101), .Z(
        n15094) );
  INV_X1 U16898 ( .A(n15105), .ZN(n15093) );
  AOI211_X1 U16899 ( .C1(n15095), .C2(n15094), .A(n15142), .B(n15093), .ZN(
        n15099) );
  NAND2_X1 U16900 ( .A1(n15680), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n15097) );
  OAI211_X1 U16901 ( .C1(n15699), .C2(n15106), .A(n15097), .B(n15096), .ZN(
        n15098) );
  OR3_X1 U16902 ( .A1(n15100), .A2(n15099), .A3(n15098), .ZN(P1_U3259) );
  XNOR2_X1 U16903 ( .A(n15123), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n15103) );
  NOR2_X1 U16904 ( .A1(n15104), .A2(n15103), .ZN(n15122) );
  AOI211_X1 U16905 ( .C1(n15104), .C2(n15103), .A(n15102), .B(n15122), .ZN(
        n15115) );
  MUX2_X1 U16906 ( .A(n15107), .B(P1_REG2_REG_17__SCAN_IN), .S(n15120), .Z(
        n15108) );
  NAND2_X1 U16907 ( .A1(n15108), .A2(n15109), .ZN(n15119) );
  OAI211_X1 U16908 ( .C1(n15109), .C2(n15108), .A(n15724), .B(n15119), .ZN(
        n15113) );
  INV_X1 U16909 ( .A(n15110), .ZN(n15111) );
  AOI21_X1 U16910 ( .B1(n15680), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n15111), 
        .ZN(n15112) );
  OAI211_X1 U16911 ( .C1(n15699), .C2(n15120), .A(n15113), .B(n15112), .ZN(
        n15114) );
  OR2_X1 U16912 ( .A1(n15115), .A2(n15114), .ZN(P1_U3260) );
  NOR2_X1 U16913 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n15116), .ZN(n15118) );
  NOR2_X1 U16914 ( .A1(n15699), .A2(n15131), .ZN(n15117) );
  AOI211_X1 U16915 ( .C1(n15680), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n15118), 
        .B(n15117), .ZN(n15130) );
  OAI21_X1 U16916 ( .B1(n15107), .B2(n15120), .A(n15119), .ZN(n15136) );
  XNOR2_X1 U16917 ( .A(n15131), .B(n15136), .ZN(n15121) );
  NAND2_X1 U16918 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n15121), .ZN(n15139) );
  OAI211_X1 U16919 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n15121), .A(n15724), 
        .B(n15139), .ZN(n15129) );
  INV_X1 U16920 ( .A(n15124), .ZN(n15127) );
  INV_X1 U16921 ( .A(n15134), .ZN(n15126) );
  OAI211_X1 U16922 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n15127), .A(n15723), 
        .B(n15126), .ZN(n15128) );
  NAND3_X1 U16923 ( .A1(n15130), .A2(n15129), .A3(n15128), .ZN(P1_U3261) );
  NOR2_X1 U16924 ( .A1(n15132), .A2(n15131), .ZN(n15133) );
  INV_X1 U16925 ( .A(n15145), .ZN(n15143) );
  NAND2_X1 U16926 ( .A1(n15137), .A2(n15136), .ZN(n15138) );
  NAND2_X1 U16927 ( .A1(n15139), .A2(n15138), .ZN(n15141) );
  XNOR2_X1 U16928 ( .A(n15141), .B(n15140), .ZN(n15144) );
  NAND2_X1 U16929 ( .A1(n15447), .A2(n15174), .ZN(n15155) );
  AOI21_X1 U16930 ( .B1(n15150), .B2(P1_B_REG_SCAN_IN), .A(n15411), .ZN(n15178) );
  NAND2_X1 U16931 ( .A1(n15178), .A2(n15151), .ZN(n15445) );
  NOR2_X1 U16932 ( .A1(n15445), .A2(n15764), .ZN(n15157) );
  NOR2_X1 U16933 ( .A1(n15148), .A2(n15418), .ZN(n15153) );
  AOI211_X1 U16934 ( .C1(n15764), .C2(P1_REG2_REG_31__SCAN_IN), .A(n15157), 
        .B(n15153), .ZN(n15154) );
  OAI21_X1 U16935 ( .B1(n15304), .B2(n15444), .A(n15154), .ZN(P1_U3263) );
  OAI211_X1 U16936 ( .C1(n15447), .C2(n15174), .A(n10870), .B(n15155), .ZN(
        n15446) );
  NOR2_X1 U16937 ( .A1(n6544), .A2(n15156), .ZN(n15158) );
  AOI211_X1 U16938 ( .C1(n15159), .C2(n15730), .A(n15158), .B(n15157), .ZN(
        n15160) );
  OAI21_X1 U16939 ( .B1(n15446), .B2(n15304), .A(n15160), .ZN(P1_U3264) );
  NAND2_X1 U16940 ( .A1(n15191), .A2(n15204), .ZN(n15190) );
  NAND2_X1 U16941 ( .A1(n15190), .A2(n7985), .ZN(n15163) );
  XNOR2_X1 U16942 ( .A(n15163), .B(n15168), .ZN(n15448) );
  INV_X1 U16943 ( .A(n15448), .ZN(n15189) );
  NAND2_X1 U16944 ( .A1(n15164), .A2(n15169), .ZN(n15173) );
  OR2_X1 U16945 ( .A1(n15469), .A2(n15213), .ZN(n15200) );
  AND2_X1 U16946 ( .A1(n15165), .A2(n15200), .ZN(n15166) );
  NAND3_X1 U16947 ( .A1(n15201), .A2(n15166), .A3(n15168), .ZN(n15172) );
  INV_X1 U16948 ( .A(n15166), .ZN(n15167) );
  NAND2_X1 U16949 ( .A1(n15167), .A2(n15169), .ZN(n15170) );
  MUX2_X1 U16950 ( .A(n15170), .B(n15169), .S(n15168), .Z(n15171) );
  OAI211_X1 U16951 ( .C1(n15201), .C2(n15173), .A(n15172), .B(n15171), .ZN(
        n15454) );
  AOI211_X1 U16952 ( .C1(n15175), .C2(n15196), .A(n15742), .B(n15174), .ZN(
        n15453) );
  NAND2_X1 U16953 ( .A1(n15453), .A2(n15732), .ZN(n15186) );
  INV_X1 U16954 ( .A(n15176), .ZN(n15184) );
  NAND2_X1 U16955 ( .A1(n15178), .A2(n15177), .ZN(n15450) );
  INV_X1 U16956 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n15179) );
  OAI22_X1 U16957 ( .A1(n15450), .A2(n15180), .B1(n15179), .B2(n6544), .ZN(
        n15183) );
  NAND2_X1 U16958 ( .A1(n15181), .A2(n15426), .ZN(n15449) );
  NOR2_X1 U16959 ( .A1(n15449), .A2(n15764), .ZN(n15182) );
  AOI211_X1 U16960 ( .C1(n15760), .C2(n15184), .A(n15183), .B(n15182), .ZN(
        n15185) );
  OAI211_X1 U16961 ( .C1(n15451), .C2(n15418), .A(n15186), .B(n15185), .ZN(
        n15187) );
  AOI21_X1 U16962 ( .B1(n15383), .B2(n15454), .A(n15187), .ZN(n15188) );
  OAI21_X1 U16963 ( .B1(n15189), .B2(n15333), .A(n15188), .ZN(P1_U3356) );
  OAI21_X1 U16964 ( .B1(n15191), .B2(n15204), .A(n15190), .ZN(n15460) );
  INV_X1 U16965 ( .A(n15460), .ZN(n15208) );
  AOI22_X1 U16966 ( .A1(n15192), .A2(n15760), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n15764), .ZN(n15193) );
  OAI21_X1 U16967 ( .B1(n15194), .B2(n15764), .A(n15193), .ZN(n15199) );
  AOI21_X1 U16968 ( .B1(n15462), .B2(n15195), .A(n15742), .ZN(n15197) );
  NAND2_X1 U16969 ( .A1(n15197), .A2(n15196), .ZN(n15464) );
  NOR2_X1 U16970 ( .A1(n15464), .A2(n15304), .ZN(n15198) );
  AOI211_X1 U16971 ( .C1(n15730), .C2(n15462), .A(n15199), .B(n15198), .ZN(
        n15207) );
  NAND2_X1 U16972 ( .A1(n15203), .A2(n15202), .ZN(n15458) );
  NAND2_X1 U16973 ( .A1(n15205), .A2(n15204), .ZN(n15459) );
  NAND3_X1 U16974 ( .A1(n15458), .A2(n15383), .A3(n15459), .ZN(n15206) );
  OAI211_X1 U16975 ( .C1(n15208), .C2(n15333), .A(n15207), .B(n15206), .ZN(
        P1_U3265) );
  NAND3_X1 U16976 ( .A1(n15209), .A2(n7635), .A3(n15210), .ZN(n15211) );
  NAND2_X1 U16977 ( .A1(n12737), .A2(n15211), .ZN(n15214) );
  AOI222_X1 U16978 ( .A1(n15214), .A2(n15754), .B1(n15213), .B2(n15746), .C1(
        n15212), .C2(n15426), .ZN(n15478) );
  INV_X1 U16979 ( .A(n15231), .ZN(n15215) );
  AOI21_X1 U16980 ( .B1(n15215), .B2(n15222), .A(n15742), .ZN(n15218) );
  INV_X1 U16981 ( .A(n15216), .ZN(n15217) );
  NAND2_X1 U16982 ( .A1(n15218), .A2(n15217), .ZN(n15475) );
  INV_X1 U16983 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n15219) );
  OAI22_X1 U16984 ( .A1(n15220), .A2(n15393), .B1(n15219), .B2(n6544), .ZN(
        n15221) );
  AOI21_X1 U16985 ( .B1(n15222), .B2(n15730), .A(n15221), .ZN(n15223) );
  OAI21_X1 U16986 ( .B1(n15475), .B2(n15304), .A(n15223), .ZN(n15224) );
  INV_X1 U16987 ( .A(n15224), .ZN(n15227) );
  OR2_X1 U16988 ( .A1(n15225), .A2(n7635), .ZN(n15474) );
  NAND3_X1 U16989 ( .A1(n15474), .A2(n15383), .A3(n15473), .ZN(n15226) );
  OAI211_X1 U16990 ( .C1(n15478), .C2(n15764), .A(n15227), .B(n15226), .ZN(
        P1_U3267) );
  XNOR2_X1 U16991 ( .A(n15228), .B(n15235), .ZN(n15485) );
  NAND2_X1 U16992 ( .A1(n15250), .A2(n15482), .ZN(n15229) );
  NAND2_X1 U16993 ( .A1(n15229), .A2(n10870), .ZN(n15230) );
  NOR2_X1 U16994 ( .A1(n15231), .A2(n15230), .ZN(n15480) );
  INV_X1 U16995 ( .A(n15482), .ZN(n15234) );
  AOI22_X1 U16996 ( .A1(n15232), .A2(n15760), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n15764), .ZN(n15233) );
  OAI21_X1 U16997 ( .B1(n15234), .B2(n15418), .A(n15233), .ZN(n15239) );
  OAI21_X1 U16998 ( .B1(n15236), .B2(n15235), .A(n15209), .ZN(n15237) );
  NAND2_X1 U16999 ( .A1(n15237), .A2(n15754), .ZN(n15484) );
  AOI21_X1 U17000 ( .B1(n15484), .B2(n15479), .A(n15764), .ZN(n15238) );
  AOI211_X1 U17001 ( .C1(n15480), .C2(n15732), .A(n15239), .B(n15238), .ZN(
        n15240) );
  OAI21_X1 U17002 ( .B1(n15423), .B2(n15485), .A(n15240), .ZN(P1_U3268) );
  XNOR2_X1 U17003 ( .A(n15241), .B(n15244), .ZN(n15490) );
  INV_X1 U17004 ( .A(n15242), .ZN(n15247) );
  NOR3_X1 U17005 ( .A1(n15243), .A2(n15245), .A3(n15244), .ZN(n15246) );
  OAI21_X1 U17006 ( .B1(n15247), .B2(n15246), .A(n15754), .ZN(n15249) );
  NAND2_X1 U17007 ( .A1(n15249), .A2(n15248), .ZN(n15486) );
  AOI21_X1 U17008 ( .B1(n6578), .B2(n15488), .A(n15742), .ZN(n15251) );
  AND2_X1 U17009 ( .A1(n15251), .A2(n15250), .ZN(n15487) );
  NAND2_X1 U17010 ( .A1(n15487), .A2(n15732), .ZN(n15254) );
  AOI22_X1 U17011 ( .A1(n15252), .A2(n15760), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n15764), .ZN(n15253) );
  OAI211_X1 U17012 ( .C1(n15255), .C2(n15418), .A(n15254), .B(n15253), .ZN(
        n15256) );
  AOI21_X1 U17013 ( .B1(n15486), .B2(n6544), .A(n15256), .ZN(n15257) );
  OAI21_X1 U17014 ( .B1(n15423), .B2(n15490), .A(n15257), .ZN(P1_U3269) );
  XOR2_X1 U17015 ( .A(n15259), .B(n15258), .Z(n15497) );
  AOI21_X1 U17016 ( .B1(n15260), .B2(n15259), .A(n15243), .ZN(n15261) );
  INV_X1 U17017 ( .A(n15261), .ZN(n15495) );
  OAI211_X1 U17018 ( .C1(n15270), .C2(n15493), .A(n10870), .B(n6578), .ZN(
        n15492) );
  OAI21_X1 U17019 ( .B1(n15262), .B2(n15393), .A(n15491), .ZN(n15263) );
  MUX2_X1 U17020 ( .A(P1_REG2_REG_23__SCAN_IN), .B(n15263), .S(n6544), .Z(
        n15264) );
  AOI21_X1 U17021 ( .B1(n15265), .B2(n15730), .A(n15264), .ZN(n15266) );
  OAI21_X1 U17022 ( .B1(n15492), .B2(n15304), .A(n15266), .ZN(n15267) );
  AOI21_X1 U17023 ( .B1(n15495), .B2(n15313), .A(n15267), .ZN(n15268) );
  OAI21_X1 U17024 ( .B1(n15497), .B2(n15423), .A(n15268), .ZN(P1_U3270) );
  XNOR2_X1 U17025 ( .A(n15269), .B(n15280), .ZN(n15504) );
  OAI21_X1 U17026 ( .B1(n15286), .B2(n15277), .A(n10870), .ZN(n15271) );
  NOR2_X1 U17027 ( .A1(n15271), .A2(n15270), .ZN(n15498) );
  INV_X1 U17028 ( .A(n15272), .ZN(n15273) );
  AOI22_X1 U17029 ( .A1(n15273), .A2(n15760), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n15764), .ZN(n15276) );
  OAI22_X1 U17030 ( .A1(n15274), .A2(n15411), .B1(n12727), .B2(n15758), .ZN(
        n15499) );
  NAND2_X1 U17031 ( .A1(n15499), .A2(n6544), .ZN(n15275) );
  OAI211_X1 U17032 ( .C1(n15277), .C2(n15418), .A(n15276), .B(n15275), .ZN(
        n15278) );
  AOI21_X1 U17033 ( .B1(n15498), .B2(n15732), .A(n15278), .ZN(n15283) );
  OAI21_X1 U17034 ( .B1(n15281), .B2(n15280), .A(n15279), .ZN(n15501) );
  NAND2_X1 U17035 ( .A1(n15501), .A2(n15383), .ZN(n15282) );
  OAI211_X1 U17036 ( .C1(n15504), .C2(n15333), .A(n15283), .B(n15282), .ZN(
        P1_U3271) );
  XNOR2_X1 U17037 ( .A(n15285), .B(n15284), .ZN(n15509) );
  AOI211_X1 U17038 ( .C1(n15507), .C2(n15302), .A(n15742), .B(n15286), .ZN(
        n15506) );
  OAI22_X1 U17039 ( .A1(n15288), .A2(n15418), .B1(n15287), .B2(n6544), .ZN(
        n15296) );
  XNOR2_X1 U17040 ( .A(n15290), .B(n15289), .ZN(n15292) );
  OAI21_X1 U17041 ( .B1(n15292), .B2(n15829), .A(n15291), .ZN(n15505) );
  AOI21_X1 U17042 ( .B1(n15293), .B2(n15760), .A(n15505), .ZN(n15294) );
  NOR2_X1 U17043 ( .A1(n15294), .A2(n15764), .ZN(n15295) );
  AOI211_X1 U17044 ( .C1(n15506), .C2(n15732), .A(n15296), .B(n15295), .ZN(
        n15297) );
  OAI21_X1 U17045 ( .B1(n15509), .B2(n15423), .A(n15297), .ZN(P1_U3272) );
  OAI21_X1 U17046 ( .B1(n7447), .B2(n6587), .A(n6723), .ZN(n15516) );
  OAI21_X1 U17047 ( .B1(n15300), .B2(n15299), .A(n15298), .ZN(n15301) );
  INV_X1 U17048 ( .A(n15301), .ZN(n15514) );
  AOI21_X1 U17049 ( .B1(n15318), .B2(n15305), .A(n15742), .ZN(n15303) );
  NAND2_X1 U17050 ( .A1(n15303), .A2(n15302), .ZN(n15511) );
  NOR2_X1 U17051 ( .A1(n15511), .A2(n15304), .ZN(n15312) );
  NAND2_X1 U17052 ( .A1(n15305), .A2(n15730), .ZN(n15309) );
  OAI22_X1 U17053 ( .A1(n15510), .A2(n15764), .B1(n15306), .B2(n15393), .ZN(
        n15307) );
  INV_X1 U17054 ( .A(n15307), .ZN(n15308) );
  OAI211_X1 U17055 ( .C1(n6544), .C2(n15310), .A(n15309), .B(n15308), .ZN(
        n15311) );
  AOI211_X1 U17056 ( .C1(n15514), .C2(n15313), .A(n15312), .B(n15311), .ZN(
        n15314) );
  OAI21_X1 U17057 ( .B1(n15423), .B2(n15516), .A(n15314), .ZN(P1_U3273) );
  AOI21_X1 U17058 ( .B1(n15317), .B2(n15316), .A(n15315), .ZN(n15523) );
  INV_X1 U17059 ( .A(n15343), .ZN(n15320) );
  INV_X1 U17060 ( .A(n15318), .ZN(n15319) );
  AOI211_X1 U17061 ( .C1(n15519), .C2(n15320), .A(n15742), .B(n15319), .ZN(
        n15517) );
  OAI22_X1 U17062 ( .A1(n15322), .A2(n15411), .B1(n15321), .B2(n15758), .ZN(
        n15518) );
  AOI21_X1 U17063 ( .B1(n15323), .B2(n15760), .A(n15518), .ZN(n15324) );
  NOR2_X1 U17064 ( .A1(n15324), .A2(n15764), .ZN(n15325) );
  AOI21_X1 U17065 ( .B1(n15764), .B2(P1_REG2_REG_19__SCAN_IN), .A(n15325), 
        .ZN(n15326) );
  OAI21_X1 U17066 ( .B1(n15327), .B2(n15418), .A(n15326), .ZN(n15328) );
  AOI21_X1 U17067 ( .B1(n15517), .B2(n15732), .A(n15328), .ZN(n15332) );
  XNOR2_X1 U17068 ( .A(n15330), .B(n15329), .ZN(n15520) );
  NAND2_X1 U17069 ( .A1(n15520), .A2(n15383), .ZN(n15331) );
  OAI211_X1 U17070 ( .C1(n15523), .C2(n15333), .A(n15332), .B(n15331), .ZN(
        P1_U3274) );
  XNOR2_X1 U17071 ( .A(n15335), .B(n15334), .ZN(n15528) );
  NOR2_X1 U17072 ( .A1(n15409), .A2(n15355), .ZN(n15338) );
  OAI21_X1 U17073 ( .B1(n15338), .B2(n15337), .A(n15336), .ZN(n15339) );
  XNOR2_X1 U17074 ( .A(n15339), .B(n12720), .ZN(n15342) );
  OAI222_X1 U17075 ( .A1(n15342), .A2(n15829), .B1(n15411), .B2(n15341), .C1(
        n15758), .C2(n15340), .ZN(n15526) );
  NAND2_X1 U17076 ( .A1(n15526), .A2(n6544), .ZN(n15351) );
  OAI21_X1 U17077 ( .B1(n15363), .B2(n15345), .A(n10870), .ZN(n15344) );
  NOR2_X1 U17078 ( .A1(n15344), .A2(n15343), .ZN(n15524) );
  NOR2_X1 U17079 ( .A1(n15345), .A2(n15418), .ZN(n15349) );
  OAI22_X1 U17080 ( .A1(n6544), .A2(n15347), .B1(n15346), .B2(n15393), .ZN(
        n15348) );
  AOI211_X1 U17081 ( .C1(n15524), .C2(n15732), .A(n15349), .B(n15348), .ZN(
        n15350) );
  OAI211_X1 U17082 ( .C1(n15528), .C2(n15423), .A(n15351), .B(n15350), .ZN(
        P1_U3275) );
  XNOR2_X1 U17083 ( .A(n15352), .B(n15357), .ZN(n15534) );
  AND2_X1 U17084 ( .A1(n15409), .A2(n15353), .ZN(n15356) );
  OAI21_X1 U17085 ( .B1(n15356), .B2(n15355), .A(n15354), .ZN(n15358) );
  XNOR2_X1 U17086 ( .A(n15358), .B(n15357), .ZN(n15360) );
  AOI22_X1 U17087 ( .A1(n15360), .A2(n15754), .B1(n15746), .B2(n15359), .ZN(
        n15533) );
  INV_X1 U17088 ( .A(n15533), .ZN(n15362) );
  NOR2_X1 U17089 ( .A1(n15361), .A2(n15758), .ZN(n15530) );
  OAI21_X1 U17090 ( .B1(n15362), .B2(n15530), .A(n6544), .ZN(n15368) );
  AOI211_X1 U17091 ( .C1(n15531), .C2(n15377), .A(n15742), .B(n15363), .ZN(
        n15529) );
  AOI22_X1 U17092 ( .A1(n15764), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n15364), 
        .B2(n15760), .ZN(n15365) );
  OAI21_X1 U17093 ( .B1(n7824), .B2(n15418), .A(n15365), .ZN(n15366) );
  AOI21_X1 U17094 ( .B1(n15529), .B2(n15732), .A(n15366), .ZN(n15367) );
  OAI211_X1 U17095 ( .C1(n15534), .C2(n15423), .A(n15368), .B(n15367), .ZN(
        P1_U3276) );
  NAND2_X1 U17096 ( .A1(n15409), .A2(n15408), .ZN(n15407) );
  NAND2_X1 U17097 ( .A1(n15407), .A2(n15369), .ZN(n15389) );
  NAND2_X1 U17098 ( .A1(n15389), .A2(n15396), .ZN(n15388) );
  NAND2_X1 U17099 ( .A1(n15388), .A2(n15370), .ZN(n15371) );
  XNOR2_X1 U17100 ( .A(n15371), .B(n15376), .ZN(n15373) );
  AOI21_X1 U17101 ( .B1(n15373), .B2(n15754), .A(n15372), .ZN(n15539) );
  OAI21_X1 U17102 ( .B1(n15376), .B2(n15375), .A(n15374), .ZN(n15535) );
  INV_X1 U17103 ( .A(n15377), .ZN(n15378) );
  AOI211_X1 U17104 ( .C1(n15537), .C2(n15385), .A(n15742), .B(n15378), .ZN(
        n15536) );
  NAND2_X1 U17105 ( .A1(n15536), .A2(n15732), .ZN(n15381) );
  AOI22_X1 U17106 ( .A1(n15764), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n15379), 
        .B2(n15760), .ZN(n15380) );
  OAI211_X1 U17107 ( .C1(n7825), .C2(n15418), .A(n15381), .B(n15380), .ZN(
        n15382) );
  AOI21_X1 U17108 ( .B1(n15383), .B2(n15535), .A(n15382), .ZN(n15384) );
  OAI21_X1 U17109 ( .B1(n15539), .B2(n15764), .A(n15384), .ZN(P1_U3277) );
  INV_X1 U17110 ( .A(n15414), .ZN(n15387) );
  INV_X1 U17111 ( .A(n15385), .ZN(n15386) );
  AOI211_X1 U17112 ( .C1(n15543), .C2(n15387), .A(n15742), .B(n15386), .ZN(
        n15542) );
  OAI211_X1 U17113 ( .C1(n15389), .C2(n15396), .A(n15388), .B(n15754), .ZN(
        n15391) );
  NAND2_X1 U17114 ( .A1(n15391), .A2(n15390), .ZN(n15541) );
  AOI21_X1 U17115 ( .B1(n15542), .B2(n6539), .A(n15541), .ZN(n15401) );
  OAI22_X1 U17116 ( .A1(n6544), .A2(n15717), .B1(n15394), .B2(n15393), .ZN(
        n15399) );
  NOR2_X1 U17117 ( .A1(n15408), .A2(n15402), .ZN(n15403) );
  NOR2_X1 U17118 ( .A1(n15403), .A2(n15395), .ZN(n15397) );
  XNOR2_X1 U17119 ( .A(n15397), .B(n15396), .ZN(n15545) );
  NOR2_X1 U17120 ( .A1(n15545), .A2(n15423), .ZN(n15398) );
  AOI211_X1 U17121 ( .C1(n15730), .C2(n15543), .A(n15399), .B(n15398), .ZN(
        n15400) );
  OAI21_X1 U17122 ( .B1(n15401), .B2(n15764), .A(n15400), .ZN(P1_U3278) );
  INV_X1 U17123 ( .A(n15402), .ZN(n15406) );
  INV_X1 U17124 ( .A(n15403), .ZN(n15404) );
  OAI21_X1 U17125 ( .B1(n15406), .B2(n15405), .A(n15404), .ZN(n15551) );
  OAI211_X1 U17126 ( .C1(n15409), .C2(n15408), .A(n15754), .B(n15407), .ZN(
        n15550) );
  INV_X1 U17127 ( .A(n15550), .ZN(n15413) );
  OAI22_X1 U17128 ( .A1(n15412), .A2(n15411), .B1(n15758), .B2(n15410), .ZN(
        n15547) );
  OAI21_X1 U17129 ( .B1(n15413), .B2(n15547), .A(n6544), .ZN(n15422) );
  AOI211_X1 U17130 ( .C1(n15548), .C2(n15415), .A(n15742), .B(n15414), .ZN(
        n15546) );
  AOI22_X1 U17131 ( .A1(n15764), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n15416), 
        .B2(n15760), .ZN(n15417) );
  OAI21_X1 U17132 ( .B1(n15419), .B2(n15418), .A(n15417), .ZN(n15420) );
  AOI21_X1 U17133 ( .B1(n15546), .B2(n15732), .A(n15420), .ZN(n15421) );
  OAI211_X1 U17134 ( .C1(n15551), .C2(n15423), .A(n15422), .B(n15421), .ZN(
        P1_U3279) );
  XNOR2_X1 U17135 ( .A(n15424), .B(n15429), .ZN(n15437) );
  AOI22_X1 U17136 ( .A1(n15426), .A2(n15751), .B1(n15746), .B2(n15425), .ZN(
        n15432) );
  OAI21_X1 U17137 ( .B1(n15429), .B2(n15428), .A(n15427), .ZN(n15430) );
  NAND2_X1 U17138 ( .A1(n15430), .A2(n15754), .ZN(n15431) );
  OAI211_X1 U17139 ( .C1(n15437), .C2(n15433), .A(n15432), .B(n15431), .ZN(
        n15781) );
  MUX2_X1 U17140 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n15781), .S(n6544), .Z(
        n15434) );
  INV_X1 U17141 ( .A(n15434), .ZN(n15443) );
  OAI211_X1 U17142 ( .C1(n15739), .C2(n15780), .A(n10870), .B(n15435), .ZN(
        n15779) );
  INV_X1 U17143 ( .A(n15779), .ZN(n15436) );
  AOI22_X1 U17144 ( .A1(n15732), .A2(n15436), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n15760), .ZN(n15442) );
  INV_X1 U17145 ( .A(n15437), .ZN(n15783) );
  INV_X1 U17146 ( .A(n15438), .ZN(n15761) );
  NAND2_X1 U17147 ( .A1(n15783), .A2(n15761), .ZN(n15441) );
  NAND2_X1 U17148 ( .A1(n15730), .A2(n15439), .ZN(n15440) );
  NAND4_X1 U17149 ( .A1(n15443), .A2(n15442), .A3(n15441), .A4(n15440), .ZN(
        P1_U3291) );
  OAI211_X1 U17150 ( .C1(n15148), .C2(n15827), .A(n15444), .B(n15445), .ZN(
        n15563) );
  MUX2_X1 U17151 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15563), .S(n15850), .Z(
        P1_U3559) );
  OAI211_X1 U17152 ( .C1(n15447), .C2(n15827), .A(n15446), .B(n15445), .ZN(
        n15564) );
  MUX2_X1 U17153 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15564), .S(n15850), .Z(
        P1_U3558) );
  NAND2_X1 U17154 ( .A1(n15448), .A2(n15754), .ZN(n15457) );
  OAI211_X1 U17155 ( .C1(n15451), .C2(n15827), .A(n15450), .B(n15449), .ZN(
        n15452) );
  NAND3_X1 U17156 ( .A1(n15457), .A2(n15456), .A3(n15455), .ZN(n15565) );
  MUX2_X1 U17157 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n15565), .S(n15850), .Z(
        P1_U3557) );
  NAND3_X1 U17158 ( .A1(n15459), .A2(n15458), .A3(n15835), .ZN(n15467) );
  NAND2_X1 U17159 ( .A1(n15460), .A2(n15754), .ZN(n15466) );
  AOI21_X1 U17160 ( .B1(n15462), .B2(n15813), .A(n15461), .ZN(n15463) );
  MUX2_X1 U17161 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15566), .S(n15850), .Z(
        P1_U3556) );
  NAND2_X1 U17162 ( .A1(n15469), .A2(n15813), .ZN(n15471) );
  MUX2_X1 U17163 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15567), .S(n15850), .Z(
        P1_U3555) );
  NAND3_X1 U17164 ( .A1(n15474), .A2(n15835), .A3(n15473), .ZN(n15476) );
  NAND4_X1 U17165 ( .A1(n15478), .A2(n15477), .A3(n15476), .A4(n15475), .ZN(
        n15568) );
  MUX2_X1 U17166 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15568), .S(n15850), .Z(
        P1_U3554) );
  INV_X1 U17167 ( .A(n15479), .ZN(n15481) );
  AOI211_X1 U17168 ( .C1(n15813), .C2(n15482), .A(n15481), .B(n15480), .ZN(
        n15483) );
  OAI211_X1 U17169 ( .C1(n15801), .C2(n15485), .A(n15484), .B(n15483), .ZN(
        n15569) );
  MUX2_X1 U17170 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15569), .S(n15850), .Z(
        P1_U3553) );
  AOI211_X1 U17171 ( .C1(n15813), .C2(n15488), .A(n15487), .B(n15486), .ZN(
        n15489) );
  OAI21_X1 U17172 ( .B1(n15801), .B2(n15490), .A(n15489), .ZN(n15570) );
  MUX2_X1 U17173 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15570), .S(n15850), .Z(
        P1_U3552) );
  OAI211_X1 U17174 ( .C1(n15493), .C2(n15827), .A(n15492), .B(n15491), .ZN(
        n15494) );
  AOI21_X1 U17175 ( .B1(n15495), .B2(n15754), .A(n15494), .ZN(n15496) );
  OAI21_X1 U17176 ( .B1(n15801), .B2(n15497), .A(n15496), .ZN(n15571) );
  MUX2_X1 U17177 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15571), .S(n15850), .Z(
        P1_U3551) );
  AOI211_X1 U17178 ( .C1(n15813), .C2(n15500), .A(n15499), .B(n15498), .ZN(
        n15503) );
  NAND2_X1 U17179 ( .A1(n15501), .A2(n15835), .ZN(n15502) );
  OAI211_X1 U17180 ( .C1(n15504), .C2(n15829), .A(n15503), .B(n15502), .ZN(
        n15572) );
  MUX2_X1 U17181 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15572), .S(n15850), .Z(
        P1_U3550) );
  AOI211_X1 U17182 ( .C1(n15813), .C2(n15507), .A(n15506), .B(n15505), .ZN(
        n15508) );
  OAI21_X1 U17183 ( .B1(n15801), .B2(n15509), .A(n15508), .ZN(n15573) );
  MUX2_X1 U17184 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15573), .S(n15850), .Z(
        P1_U3549) );
  OAI211_X1 U17185 ( .C1(n15512), .C2(n15827), .A(n15511), .B(n15510), .ZN(
        n15513) );
  AOI21_X1 U17186 ( .B1(n15514), .B2(n15754), .A(n15513), .ZN(n15515) );
  OAI21_X1 U17187 ( .B1(n15801), .B2(n15516), .A(n15515), .ZN(n15574) );
  MUX2_X1 U17188 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15574), .S(n15850), .Z(
        P1_U3548) );
  AOI211_X1 U17189 ( .C1(n15813), .C2(n15519), .A(n15518), .B(n15517), .ZN(
        n15522) );
  NAND2_X1 U17190 ( .A1(n15520), .A2(n15835), .ZN(n15521) );
  OAI211_X1 U17191 ( .C1(n15523), .C2(n15829), .A(n15522), .B(n15521), .ZN(
        n15575) );
  MUX2_X1 U17192 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15575), .S(n15850), .Z(
        P1_U3547) );
  NOR3_X1 U17193 ( .A1(n15526), .A2(n15525), .A3(n15524), .ZN(n15527) );
  OAI21_X1 U17194 ( .B1(n15801), .B2(n15528), .A(n15527), .ZN(n15576) );
  MUX2_X1 U17195 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15576), .S(n15850), .Z(
        P1_U3546) );
  AOI211_X1 U17196 ( .C1(n15813), .C2(n15531), .A(n15530), .B(n15529), .ZN(
        n15532) );
  OAI211_X1 U17197 ( .C1(n15801), .C2(n15534), .A(n15533), .B(n15532), .ZN(
        n15577) );
  MUX2_X1 U17198 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15577), .S(n15850), .Z(
        P1_U3545) );
  INV_X1 U17199 ( .A(n15535), .ZN(n15540) );
  AOI21_X1 U17200 ( .B1(n15813), .B2(n15537), .A(n15536), .ZN(n15538) );
  OAI211_X1 U17201 ( .C1(n15801), .C2(n15540), .A(n15539), .B(n15538), .ZN(
        n15578) );
  MUX2_X1 U17202 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15578), .S(n15850), .Z(
        P1_U3544) );
  AOI211_X1 U17203 ( .C1(n15813), .C2(n15543), .A(n15542), .B(n15541), .ZN(
        n15544) );
  OAI21_X1 U17204 ( .B1(n15801), .B2(n15545), .A(n15544), .ZN(n15579) );
  MUX2_X1 U17205 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15579), .S(n15850), .Z(
        P1_U3543) );
  AOI211_X1 U17206 ( .C1(n15813), .C2(n15548), .A(n15547), .B(n15546), .ZN(
        n15549) );
  OAI211_X1 U17207 ( .C1(n15801), .C2(n15551), .A(n15550), .B(n15549), .ZN(
        n15580) );
  MUX2_X1 U17208 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15580), .S(n15850), .Z(
        P1_U3542) );
  AOI21_X1 U17209 ( .B1(n15813), .B2(n15553), .A(n15552), .ZN(n15554) );
  OAI211_X1 U17210 ( .C1(n15801), .C2(n15556), .A(n15555), .B(n15554), .ZN(
        n15581) );
  MUX2_X1 U17211 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n15581), .S(n15850), .Z(
        P1_U3541) );
  INV_X1 U17212 ( .A(n15557), .ZN(n15562) );
  AOI21_X1 U17213 ( .B1(n15813), .B2(n15559), .A(n15558), .ZN(n15560) );
  OAI211_X1 U17214 ( .C1(n15801), .C2(n15562), .A(n15561), .B(n15560), .ZN(
        n15582) );
  MUX2_X1 U17215 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n15582), .S(n15850), .Z(
        P1_U3539) );
  MUX2_X1 U17216 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15563), .S(n15838), .Z(
        P1_U3527) );
  MUX2_X1 U17217 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15564), .S(n15838), .Z(
        P1_U3526) );
  MUX2_X1 U17218 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n15565), .S(n15838), .Z(
        P1_U3525) );
  MUX2_X1 U17219 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n15566), .S(n15838), .Z(
        P1_U3524) );
  MUX2_X1 U17220 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15568), .S(n15838), .Z(
        P1_U3522) );
  MUX2_X1 U17221 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15569), .S(n15838), .Z(
        P1_U3521) );
  MUX2_X1 U17222 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15570), .S(n15838), .Z(
        P1_U3520) );
  MUX2_X1 U17223 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15571), .S(n15838), .Z(
        P1_U3519) );
  MUX2_X1 U17224 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15572), .S(n15838), .Z(
        P1_U3518) );
  MUX2_X1 U17225 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15573), .S(n15838), .Z(
        P1_U3517) );
  MUX2_X1 U17226 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15574), .S(n15838), .Z(
        P1_U3516) );
  MUX2_X1 U17227 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15575), .S(n15838), .Z(
        P1_U3515) );
  MUX2_X1 U17228 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15576), .S(n15838), .Z(
        P1_U3513) );
  MUX2_X1 U17229 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15577), .S(n15838), .Z(
        P1_U3510) );
  MUX2_X1 U17230 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15578), .S(n15838), .Z(
        P1_U3507) );
  MUX2_X1 U17231 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15579), .S(n15838), .Z(
        P1_U3504) );
  MUX2_X1 U17232 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15580), .S(n15838), .Z(
        P1_U3501) );
  MUX2_X1 U17233 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n15581), .S(n15838), .Z(
        P1_U3498) );
  MUX2_X1 U17234 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n15582), .S(n15838), .Z(
        P1_U3492) );
  INV_X1 U17235 ( .A(n15583), .ZN(n15590) );
  NOR4_X1 U17236 ( .A1(n15586), .A2(P1_IR_REG_30__SCAN_IN), .A3(n15585), .A4(
        P1_U3086), .ZN(n15587) );
  AOI21_X1 U17237 ( .B1(n15588), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n15587), 
        .ZN(n15589) );
  OAI21_X1 U17238 ( .B1(n15590), .B2(n15595), .A(n15589), .ZN(P1_U3324) );
  OAI222_X1 U17239 ( .A1(n15597), .A2(n15593), .B1(n15595), .B2(n15592), .C1(
        n15591), .C2(P1_U3086), .ZN(P1_U3326) );
  OAI222_X1 U17240 ( .A1(n15597), .A2(n15596), .B1(n15595), .B2(n15594), .C1(
        P1_U3086), .C2(n15674), .ZN(P1_U3328) );
  MUX2_X1 U17241 ( .A(n15599), .B(n15598), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  MUX2_X1 U17242 ( .A(n15600), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XOR2_X1 U17243 ( .A(n15602), .B(n15601), .Z(SUB_1596_U53) );
  XOR2_X1 U17244 ( .A(n15603), .B(n15604), .Z(SUB_1596_U59) );
  XOR2_X1 U17245 ( .A(n15605), .B(n15606), .Z(SUB_1596_U57) );
  XOR2_X1 U17246 ( .A(n15607), .B(n15608), .Z(SUB_1596_U56) );
  XOR2_X1 U17247 ( .A(n15609), .B(P2_ADDR_REG_8__SCAN_IN), .Z(SUB_1596_U55) );
  NAND2_X1 U17248 ( .A1(n15613), .A2(n15612), .ZN(n15616) );
  NAND2_X1 U17249 ( .A1(P3_ADDR_REG_14__SCAN_IN), .A2(n15614), .ZN(n15615) );
  NAND2_X1 U17250 ( .A1(n15616), .A2(n15615), .ZN(n15626) );
  XNOR2_X1 U17251 ( .A(P3_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n15625) );
  XNOR2_X1 U17252 ( .A(n15626), .B(n15625), .ZN(n15617) );
  INV_X1 U17253 ( .A(n15617), .ZN(n15618) );
  NAND2_X1 U17254 ( .A1(n15619), .A2(n15618), .ZN(n15623) );
  INV_X1 U17255 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15621) );
  OAI21_X1 U17256 ( .B1(n15622), .B2(n15621), .A(n15624), .ZN(SUB_1596_U65) );
  NAND2_X1 U17257 ( .A1(n15626), .A2(n15625), .ZN(n15629) );
  INV_X1 U17258 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15627) );
  NAND2_X1 U17259 ( .A1(n15627), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n15628) );
  NAND2_X1 U17260 ( .A1(n15629), .A2(n15628), .ZN(n15640) );
  XNOR2_X1 U17261 ( .A(n15636), .B(P1_ADDR_REG_16__SCAN_IN), .ZN(n15630) );
  XNOR2_X1 U17262 ( .A(n15640), .B(n15630), .ZN(n15631) );
  NAND2_X1 U17263 ( .A1(n15633), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n15634) );
  NAND2_X1 U17264 ( .A1(n15635), .A2(n15634), .ZN(SUB_1596_U64) );
  NAND2_X1 U17265 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n15636), .ZN(n15639) );
  INV_X1 U17266 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n15637) );
  AND2_X1 U17267 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n15637), .ZN(n15638) );
  AOI21_X1 U17268 ( .B1(n15640), .B2(n15639), .A(n15638), .ZN(n15649) );
  INV_X1 U17269 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n15641) );
  XNOR2_X1 U17270 ( .A(n15649), .B(n15641), .ZN(n15648) );
  XNOR2_X1 U17271 ( .A(n15648), .B(P3_ADDR_REG_17__SCAN_IN), .ZN(n15642) );
  INV_X1 U17272 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15646) );
  XNOR2_X1 U17273 ( .A(n15647), .B(n15646), .ZN(SUB_1596_U63) );
  INV_X1 U17274 ( .A(n15642), .ZN(n15643) );
  AND2_X1 U17275 ( .A1(n15644), .A2(n15643), .ZN(n15645) );
  NAND2_X1 U17276 ( .A1(n15648), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n15651) );
  OR2_X1 U17277 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n15649), .ZN(n15650) );
  NAND2_X1 U17278 ( .A1(n15651), .A2(n15650), .ZN(n15657) );
  XNOR2_X1 U17279 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n15652) );
  XNOR2_X1 U17280 ( .A(n15657), .B(n15652), .ZN(n15654) );
  INV_X1 U17281 ( .A(n15654), .ZN(n15653) );
  INV_X1 U17282 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n15656) );
  INV_X1 U17283 ( .A(n15657), .ZN(n15660) );
  INV_X1 U17284 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15658) );
  OR2_X1 U17285 ( .A1(n15658), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n15659) );
  AOI22_X1 U17286 ( .A1(n15660), .A2(n15659), .B1(P1_ADDR_REG_18__SCAN_IN), 
        .B2(n15658), .ZN(n15664) );
  XNOR2_X1 U17287 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n15662) );
  XNOR2_X1 U17288 ( .A(n15661), .B(n15662), .ZN(n15663) );
  XNOR2_X1 U17289 ( .A(n15664), .B(n15663), .ZN(n15665) );
  AOI21_X1 U17290 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15666) );
  OAI21_X1 U17291 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n15666), 
        .ZN(U28) );
  AOI21_X1 U17292 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n15667) );
  OAI21_X1 U17293 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n15667), 
        .ZN(U29) );
  AND2_X1 U17294 ( .A1(n15669), .A2(n15668), .ZN(n15671) );
  XNOR2_X1 U17295 ( .A(n15671), .B(n15670), .ZN(SUB_1596_U61) );
  INV_X1 U17296 ( .A(n15672), .ZN(n15679) );
  NAND2_X1 U17297 ( .A1(n15674), .A2(n15673), .ZN(n15677) );
  NAND2_X1 U17298 ( .A1(n15675), .A2(n15677), .ZN(n15676) );
  MUX2_X1 U17299 ( .A(n15677), .B(n15676), .S(P1_IR_REG_0__SCAN_IN), .Z(n15678) );
  NAND2_X1 U17300 ( .A1(n15679), .A2(n15678), .ZN(n15682) );
  AOI22_X1 U17301 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n15680), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n15681) );
  OAI21_X1 U17302 ( .B1(n15683), .B2(n15682), .A(n15681), .ZN(P1_U3243) );
  MUX2_X1 U17303 ( .A(n11514), .B(P1_REG2_REG_4__SCAN_IN), .S(n15684), .Z(
        n15685) );
  NAND3_X1 U17304 ( .A1(n15687), .A2(n15686), .A3(n15685), .ZN(n15688) );
  NAND3_X1 U17305 ( .A1(n15724), .A2(n15689), .A3(n15688), .ZN(n15697) );
  INV_X1 U17306 ( .A(n15690), .ZN(n15693) );
  NAND3_X1 U17307 ( .A1(n15693), .A2(n15692), .A3(n15691), .ZN(n15694) );
  NAND3_X1 U17308 ( .A1(n15723), .A2(n15695), .A3(n15694), .ZN(n15696) );
  OAI211_X1 U17309 ( .C1(n15699), .C2(n15698), .A(n15697), .B(n15696), .ZN(
        n15700) );
  NOR2_X1 U17310 ( .A1(n15701), .A2(n15700), .ZN(n15703) );
  NAND2_X1 U17311 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n15702) );
  OAI211_X1 U17312 ( .C1(n15728), .C2(n15704), .A(n15703), .B(n15702), .ZN(
        P1_U3247) );
  OAI21_X1 U17313 ( .B1(n15707), .B2(n15706), .A(n15705), .ZN(n15712) );
  XNOR2_X1 U17314 ( .A(n15709), .B(n15708), .ZN(n15711) );
  AOI222_X1 U17315 ( .A1(n15712), .A2(n15724), .B1(n15723), .B2(n15711), .C1(
        n15710), .C2(n15720), .ZN(n15714) );
  OAI211_X1 U17316 ( .C1(n15715), .C2(n15728), .A(n15714), .B(n15713), .ZN(
        P1_U3255) );
  OAI21_X1 U17317 ( .B1(n15718), .B2(n15717), .A(n15716), .ZN(n15725) );
  XNOR2_X1 U17318 ( .A(n15719), .B(P1_REG1_REG_15__SCAN_IN), .ZN(n15722) );
  AOI222_X1 U17319 ( .A1(n15725), .A2(n15724), .B1(n15723), .B2(n15722), .C1(
        n15721), .C2(n15720), .ZN(n15727) );
  OAI211_X1 U17320 ( .C1(n15627), .C2(n15728), .A(n15727), .B(n15726), .ZN(
        P1_U3258) );
  AOI222_X1 U17321 ( .A1(n15731), .A2(n15730), .B1(P1_REG2_REG_6__SCAN_IN), 
        .B2(n15764), .C1(n15760), .C2(n15729), .ZN(n15736) );
  AOI22_X1 U17322 ( .A1(n15734), .A2(n15761), .B1(n15733), .B2(n15732), .ZN(
        n15735) );
  OAI211_X1 U17323 ( .C1(n15764), .C2(n15737), .A(n15736), .B(n15735), .ZN(
        P1_U3287) );
  XNOR2_X1 U17324 ( .A(n15750), .B(n15738), .ZN(n15777) );
  INV_X1 U17325 ( .A(n15739), .ZN(n15741) );
  NAND2_X1 U17326 ( .A1(n15744), .A2(n8869), .ZN(n15740) );
  NAND2_X1 U17327 ( .A1(n15741), .A2(n15740), .ZN(n15752) );
  OR2_X1 U17328 ( .A1(n15752), .A2(n15742), .ZN(n15774) );
  NAND2_X1 U17329 ( .A1(n15744), .A2(n15743), .ZN(n15747) );
  NAND2_X1 U17330 ( .A1(n15746), .A2(n15745), .ZN(n15772) );
  OAI211_X1 U17331 ( .C1(n15774), .C2(n15748), .A(n15747), .B(n15772), .ZN(
        n15759) );
  OAI21_X1 U17332 ( .B1(n15750), .B2(n15749), .A(n15754), .ZN(n15757) );
  XNOR2_X1 U17333 ( .A(n15752), .B(n15751), .ZN(n15755) );
  AOI21_X1 U17334 ( .B1(n15755), .B2(n15754), .A(n15753), .ZN(n15756) );
  AOI21_X1 U17335 ( .B1(n15758), .B2(n15757), .A(n15756), .ZN(n15775) );
  AOI211_X1 U17336 ( .C1(n15792), .C2(n15777), .A(n15759), .B(n15775), .ZN(
        n15763) );
  AOI22_X1 U17337 ( .A1(n15761), .A2(n15777), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n15760), .ZN(n15762) );
  OAI221_X1 U17338 ( .B1(n15764), .B2(n15763), .C1(n6544), .C2(n10679), .A(
        n15762), .ZN(P1_U3292) );
  NOR2_X1 U17339 ( .A1(n15770), .A2(n15765), .ZN(P1_U3294) );
  AND2_X1 U17340 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15771), .ZN(P1_U3295) );
  AND2_X1 U17341 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15771), .ZN(P1_U3296) );
  AND2_X1 U17342 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15771), .ZN(P1_U3297) );
  NOR2_X1 U17343 ( .A1(n15770), .A2(n15766), .ZN(P1_U3298) );
  AND2_X1 U17344 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15771), .ZN(P1_U3299) );
  AND2_X1 U17345 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15771), .ZN(P1_U3300) );
  AND2_X1 U17346 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15771), .ZN(P1_U3301) );
  AND2_X1 U17347 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15771), .ZN(P1_U3302) );
  AND2_X1 U17348 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15771), .ZN(P1_U3303) );
  NOR2_X1 U17349 ( .A1(n15770), .A2(n15767), .ZN(P1_U3304) );
  AND2_X1 U17350 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15771), .ZN(P1_U3305) );
  AND2_X1 U17351 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15771), .ZN(P1_U3306) );
  AND2_X1 U17352 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15771), .ZN(P1_U3307) );
  AND2_X1 U17353 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15771), .ZN(P1_U3308) );
  AND2_X1 U17354 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15771), .ZN(P1_U3309) );
  AND2_X1 U17355 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15771), .ZN(P1_U3310) );
  AND2_X1 U17356 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15771), .ZN(P1_U3311) );
  AND2_X1 U17357 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15771), .ZN(P1_U3312) );
  AND2_X1 U17358 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15771), .ZN(P1_U3313) );
  AND2_X1 U17359 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15771), .ZN(P1_U3314) );
  AND2_X1 U17360 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15771), .ZN(P1_U3315) );
  AND2_X1 U17361 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15771), .ZN(P1_U3316) );
  NOR2_X1 U17362 ( .A1(n15770), .A2(n15768), .ZN(P1_U3317) );
  AND2_X1 U17363 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15771), .ZN(P1_U3318) );
  AND2_X1 U17364 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15771), .ZN(P1_U3319) );
  NOR2_X1 U17365 ( .A1(n15770), .A2(n15769), .ZN(P1_U3320) );
  AND2_X1 U17366 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15771), .ZN(P1_U3321) );
  AND2_X1 U17367 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15771), .ZN(P1_U3322) );
  AND2_X1 U17368 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15771), .ZN(P1_U3323) );
  NAND3_X1 U17369 ( .A1(n15774), .A2(n15773), .A3(n15772), .ZN(n15776) );
  AOI211_X1 U17370 ( .C1(n15835), .C2(n15777), .A(n15776), .B(n15775), .ZN(
        n15839) );
  INV_X1 U17371 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n15778) );
  AOI22_X1 U17372 ( .A1(n15838), .A2(n15839), .B1(n15778), .B2(n15836), .ZN(
        P1_U3462) );
  OAI21_X1 U17373 ( .B1(n15780), .B2(n15827), .A(n15779), .ZN(n15782) );
  AOI211_X1 U17374 ( .C1(n7453), .C2(n15783), .A(n15782), .B(n15781), .ZN(
        n15841) );
  INV_X1 U17375 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n15784) );
  AOI22_X1 U17376 ( .A1(n15838), .A2(n15841), .B1(n15784), .B2(n15836), .ZN(
        P1_U3465) );
  INV_X1 U17377 ( .A(n15788), .ZN(n15791) );
  AOI21_X1 U17378 ( .B1(n15813), .B2(n15786), .A(n15785), .ZN(n15787) );
  OAI21_X1 U17379 ( .B1(n15788), .B2(n15815), .A(n15787), .ZN(n15789) );
  AOI211_X1 U17380 ( .C1(n15792), .C2(n15791), .A(n15790), .B(n15789), .ZN(
        n15843) );
  INV_X1 U17381 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n15793) );
  AOI22_X1 U17382 ( .A1(n15838), .A2(n15843), .B1(n15793), .B2(n15836), .ZN(
        P1_U3468) );
  INV_X1 U17383 ( .A(n15794), .ZN(n15796) );
  OAI211_X1 U17384 ( .C1(n15801), .C2(n15797), .A(n15796), .B(n15795), .ZN(
        n15799) );
  NOR2_X1 U17385 ( .A1(n15799), .A2(n15798), .ZN(n15844) );
  INV_X1 U17386 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n15800) );
  AOI22_X1 U17387 ( .A1(n15838), .A2(n15844), .B1(n15800), .B2(n15836), .ZN(
        P1_U3471) );
  NOR2_X1 U17388 ( .A1(n15802), .A2(n15801), .ZN(n15809) );
  INV_X1 U17389 ( .A(n15803), .ZN(n15805) );
  NAND2_X1 U17390 ( .A1(n15805), .A2(n15804), .ZN(n15806) );
  NOR4_X1 U17391 ( .A1(n15809), .A2(n15808), .A3(n15807), .A4(n15806), .ZN(
        n15845) );
  INV_X1 U17392 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15810) );
  AOI22_X1 U17393 ( .A1(n15838), .A2(n15845), .B1(n15810), .B2(n15836), .ZN(
        P1_U3474) );
  AOI21_X1 U17394 ( .B1(n15813), .B2(n15812), .A(n15811), .ZN(n15814) );
  OAI21_X1 U17395 ( .B1(n15816), .B2(n15815), .A(n15814), .ZN(n15817) );
  NOR2_X1 U17396 ( .A1(n15818), .A2(n15817), .ZN(n15846) );
  INV_X1 U17397 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15819) );
  AOI22_X1 U17398 ( .A1(n15838), .A2(n15846), .B1(n15819), .B2(n15836), .ZN(
        P1_U3480) );
  OAI21_X1 U17399 ( .B1(n15821), .B2(n15827), .A(n15820), .ZN(n15823) );
  AOI211_X1 U17400 ( .C1(n15835), .C2(n15824), .A(n15823), .B(n15822), .ZN(
        n15847) );
  AOI22_X1 U17401 ( .A1(n15838), .A2(n15847), .B1(n15825), .B2(n15836), .ZN(
        P1_U3483) );
  OAI21_X1 U17402 ( .B1(n15828), .B2(n15827), .A(n15826), .ZN(n15833) );
  NOR3_X1 U17403 ( .A1(n15831), .A2(n15830), .A3(n15829), .ZN(n15832) );
  AOI211_X1 U17404 ( .C1(n15835), .C2(n15834), .A(n15833), .B(n15832), .ZN(
        n15849) );
  INV_X1 U17405 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n15837) );
  AOI22_X1 U17406 ( .A1(n15838), .A2(n15849), .B1(n15837), .B2(n15836), .ZN(
        P1_U3489) );
  AOI22_X1 U17407 ( .A1(n15850), .A2(n15839), .B1(n8862), .B2(n15848), .ZN(
        P1_U3529) );
  AOI22_X1 U17408 ( .A1(n15850), .A2(n15841), .B1(n15840), .B2(n15848), .ZN(
        P1_U3530) );
  AOI22_X1 U17409 ( .A1(n15850), .A2(n15843), .B1(n15842), .B2(n15848), .ZN(
        P1_U3531) );
  AOI22_X1 U17410 ( .A1(n15850), .A2(n15844), .B1(n10668), .B2(n15848), .ZN(
        P1_U3532) );
  AOI22_X1 U17411 ( .A1(n15850), .A2(n15845), .B1(n10669), .B2(n15848), .ZN(
        P1_U3533) );
  AOI22_X1 U17412 ( .A1(n15850), .A2(n15846), .B1(n10671), .B2(n15848), .ZN(
        P1_U3535) );
  AOI22_X1 U17413 ( .A1(n15850), .A2(n15847), .B1(n10746), .B2(n15848), .ZN(
        P1_U3536) );
  AOI22_X1 U17414 ( .A1(n15850), .A2(n15849), .B1(n11070), .B2(n15848), .ZN(
        P1_U3538) );
  NOR2_X1 U17415 ( .A1(n15851), .A2(P2_U3947), .ZN(P2_U3087) );
  OAI21_X1 U17416 ( .B1(n15854), .B2(n15853), .A(n15852), .ZN(n15859) );
  NAND2_X1 U17417 ( .A1(n15894), .A2(n15855), .ZN(n15858) );
  OR2_X1 U17418 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15856), .ZN(n15857) );
  OAI211_X1 U17419 ( .C1(n15873), .C2(n15859), .A(n15858), .B(n15857), .ZN(
        n15860) );
  INV_X1 U17420 ( .A(n15860), .ZN(n15865) );
  OAI211_X1 U17421 ( .C1(n15863), .C2(n15862), .A(n15892), .B(n15861), .ZN(
        n15864) );
  OAI211_X1 U17422 ( .C1(n15900), .C2(n16027), .A(n15865), .B(n15864), .ZN(
        P2_U3217) );
  OAI21_X1 U17423 ( .B1(n15868), .B2(n15867), .A(n15866), .ZN(n15872) );
  NAND2_X1 U17424 ( .A1(n15894), .A2(n15869), .ZN(n15871) );
  OAI211_X1 U17425 ( .C1(n15873), .C2(n15872), .A(n15871), .B(n15870), .ZN(
        n15874) );
  INV_X1 U17426 ( .A(n15874), .ZN(n15879) );
  OAI211_X1 U17427 ( .C1(n15877), .C2(n15876), .A(n15892), .B(n15875), .ZN(
        n15878) );
  OAI211_X1 U17428 ( .C1(n15900), .C2(n15880), .A(n15879), .B(n15878), .ZN(
        P2_U3219) );
  AND2_X1 U17429 ( .A1(n15882), .A2(n15881), .ZN(n15885) );
  OAI21_X1 U17430 ( .B1(n15885), .B2(n15884), .A(n15883), .ZN(n15897) );
  INV_X1 U17431 ( .A(n15886), .ZN(n15888) );
  NAND3_X1 U17432 ( .A1(n15889), .A2(n15888), .A3(n15887), .ZN(n15890) );
  NAND2_X1 U17433 ( .A1(n15891), .A2(n15890), .ZN(n15893) );
  AOI222_X1 U17434 ( .A1(n15897), .A2(n15896), .B1(n15895), .B2(n15894), .C1(
        n15893), .C2(n15892), .ZN(n15899) );
  OAI211_X1 U17435 ( .C1(n15901), .C2(n15900), .A(n15899), .B(n15898), .ZN(
        P2_U3226) );
  NOR2_X1 U17436 ( .A1(n15911), .A2(n15902), .ZN(n15907) );
  AND2_X1 U17437 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15908), .ZN(P2_U3266) );
  AND2_X1 U17438 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15908), .ZN(P2_U3267) );
  AND2_X1 U17439 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15908), .ZN(P2_U3268) );
  AND2_X1 U17440 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15908), .ZN(P2_U3269) );
  AND2_X1 U17441 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15908), .ZN(P2_U3270) );
  AND2_X1 U17442 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15908), .ZN(P2_U3271) );
  AND2_X1 U17443 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15908), .ZN(P2_U3272) );
  AND2_X1 U17444 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15908), .ZN(P2_U3273) );
  NOR2_X1 U17445 ( .A1(n15907), .A2(n15903), .ZN(P2_U3274) );
  AND2_X1 U17446 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15908), .ZN(P2_U3275) );
  NOR2_X1 U17447 ( .A1(n15907), .A2(n15904), .ZN(P2_U3276) );
  AND2_X1 U17448 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15908), .ZN(P2_U3277) );
  AND2_X1 U17449 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15908), .ZN(P2_U3278) );
  AND2_X1 U17450 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15908), .ZN(P2_U3279) );
  AND2_X1 U17451 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15908), .ZN(P2_U3280) );
  AND2_X1 U17452 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15908), .ZN(P2_U3281) );
  AND2_X1 U17453 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15908), .ZN(P2_U3282) );
  AND2_X1 U17454 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15908), .ZN(P2_U3283) );
  AND2_X1 U17455 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15908), .ZN(P2_U3284) );
  AND2_X1 U17456 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15908), .ZN(P2_U3285) );
  NOR2_X1 U17457 ( .A1(n15907), .A2(n15905), .ZN(P2_U3286) );
  AND2_X1 U17458 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15908), .ZN(P2_U3287) );
  AND2_X1 U17459 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15908), .ZN(P2_U3288) );
  AND2_X1 U17460 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15908), .ZN(P2_U3289) );
  AND2_X1 U17461 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15908), .ZN(P2_U3290) );
  AND2_X1 U17462 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15908), .ZN(P2_U3291) );
  NOR2_X1 U17463 ( .A1(n15907), .A2(n15906), .ZN(P2_U3292) );
  AND2_X1 U17464 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15908), .ZN(P2_U3293) );
  AND2_X1 U17465 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15908), .ZN(P2_U3294) );
  AND2_X1 U17466 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15908), .ZN(P2_U3295) );
  AOI22_X1 U17467 ( .A1(n15914), .A2(n15910), .B1(n15909), .B2(n15911), .ZN(
        P2_U3416) );
  AOI22_X1 U17468 ( .A1(n15914), .A2(n15913), .B1(n15912), .B2(n15911), .ZN(
        P2_U3417) );
  INV_X1 U17469 ( .A(n15915), .ZN(n15916) );
  OAI21_X1 U17470 ( .B1(n15917), .B2(n15931), .A(n15916), .ZN(n15920) );
  INV_X1 U17471 ( .A(n15918), .ZN(n15919) );
  AOI211_X1 U17472 ( .C1(n15937), .C2(n15921), .A(n15920), .B(n15919), .ZN(
        n15939) );
  INV_X1 U17473 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15922) );
  AOI22_X1 U17474 ( .A1(n14818), .A2(n15939), .B1(n15922), .B2(n15938), .ZN(
        P2_U3436) );
  OAI21_X1 U17475 ( .B1(n15924), .B2(n15931), .A(n15923), .ZN(n15927) );
  INV_X1 U17476 ( .A(n15925), .ZN(n15926) );
  AOI211_X1 U17477 ( .C1(n15929), .C2(n15928), .A(n15927), .B(n15926), .ZN(
        n15940) );
  AOI22_X1 U17478 ( .A1(n14818), .A2(n15940), .B1(n9528), .B2(n15938), .ZN(
        P2_U3442) );
  OAI21_X1 U17479 ( .B1(n15932), .B2(n15931), .A(n15930), .ZN(n15935) );
  INV_X1 U17480 ( .A(n15933), .ZN(n15934) );
  AOI211_X1 U17481 ( .C1(n15937), .C2(n15936), .A(n15935), .B(n15934), .ZN(
        n15943) );
  AOI22_X1 U17482 ( .A1(n14818), .A2(n15943), .B1(n9557), .B2(n15938), .ZN(
        P2_U3448) );
  AOI22_X1 U17483 ( .A1(n15944), .A2(n15939), .B1(n9502), .B2(n15941), .ZN(
        P2_U3501) );
  AOI22_X1 U17484 ( .A1(n15944), .A2(n15940), .B1(n9529), .B2(n15941), .ZN(
        P2_U3503) );
  AOI22_X1 U17485 ( .A1(n15944), .A2(n15943), .B1(n15942), .B2(n15941), .ZN(
        P2_U3505) );
  NOR2_X1 U17486 ( .A1(P3_U3897), .A2(n15945), .ZN(P3_U3150) );
  AOI21_X1 U17487 ( .B1(n15947), .B2(n15994), .A(n15946), .ZN(n15948) );
  INV_X1 U17488 ( .A(n15948), .ZN(n15951) );
  AOI222_X1 U17489 ( .A1(n15951), .A2(n15995), .B1(n15950), .B2(n15958), .C1(
        n15949), .C2(n15977), .ZN(n15952) );
  OAI21_X1 U17490 ( .B1(n15995), .B2(n7586), .A(n15952), .ZN(P3_U3226) );
  INV_X1 U17491 ( .A(n15953), .ZN(n15955) );
  OAI21_X1 U17492 ( .B1(n15956), .B2(n15955), .A(n15954), .ZN(n15960) );
  AOI222_X1 U17493 ( .A1(n15995), .A2(n15960), .B1(n15959), .B2(n15958), .C1(
        n15957), .C2(n15977), .ZN(n15961) );
  OAI21_X1 U17494 ( .B1(n15995), .B2(n15962), .A(n15961), .ZN(P3_U3227) );
  XNOR2_X1 U17495 ( .A(n15965), .B(n15963), .ZN(n15971) );
  OAI21_X1 U17496 ( .B1(n15966), .B2(n15965), .A(n15964), .ZN(n16004) );
  OAI22_X1 U17497 ( .A1(n10860), .A2(n15990), .B1(n15967), .B2(n15992), .ZN(
        n15968) );
  AOI21_X1 U17498 ( .B1(n16004), .B2(n15969), .A(n15968), .ZN(n15970) );
  OAI21_X1 U17499 ( .B1(n15971), .B2(n15988), .A(n15970), .ZN(n16002) );
  INV_X1 U17500 ( .A(n16004), .ZN(n15975) );
  NOR2_X1 U17501 ( .A1(n15972), .A2(n15981), .ZN(n16003) );
  INV_X1 U17502 ( .A(n16003), .ZN(n15973) );
  OAI22_X1 U17503 ( .A1(n15975), .A2(n15974), .B1(n15983), .B2(n15973), .ZN(
        n15976) );
  AOI211_X1 U17504 ( .C1(n15977), .C2(P3_REG3_REG_2__SCAN_IN), .A(n16002), .B(
        n15976), .ZN(n15978) );
  AOI22_X1 U17505 ( .A1(n15997), .A2(n15979), .B1(n15978), .B2(n15995), .ZN(
        P3_U3231) );
  XNOR2_X1 U17506 ( .A(n15980), .B(n10905), .ZN(n16000) );
  NOR2_X1 U17507 ( .A1(n15982), .A2(n15981), .ZN(n15999) );
  INV_X1 U17508 ( .A(n15999), .ZN(n15984) );
  OAI22_X1 U17509 ( .A1(n15985), .A2(n10057), .B1(n15984), .B2(n15983), .ZN(
        n15993) );
  XNOR2_X1 U17510 ( .A(n10905), .B(n15986), .ZN(n15987) );
  OAI222_X1 U17511 ( .A1(n15992), .A2(n15991), .B1(n15990), .B2(n15989), .C1(
        n15988), .C2(n15987), .ZN(n15998) );
  AOI211_X1 U17512 ( .C1(n15994), .C2(n16000), .A(n15993), .B(n15998), .ZN(
        n15996) );
  AOI22_X1 U17513 ( .A1(n15997), .A2(n7338), .B1(n15996), .B2(n15995), .ZN(
        P3_U3232) );
  INV_X1 U17514 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n16001) );
  AOI211_X1 U17515 ( .C1(n16007), .C2(n16000), .A(n15999), .B(n15998), .ZN(
        n16019) );
  AOI22_X1 U17516 ( .A1(n16018), .A2(n16001), .B1(n16019), .B2(n16017), .ZN(
        P3_U3393) );
  INV_X1 U17517 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n16005) );
  AOI211_X1 U17518 ( .C1(n16013), .C2(n16004), .A(n16003), .B(n16002), .ZN(
        n16020) );
  AOI22_X1 U17519 ( .A1(n16018), .A2(n16005), .B1(n16020), .B2(n16017), .ZN(
        P3_U3396) );
  AOI22_X1 U17520 ( .A1(n16008), .A2(n16007), .B1(n16006), .B2(n16011), .ZN(
        n16009) );
  AND2_X1 U17521 ( .A1(n16010), .A2(n16009), .ZN(n16022) );
  AOI22_X1 U17522 ( .A1(n16018), .A2(n8210), .B1(n16022), .B2(n16017), .ZN(
        P3_U3402) );
  AOI22_X1 U17523 ( .A1(n16014), .A2(n16013), .B1(n16012), .B2(n16011), .ZN(
        n16015) );
  AND2_X1 U17524 ( .A1(n16016), .A2(n16015), .ZN(n16024) );
  AOI22_X1 U17525 ( .A1(n16018), .A2(n8145), .B1(n16024), .B2(n16017), .ZN(
        P3_U3405) );
  AOI22_X1 U17526 ( .A1(n13911), .A2(n16019), .B1(n7337), .B2(n16023), .ZN(
        P3_U3460) );
  AOI22_X1 U17527 ( .A1(n13911), .A2(n16020), .B1(n11143), .B2(n16023), .ZN(
        P3_U3461) );
  AOI22_X1 U17528 ( .A1(n13911), .A2(n16022), .B1(n16021), .B2(n16023), .ZN(
        P3_U3463) );
  AOI22_X1 U17529 ( .A1(n13911), .A2(n16024), .B1(n11200), .B2(n16023), .ZN(
        P3_U3464) );
  AND2_X1 U17530 ( .A1(n16026), .A2(n16025), .ZN(n16028) );
  XNOR2_X1 U17531 ( .A(n16028), .B(n16027), .ZN(SUB_1596_U60) );
  XOR2_X1 U17532 ( .A(n16030), .B(n16029), .Z(SUB_1596_U5) );
  NAND2_X1 U12243 ( .A1(n9697), .A2(n9696), .ZN(n14580) );
  AND2_X1 U7290 ( .A1(n6575), .A2(n7413), .ZN(n7526) );
  CLKBUF_X1 U7301 ( .A(n8174), .Z(n6551) );
  CLKBUF_X1 U7318 ( .A(n8615), .Z(n6541) );
  INV_X1 U7330 ( .A(n15419), .ZN(n15548) );
  CLKBUF_X1 U7332 ( .A(n13146), .Z(n6543) );
  NAND2_X1 U7333 ( .A1(n9783), .A2(n9782), .ZN(n14700) );
  NAND2_X1 U7347 ( .A1(n9738), .A2(n9737), .ZN(n14491) );
  NAND2_X1 U7351 ( .A1(n9213), .A2(n9212), .ZN(n15507) );
  CLKBUF_X1 U7352 ( .A(n8843), .Z(n10642) );
  OR2_X1 U7353 ( .A1(n8989), .A2(n8988), .ZN(n9013) );
  CLKBUF_X3 U7360 ( .A(n8615), .Z(n6542) );
  INV_X1 U7380 ( .A(n10860), .ZN(n8170) );
  AND2_X1 U8263 ( .A1(n9720), .A2(n9719), .ZN(n14552) );
  CLKBUF_X1 U9357 ( .A(n15392), .Z(n6539) );
  AND2_X1 U9982 ( .A1(n7945), .A2(n7946), .ZN(n16036) );
  INV_X1 U10307 ( .A(n8615), .ZN(n8069) );
endmodule

