

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881;

  INV_X2 U2375 ( .A(n3994), .ZN(U4043) );
  NAND2_X1 U2376 ( .A1(n4470), .A2(n2408), .ZN(n4022) );
  XOR2_X1 U2377 ( .A(n2390), .B(n3237), .Z(n4434) );
  NOR2_X1 U2378 ( .A1(n2851), .A2(n2850), .ZN(n2849) );
  AOI21_X1 U2379 ( .B1(n2382), .B2(n4387), .A(n2726), .ZN(n2851) );
  NAND2_X1 U2380 ( .A1(n2556), .A2(n2366), .ZN(n2369) );
  INV_X1 U2381 ( .A(n2784), .ZN(n3837) );
  NAND2_X1 U2382 ( .A1(n2356), .A2(n2355), .ZN(n2359) );
  NAND2_X1 U2384 ( .A1(n2349), .A2(n2348), .ZN(n2354) );
  INV_X1 U2385 ( .A(n2805), .ZN(n3725) );
  NAND2_X1 U2386 ( .A1(n3996), .A2(n2345), .ZN(n4010) );
  AND2_X1 U2387 ( .A1(n2194), .A2(n2192), .ZN(n2151) );
  BUF_X1 U2388 ( .A(IR_REG_0__SCAN_IN), .Z(n4603) );
  AOI21_X2 U2389 ( .B1(n3425), .B2(REG1_REG_18__SCAN_IN), .A(n4479), .ZN(n2415) );
  NOR2_X2 U2390 ( .A1(n4453), .A2(n2210), .ZN(n2407) );
  NOR2_X2 U2391 ( .A1(n2391), .A2(n4433), .ZN(n3403) );
  NOR2_X1 U2392 ( .A1(n4444), .A2(n4766), .ZN(n4443) );
  XNOR2_X1 U2393 ( .A(n2400), .B(n2399), .ZN(n4444) );
  NOR2_X2 U2394 ( .A1(n2849), .A2(n2135), .ZN(n2386) );
  NAND4_X1 U2395 ( .A1(n2665), .A2(n2664), .A3(n2663), .A4(n2662), .ZN(n2688)
         );
  AND2_X1 U2396 ( .A1(n2585), .A2(n2584), .ZN(n2681) );
  NAND4_X2 U2397 ( .A1(n2684), .A2(n2685), .A3(n2683), .A4(n2687), .ZN(n2762)
         );
  NAND2_X2 U2399 ( .A1(n2700), .A2(n3556), .ZN(n2741) );
  INV_X1 U2400 ( .A(n4208), .ZN(n2981) );
  BUF_X2 U2401 ( .A(n2680), .Z(n3489) );
  INV_X1 U2402 ( .A(n2584), .ZN(n2586) );
  INV_X1 U2404 ( .A(IR_REG_23__SCAN_IN), .ZN(n4692) );
  MUX2_X1 U2405 ( .A(n4772), .B(n4344), .S(n4577), .Z(n4246) );
  MUX2_X1 U2406 ( .A(n4345), .B(n4344), .S(n4565), .Z(n4349) );
  NAND2_X1 U2407 ( .A1(n3942), .A2(n3946), .ZN(n3917) );
  AOI21_X1 U2408 ( .B1(n3776), .B2(n3775), .A(n3774), .ZN(n3777) );
  NAND2_X1 U2409 ( .A1(n3649), .A2(n3648), .ZN(n3651) );
  NAND2_X1 U2410 ( .A1(n2280), .A2(n2281), .ZN(n3674) );
  OR2_X1 U2411 ( .A1(n3379), .A2(n3528), .ZN(n3649) );
  AOI21_X1 U2412 ( .B1(n3318), .B2(n3317), .A(n3316), .ZN(n3354) );
  OAI21_X1 U2413 ( .B1(n3101), .B2(n3029), .A(n3579), .ZN(n3069) );
  AND3_X2 U2414 ( .A1(n2205), .A2(n2204), .A3(n2164), .ZN(n2390) );
  NAND2_X1 U2415 ( .A1(n2172), .A2(n3569), .ZN(n3101) );
  INV_X2 U2416 ( .A(n4505), .ZN(n4396) );
  NAND3_X2 U2417 ( .A1(n2796), .A2(n3629), .A3(n4382), .ZN(n3949) );
  AOI21_X1 U2418 ( .B1(n3570), .B2(n3025), .A(n2140), .ZN(n2223) );
  AND2_X1 U2419 ( .A1(n2865), .A2(n2864), .ZN(n2868) );
  CLKBUF_X3 U2420 ( .A(n2784), .Z(n3825) );
  AND2_X2 U2421 ( .A1(n3843), .A2(n4551), .ZN(n3830) );
  AND2_X2 U2422 ( .A1(n2741), .A2(n2740), .ZN(n3843) );
  NAND4_X1 U2423 ( .A1(n2636), .A2(n2635), .A3(n2634), .A4(n2633), .ZN(n4208)
         );
  INV_X4 U2424 ( .A(n2679), .ZN(n3488) );
  NAND2_X1 U2425 ( .A1(n2514), .A2(n2517), .ZN(n2584) );
  XNOR2_X1 U2426 ( .A(n2518), .B(n3884), .ZN(n2585) );
  NAND2_X1 U2427 ( .A1(n2171), .A2(n2512), .ZN(n2514) );
  NAND2_X1 U2428 ( .A1(n2517), .A2(n2522), .ZN(n2518) );
  NOR2_X1 U2429 ( .A1(n2149), .A2(n2481), .ZN(n2270) );
  OR2_X1 U2430 ( .A1(n2480), .A2(n2479), .ZN(n2481) );
  AND2_X1 U2431 ( .A1(n2229), .A2(n2420), .ZN(n2183) );
  INV_X1 U2432 ( .A(n2333), .ZN(n2134) );
  AND4_X1 U2433 ( .A1(n2320), .A2(n2318), .A3(n2335), .A4(n2319), .ZN(n2229)
         );
  AND2_X1 U2434 ( .A1(n2317), .A2(n2337), .ZN(n2320) );
  NOR2_X2 U2435 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2343)
         );
  NOR2_X1 U2436 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2335)
         );
  INV_X1 U2437 ( .A(IR_REG_24__SCAN_IN), .ZN(n4691) );
  AND2_X1 U2438 ( .A1(n4386), .A2(REG1_REG_9__SCAN_IN), .ZN(n2135) );
  NAND2_X1 U2439 ( .A1(n2371), .A2(n2370), .ZN(n2569) );
  XNOR2_X1 U2440 ( .A(n2346), .B(IR_REG_2__SCAN_IN), .ZN(n4391) );
  INV_X1 U2441 ( .A(n3830), .ZN(n3838) );
  INV_X1 U2442 ( .A(n3925), .ZN(n2306) );
  INV_X1 U2443 ( .A(n3384), .ZN(n2283) );
  NOR2_X1 U2444 ( .A1(n2143), .A2(n2165), .ZN(n2278) );
  OAI21_X1 U2445 ( .B1(n2682), .B2(n2447), .A(n2217), .ZN(n2863) );
  NAND2_X1 U2446 ( .A1(n2682), .A2(DATAI_1_), .ZN(n2217) );
  NAND2_X1 U2447 ( .A1(n2584), .A2(n2583), .ZN(n2670) );
  NAND2_X1 U2448 ( .A1(n4026), .A2(n2201), .ZN(n4485) );
  NAND2_X1 U2449 ( .A1(n3427), .A2(n2202), .ZN(n2201) );
  INV_X1 U2450 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2202) );
  NOR2_X1 U2451 ( .A1(n4485), .A2(n4486), .ZN(n4484) );
  CLKBUF_X1 U2452 ( .A(n2670), .Z(n2638) );
  AND2_X1 U2453 ( .A1(n3466), .A2(n2920), .ZN(n3485) );
  NAND2_X1 U2454 ( .A1(n2243), .A2(n2242), .ZN(n4095) );
  AOI21_X1 U2455 ( .B1(n2244), .B2(n2142), .A(n2162), .ZN(n2242) );
  AOI21_X1 U2456 ( .B1(n2226), .B2(n2228), .A(n2161), .ZN(n2224) );
  NAND2_X1 U2457 ( .A1(n2291), .A2(n2289), .ZN(n3888) );
  NAND2_X1 U2458 ( .A1(n3815), .A2(n2290), .ZN(n2289) );
  AOI21_X1 U2459 ( .B1(n3818), .B2(n2294), .A(n2292), .ZN(n2291) );
  AND2_X1 U2460 ( .A1(n2299), .A2(n2308), .ZN(n2290) );
  OAI22_X1 U2461 ( .A1(n2239), .A2(n3180), .B1(n3231), .B2(n3270), .ZN(n2238)
         );
  NAND2_X1 U2462 ( .A1(n3117), .A2(n3118), .ZN(n2239) );
  NOR2_X1 U2463 ( .A1(n2241), .A2(n3180), .ZN(n2240) );
  INV_X1 U2464 ( .A(n3117), .ZN(n2241) );
  NAND2_X1 U2465 ( .A1(n2454), .A2(n2453), .ZN(n2455) );
  INV_X1 U2466 ( .A(n2463), .ZN(n2191) );
  NOR2_X1 U2467 ( .A1(n4458), .A2(n2203), .ZN(n2476) );
  AND2_X1 U2468 ( .A1(n3376), .A2(REG2_REG_15__SCAN_IN), .ZN(n2203) );
  AND2_X1 U2469 ( .A1(n3463), .A2(n3462), .ZN(n3875) );
  INV_X1 U2470 ( .A(n2240), .ZN(n2233) );
  INV_X1 U2471 ( .A(n2238), .ZN(n2235) );
  NOR2_X1 U2472 ( .A1(n2238), .A2(n3519), .ZN(n2236) );
  NAND2_X1 U2473 ( .A1(n3119), .A2(n2240), .ZN(n2237) );
  NAND2_X1 U2474 ( .A1(n2983), .A2(n3154), .ZN(n3567) );
  NAND2_X1 U2475 ( .A1(n2979), .A2(n2978), .ZN(n2231) );
  NAND2_X1 U2476 ( .A1(n2960), .A2(n4212), .ZN(n3558) );
  NAND2_X1 U2477 ( .A1(n4314), .A2(n3393), .ZN(n2176) );
  NAND2_X1 U2478 ( .A1(n2271), .A2(n4613), .ZN(n2440) );
  INV_X1 U2479 ( .A(IR_REG_6__SCAN_IN), .ZN(n2334) );
  INV_X1 U2480 ( .A(IR_REG_2__SCAN_IN), .ZN(n2314) );
  NAND2_X1 U2481 ( .A1(n2193), .A2(n2326), .ZN(n2192) );
  INV_X1 U2482 ( .A(IR_REG_1__SCAN_IN), .ZN(n2193) );
  INV_X1 U2483 ( .A(n3935), .ZN(n2308) );
  NAND2_X1 U2484 ( .A1(n2266), .A2(n3799), .ZN(n2264) );
  NAND2_X1 U2485 ( .A1(n2688), .A2(n2784), .ZN(n2251) );
  INV_X1 U2486 ( .A(n3136), .ZN(n2259) );
  INV_X1 U2487 ( .A(n2261), .ZN(n2260) );
  INV_X1 U2488 ( .A(n2258), .ZN(n2257) );
  OAI21_X1 U2489 ( .B1(n3061), .B2(n2259), .A(n3204), .ZN(n2258) );
  INV_X1 U2490 ( .A(n3210), .ZN(n3206) );
  OR2_X1 U2491 ( .A1(n2615), .A2(n4660), .ZN(n2622) );
  AND2_X1 U2492 ( .A1(n2275), .A2(n2163), .ZN(n2272) );
  NAND2_X1 U2493 ( .A1(n2278), .A2(n2277), .ZN(n2276) );
  NAND2_X1 U2494 ( .A1(n3943), .A2(n3944), .ZN(n3942) );
  AOI21_X1 U2495 ( .B1(n2150), .B2(n3298), .A(n2287), .ZN(n2286) );
  NOR2_X1 U2496 ( .A1(n3296), .A2(n2288), .ZN(n2287) );
  NOR2_X1 U2497 ( .A1(n3956), .A2(n2269), .ZN(n2266) );
  OR2_X1 U2498 ( .A1(n3917), .A2(n3799), .ZN(n2267) );
  AOI21_X1 U2499 ( .B1(n2762), .B2(n3830), .A(n2775), .ZN(n2776) );
  XNOR2_X1 U2500 ( .A(n2774), .B(n2805), .ZN(n2778) );
  NAND2_X1 U2501 ( .A1(n2306), .A2(n2157), .ZN(n2304) );
  NAND2_X1 U2502 ( .A1(n2305), .A2(n3817), .ZN(n2303) );
  NAND2_X1 U2503 ( .A1(n3818), .A2(n3817), .ZN(n2297) );
  NAND2_X1 U2504 ( .A1(n3815), .A2(n2308), .ZN(n2307) );
  NOR2_X1 U2505 ( .A1(n3684), .A2(n3683), .ZN(n3720) );
  NAND2_X1 U2506 ( .A1(n2551), .A2(n2458), .ZN(n2459) );
  NAND2_X1 U2507 ( .A1(n2467), .A2(n2197), .ZN(n2468) );
  NAND2_X1 U2508 ( .A1(n4386), .A2(REG2_REG_9__SCAN_IN), .ZN(n2197) );
  OR2_X1 U2509 ( .A1(n4424), .A2(n4764), .ZN(n2207) );
  NAND2_X1 U2510 ( .A1(n2470), .A2(n4427), .ZN(n2471) );
  OAI22_X1 U2511 ( .A1(n3401), .A2(n2195), .B1(n3300), .B2(
        REG2_REG_13__SCAN_IN), .ZN(n2473) );
  NOR2_X1 U2512 ( .A1(n3408), .A2(n2196), .ZN(n2195) );
  INV_X1 U2513 ( .A(REG2_REG_13__SCAN_IN), .ZN(n2196) );
  XNOR2_X1 U2514 ( .A(n2476), .B(n3414), .ZN(n4469) );
  NAND2_X1 U2515 ( .A1(n4469), .A2(n4468), .ZN(n4467) );
  OR2_X1 U2516 ( .A1(n3486), .A2(n3848), .ZN(n4033) );
  AND2_X1 U2517 ( .A1(n3860), .A2(n2248), .ZN(n2247) );
  OR2_X1 U2518 ( .A1(n3861), .A2(n2249), .ZN(n2248) );
  OR2_X1 U2519 ( .A1(n4156), .A2(n2187), .ZN(n3858) );
  NOR2_X1 U2520 ( .A1(n3547), .A2(n4134), .ZN(n4154) );
  OR2_X1 U2521 ( .A1(n3328), .A2(n2648), .ZN(n3417) );
  OR2_X1 U2522 ( .A1(n3730), .A2(n4314), .ZN(n3704) );
  OAI21_X1 U2523 ( .B1(n3123), .B2(n3122), .A(n3574), .ZN(n3184) );
  AND2_X1 U2524 ( .A1(n2586), .A2(n2585), .ZN(n2680) );
  AND2_X1 U2525 ( .A1(n2734), .A2(n2733), .ZN(n2954) );
  AND2_X1 U2526 ( .A1(n2750), .A2(n2759), .ZN(n2953) );
  NOR2_X1 U2527 ( .A1(n4064), .A2(n4053), .ZN(n4226) );
  OR2_X1 U2528 ( .A1(n4062), .A2(n4237), .ZN(n4064) );
  NAND2_X1 U2529 ( .A1(n4086), .A2(n4048), .ZN(n4062) );
  AND2_X1 U2530 ( .A1(n4103), .A2(n4088), .ZN(n4086) );
  NOR2_X1 U2531 ( .A1(n2137), .A2(n3768), .ZN(n4195) );
  INV_X1 U2532 ( .A(n3685), .ZN(n4314) );
  OR2_X1 U2533 ( .A1(n3366), .A2(n3323), .ZN(n3367) );
  NAND2_X1 U2534 ( .A1(n3243), .A2(n3290), .ZN(n3366) );
  AND2_X1 U2535 ( .A1(n3409), .A2(n2694), .ZN(n4297) );
  NAND2_X1 U2536 ( .A1(n3364), .A2(n4557), .ZN(n4549) );
  NAND2_X1 U2537 ( .A1(n2530), .A2(n2529), .ZN(n2718) );
  AND2_X1 U2538 ( .A1(n2740), .A2(n2752), .ZN(n2759) );
  NAND2_X1 U2539 ( .A1(n2511), .A2(IR_REG_31__SCAN_IN), .ZN(n2512) );
  OAI21_X1 U2540 ( .B1(n2513), .B2(n2483), .A(IR_REG_29__SCAN_IN), .ZN(n2171)
         );
  OAI21_X1 U2541 ( .B1(n2440), .B2(IR_REG_22__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2432) );
  NAND2_X1 U2542 ( .A1(n2411), .A2(n2522), .ZN(n2412) );
  INV_X1 U2543 ( .A(IR_REG_19__SCAN_IN), .ZN(n4685) );
  OR2_X1 U2544 ( .A1(n2340), .A2(IR_REG_9__SCAN_IN), .ZN(n2384) );
  INV_X1 U2545 ( .A(n2326), .ZN(n2522) );
  AOI21_X1 U2546 ( .B1(n3888), .B2(n3887), .A(n2310), .ZN(n3847) );
  INV_X1 U2547 ( .A(n3353), .ZN(n3662) );
  INV_X1 U2548 ( .A(n4384), .ZN(n3627) );
  OAI21_X1 U2549 ( .B1(n4090), .B2(n2679), .A(n2925), .ZN(n4249) );
  NAND2_X1 U2550 ( .A1(n2450), .A2(n2449), .ZN(n4017) );
  INV_X1 U2551 ( .A(n4390), .ZN(n2550) );
  XNOR2_X1 U2552 ( .A(n2468), .B(n4520), .ZN(n4420) );
  NAND2_X1 U2553 ( .A1(n4420), .A2(REG2_REG_10__SCAN_IN), .ZN(n4419) );
  XNOR2_X1 U2554 ( .A(n2471), .B(n4517), .ZN(n4440) );
  NAND2_X1 U2555 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4440), .ZN(n4439) );
  NOR2_X1 U2556 ( .A1(n4480), .A2(n4481), .ZN(n4479) );
  NAND2_X1 U2557 ( .A1(n2216), .A2(n4474), .ZN(n2215) );
  NAND2_X1 U2558 ( .A1(n4480), .A2(n4481), .ZN(n2216) );
  OAI21_X1 U2559 ( .B1(n4490), .B2(n4511), .A(n2213), .ZN(n2212) );
  AOI21_X1 U2560 ( .B1(n4483), .B2(ADDR_REG_18__SCAN_IN), .A(n4482), .ZN(n2213) );
  XNOR2_X1 U2561 ( .A(n2199), .B(n2198), .ZN(n2495) );
  INV_X1 U2562 ( .A(n2478), .ZN(n2198) );
  NOR2_X1 U2563 ( .A1(n4484), .A2(n2200), .ZN(n2199) );
  AND2_X1 U2564 ( .A1(n2540), .A2(n4007), .ZN(n4488) );
  INV_X1 U2565 ( .A(n4502), .ZN(n4162) );
  INV_X1 U2566 ( .A(n2689), .ZN(n3518) );
  INV_X1 U2567 ( .A(n2740), .ZN(n2744) );
  INV_X1 U2568 ( .A(n3905), .ZN(n2277) );
  NAND2_X1 U2569 ( .A1(n3963), .A2(n2277), .ZN(n2275) );
  INV_X1 U2570 ( .A(n2156), .ZN(n2305) );
  AND2_X1 U2571 ( .A1(n3549), .A2(n4111), .ZN(n3876) );
  OAI21_X1 U2572 ( .B1(n2569), .B2(n2376), .A(n2377), .ZN(n2381) );
  AND2_X1 U2573 ( .A1(n3376), .A2(REG1_REG_15__SCAN_IN), .ZN(n2210) );
  NOR2_X1 U2574 ( .A1(n3863), .A2(n2245), .ZN(n2244) );
  INV_X1 U2575 ( .A(n2247), .ZN(n2245) );
  INV_X1 U2576 ( .A(n2227), .ZN(n2226) );
  OAI21_X1 U2577 ( .B1(n3746), .B2(n2228), .A(n3853), .ZN(n2227) );
  NAND2_X1 U2578 ( .A1(n4295), .A2(n3855), .ZN(n3853) );
  INV_X1 U2579 ( .A(n3755), .ZN(n2228) );
  NAND2_X1 U2580 ( .A1(n3567), .A2(n3564), .ZN(n2230) );
  NAND2_X1 U2581 ( .A1(n2677), .A2(REG2_REG_1__SCAN_IN), .ZN(n2687) );
  OR2_X1 U2582 ( .A1(n2679), .A2(n2678), .ZN(n2684) );
  NAND2_X1 U2583 ( .A1(n2680), .A2(REG1_REG_1__SCAN_IN), .ZN(n2685) );
  AND2_X1 U2584 ( .A1(n4131), .A2(n4130), .ZN(n4171) );
  AND2_X1 U2585 ( .A1(n4493), .A2(n2888), .ZN(n2879) );
  OR2_X1 U2586 ( .A1(n2718), .A2(n2715), .ZN(n2734) );
  INV_X1 U2587 ( .A(IR_REG_25__SCAN_IN), .ZN(n2423) );
  AND4_X1 U2588 ( .A1(n2419), .A2(n2418), .A3(n2417), .A4(n2416), .ZN(n2420)
         );
  INV_X1 U2589 ( .A(n2480), .ZN(n2425) );
  INV_X1 U2590 ( .A(IR_REG_18__SCAN_IN), .ZN(n4686) );
  NAND2_X1 U2591 ( .A1(n2311), .A2(n2322), .ZN(n2323) );
  INV_X1 U2592 ( .A(IR_REG_17__SCAN_IN), .ZN(n2328) );
  INV_X1 U2593 ( .A(IR_REG_13__SCAN_IN), .ZN(n4602) );
  INV_X1 U2594 ( .A(IR_REG_7__SCAN_IN), .ZN(n2373) );
  AOI21_X1 U2595 ( .B1(n2300), .B2(n3976), .A(n3975), .ZN(n2299) );
  INV_X1 U2596 ( .A(n2304), .ZN(n2300) );
  NOR2_X1 U2597 ( .A1(n2295), .A2(n2293), .ZN(n2292) );
  NOR2_X1 U2598 ( .A1(n2302), .A2(n2296), .ZN(n2295) );
  INV_X1 U2599 ( .A(n2299), .ZN(n2293) );
  INV_X1 U2600 ( .A(n3976), .ZN(n2296) );
  AND2_X1 U2601 ( .A1(n2299), .A2(n3817), .ZN(n2294) );
  AND2_X1 U2602 ( .A1(n3072), .A2(REG3_REG_10__SCAN_IN), .ZN(n3074) );
  NAND2_X1 U2603 ( .A1(n2907), .A2(REG3_REG_7__SCAN_IN), .ZN(n2615) );
  OAI21_X1 U2604 ( .B1(n3818), .B2(n2305), .A(n3817), .ZN(n3934) );
  INV_X1 U2605 ( .A(n3843), .ZN(n3835) );
  AND2_X1 U2606 ( .A1(n3309), .A2(n3308), .ZN(n3384) );
  NAND2_X1 U2607 ( .A1(n3074), .A2(REG3_REG_11__SCAN_IN), .ZN(n2656) );
  INV_X1 U2608 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2600) );
  INV_X1 U2609 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2601) );
  OR3_X1 U2610 ( .A1(n2656), .A2(n2601), .A3(n2600), .ZN(n2602) );
  INV_X1 U2611 ( .A(n4212), .ZN(n2948) );
  NOR2_X1 U2612 ( .A1(n2905), .A2(n2904), .ZN(n2907) );
  INV_X1 U2613 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2904) );
  NOR2_X1 U2614 ( .A1(n2602), .A2(n4658), .ZN(n3326) );
  AND3_X1 U2615 ( .A1(n2877), .A2(n2954), .A3(n2951), .ZN(n2796) );
  XNOR2_X1 U2616 ( .A(n2452), .B(n2550), .ZN(n2545) );
  XNOR2_X1 U2617 ( .A(n2455), .B(n2498), .ZN(n4404) );
  OAI21_X1 U2618 ( .B1(n2461), .B2(n2191), .A(n2189), .ZN(n2465) );
  INV_X1 U2619 ( .A(n2190), .ZN(n2189) );
  XNOR2_X1 U2620 ( .A(n2381), .B(n3026), .ZN(n2727) );
  NOR2_X1 U2621 ( .A1(n2847), .A2(n2846), .ZN(n2845) );
  OR2_X1 U2622 ( .A1(n4416), .A2(n4764), .ZN(n2209) );
  NAND2_X1 U2623 ( .A1(n2387), .A2(n2206), .ZN(n2204) );
  INV_X1 U2624 ( .A(n4424), .ZN(n2206) );
  NOR2_X1 U2625 ( .A1(n2313), .A2(n2397), .ZN(n2400) );
  INV_X1 U2626 ( .A(n2396), .ZN(n2397) );
  XNOR2_X1 U2627 ( .A(n2407), .B(n3414), .ZN(n4472) );
  NAND2_X1 U2628 ( .A1(n4472), .A2(n4471), .ZN(n4470) );
  NAND2_X1 U2629 ( .A1(n4467), .A2(n2477), .ZN(n4027) );
  AND2_X1 U2630 ( .A1(n3425), .A2(REG2_REG_18__SCAN_IN), .ZN(n2200) );
  INV_X1 U2631 ( .A(n4248), .ZN(n4048) );
  AND2_X1 U2632 ( .A1(n3875), .A2(n2169), .ZN(n2168) );
  NAND2_X1 U2633 ( .A1(n3874), .A2(n2170), .ZN(n2169) );
  NAND2_X1 U2634 ( .A1(n4139), .A2(n4161), .ZN(n2249) );
  INV_X1 U2635 ( .A(n4144), .ZN(n4138) );
  OR2_X1 U2636 ( .A1(n4152), .A2(n4154), .ZN(n2250) );
  NAND2_X1 U2637 ( .A1(n4193), .A2(n4283), .ZN(n4173) );
  AND2_X1 U2638 ( .A1(n2682), .A2(DATAI_20_), .ZN(n4196) );
  NAND2_X1 U2639 ( .A1(n3907), .A2(n3968), .ZN(n3755) );
  NOR2_X1 U2640 ( .A1(n3417), .A2(n2580), .ZN(n3419) );
  AOI22_X1 U2641 ( .A1(n3745), .A2(n3744), .B1(n3743), .B2(n3742), .ZN(n3747)
         );
  NAND2_X1 U2642 ( .A1(n3747), .A2(n3746), .ZN(n3756) );
  NAND2_X1 U2643 ( .A1(n3707), .A2(n3706), .ZN(n4185) );
  AND2_X1 U2644 ( .A1(n3690), .A2(n3698), .ZN(n3644) );
  AND2_X1 U2645 ( .A1(n3410), .A2(n3411), .ZN(n3531) );
  INV_X1 U2646 ( .A(n2236), .ZN(n2234) );
  AOI21_X1 U2647 ( .B1(n2236), .B2(n2233), .A(n2148), .ZN(n2232) );
  NAND2_X1 U2648 ( .A1(n3184), .A2(n3589), .ZN(n3185) );
  NAND2_X1 U2649 ( .A1(n2237), .A2(n2236), .ZN(n3236) );
  NAND2_X1 U2650 ( .A1(n2237), .A2(n2235), .ZN(n3182) );
  NAND2_X1 U2651 ( .A1(n3070), .A2(n3578), .ZN(n3123) );
  AND2_X1 U2652 ( .A1(n2592), .A2(n2591), .ZN(n3211) );
  NAND2_X1 U2653 ( .A1(n3027), .A2(n3577), .ZN(n2172) );
  NAND2_X1 U2654 ( .A1(n2829), .A2(REG3_REG_5__SCAN_IN), .ZN(n2905) );
  OAI21_X1 U2655 ( .B1(n3153), .B2(n2987), .A(n3567), .ZN(n3004) );
  AND4_X1 U2656 ( .A1(n2812), .A2(n2811), .A3(n2810), .A4(n2809), .ZN(n2989)
         );
  INV_X1 U2657 ( .A(n2997), .ZN(n3000) );
  NAND2_X1 U2658 ( .A1(n3151), .A2(n3154), .ZN(n2185) );
  AND2_X1 U2659 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2829) );
  INV_X1 U2660 ( .A(n2230), .ZN(n3152) );
  NAND2_X1 U2661 ( .A1(n2986), .A2(n3563), .ZN(n3153) );
  AND2_X1 U2662 ( .A1(n2832), .A2(n2831), .ZN(n3155) );
  NAND2_X1 U2663 ( .A1(n2958), .A2(n3529), .ZN(n2986) );
  NOR2_X1 U2664 ( .A1(n2964), .A2(n2977), .ZN(n3151) );
  OR2_X1 U2665 ( .A1(n2443), .A2(IR_REG_27__SCAN_IN), .ZN(n2219) );
  NAND2_X1 U2666 ( .A1(n2689), .A2(n3553), .ZN(n2693) );
  OR2_X1 U2667 ( .A1(n2689), .A2(n3553), .ZN(n2872) );
  AND2_X1 U2668 ( .A1(n4118), .A2(n4105), .ZN(n4103) );
  NOR2_X1 U2669 ( .A1(n4143), .A2(n4265), .ZN(n4118) );
  INV_X1 U2670 ( .A(n4120), .ZN(n4265) );
  OR2_X1 U2671 ( .A1(n4279), .A2(n4138), .ZN(n4143) );
  AND2_X1 U2672 ( .A1(n4195), .A2(n4292), .ZN(n4193) );
  INV_X1 U2673 ( .A(n2176), .ZN(n2175) );
  INV_X1 U2674 ( .A(n3388), .ZN(n4331) );
  NOR2_X1 U2675 ( .A1(n3367), .A2(n3660), .ZN(n3652) );
  INV_X1 U2676 ( .A(n3323), .ZN(n3368) );
  NOR2_X1 U2677 ( .A1(n3191), .A2(n3260), .ZN(n3243) );
  NAND2_X1 U2678 ( .A1(n2188), .A2(n3231), .ZN(n3191) );
  AND2_X1 U2679 ( .A1(n3106), .A2(n3105), .ZN(n3107) );
  NAND2_X1 U2680 ( .A1(n3107), .A2(n3145), .ZN(n3086) );
  NOR2_X1 U2681 ( .A1(n3011), .A2(n3020), .ZN(n3106) );
  NAND2_X1 U2682 ( .A1(n3151), .A2(n2184), .ZN(n3011) );
  NOR2_X1 U2683 ( .A1(n3000), .A2(n2984), .ZN(n2184) );
  INV_X1 U2684 ( .A(n4549), .ZN(n4543) );
  AND2_X1 U2685 ( .A1(n2695), .A2(n4491), .ZN(n4326) );
  INV_X1 U2686 ( .A(n4321), .ZN(n4330) );
  INV_X1 U2687 ( .A(IR_REG_20__SCAN_IN), .ZN(n2524) );
  NAND2_X1 U2688 ( .A1(n2523), .A2(n2522), .ZN(n2525) );
  INV_X1 U2689 ( .A(IR_REG_16__SCAN_IN), .ZN(n2405) );
  INV_X1 U2690 ( .A(IR_REG_15__SCAN_IN), .ZN(n2322) );
  OR2_X1 U2691 ( .A1(n2372), .A2(n2336), .ZN(n2340) );
  NOR2_X1 U2692 ( .A1(n2333), .A2(IR_REG_5__SCAN_IN), .ZN(n2367) );
  INV_X1 U2693 ( .A(n2343), .ZN(n2344) );
  NAND2_X1 U2694 ( .A1(n2152), .A2(n4603), .ZN(n2194) );
  NAND2_X1 U2695 ( .A1(n3062), .A2(n3061), .ZN(n3137) );
  AOI21_X1 U2696 ( .B1(n2138), .B2(n2282), .A(n2166), .ZN(n2281) );
  NAND2_X1 U2697 ( .A1(n3297), .A2(n2138), .ZN(n2280) );
  INV_X1 U2698 ( .A(n2154), .ZN(n2282) );
  NAND2_X1 U2699 ( .A1(n2265), .A2(n2159), .ZN(n3898) );
  NOR2_X1 U2700 ( .A1(n3895), .A2(n3896), .ZN(n3809) );
  INV_X1 U2701 ( .A(n2273), .ZN(n3904) );
  OAI21_X1 U2702 ( .B1(n3777), .B2(n2274), .A(n2279), .ZN(n2273) );
  INV_X1 U2703 ( .A(n2278), .ZN(n2274) );
  AND2_X1 U2704 ( .A1(n4033), .A2(n3478), .ZN(n4065) );
  NAND2_X1 U2705 ( .A1(n3137), .A2(n3136), .ZN(n3205) );
  AND2_X1 U2706 ( .A1(n2146), .A2(n2251), .ZN(n2769) );
  INV_X1 U2707 ( .A(n2863), .ZN(n2888) );
  NAND2_X1 U2708 ( .A1(n3934), .A2(n2307), .ZN(n3927) );
  NAND2_X1 U2709 ( .A1(n2898), .A2(n2897), .ZN(n2928) );
  OR2_X1 U2710 ( .A1(n3722), .A2(n3721), .ZN(n3723) );
  NAND2_X1 U2711 ( .A1(n2821), .A2(n2820), .ZN(n2898) );
  NAND2_X1 U2712 ( .A1(n2256), .A2(n2255), .ZN(n3209) );
  AOI22_X1 U2713 ( .A1(n2260), .A2(n2262), .B1(n2257), .B2(n2259), .ZN(n2255)
         );
  INV_X1 U2714 ( .A(n2745), .ZN(n4493) );
  NAND2_X1 U2715 ( .A1(n2284), .A2(n2286), .ZN(n3385) );
  NAND2_X1 U2716 ( .A1(n2285), .A2(n2154), .ZN(n2284) );
  INV_X1 U2717 ( .A(n3297), .ZN(n2285) );
  NAND2_X1 U2718 ( .A1(n2267), .A2(n2268), .ZN(n3955) );
  INV_X1 U2719 ( .A(n3991), .ZN(n3270) );
  INV_X1 U2720 ( .A(n2795), .ZN(n2792) );
  AOI21_X1 U2721 ( .B1(n2927), .B2(n2254), .A(n2145), .ZN(n2252) );
  INV_X1 U2722 ( .A(n2897), .ZN(n2254) );
  NAND2_X1 U2723 ( .A1(n2298), .A2(n2304), .ZN(n3979) );
  NAND2_X1 U2724 ( .A1(n2141), .A2(n2307), .ZN(n2298) );
  NAND2_X1 U2725 ( .A1(n2828), .A2(n2827), .ZN(n3985) );
  NAND2_X1 U2726 ( .A1(n3472), .A2(n3471), .ZN(n4080) );
  OAI21_X1 U2727 ( .B1(n3937), .B2(n2679), .A(n2843), .ZN(n3862) );
  NAND2_X1 U2728 ( .A1(n3458), .A2(n3457), .ZN(n4266) );
  NAND2_X1 U2729 ( .A1(n3436), .A2(n3435), .ZN(n4288) );
  INV_X1 U2730 ( .A(n4316), .ZN(n3743) );
  NAND4_X1 U2731 ( .A1(n2607), .A2(n2606), .A3(n2605), .A4(n2604), .ZN(n3353)
         );
  INV_X1 U2732 ( .A(n2989), .ZN(n2983) );
  AND3_X1 U2733 ( .A1(n2673), .A2(n2672), .A3(n2671), .ZN(n2675) );
  OR2_X1 U2734 ( .A1(n2670), .A2(n4206), .ZN(n2673) );
  OR2_X1 U2735 ( .A1(n2740), .A2(n4509), .ZN(n3994) );
  AND2_X1 U2736 ( .A1(n2490), .A2(n2488), .ZN(n2540) );
  NAND2_X1 U2737 ( .A1(n3995), .A2(n4006), .ZN(n4015) );
  XNOR2_X1 U2738 ( .A(n2459), .B(n2564), .ZN(n2562) );
  NAND2_X1 U2739 ( .A1(n2461), .A2(n2460), .ZN(n2576) );
  NAND2_X1 U2740 ( .A1(n2576), .A2(n2463), .ZN(n2574) );
  XNOR2_X1 U2741 ( .A(n2465), .B(n3026), .ZN(n2724) );
  NAND2_X1 U2742 ( .A1(n4419), .A2(n2469), .ZN(n4428) );
  NAND2_X1 U2743 ( .A1(n2205), .A2(n2204), .ZN(n4423) );
  NAND2_X1 U2744 ( .A1(n2472), .A2(n4439), .ZN(n3401) );
  XNOR2_X1 U2745 ( .A(n2473), .B(n2399), .ZN(n4447) );
  NOR2_X1 U2746 ( .A1(n4447), .A2(n4794), .ZN(n4446) );
  AND2_X1 U2747 ( .A1(n3494), .A2(n3493), .ZN(n4241) );
  OR2_X1 U2748 ( .A1(n3485), .A2(n2921), .ZN(n4090) );
  OR2_X1 U2749 ( .A1(n4152), .A2(n2142), .ZN(n2246) );
  NAND2_X1 U2750 ( .A1(n4193), .A2(n2186), .ZN(n4279) );
  NOR2_X1 U2751 ( .A1(n4161), .A2(n2187), .ZN(n2186) );
  NOR3_X1 U2752 ( .A1(n3367), .A2(n4325), .A3(n3660), .ZN(n3653) );
  INV_X1 U2753 ( .A(n4328), .ZN(n3730) );
  INV_X1 U2754 ( .A(n3262), .ZN(n3343) );
  INV_X1 U2755 ( .A(n3202), .ZN(n3230) );
  AND2_X1 U2756 ( .A1(n4505), .A2(n2976), .ZN(n4192) );
  NAND2_X1 U2757 ( .A1(n3110), .A2(n3025), .ZN(n3082) );
  AND2_X1 U2758 ( .A1(n4505), .A2(n3627), .ZN(n3749) );
  OR2_X1 U2759 ( .A1(n2689), .A2(n2690), .ZN(n2691) );
  NAND2_X2 U2760 ( .A1(n2955), .A2(n4162), .ZN(n4505) );
  AND2_X2 U2761 ( .A1(n4536), .A2(n2760), .ZN(n4502) );
  INV_X2 U2762 ( .A(n4574), .ZN(n4577) );
  NAND2_X1 U2763 ( .A1(n4225), .A2(n2180), .ZN(n4397) );
  AOI21_X1 U2764 ( .B1(n4562), .B2(n4234), .A(n4233), .ZN(n4235) );
  AND2_X1 U2765 ( .A1(n4064), .A2(n4063), .ZN(n4347) );
  AND2_X1 U2766 ( .A1(n4565), .A2(n4562), .ZN(n4346) );
  INV_X1 U2767 ( .A(n4509), .ZN(n2752) );
  INV_X1 U2768 ( .A(IR_REG_30__SCAN_IN), .ZN(n3884) );
  XNOR2_X1 U2769 ( .A(n2426), .B(IR_REG_26__SCAN_IN), .ZN(n2530) );
  NAND2_X1 U2770 ( .A1(n2434), .A2(IR_REG_31__SCAN_IN), .ZN(n2426) );
  XNOR2_X1 U2771 ( .A(n2422), .B(IR_REG_24__SCAN_IN), .ZN(n2534) );
  NAND2_X1 U2772 ( .A1(n2421), .A2(IR_REG_31__SCAN_IN), .ZN(n2422) );
  INV_X1 U2773 ( .A(n2758), .ZN(n3556) );
  AND2_X1 U2774 ( .A1(n2523), .A2(n2413), .ZN(n4384) );
  AND2_X1 U2775 ( .A1(n2339), .A2(n2388), .ZN(n4518) );
  AND2_X1 U2776 ( .A1(n2357), .A2(n2353), .ZN(n4390) );
  OR2_X1 U2777 ( .A1(n2343), .A2(n2326), .ZN(n2346) );
  INV_X1 U2778 ( .A(n2212), .ZN(n2211) );
  OR2_X1 U2779 ( .A1(n4479), .A2(n2215), .ZN(n2214) );
  OAI21_X1 U2780 ( .B1(n4397), .B2(n4174), .A(n2177), .ZN(U3261) );
  AND2_X1 U2781 ( .A1(n2179), .A2(n2178), .ZN(n2177) );
  NAND2_X1 U2782 ( .A1(n4505), .A2(n4398), .ZN(n2178) );
  OR2_X1 U2783 ( .A1(n4505), .A2(n4809), .ZN(n2179) );
  NAND3_X4 U2784 ( .A1(n2219), .A2(n2218), .A3(n2436), .ZN(n2682) );
  OR2_X1 U2785 ( .A1(n3367), .A2(n2174), .ZN(n2137) );
  AND2_X1 U2786 ( .A1(n2286), .A2(n2283), .ZN(n2138) );
  AND2_X1 U2787 ( .A1(n2134), .A2(n2229), .ZN(n2139) );
  NAND2_X1 U2788 ( .A1(n2271), .A2(n2425), .ZN(n2434) );
  AND2_X1 U2789 ( .A1(n3211), .A2(n3145), .ZN(n2140) );
  AND2_X1 U2790 ( .A1(n2297), .A2(n2301), .ZN(n2141) );
  OR2_X1 U2791 ( .A1(n4154), .A2(n3861), .ZN(n2142) );
  AND2_X1 U2792 ( .A1(n3779), .A2(n3778), .ZN(n2143) );
  INV_X1 U2793 ( .A(n2133), .ZN(n3445) );
  INV_X1 U2794 ( .A(n3299), .ZN(n2288) );
  AND2_X1 U2795 ( .A1(n2267), .A2(n2266), .ZN(n2144) );
  AND2_X1 U2796 ( .A1(n2931), .A2(n2930), .ZN(n2145) );
  NAND2_X1 U2797 ( .A1(n2246), .A2(n2247), .ZN(n4116) );
  NAND2_X1 U2798 ( .A1(n2534), .A2(n2431), .ZN(n2740) );
  NAND2_X1 U2799 ( .A1(n2745), .A2(n3843), .ZN(n2146) );
  NAND2_X1 U2800 ( .A1(n2183), .A2(n2134), .ZN(n2482) );
  NAND2_X1 U2801 ( .A1(n2151), .A2(n2344), .ZN(n2447) );
  INV_X1 U2802 ( .A(IR_REG_31__SCAN_IN), .ZN(n2326) );
  OR2_X1 U2803 ( .A1(n2257), .A2(n2260), .ZN(n2147) );
  AND2_X1 U2804 ( .A1(n3343), .A2(n3271), .ZN(n2148) );
  NAND2_X1 U2805 ( .A1(n2485), .A2(n2511), .ZN(n2149) );
  NAND2_X1 U2806 ( .A1(n3296), .A2(n2288), .ZN(n2150) );
  NAND2_X1 U2807 ( .A1(n2675), .A2(n2674), .ZN(n2866) );
  AND2_X1 U2808 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2152)
         );
  AND2_X1 U2809 ( .A1(n3028), .A2(n3579), .ZN(n3570) );
  AND2_X1 U2810 ( .A1(n2250), .A2(n2249), .ZN(n2153) );
  INV_X1 U2811 ( .A(IR_REG_27__SCAN_IN), .ZN(n2435) );
  INV_X1 U2812 ( .A(IR_REG_28__SCAN_IN), .ZN(n2485) );
  INV_X1 U2813 ( .A(IR_REG_26__SCAN_IN), .ZN(n2181) );
  INV_X2 U2814 ( .A(n2670), .ZN(n2677) );
  NAND2_X2 U2815 ( .A1(n2586), .A2(n2583), .ZN(n2679) );
  INV_X1 U2816 ( .A(IR_REG_22__SCAN_IN), .ZN(n2437) );
  OR2_X1 U2817 ( .A1(n3299), .A2(n3298), .ZN(n2154) );
  INV_X1 U2818 ( .A(IR_REG_11__SCAN_IN), .ZN(n2337) );
  NAND2_X1 U2819 ( .A1(n2225), .A2(n2224), .ZN(n4190) );
  NAND2_X1 U2820 ( .A1(n3756), .A2(n3755), .ZN(n3854) );
  NAND2_X1 U2821 ( .A1(n3297), .A2(n3296), .ZN(n2155) );
  OR2_X1 U2822 ( .A1(n3811), .A2(n3810), .ZN(n2156) );
  AND2_X1 U2823 ( .A1(n3824), .A2(n3823), .ZN(n2157) );
  OR3_X1 U2824 ( .A1(n3367), .A2(n4325), .A3(n2176), .ZN(n2158) );
  INV_X1 U2825 ( .A(n2984), .ZN(n3154) );
  AND2_X1 U2826 ( .A1(n3809), .A2(n2264), .ZN(n2159) );
  AND2_X1 U2827 ( .A1(n4331), .A2(n3393), .ZN(n2160) );
  INV_X1 U2828 ( .A(IR_REG_21__SCAN_IN), .ZN(n4613) );
  INV_X1 U2829 ( .A(n3907), .ZN(n3990) );
  AND2_X1 U2830 ( .A1(n3950), .A2(n3908), .ZN(n2161) );
  INV_X1 U2831 ( .A(n2302), .ZN(n2301) );
  AND3_X1 U2832 ( .A1(n2646), .A2(n2645), .A3(n2644), .ZN(n3950) );
  INV_X1 U2833 ( .A(n3950), .ZN(n4295) );
  INV_X1 U2834 ( .A(n2269), .ZN(n2268) );
  NOR2_X1 U2835 ( .A1(n3798), .A2(n3797), .ZN(n2269) );
  NOR2_X1 U2836 ( .A1(n2331), .A2(n2323), .ZN(n2325) );
  NOR2_X1 U2837 ( .A1(n3862), .A2(n4265), .ZN(n2162) );
  OR2_X1 U2838 ( .A1(n3785), .A2(n3784), .ZN(n2163) );
  NAND2_X1 U2839 ( .A1(n4518), .A2(REG1_REG_11__SCAN_IN), .ZN(n2164) );
  XNOR2_X1 U2840 ( .A(n2525), .B(n2524), .ZN(n2700) );
  OR2_X1 U2841 ( .A1(n3111), .A2(n3570), .ZN(n3110) );
  INV_X1 U2842 ( .A(n3766), .ZN(n3968) );
  INV_X1 U2843 ( .A(n3408), .ZN(n3300) );
  AND2_X1 U2844 ( .A1(n3749), .A2(n4562), .ZN(n4399) );
  INV_X1 U2845 ( .A(n3706), .ZN(n2170) );
  OAI21_X1 U2846 ( .B1(n3119), .B2(n3118), .A(n3117), .ZN(n3181) );
  NOR2_X1 U2847 ( .A1(n2482), .A2(n2481), .ZN(n2486) );
  AND2_X1 U2848 ( .A1(n3782), .A2(n3781), .ZN(n2165) );
  AND2_X1 U2849 ( .A1(n3307), .A2(n3306), .ZN(n2166) );
  NAND2_X1 U2850 ( .A1(n2762), .A2(n2888), .ZN(n3554) );
  NAND2_X1 U2851 ( .A1(n2231), .A2(n2982), .ZN(n3156) );
  INV_X1 U2852 ( .A(n2188), .ZN(n3124) );
  NOR2_X1 U2853 ( .A1(n3086), .A2(n3200), .ZN(n2188) );
  INV_X1 U2854 ( .A(n3963), .ZN(n2279) );
  INV_X1 U2855 ( .A(n3741), .ZN(n3742) );
  AND2_X1 U2856 ( .A1(n2209), .A2(n2208), .ZN(n2167) );
  NAND2_X1 U2857 ( .A1(n2682), .A2(DATAI_21_), .ZN(n4283) );
  INV_X1 U2858 ( .A(n4283), .ZN(n2187) );
  AND2_X1 U2859 ( .A1(n2540), .A2(n4003), .ZN(n4474) );
  NAND2_X1 U2860 ( .A1(n2182), .A2(IR_REG_31__SCAN_IN), .ZN(n2443) );
  AND2_X1 U2861 ( .A1(n2486), .A2(n2485), .ZN(n2513) );
  INV_X1 U2862 ( .A(n2585), .ZN(n2583) );
  OAI21_X2 U2863 ( .B1(n3707), .B2(n3464), .A(n2168), .ZN(n4112) );
  NAND2_X1 U2864 ( .A1(n4112), .A2(n3876), .ZN(n4097) );
  NAND2_X1 U2865 ( .A1(n2173), .A2(n3410), .ZN(n3379) );
  NAND2_X1 U2866 ( .A1(n3413), .A2(n3531), .ZN(n2173) );
  NAND3_X1 U2867 ( .A1(n3698), .A2(n2175), .A3(n3741), .ZN(n2174) );
  OR2_X1 U2868 ( .A1(n4226), .A2(n4229), .ZN(n2180) );
  NAND4_X1 U2869 ( .A1(n2425), .A2(n2183), .A3(n2134), .A4(n2181), .ZN(n2182)
         );
  NAND2_X1 U2870 ( .A1(n2185), .A2(n3000), .ZN(n2993) );
  OAI211_X1 U2871 ( .C1(n3151), .C2(n3154), .A(n2185), .B(n4562), .ZN(n4533)
         );
  OAI21_X1 U2872 ( .B1(n2460), .B2(n2191), .A(n2464), .ZN(n2190) );
  MUX2_X1 U2873 ( .A(n2448), .B(REG2_REG_1__SCAN_IN), .S(n2447), .Z(n3995) );
  NOR2_X1 U2874 ( .A1(n2474), .A2(n4446), .ZN(n4459) );
  AOI21_X1 U2875 ( .B1(n2495), .B2(n4488), .A(n2494), .ZN(n2496) );
  NAND2_X1 U2876 ( .A1(n4027), .A2(n4028), .ZN(n4026) );
  INV_X1 U2877 ( .A(n2209), .ZN(n4415) );
  INV_X1 U2878 ( .A(n2387), .ZN(n2208) );
  NAND3_X1 U2879 ( .A1(n2214), .A2(n4489), .A3(n2211), .ZN(U3258) );
  NAND2_X1 U2880 ( .A1(n2443), .A2(IR_REG_28__SCAN_IN), .ZN(n2218) );
  NOR2_X2 U2881 ( .A1(n3375), .A2(n2160), .ZN(n3643) );
  NOR2_X2 U2882 ( .A1(n3319), .A2(n3531), .ZN(n3375) );
  OAI22_X2 U2883 ( .A1(n2221), .A2(n2220), .B1(n3662), .B2(n3368), .ZN(n3319)
         );
  NOR2_X1 U2884 ( .A1(n3353), .A2(n3323), .ZN(n2220) );
  INV_X1 U2885 ( .A(n3354), .ZN(n2221) );
  NAND2_X1 U2886 ( .A1(n2222), .A2(n2223), .ZN(n3085) );
  NAND2_X1 U2887 ( .A1(n3111), .A2(n3025), .ZN(n2222) );
  NAND2_X1 U2888 ( .A1(n3747), .A2(n2226), .ZN(n2225) );
  NAND3_X1 U2889 ( .A1(n2231), .A2(n2982), .A3(n2230), .ZN(n3158) );
  OAI21_X1 U2890 ( .B1(n3119), .B2(n2234), .A(n2232), .ZN(n3318) );
  NAND2_X1 U2891 ( .A1(n4152), .A2(n2244), .ZN(n2243) );
  INV_X1 U2892 ( .A(n2250), .ZN(n4151) );
  NAND3_X1 U2893 ( .A1(n2146), .A2(n2743), .A3(n2251), .ZN(n2767) );
  NAND2_X1 U2894 ( .A1(n2253), .A2(n2252), .ZN(n3047) );
  NAND3_X1 U2895 ( .A1(n2821), .A2(n2820), .A3(n2927), .ZN(n2253) );
  NAND2_X1 U2896 ( .A1(n3062), .A2(n2147), .ZN(n2256) );
  OAI21_X1 U2897 ( .B1(n3061), .B2(n2262), .A(n3203), .ZN(n2261) );
  NAND2_X1 U2898 ( .A1(n3136), .A2(n2263), .ZN(n2262) );
  INV_X1 U2899 ( .A(n3204), .ZN(n2263) );
  NAND2_X1 U2900 ( .A1(n3917), .A2(n2266), .ZN(n2265) );
  INV_X1 U2901 ( .A(n2482), .ZN(n2271) );
  NAND2_X1 U2902 ( .A1(n2271), .A2(n2270), .ZN(n2517) );
  OAI21_X1 U2903 ( .B1(n3777), .B2(n2276), .A(n2272), .ZN(n3943) );
  NOR2_X1 U2904 ( .A1(n3777), .A2(n2143), .ZN(n3965) );
  NAND2_X1 U2905 ( .A1(n2306), .A2(n2303), .ZN(n2302) );
  NAND2_X1 U2906 ( .A1(n2868), .A2(n2867), .ZN(n2950) );
  INV_X1 U2907 ( .A(n2867), .ZN(n3530) );
  NAND2_X1 U2908 ( .A1(n2700), .A2(n4491), .ZN(n4551) );
  INV_X1 U2909 ( .A(n2700), .ZN(n2695) );
  OAI21_X2 U2910 ( .B1(n4169), .B2(n3859), .A(n3858), .ZN(n4152) );
  AOI21_X2 U2911 ( .B1(n4190), .B2(n3857), .A(n3856), .ZN(n4169) );
  NOR2_X2 U2912 ( .A1(n3870), .A2(n3869), .ZN(n4050) );
  AND2_X1 U2913 ( .A1(n2156), .A2(n3814), .ZN(n2309) );
  AND2_X1 U2914 ( .A1(n3841), .A2(n3840), .ZN(n2310) );
  AND2_X1 U2915 ( .A1(n2321), .A2(n2405), .ZN(n2311) );
  AND2_X1 U2916 ( .A1(n2351), .A2(n2315), .ZN(n2312) );
  MUX2_X1 U2917 ( .A(n3627), .B(n3416), .S(n2682), .Z(n3908) );
  NAND2_X1 U2918 ( .A1(n3158), .A2(n2985), .ZN(n2999) );
  NOR2_X1 U2919 ( .A1(n3403), .A2(n3402), .ZN(n2313) );
  INV_X1 U2920 ( .A(IR_REG_5__SCAN_IN), .ZN(n2317) );
  NAND2_X1 U2921 ( .A1(n2773), .A2(n2772), .ZN(n2774) );
  NAND2_X1 U2922 ( .A1(n2989), .A2(n2984), .ZN(n3564) );
  INV_X1 U2923 ( .A(IR_REG_29__SCAN_IN), .ZN(n2511) );
  OR2_X1 U2924 ( .A1(n4158), .A2(n4144), .ZN(n3860) );
  AND2_X1 U2925 ( .A1(n3355), .A2(n3320), .ZN(n3595) );
  NAND4_X1 U2926 ( .A1(n2687), .A2(n2686), .A3(n2685), .A4(n2684), .ZN(n2870)
         );
  INV_X1 U2927 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4658) );
  OR2_X1 U2928 ( .A1(n3283), .A2(n3282), .ZN(n3296) );
  INV_X1 U2929 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2621) );
  NAND2_X1 U2930 ( .A1(n3438), .A2(n2581), .ZN(n3440) );
  INV_X1 U2931 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4660) );
  AND2_X1 U2932 ( .A1(n2682), .A2(DATAI_27_), .ZN(n4248) );
  OR2_X1 U2933 ( .A1(n3440), .A2(n4862), .ZN(n3450) );
  NAND2_X1 U2934 ( .A1(n3002), .A2(n3001), .ZN(n3023) );
  INV_X1 U2935 ( .A(n3957), .ZN(n4161) );
  AND2_X1 U2936 ( .A1(n3591), .A2(n3590), .ZN(n3519) );
  INV_X1 U2937 ( .A(n4497), .ZN(n4327) );
  INV_X1 U2938 ( .A(n3056), .ZN(n3105) );
  OR2_X1 U2939 ( .A1(n3450), .A2(n3899), .ZN(n3452) );
  NOR2_X1 U2940 ( .A1(n3452), .A2(n4661), .ZN(n3466) );
  AND2_X1 U2941 ( .A1(n3728), .A2(n3727), .ZN(n3776) );
  NOR2_X1 U2942 ( .A1(n2622), .A2(n2621), .ZN(n3072) );
  AND2_X1 U2943 ( .A1(n3419), .A2(REG3_REG_19__SCAN_IN), .ZN(n3438) );
  INV_X1 U2944 ( .A(n4266), .ZN(n4158) );
  INV_X1 U2945 ( .A(n4325), .ZN(n3698) );
  OR2_X1 U2946 ( .A1(n2838), .A2(n3466), .ZN(n3937) );
  NOR2_X1 U2947 ( .A1(n2401), .A2(n4443), .ZN(n4455) );
  AOI21_X1 U2948 ( .B1(n4450), .B2(n4384), .A(n2491), .ZN(n2492) );
  OR2_X1 U2949 ( .A1(n4037), .A2(n3510), .ZN(n4057) );
  AND2_X1 U2950 ( .A1(n3631), .A2(n3556), .ZN(n2735) );
  INV_X1 U2951 ( .A(n3862), .ZN(n4142) );
  AND2_X1 U2952 ( .A1(n2630), .A2(n2629), .ZN(n4316) );
  INV_X1 U2953 ( .A(n4320), .ZN(n3690) );
  OR2_X1 U2954 ( .A1(n2718), .A2(D_REG_1__SCAN_IN), .ZN(n2951) );
  INV_X1 U2955 ( .A(n4326), .ZN(n4315) );
  INV_X1 U2956 ( .A(n3340), .ZN(n3290) );
  AND2_X1 U2957 ( .A1(n2700), .A2(n4384), .ZN(n4494) );
  AND2_X1 U2958 ( .A1(n2378), .A2(n2375), .ZN(n3024) );
  AND2_X1 U2959 ( .A1(n3487), .A2(n3486), .ZN(n3892) );
  AND2_X1 U2960 ( .A1(n3424), .A2(n3423), .ZN(n3907) );
  INV_X1 U2961 ( .A(n3211), .ZN(n3083) );
  AND2_X1 U2962 ( .A1(n2540), .A2(n2763), .ZN(n4450) );
  AND2_X1 U2963 ( .A1(n4382), .A2(n2735), .ZN(n4321) );
  INV_X1 U2964 ( .A(n4132), .ZN(n4170) );
  NOR2_X1 U2965 ( .A1(n3645), .A2(n3644), .ZN(n3647) );
  INV_X1 U2966 ( .A(n4297), .ZN(n4495) );
  AND2_X1 U2967 ( .A1(n4577), .A2(n4562), .ZN(n4244) );
  INV_X1 U2968 ( .A(n4196), .ZN(n4292) );
  INV_X1 U2969 ( .A(n4551), .ZN(n4562) );
  AND2_X1 U2970 ( .A1(n4494), .A2(n2692), .ZN(n4536) );
  INV_X1 U2971 ( .A(n2692), .ZN(n3631) );
  AND2_X1 U2972 ( .A1(n2490), .A2(n2489), .ZN(n4483) );
  NAND2_X1 U2973 ( .A1(n2796), .A2(n2739), .ZN(n3988) );
  NAND2_X1 U2974 ( .A1(n3484), .A2(n3483), .ZN(n4247) );
  OAI211_X1 U2975 ( .C1(n3445), .C2(n3444), .A(n3443), .B(n3442), .ZN(n4156)
         );
  INV_X1 U2976 ( .A(n4474), .ZN(n4478) );
  OR2_X1 U2977 ( .A1(n2394), .A2(n2393), .ZN(n3408) );
  INV_X1 U2978 ( .A(n4450), .ZN(n4490) );
  INV_X1 U2979 ( .A(n4192), .ZN(n4182) );
  INV_X1 U2980 ( .A(n4399), .ZN(n4174) );
  INV_X1 U2981 ( .A(n4244), .ZN(n4313) );
  OR2_X1 U2982 ( .A1(n2878), .A2(n2952), .ZN(n4574) );
  INV_X1 U2983 ( .A(n4346), .ZN(n4378) );
  OR2_X1 U2984 ( .A1(n2878), .A2(n2877), .ZN(n4563) );
  INV_X1 U2985 ( .A(n4507), .ZN(n4508) );
  AND2_X1 U2986 ( .A1(n2342), .A2(n2384), .ZN(n4386) );
  NAND2_X1 U2987 ( .A1(n2497), .A2(n2496), .ZN(U3259) );
  INV_X2 U2988 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND2_X1 U2989 ( .A1(n2343), .A2(n2314), .ZN(n2350) );
  INV_X1 U2990 ( .A(n2350), .ZN(n2316) );
  INV_X1 U2991 ( .A(IR_REG_3__SCAN_IN), .ZN(n2351) );
  INV_X1 U2992 ( .A(IR_REG_4__SCAN_IN), .ZN(n2315) );
  NAND2_X1 U2993 ( .A1(n2316), .A2(n2312), .ZN(n2333) );
  NOR2_X1 U2994 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2319)
         );
  NOR2_X1 U2995 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2318)
         );
  NAND2_X1 U2996 ( .A1(n2139), .A2(n4602), .ZN(n2331) );
  INV_X1 U2997 ( .A(IR_REG_14__SCAN_IN), .ZN(n2321) );
  NAND2_X1 U2998 ( .A1(n2325), .A2(n2328), .ZN(n2409) );
  NAND2_X1 U2999 ( .A1(n2409), .A2(IR_REG_31__SCAN_IN), .ZN(n2324) );
  XNOR2_X1 U3000 ( .A(n2324), .B(IR_REG_18__SCAN_IN), .ZN(n3425) );
  INV_X1 U3001 ( .A(n3425), .ZN(n4511) );
  INV_X1 U3002 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4769) );
  AOI22_X1 U3003 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4511), .B1(n3425), .B2(
        n4769), .ZN(n4481) );
  INV_X1 U3004 ( .A(n2325), .ZN(n2327) );
  NAND2_X1 U3005 ( .A1(n2327), .A2(n2522), .ZN(n2329) );
  MUX2_X1 U3006 ( .A(n2329), .B(IR_REG_31__SCAN_IN), .S(n2328), .Z(n2330) );
  NAND2_X1 U3007 ( .A1(n2330), .A2(n2409), .ZN(n3427) );
  INV_X1 U3008 ( .A(n3427), .ZN(n4385) );
  OR2_X1 U3009 ( .A1(n2331), .A2(IR_REG_14__SCAN_IN), .ZN(n2332) );
  NAND2_X1 U3010 ( .A1(n2332), .A2(IR_REG_31__SCAN_IN), .ZN(n2403) );
  XNOR2_X1 U3011 ( .A(n2403), .B(IR_REG_15__SCAN_IN), .ZN(n3376) );
  NAND2_X1 U3012 ( .A1(n2367), .A2(n2334), .ZN(n2372) );
  INV_X1 U3013 ( .A(n2335), .ZN(n2336) );
  OAI21_X1 U3014 ( .B1(n2384), .B2(IR_REG_10__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2338) );
  OR2_X1 U3015 ( .A1(n2338), .A2(n2337), .ZN(n2339) );
  NAND2_X1 U3016 ( .A1(n2338), .A2(n2337), .ZN(n2388) );
  NAND2_X1 U3017 ( .A1(n2340), .A2(n2522), .ZN(n2341) );
  INV_X1 U3018 ( .A(IR_REG_9__SCAN_IN), .ZN(n4601) );
  MUX2_X1 U3019 ( .A(n2341), .B(IR_REG_31__SCAN_IN), .S(n4601), .Z(n2342) );
  XNOR2_X1 U3020 ( .A(n2447), .B(REG1_REG_1__SCAN_IN), .ZN(n3998) );
  AND2_X1 U3021 ( .A1(REG1_REG_0__SCAN_IN), .A2(n4603), .ZN(n3997) );
  NAND2_X1 U3022 ( .A1(n3998), .A2(n3997), .ZN(n3996) );
  INV_X1 U3023 ( .A(n2447), .ZN(n4392) );
  NAND2_X1 U3024 ( .A1(n4392), .A2(REG1_REG_1__SCAN_IN), .ZN(n2345) );
  INV_X1 U3025 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2347) );
  XNOR2_X1 U3026 ( .A(n4391), .B(n2347), .ZN(n4011) );
  NAND2_X1 U3027 ( .A1(n4010), .A2(n4011), .ZN(n2349) );
  NAND2_X1 U3028 ( .A1(n2136), .A2(REG1_REG_2__SCAN_IN), .ZN(n2348) );
  NAND2_X1 U3029 ( .A1(n2350), .A2(IR_REG_31__SCAN_IN), .ZN(n2352) );
  NAND2_X1 U3030 ( .A1(n2352), .A2(n2351), .ZN(n2357) );
  OR2_X1 U3031 ( .A1(n2352), .A2(n2351), .ZN(n2353) );
  XNOR2_X1 U3032 ( .A(n2354), .B(n2550), .ZN(n2544) );
  NAND2_X1 U3033 ( .A1(n2544), .A2(REG1_REG_3__SCAN_IN), .ZN(n2356) );
  NAND2_X1 U3034 ( .A1(n2354), .A2(n4390), .ZN(n2355) );
  NAND2_X1 U3035 ( .A1(n2357), .A2(IR_REG_31__SCAN_IN), .ZN(n2358) );
  XNOR2_X1 U3036 ( .A(n2358), .B(IR_REG_4__SCAN_IN), .ZN(n4406) );
  INV_X1 U3037 ( .A(n4406), .ZN(n2498) );
  XNOR2_X1 U3038 ( .A(n2359), .B(n2498), .ZN(n4401) );
  NAND2_X1 U3039 ( .A1(n4401), .A2(REG1_REG_4__SCAN_IN), .ZN(n2361) );
  NAND2_X1 U3040 ( .A1(n2359), .A2(n4406), .ZN(n2360) );
  NAND2_X1 U3041 ( .A1(n2361), .A2(n2360), .ZN(n2557) );
  INV_X1 U3042 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2365) );
  INV_X1 U3043 ( .A(n2367), .ZN(n2364) );
  NAND2_X1 U3044 ( .A1(n2333), .A2(IR_REG_31__SCAN_IN), .ZN(n2362) );
  MUX2_X1 U3045 ( .A(IR_REG_31__SCAN_IN), .B(n2362), .S(IR_REG_5__SCAN_IN), 
        .Z(n2363) );
  NAND2_X1 U3046 ( .A1(n2364), .A2(n2363), .ZN(n2900) );
  MUX2_X1 U3047 ( .A(n2365), .B(REG1_REG_5__SCAN_IN), .S(n2900), .Z(n2558) );
  NAND2_X1 U3048 ( .A1(n2557), .A2(n2558), .ZN(n2556) );
  INV_X1 U3049 ( .A(n2900), .ZN(n4389) );
  NAND2_X1 U3050 ( .A1(n4389), .A2(REG1_REG_5__SCAN_IN), .ZN(n2366) );
  OR2_X1 U3051 ( .A1(n2367), .A2(n2483), .ZN(n2368) );
  XNOR2_X1 U3052 ( .A(n2368), .B(IR_REG_6__SCAN_IN), .ZN(n4388) );
  INV_X1 U3053 ( .A(n4388), .ZN(n2564) );
  XNOR2_X1 U3054 ( .A(n2369), .B(n2564), .ZN(n2561) );
  NAND2_X1 U3055 ( .A1(n2561), .A2(REG1_REG_6__SCAN_IN), .ZN(n2371) );
  NAND2_X1 U3056 ( .A1(n2369), .A2(n4388), .ZN(n2370) );
  NAND2_X1 U3057 ( .A1(n2372), .A2(n2522), .ZN(n2374) );
  NAND2_X1 U3058 ( .A1(n2374), .A2(n2373), .ZN(n2378) );
  OR2_X1 U3059 ( .A1(n2374), .A2(n2373), .ZN(n2375) );
  AND2_X1 U3060 ( .A1(n3024), .A2(REG1_REG_7__SCAN_IN), .ZN(n2376) );
  OR2_X1 U3061 ( .A1(n3024), .A2(REG1_REG_7__SCAN_IN), .ZN(n2377) );
  INV_X1 U3062 ( .A(n2381), .ZN(n2382) );
  NAND2_X1 U3063 ( .A1(n2378), .A2(IR_REG_31__SCAN_IN), .ZN(n2380) );
  INV_X1 U3064 ( .A(IR_REG_8__SCAN_IN), .ZN(n2379) );
  XNOR2_X1 U3065 ( .A(n2380), .B(n2379), .ZN(n3026) );
  INV_X1 U3066 ( .A(n3026), .ZN(n4387) );
  INV_X1 U3067 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2728) );
  NOR2_X1 U3068 ( .A1(n2727), .A2(n2728), .ZN(n2726) );
  INV_X1 U3069 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2383) );
  MUX2_X1 U3070 ( .A(n2383), .B(REG1_REG_9__SCAN_IN), .S(n4386), .Z(n2850) );
  NAND2_X1 U3071 ( .A1(n2384), .A2(IR_REG_31__SCAN_IN), .ZN(n2385) );
  XNOR2_X1 U3072 ( .A(n2385), .B(IR_REG_10__SCAN_IN), .ZN(n3120) );
  INV_X1 U3073 ( .A(n3120), .ZN(n4520) );
  NOR2_X1 U3074 ( .A1(n2386), .A2(n4520), .ZN(n2387) );
  INV_X1 U3075 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4764) );
  XNOR2_X1 U3076 ( .A(n4520), .B(n2386), .ZN(n4416) );
  INV_X1 U3077 ( .A(n4518), .ZN(n4432) );
  INV_X1 U3078 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4575) );
  AOI22_X1 U3079 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4432), .B1(n4518), .B2(
        n4575), .ZN(n4424) );
  NAND2_X1 U3080 ( .A1(n2388), .A2(IR_REG_31__SCAN_IN), .ZN(n2389) );
  XNOR2_X1 U3081 ( .A(n2389), .B(IR_REG_12__SCAN_IN), .ZN(n3237) );
  INV_X1 U3082 ( .A(n3237), .ZN(n4517) );
  NOR2_X1 U3083 ( .A1(n2390), .A2(n4517), .ZN(n2391) );
  INV_X1 U3084 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4435) );
  NOR2_X1 U3085 ( .A1(n4435), .A2(n4434), .ZN(n4433) );
  INV_X1 U3086 ( .A(IR_REG_31__SCAN_IN), .ZN(n2483) );
  NOR2_X1 U3087 ( .A1(n2139), .A2(n2483), .ZN(n2392) );
  MUX2_X1 U3088 ( .A(n2483), .B(n2392), .S(IR_REG_13__SCAN_IN), .Z(n2394) );
  INV_X1 U3089 ( .A(n2331), .ZN(n2393) );
  NAND2_X1 U3090 ( .A1(n3300), .A2(REG1_REG_13__SCAN_IN), .ZN(n2396) );
  INV_X1 U3091 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3640) );
  NAND2_X1 U3092 ( .A1(n3408), .A2(n3640), .ZN(n2395) );
  NAND2_X1 U3093 ( .A1(n2396), .A2(n2395), .ZN(n3402) );
  NAND2_X1 U3094 ( .A1(n2331), .A2(IR_REG_31__SCAN_IN), .ZN(n2398) );
  XNOR2_X1 U3095 ( .A(n2398), .B(IR_REG_14__SCAN_IN), .ZN(n4514) );
  NOR2_X1 U3096 ( .A1(n2400), .A2(n2399), .ZN(n2401) );
  INV_X1 U3097 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4766) );
  INV_X1 U3098 ( .A(n4514), .ZN(n2399) );
  INV_X1 U3099 ( .A(n3376), .ZN(n4513) );
  INV_X1 U3100 ( .A(REG1_REG_15__SCAN_IN), .ZN(n2402) );
  AOI22_X1 U3101 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4513), .B1(n3376), .B2(
        n2402), .ZN(n4454) );
  NOR2_X1 U3102 ( .A1(n4455), .A2(n4454), .ZN(n4453) );
  NAND2_X1 U3103 ( .A1(n2403), .A2(n2322), .ZN(n2404) );
  NAND2_X1 U3104 ( .A1(n2404), .A2(n2522), .ZN(n2406) );
  XNOR2_X1 U3105 ( .A(n2406), .B(n2405), .ZN(n4512) );
  NAND2_X1 U3106 ( .A1(n2407), .A2(n4512), .ZN(n2408) );
  INV_X1 U3107 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4471) );
  XNOR2_X1 U3108 ( .A(n3427), .B(REG1_REG_17__SCAN_IN), .ZN(n4023) );
  NAND2_X1 U3109 ( .A1(n4022), .A2(n4023), .ZN(n4021) );
  OAI21_X1 U3110 ( .B1(n4385), .B2(REG1_REG_17__SCAN_IN), .A(n4021), .ZN(n4480) );
  INV_X1 U3111 ( .A(n2409), .ZN(n2410) );
  NAND2_X1 U3112 ( .A1(n2410), .A2(n4686), .ZN(n2411) );
  NAND2_X1 U3113 ( .A1(n2412), .A2(n4685), .ZN(n2523) );
  OR2_X1 U3114 ( .A1(n2412), .A2(n4685), .ZN(n2413) );
  XNOR2_X1 U3115 ( .A(n3627), .B(REG1_REG_19__SCAN_IN), .ZN(n2414) );
  XNOR2_X1 U3116 ( .A(n2415), .B(n2414), .ZN(n2444) );
  NOR2_X1 U3117 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2419)
         );
  NOR2_X1 U3118 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2418)
         );
  NOR2_X1 U3119 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2417)
         );
  NOR2_X1 U3120 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2416)
         );
  NAND2_X1 U3121 ( .A1(n2432), .A2(n4692), .ZN(n2421) );
  NAND4_X1 U3122 ( .A1(n4692), .A2(n4613), .A3(n4691), .A4(n2437), .ZN(n2427)
         );
  INV_X1 U3123 ( .A(n2427), .ZN(n2424) );
  NAND2_X1 U3124 ( .A1(n2424), .A2(n2423), .ZN(n2480) );
  INV_X1 U3125 ( .A(n2530), .ZN(n2535) );
  OR2_X1 U3126 ( .A1(n2482), .A2(n2427), .ZN(n2428) );
  NAND2_X1 U3127 ( .A1(n2428), .A2(n2522), .ZN(n2429) );
  MUX2_X1 U3128 ( .A(IR_REG_31__SCAN_IN), .B(n2429), .S(IR_REG_25__SCAN_IN), 
        .Z(n2430) );
  NAND2_X1 U3129 ( .A1(n2430), .A2(n2434), .ZN(n2531) );
  NOR2_X1 U3130 ( .A1(n2535), .A2(n2531), .ZN(n2431) );
  XNOR2_X1 U3131 ( .A(n2432), .B(n4692), .ZN(n2824) );
  NAND2_X1 U3132 ( .A1(n2824), .A2(STATE_REG_SCAN_IN), .ZN(n4509) );
  OR2_X1 U3133 ( .A1(n2824), .A2(U3149), .ZN(n3633) );
  INV_X1 U3134 ( .A(n3633), .ZN(n2433) );
  OR2_X1 U3135 ( .A1(n2759), .A2(n2433), .ZN(n2490) );
  NAND2_X1 U3136 ( .A1(n2485), .A2(IR_REG_27__SCAN_IN), .ZN(n2436) );
  NAND2_X1 U3137 ( .A1(n2440), .A2(n2522), .ZN(n2438) );
  XNOR2_X1 U3138 ( .A(n2437), .B(n2438), .ZN(n2692) );
  NAND2_X1 U3139 ( .A1(n2482), .A2(IR_REG_31__SCAN_IN), .ZN(n2439) );
  MUX2_X1 U3140 ( .A(IR_REG_31__SCAN_IN), .B(n2439), .S(IR_REG_21__SCAN_IN), 
        .Z(n2441) );
  NAND2_X1 U3141 ( .A1(n2441), .A2(n2440), .ZN(n2758) );
  NAND2_X1 U3142 ( .A1(n2824), .A2(n2735), .ZN(n2442) );
  AND2_X1 U3143 ( .A1(n2682), .A2(n2442), .ZN(n2488) );
  XNOR2_X1 U3144 ( .A(n2443), .B(IR_REG_27__SCAN_IN), .ZN(n4383) );
  INV_X1 U3145 ( .A(n4383), .ZN(n4003) );
  NAND2_X1 U3146 ( .A1(n2444), .A2(n4474), .ZN(n2497) );
  INV_X1 U3147 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2445) );
  MUX2_X1 U31480 ( .A(n2445), .B(REG2_REG_19__SCAN_IN), .S(n4384), .Z(n2478)
         );
  NAND2_X1 U31490 ( .A1(REG2_REG_18__SCAN_IN), .A2(n3425), .ZN(n2446) );
  OAI21_X1 U3150 ( .B1(REG2_REG_18__SCAN_IN), .B2(n3425), .A(n2446), .ZN(n4486) );
  NAND2_X1 U3151 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4518), .ZN(n2470) );
  INV_X1 U3152 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4791) );
  AOI22_X1 U3153 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4518), .B1(n4432), .B2(
        n4791), .ZN(n4429) );
  INV_X1 U3154 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3089) );
  INV_X1 U3155 ( .A(n4386), .ZN(n2855) );
  INV_X1 U3156 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2448) );
  AND2_X1 U3157 ( .A1(REG2_REG_0__SCAN_IN), .A2(n4603), .ZN(n4006) );
  NAND2_X1 U3158 ( .A1(n4392), .A2(REG2_REG_1__SCAN_IN), .ZN(n4014) );
  NAND2_X1 U3159 ( .A1(n4015), .A2(n4014), .ZN(n2450) );
  INV_X1 U3160 ( .A(REG2_REG_2__SCAN_IN), .ZN(n4206) );
  MUX2_X1 U3161 ( .A(REG2_REG_2__SCAN_IN), .B(n4206), .S(n2136), .Z(n2449) );
  NAND2_X1 U3162 ( .A1(n2136), .A2(REG2_REG_2__SCAN_IN), .ZN(n2451) );
  NAND2_X1 U3163 ( .A1(n4017), .A2(n2451), .ZN(n2452) );
  NAND2_X1 U3164 ( .A1(n2545), .A2(REG2_REG_3__SCAN_IN), .ZN(n2454) );
  NAND2_X1 U3165 ( .A1(n2452), .A2(n4390), .ZN(n2453) );
  NAND2_X1 U3166 ( .A1(n4404), .A2(REG2_REG_4__SCAN_IN), .ZN(n2457) );
  NAND2_X1 U3167 ( .A1(n2455), .A2(n4406), .ZN(n2456) );
  NAND2_X1 U3168 ( .A1(n2457), .A2(n2456), .ZN(n2553) );
  INV_X1 U3169 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2992) );
  MUX2_X1 U3170 ( .A(n2992), .B(REG2_REG_5__SCAN_IN), .S(n2900), .Z(n2552) );
  NAND2_X1 U3171 ( .A1(n2553), .A2(n2552), .ZN(n2551) );
  NAND2_X1 U3172 ( .A1(n4389), .A2(REG2_REG_5__SCAN_IN), .ZN(n2458) );
  NAND2_X1 U3173 ( .A1(n2562), .A2(REG2_REG_6__SCAN_IN), .ZN(n2461) );
  NAND2_X1 U3174 ( .A1(n2459), .A2(n4388), .ZN(n2460) );
  INV_X1 U3175 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2462) );
  MUX2_X1 U3176 ( .A(REG2_REG_7__SCAN_IN), .B(n2462), .S(n3024), .Z(n2463) );
  NAND2_X1 U3177 ( .A1(n3024), .A2(REG2_REG_7__SCAN_IN), .ZN(n2464) );
  AND2_X1 U3178 ( .A1(n2465), .A2(n4387), .ZN(n2466) );
  AOI21_X1 U3179 ( .B1(n2724), .B2(REG2_REG_8__SCAN_IN), .A(n2466), .ZN(n2847)
         );
  MUX2_X1 U3180 ( .A(n3089), .B(REG2_REG_9__SCAN_IN), .S(n4386), .Z(n2846) );
  INV_X1 U3181 ( .A(n2845), .ZN(n2467) );
  NAND2_X1 U3182 ( .A1(n3120), .A2(n2468), .ZN(n2469) );
  NAND2_X1 U3183 ( .A1(n4429), .A2(n4428), .ZN(n4427) );
  NAND2_X1 U3184 ( .A1(n3237), .A2(n2471), .ZN(n2472) );
  NOR2_X1 U3185 ( .A1(n2399), .A2(n2473), .ZN(n2474) );
  INV_X1 U3186 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4794) );
  INV_X1 U3187 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2475) );
  AOI22_X1 U3188 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4513), .B1(n3376), .B2(
        n2475), .ZN(n4460) );
  NOR2_X1 U3189 ( .A1(n4459), .A2(n4460), .ZN(n4458) );
  NAND2_X1 U3190 ( .A1(n2476), .A2(n4512), .ZN(n2477) );
  INV_X1 U3191 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4468) );
  XNOR2_X1 U3192 ( .A(n3427), .B(REG2_REG_17__SCAN_IN), .ZN(n4028) );
  NAND2_X1 U3193 ( .A1(n2181), .A2(n2435), .ZN(n2479) );
  NOR2_X1 U3194 ( .A1(n2486), .A2(n2483), .ZN(n2484) );
  MUX2_X1 U3195 ( .A(n2483), .B(n2484), .S(IR_REG_28__SCAN_IN), .Z(n2487) );
  NOR2_X1 U3196 ( .A1(n2487), .A2(n2513), .ZN(n4382) );
  AND2_X1 U3197 ( .A1(n4382), .A2(n4383), .ZN(n4007) );
  INV_X1 U3198 ( .A(n2488), .ZN(n2489) );
  INV_X1 U3199 ( .A(n4483), .ZN(n4465) );
  INV_X1 U3200 ( .A(ADDR_REG_19__SCAN_IN), .ZN(n4812) );
  NAND2_X1 U3201 ( .A1(n4483), .A2(ADDR_REG_19__SCAN_IN), .ZN(n2493) );
  INV_X1 U3202 ( .A(n4382), .ZN(n2763) );
  NAND2_X1 U3203 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3906) );
  INV_X1 U3204 ( .A(n3906), .ZN(n2491) );
  NAND2_X1 U3205 ( .A1(n2493), .A2(n2492), .ZN(n2494) );
  INV_X1 U3206 ( .A(DATAI_4_), .ZN(n2499) );
  MUX2_X1 U3207 ( .A(n2499), .B(n2498), .S(STATE_REG_SCAN_IN), .Z(n2500) );
  INV_X1 U3208 ( .A(n2500), .ZN(U3348) );
  NAND2_X1 U3209 ( .A1(U3149), .A2(DATAI_25_), .ZN(n2501) );
  OAI21_X1 U32100 ( .B1(n2531), .B2(U3149), .A(n2501), .ZN(U3327) );
  INV_X1 U32110 ( .A(DATAI_21_), .ZN(n4632) );
  NAND2_X1 U32120 ( .A1(n3556), .A2(STATE_REG_SCAN_IN), .ZN(n2502) );
  OAI21_X1 U32130 ( .B1(STATE_REG_SCAN_IN), .B2(n4632), .A(n2502), .ZN(U3331)
         );
  INV_X1 U32140 ( .A(DATAI_26_), .ZN(n2504) );
  NAND2_X1 U32150 ( .A1(n2530), .A2(STATE_REG_SCAN_IN), .ZN(n2503) );
  OAI21_X1 U32160 ( .B1(STATE_REG_SCAN_IN), .B2(n2504), .A(n2503), .ZN(U3326)
         );
  INV_X1 U32170 ( .A(DATAI_13_), .ZN(n2506) );
  NAND2_X1 U32180 ( .A1(n3300), .A2(STATE_REG_SCAN_IN), .ZN(n2505) );
  OAI21_X1 U32190 ( .B1(STATE_REG_SCAN_IN), .B2(n2506), .A(n2505), .ZN(U3339)
         );
  INV_X1 U32200 ( .A(DATAI_7_), .ZN(n2507) );
  INV_X1 U32210 ( .A(n3024), .ZN(n2571) );
  MUX2_X1 U32220 ( .A(n2507), .B(n2571), .S(STATE_REG_SCAN_IN), .Z(n2508) );
  INV_X1 U32230 ( .A(n2508), .ZN(U3345) );
  INV_X1 U32240 ( .A(DATAI_22_), .ZN(n2510) );
  NAND2_X1 U32250 ( .A1(n3631), .A2(STATE_REG_SCAN_IN), .ZN(n2509) );
  OAI21_X1 U32260 ( .B1(STATE_REG_SCAN_IN), .B2(n2510), .A(n2509), .ZN(U3330)
         );
  INV_X1 U32270 ( .A(DATAI_29_), .ZN(n2516) );
  NAND2_X1 U32280 ( .A1(n2586), .A2(STATE_REG_SCAN_IN), .ZN(n2515) );
  OAI21_X1 U32290 ( .B1(STATE_REG_SCAN_IN), .B2(n2516), .A(n2515), .ZN(U3323)
         );
  INV_X1 U32300 ( .A(DATAI_30_), .ZN(n4629) );
  NAND2_X1 U32310 ( .A1(n2583), .A2(STATE_REG_SCAN_IN), .ZN(n2519) );
  OAI21_X1 U32320 ( .B1(STATE_REG_SCAN_IN), .B2(n4629), .A(n2519), .ZN(U3322)
         );
  INV_X1 U32330 ( .A(DATAI_24_), .ZN(n2521) );
  NAND2_X1 U32340 ( .A1(n2534), .A2(STATE_REG_SCAN_IN), .ZN(n2520) );
  OAI21_X1 U32350 ( .B1(STATE_REG_SCAN_IN), .B2(n2521), .A(n2520), .ZN(U3328)
         );
  INV_X1 U32360 ( .A(DATAI_20_), .ZN(n2527) );
  NAND2_X1 U32370 ( .A1(n2695), .A2(STATE_REG_SCAN_IN), .ZN(n2526) );
  OAI21_X1 U32380 ( .B1(STATE_REG_SCAN_IN), .B2(n2527), .A(n2526), .ZN(U3332)
         );
  NAND2_X1 U32390 ( .A1(n2531), .A2(B_REG_SCAN_IN), .ZN(n2528) );
  MUX2_X1 U32400 ( .A(n2528), .B(B_REG_SCAN_IN), .S(n2534), .Z(n2529) );
  NAND2_X1 U32410 ( .A1(n2718), .A2(n2759), .ZN(n4507) );
  INV_X1 U32420 ( .A(D_REG_1__SCAN_IN), .ZN(n2533) );
  NAND2_X1 U32430 ( .A1(n2535), .A2(n2531), .ZN(n2733) );
  INV_X1 U32440 ( .A(n2733), .ZN(n2532) );
  AOI22_X1 U32450 ( .A1(n4507), .A2(n2533), .B1(n2532), .B2(n2752), .ZN(U3459)
         );
  INV_X1 U32460 ( .A(D_REG_0__SCAN_IN), .ZN(n2719) );
  INV_X1 U32470 ( .A(n2534), .ZN(n2536) );
  NAND2_X1 U32480 ( .A1(n2536), .A2(n2535), .ZN(n2721) );
  INV_X1 U32490 ( .A(n2721), .ZN(n2537) );
  AOI22_X1 U32500 ( .A1(n4507), .A2(n2719), .B1(n2537), .B2(n2752), .ZN(U3458)
         );
  INV_X1 U32510 ( .A(n4603), .ZN(n4669) );
  INV_X1 U32520 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2742) );
  INV_X1 U32530 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4780) );
  NAND2_X1 U32540 ( .A1(n4383), .A2(n4780), .ZN(n2538) );
  NAND2_X1 U32550 ( .A1(n4382), .A2(n2538), .ZN(n4005) );
  AOI21_X1 U32560 ( .B1(n2742), .B2(n4003), .A(n4005), .ZN(n2539) );
  XOR2_X1 U32570 ( .A(n4669), .B(n2539), .Z(n2543) );
  INV_X1 U32580 ( .A(n2540), .ZN(n2542) );
  AOI22_X1 U32590 ( .A1(n4483), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n2541) );
  OAI21_X1 U32600 ( .B1(n2543), .B2(n2542), .A(n2541), .ZN(U3240) );
  XOR2_X1 U32610 ( .A(n2544), .B(REG1_REG_3__SCAN_IN), .Z(n2547) );
  INV_X1 U32620 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2965) );
  XNOR2_X1 U32630 ( .A(n2545), .B(n2965), .ZN(n2546) );
  AOI22_X1 U32640 ( .A1(n4474), .A2(n2547), .B1(n4488), .B2(n2546), .ZN(n2549)
         );
  AOI22_X1 U32650 ( .A1(n4483), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n2548) );
  OAI211_X1 U32660 ( .C1(n2550), .C2(n4490), .A(n2549), .B(n2548), .ZN(U3243)
         );
  AND2_X1 U32670 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n2914) );
  INV_X1 U32680 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n4823) );
  OAI211_X1 U32690 ( .C1(n2553), .C2(n2552), .A(n4488), .B(n2551), .ZN(n2554)
         );
  OAI21_X1 U32700 ( .B1(n4465), .B2(n4823), .A(n2554), .ZN(n2555) );
  NOR2_X1 U32710 ( .A1(n2914), .A2(n2555), .ZN(n2560) );
  OAI211_X1 U32720 ( .C1(n2558), .C2(n2557), .A(n4474), .B(n2556), .ZN(n2559)
         );
  OAI211_X1 U32730 ( .C1(n4490), .C2(n2900), .A(n2560), .B(n2559), .ZN(U3245)
         );
  XNOR2_X1 U32740 ( .A(n2561), .B(REG1_REG_6__SCAN_IN), .ZN(n2568) );
  XOR2_X1 U32750 ( .A(REG2_REG_6__SCAN_IN), .B(n2562), .Z(n2566) );
  NOR2_X1 U32760 ( .A1(STATE_REG_SCAN_IN), .A2(n2904), .ZN(n2944) );
  AOI21_X1 U32770 ( .B1(n4483), .B2(ADDR_REG_6__SCAN_IN), .A(n2944), .ZN(n2563) );
  OAI21_X1 U32780 ( .B1(n4490), .B2(n2564), .A(n2563), .ZN(n2565) );
  AOI21_X1 U32790 ( .B1(n4488), .B2(n2566), .A(n2565), .ZN(n2567) );
  OAI21_X1 U32800 ( .B1(n2568), .B2(n4478), .A(n2567), .ZN(U3246) );
  NOR2_X1 U32810 ( .A1(n4483), .A2(U4043), .ZN(U3148) );
  INV_X1 U32820 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4571) );
  MUX2_X1 U32830 ( .A(n4571), .B(REG1_REG_7__SCAN_IN), .S(n3024), .Z(n2570) );
  XOR2_X1 U32840 ( .A(n2570), .B(n2569), .Z(n2579) );
  NOR2_X1 U32850 ( .A1(STATE_REG_SCAN_IN), .A2(n4585), .ZN(n3066) );
  NOR2_X1 U32860 ( .A1(n4490), .A2(n2571), .ZN(n2572) );
  AOI211_X1 U32870 ( .C1(n4483), .C2(ADDR_REG_7__SCAN_IN), .A(n3066), .B(n2572), .ZN(n2578) );
  MUX2_X1 U32880 ( .A(n2462), .B(REG2_REG_7__SCAN_IN), .S(n3024), .Z(n2573) );
  INV_X1 U32890 ( .A(n2573), .ZN(n2575) );
  OAI211_X1 U32900 ( .C1(n2576), .C2(n2575), .A(n2574), .B(n4488), .ZN(n2577)
         );
  OAI211_X1 U32910 ( .C1(n2579), .C2(n4478), .A(n2578), .B(n2577), .ZN(U3247)
         );
  INV_X1 U32920 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n4848) );
  INV_X1 U32930 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4753) );
  NAND2_X1 U32940 ( .A1(n3326), .A2(REG3_REG_15__SCAN_IN), .ZN(n3328) );
  INV_X1 U32950 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2648) );
  NAND2_X1 U32960 ( .A1(REG3_REG_17__SCAN_IN), .A2(REG3_REG_18__SCAN_IN), .ZN(
        n2580) );
  AND2_X1 U32970 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_20__SCAN_IN), .ZN(
        n2581) );
  INV_X1 U32980 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4862) );
  NAND2_X1 U32990 ( .A1(n3440), .A2(n4862), .ZN(n2582) );
  NAND2_X1 U33000 ( .A1(n3450), .A2(n2582), .ZN(n4163) );
  OR2_X1 U33010 ( .A1(n4163), .A2(n2679), .ZN(n2588) );
  AOI22_X1 U33020 ( .A1(n2677), .A2(REG2_REG_22__SCAN_IN), .B1(n3489), .B2(
        REG1_REG_22__SCAN_IN), .ZN(n2587) );
  OAI211_X1 U33030 ( .C1(n3445), .C2(n4753), .A(n2588), .B(n2587), .ZN(n4139)
         );
  NAND2_X1 U33040 ( .A1(n4139), .A2(U4043), .ZN(n2589) );
  OAI21_X1 U33050 ( .B1(U4043), .B2(n4848), .A(n2589), .ZN(U3572) );
  INV_X1 U33060 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n4832) );
  AOI22_X1 U33070 ( .A1(n2677), .A2(REG2_REG_8__SCAN_IN), .B1(n3489), .B2(
        REG1_REG_8__SCAN_IN), .ZN(n2592) );
  NAND2_X1 U33080 ( .A1(n2615), .A2(n4660), .ZN(n2590) );
  AND2_X1 U33090 ( .A1(n2622), .A2(n2590), .ZN(n3148) );
  AOI22_X1 U33100 ( .A1(n3488), .A2(n3148), .B1(n2133), .B2(
        REG0_REG_8__SCAN_IN), .ZN(n2591) );
  NAND2_X1 U33110 ( .A1(n3083), .A2(U4043), .ZN(n2593) );
  OAI21_X1 U33120 ( .B1(U4043), .B2(n4832), .A(n2593), .ZN(U3558) );
  INV_X1 U33130 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n4842) );
  NAND2_X1 U33140 ( .A1(n2677), .A2(REG2_REG_14__SCAN_IN), .ZN(n2598) );
  AND2_X1 U33150 ( .A1(n2602), .A2(n4658), .ZN(n2594) );
  NOR2_X1 U33160 ( .A1(n3326), .A2(n2594), .ZN(n3396) );
  NAND2_X1 U33170 ( .A1(n3488), .A2(n3396), .ZN(n2597) );
  NAND2_X1 U33180 ( .A1(n3489), .A2(REG1_REG_14__SCAN_IN), .ZN(n2596) );
  NAND2_X1 U33190 ( .A1(n2133), .A2(REG0_REG_14__SCAN_IN), .ZN(n2595) );
  NAND4_X1 U33200 ( .A1(n2598), .A2(n2597), .A3(n2596), .A4(n2595), .ZN(n3388)
         );
  NAND2_X1 U33210 ( .A1(n3388), .A2(U4043), .ZN(n2599) );
  OAI21_X1 U33220 ( .B1(U4043), .B2(n4842), .A(n2599), .ZN(U3564) );
  INV_X1 U33230 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n4843) );
  NAND2_X1 U33240 ( .A1(n2677), .A2(REG2_REG_13__SCAN_IN), .ZN(n2607) );
  OAI21_X1 U33250 ( .B1(n2656), .B2(n2601), .A(n2600), .ZN(n2603) );
  AND2_X1 U33260 ( .A1(n2603), .A2(n2602), .ZN(n3370) );
  NAND2_X1 U33270 ( .A1(n3488), .A2(n3370), .ZN(n2606) );
  NAND2_X1 U33280 ( .A1(n3489), .A2(REG1_REG_13__SCAN_IN), .ZN(n2605) );
  NAND2_X1 U33290 ( .A1(n2133), .A2(REG0_REG_13__SCAN_IN), .ZN(n2604) );
  NAND2_X1 U33300 ( .A1(n3353), .A2(U4043), .ZN(n2608) );
  OAI21_X1 U33310 ( .B1(U4043), .B2(n4843), .A(n2608), .ZN(U3563) );
  INV_X1 U33320 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n4840) );
  NAND2_X1 U33330 ( .A1(n2677), .A2(REG2_REG_12__SCAN_IN), .ZN(n2612) );
  XNOR2_X1 U33340 ( .A(n2656), .B(REG3_REG_12__SCAN_IN), .ZN(n3293) );
  NAND2_X1 U33350 ( .A1(n3488), .A2(n3293), .ZN(n2611) );
  NAND2_X1 U33360 ( .A1(n3489), .A2(REG1_REG_12__SCAN_IN), .ZN(n2610) );
  NAND2_X1 U33370 ( .A1(n2133), .A2(REG0_REG_12__SCAN_IN), .ZN(n2609) );
  NAND4_X1 U33380 ( .A1(n2612), .A2(n2611), .A3(n2610), .A4(n2609), .ZN(n3362)
         );
  NAND2_X1 U33390 ( .A1(n3362), .A2(U4043), .ZN(n2613) );
  OAI21_X1 U33400 ( .B1(U4043), .B2(n4840), .A(n2613), .ZN(U3562) );
  INV_X1 U33410 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n4829) );
  NAND2_X1 U33420 ( .A1(n2677), .A2(REG2_REG_7__SCAN_IN), .ZN(n2619) );
  OR2_X1 U33430 ( .A1(n2907), .A2(REG3_REG_7__SCAN_IN), .ZN(n2614) );
  AND2_X1 U33440 ( .A1(n2615), .A2(n2614), .ZN(n3046) );
  NAND2_X1 U33450 ( .A1(n3488), .A2(n3046), .ZN(n2618) );
  NAND2_X1 U33460 ( .A1(n3489), .A2(REG1_REG_7__SCAN_IN), .ZN(n2617) );
  NAND2_X1 U33470 ( .A1(n2133), .A2(REG0_REG_7__SCAN_IN), .ZN(n2616) );
  NAND4_X1 U33480 ( .A1(n2619), .A2(n2618), .A3(n2617), .A4(n2616), .ZN(n3058)
         );
  NAND2_X1 U33490 ( .A1(n3058), .A2(U4043), .ZN(n2620) );
  OAI21_X1 U33500 ( .B1(U4043), .B2(n4829), .A(n2620), .ZN(U3557) );
  INV_X1 U33510 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n4833) );
  NAND2_X1 U33520 ( .A1(n2677), .A2(REG2_REG_9__SCAN_IN), .ZN(n2627) );
  AND2_X1 U3353 ( .A1(n2622), .A2(n2621), .ZN(n2623) );
  NOR2_X1 U33540 ( .A1(n3072), .A2(n2623), .ZN(n3215) );
  NAND2_X1 U3355 ( .A1(n3488), .A2(n3215), .ZN(n2626) );
  NAND2_X1 U3356 ( .A1(n3489), .A2(REG1_REG_9__SCAN_IN), .ZN(n2625) );
  NAND2_X1 U3357 ( .A1(n2133), .A2(REG0_REG_9__SCAN_IN), .ZN(n2624) );
  NAND4_X1 U3358 ( .A1(n2627), .A2(n2626), .A3(n2625), .A4(n2624), .ZN(n3202)
         );
  NAND2_X1 U3359 ( .A1(n3202), .A2(U4043), .ZN(n2628) );
  OAI21_X1 U3360 ( .B1(U4043), .B2(n4833), .A(n2628), .ZN(U3559) );
  INV_X1 U3361 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4845) );
  AOI22_X1 U3362 ( .A1(n2677), .A2(REG2_REG_17__SCAN_IN), .B1(n3489), .B2(
        REG1_REG_17__SCAN_IN), .ZN(n2630) );
  XNOR2_X1 U3363 ( .A(n3417), .B(REG3_REG_17__SCAN_IN), .ZN(n3732) );
  AOI22_X1 U3364 ( .A1(n3488), .A2(n3732), .B1(n2133), .B2(
        REG0_REG_17__SCAN_IN), .ZN(n2629) );
  NAND2_X1 U3365 ( .A1(n3743), .A2(U4043), .ZN(n2631) );
  OAI21_X1 U3366 ( .B1(U4043), .B2(n4845), .A(n2631), .ZN(U3567) );
  INV_X1 U3367 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n4830) );
  INV_X1 U3368 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2632) );
  NAND2_X1 U3369 ( .A1(n3488), .A2(n2632), .ZN(n2636) );
  NAND2_X1 U3370 ( .A1(n2677), .A2(REG2_REG_3__SCAN_IN), .ZN(n2635) );
  NAND2_X1 U3371 ( .A1(n2680), .A2(REG1_REG_3__SCAN_IN), .ZN(n2634) );
  NAND2_X1 U3372 ( .A1(n2133), .A2(REG0_REG_3__SCAN_IN), .ZN(n2633) );
  NAND2_X1 U3373 ( .A1(n4208), .A2(U4043), .ZN(n2637) );
  OAI21_X1 U3374 ( .B1(U4043), .B2(n4830), .A(n2637), .ZN(U3553) );
  INV_X1 U3375 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n4859) );
  INV_X1 U3376 ( .A(REG2_REG_31__SCAN_IN), .ZN(n2641) );
  NAND2_X1 U3377 ( .A1(n3489), .A2(REG1_REG_31__SCAN_IN), .ZN(n2640) );
  NAND2_X1 U3378 ( .A1(n2133), .A2(REG0_REG_31__SCAN_IN), .ZN(n2639) );
  OAI211_X1 U3379 ( .C1(n2638), .C2(n2641), .A(n2640), .B(n2639), .ZN(n4221)
         );
  NAND2_X1 U3380 ( .A1(n4221), .A2(U4043), .ZN(n2642) );
  OAI21_X1 U3381 ( .B1(U4043), .B2(n4859), .A(n2642), .ZN(U3581) );
  INV_X1 U3382 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n4849) );
  NOR2_X1 U3383 ( .A1(n3419), .A2(REG3_REG_19__SCAN_IN), .ZN(n2643) );
  NOR2_X1 U3384 ( .A1(n3438), .A2(n2643), .ZN(n3911) );
  NAND2_X1 U3385 ( .A1(n3911), .A2(n3488), .ZN(n2646) );
  AOI22_X1 U3386 ( .A1(n2677), .A2(REG2_REG_19__SCAN_IN), .B1(n3489), .B2(
        REG1_REG_19__SCAN_IN), .ZN(n2645) );
  NAND2_X1 U3387 ( .A1(n2133), .A2(REG0_REG_19__SCAN_IN), .ZN(n2644) );
  NAND2_X1 U3388 ( .A1(n4295), .A2(U4043), .ZN(n2647) );
  OAI21_X1 U3389 ( .B1(U4043), .B2(n4849), .A(n2647), .ZN(U3569) );
  INV_X1 U3390 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n4846) );
  NAND2_X1 U3391 ( .A1(n2677), .A2(REG2_REG_16__SCAN_IN), .ZN(n2653) );
  NAND2_X1 U3392 ( .A1(n3328), .A2(n2648), .ZN(n2649) );
  AND2_X1 U3393 ( .A1(n3417), .A2(n2649), .ZN(n3693) );
  NAND2_X1 U3394 ( .A1(n3488), .A2(n3693), .ZN(n2652) );
  NAND2_X1 U3395 ( .A1(n3489), .A2(REG1_REG_16__SCAN_IN), .ZN(n2651) );
  NAND2_X1 U3396 ( .A1(n2133), .A2(REG0_REG_16__SCAN_IN), .ZN(n2650) );
  NAND4_X1 U3397 ( .A1(n2653), .A2(n2652), .A3(n2651), .A4(n2650), .ZN(n4328)
         );
  NAND2_X1 U3398 ( .A1(n4328), .A2(U4043), .ZN(n2654) );
  OAI21_X1 U3399 ( .B1(U4043), .B2(n4846), .A(n2654), .ZN(U3566) );
  INV_X1 U3400 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n4839) );
  NAND2_X1 U3401 ( .A1(n2677), .A2(REG2_REG_11__SCAN_IN), .ZN(n2660) );
  OR2_X1 U3402 ( .A1(n3074), .A2(REG3_REG_11__SCAN_IN), .ZN(n2655) );
  AND2_X1 U3403 ( .A1(n2656), .A2(n2655), .ZN(n3192) );
  NAND2_X1 U3404 ( .A1(n3488), .A2(n3192), .ZN(n2659) );
  NAND2_X1 U3405 ( .A1(n3489), .A2(REG1_REG_11__SCAN_IN), .ZN(n2658) );
  NAND2_X1 U3406 ( .A1(n2133), .A2(REG0_REG_11__SCAN_IN), .ZN(n2657) );
  NAND4_X1 U3407 ( .A1(n2660), .A2(n2659), .A3(n2658), .A4(n2657), .ZN(n3262)
         );
  NAND2_X1 U3408 ( .A1(n3262), .A2(U4043), .ZN(n2661) );
  OAI21_X1 U3409 ( .B1(U4043), .B2(n4839), .A(n2661), .ZN(U3561) );
  INV_X1 U3410 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n4827) );
  NAND2_X1 U3411 ( .A1(n3488), .A2(REG3_REG_0__SCAN_IN), .ZN(n2665) );
  NAND2_X1 U3412 ( .A1(n2677), .A2(REG2_REG_0__SCAN_IN), .ZN(n2664) );
  NAND2_X1 U3413 ( .A1(n2681), .A2(REG0_REG_0__SCAN_IN), .ZN(n2663) );
  NAND2_X1 U3414 ( .A1(n2680), .A2(REG1_REG_0__SCAN_IN), .ZN(n2662) );
  INV_X1 U3415 ( .A(n2688), .ZN(n2887) );
  NAND2_X1 U3416 ( .A1(n2688), .A2(U4043), .ZN(n2666) );
  OAI21_X1 U3417 ( .B1(U4043), .B2(n4827), .A(n2666), .ZN(U3550) );
  INV_X1 U3418 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n4858) );
  NAND2_X1 U3419 ( .A1(n3489), .A2(REG1_REG_30__SCAN_IN), .ZN(n2668) );
  NAND2_X1 U3420 ( .A1(n2133), .A2(REG0_REG_30__SCAN_IN), .ZN(n2667) );
  OAI211_X1 U3421 ( .C1(n2638), .C2(n4809), .A(n2668), .B(n2667), .ZN(n4042)
         );
  NAND2_X1 U3422 ( .A1(n4042), .A2(U4043), .ZN(n2669) );
  OAI21_X1 U3423 ( .B1(U4043), .B2(n4858), .A(n2669), .ZN(U3580) );
  INV_X1 U3424 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n4826) );
  NAND2_X1 U3425 ( .A1(n2680), .A2(REG1_REG_2__SCAN_IN), .ZN(n2672) );
  NAND2_X1 U3426 ( .A1(n2681), .A2(REG0_REG_2__SCAN_IN), .ZN(n2671) );
  NAND2_X1 U3427 ( .A1(n3488), .A2(REG3_REG_2__SCAN_IN), .ZN(n2674) );
  NAND2_X1 U3428 ( .A1(n2866), .A2(U4043), .ZN(n2676) );
  OAI21_X1 U3429 ( .B1(U4043), .B2(n4826), .A(n2676), .ZN(U3552) );
  INV_X1 U3430 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2678) );
  NAND2_X1 U3431 ( .A1(n2681), .A2(REG0_REG_1__SCAN_IN), .ZN(n2683) );
  AND2_X1 U3432 ( .A1(n2863), .A2(n2683), .ZN(n2686) );
  NAND2_X1 U3433 ( .A1(n3554), .A2(n2870), .ZN(n2689) );
  MUX2_X1 U3434 ( .A(n4603), .B(DATAI_0_), .S(n2682), .Z(n2745) );
  AND2_X1 U3435 ( .A1(n2688), .A2(n2745), .ZN(n2690) );
  NAND2_X1 U3436 ( .A1(n2689), .A2(n2690), .ZN(n2865) );
  AND2_X1 U3437 ( .A1(n2865), .A2(n2691), .ZN(n2971) );
  INV_X1 U3438 ( .A(n2879), .ZN(n2881) );
  OAI21_X1 U3439 ( .B1(n2888), .B2(n4493), .A(n2881), .ZN(n2974) );
  AND2_X1 U3440 ( .A1(n2692), .A2(n2758), .ZN(n4491) );
  NOR2_X1 U3441 ( .A1(n2974), .A2(n4551), .ZN(n2704) );
  NAND2_X1 U3442 ( .A1(n2887), .A2(n2745), .ZN(n3553) );
  NAND2_X1 U3443 ( .A1(n2872), .A2(n2693), .ZN(n2699) );
  NAND2_X1 U3444 ( .A1(n2695), .A2(n3556), .ZN(n3409) );
  NAND2_X1 U3445 ( .A1(n4384), .A2(n3631), .ZN(n2694) );
  NAND2_X1 U3446 ( .A1(n2688), .A2(n4321), .ZN(n2697) );
  NAND2_X1 U3447 ( .A1(n2763), .A2(n2735), .ZN(n4497) );
  NAND2_X1 U3448 ( .A1(n2866), .A2(n4327), .ZN(n2696) );
  OAI211_X1 U3449 ( .C1(n4315), .C2(n2888), .A(n2697), .B(n2696), .ZN(n2698)
         );
  AOI21_X1 U3450 ( .B1(n2699), .B2(n4495), .A(n2698), .ZN(n2703) );
  XNOR2_X1 U3451 ( .A(n2741), .B(n3631), .ZN(n2701) );
  NAND2_X1 U3452 ( .A1(n2701), .A2(n3627), .ZN(n3364) );
  INV_X1 U3453 ( .A(n3364), .ZN(n4496) );
  NAND2_X1 U3454 ( .A1(n2971), .A2(n4496), .ZN(n2702) );
  NAND2_X1 U3455 ( .A1(n2703), .A2(n2702), .ZN(n2969) );
  AOI211_X1 U3456 ( .C1(n2971), .C2(n4536), .A(n2704), .B(n2969), .ZN(n4527)
         );
  NAND2_X1 U3457 ( .A1(n2951), .A2(n2733), .ZN(n2717) );
  NAND2_X1 U34580 ( .A1(n2700), .A2(n3627), .ZN(n2705) );
  NAND2_X1 U34590 ( .A1(n2705), .A2(n2735), .ZN(n2750) );
  INV_X1 U3460 ( .A(D_REG_18__SCAN_IN), .ZN(n4717) );
  INV_X1 U3461 ( .A(D_REG_22__SCAN_IN), .ZN(n4719) );
  INV_X1 U3462 ( .A(D_REG_27__SCAN_IN), .ZN(n4722) );
  INV_X1 U3463 ( .A(D_REG_3__SCAN_IN), .ZN(n4702) );
  NAND4_X1 U3464 ( .A1(n4717), .A2(n4719), .A3(n4722), .A4(n4702), .ZN(n2706)
         );
  NOR4_X1 U3465 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_31__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(n2706), .ZN(n4600) );
  NOR4_X1 U3466 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2708) );
  NOR3_X1 U34670 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .ZN(n2707) );
  NAND3_X1 U3468 ( .A1(n4600), .A2(n2708), .A3(n2707), .ZN(n2714) );
  NOR4_X1 U34690 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_26__SCAN_IN), .ZN(n2712) );
  NOR4_X1 U3470 ( .A1(D_REG_24__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_11__SCAN_IN), .ZN(n2711) );
  NOR4_X1 U34710 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_15__SCAN_IN), .A3(
        D_REG_19__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2710) );
  NOR4_X1 U3472 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2709) );
  NAND4_X1 U34730 ( .A1(n2712), .A2(n2711), .A3(n2710), .A4(n2709), .ZN(n2713)
         );
  NOR2_X1 U3474 ( .A1(n2714), .A2(n2713), .ZN(n2715) );
  NAND2_X1 U34750 ( .A1(n4536), .A2(n2758), .ZN(n2716) );
  NAND4_X1 U3476 ( .A1(n2717), .A2(n2953), .A3(n2734), .A4(n2716), .ZN(n2878)
         );
  INV_X1 U34770 ( .A(n2718), .ZN(n2720) );
  NAND2_X1 U3478 ( .A1(n2720), .A2(n2719), .ZN(n2722) );
  NAND2_X1 U34790 ( .A1(n2722), .A2(n2721), .ZN(n2952) );
  NAND2_X1 U3480 ( .A1(n4574), .A2(REG1_REG_1__SCAN_IN), .ZN(n2723) );
  OAI21_X1 U34810 ( .B1(n4527), .B2(n4574), .A(n2723), .ZN(U3519) );
  XNOR2_X1 U3482 ( .A(n2724), .B(REG2_REG_8__SCAN_IN), .ZN(n2732) );
  INV_X1 U34830 ( .A(n4488), .ZN(n4445) );
  INV_X1 U3484 ( .A(ADDR_REG_8__SCAN_IN), .ZN(n2725) );
  OR2_X1 U34850 ( .A1(n4660), .A2(STATE_REG_SCAN_IN), .ZN(n3143) );
  OAI21_X1 U3486 ( .B1(n4465), .B2(n2725), .A(n3143), .ZN(n2730) );
  AOI211_X1 U34870 ( .C1(n2728), .C2(n2727), .A(n4478), .B(n2726), .ZN(n2729)
         );
  AOI211_X1 U3488 ( .C1(n4450), .C2(n4387), .A(n2730), .B(n2729), .ZN(n2731)
         );
  OAI21_X1 U34890 ( .B1(n2732), .B2(n4445), .A(n2731), .ZN(U3248) );
  INV_X1 U3490 ( .A(n2952), .ZN(n2877) );
  NAND2_X1 U34910 ( .A1(n4384), .A2(n4491), .ZN(n2737) );
  INV_X1 U3492 ( .A(n2735), .ZN(n2736) );
  NAND2_X1 U34930 ( .A1(n2737), .A2(n2736), .ZN(n2738) );
  OR2_X1 U3494 ( .A1(n4326), .A2(n2738), .ZN(n2748) );
  INV_X1 U34950 ( .A(n2759), .ZN(n2756) );
  NOR2_X1 U3496 ( .A1(n2748), .A2(n2756), .ZN(n2739) );
  NOR2_X2 U34970 ( .A1(n2744), .A2(n2741), .ZN(n2784) );
  OR2_X1 U3498 ( .A1(n2740), .A2(n2742), .ZN(n2743) );
  NAND2_X1 U34990 ( .A1(n2688), .A2(n3830), .ZN(n2747) );
  AOI22_X1 U3500 ( .A1(n2784), .A2(n2745), .B1(n2744), .B2(n4603), .ZN(n2746)
         );
  NAND2_X1 U35010 ( .A1(n2747), .A2(n2746), .ZN(n2766) );
  XNOR2_X1 U3502 ( .A(n2767), .B(n2766), .ZN(n4004) );
  INV_X1 U35030 ( .A(n2796), .ZN(n2757) );
  NAND2_X1 U3504 ( .A1(n2748), .A2(n4315), .ZN(n2749) );
  NAND2_X1 U35050 ( .A1(n2757), .A2(n2749), .ZN(n2751) );
  NAND2_X1 U35060 ( .A1(n2751), .A2(n2750), .ZN(n2826) );
  INV_X1 U35070 ( .A(n2826), .ZN(n2755) );
  NAND2_X1 U35080 ( .A1(n3627), .A2(n3631), .ZN(n2768) );
  INV_X1 U35090 ( .A(n2768), .ZN(n2753) );
  NAND2_X1 U35100 ( .A1(n2753), .A2(n2752), .ZN(n2754) );
  NOR2_X1 U35110 ( .A1(n3837), .A2(n2754), .ZN(n3629) );
  NAND2_X1 U35120 ( .A1(n2757), .A2(n3629), .ZN(n2827) );
  NAND3_X1 U35130 ( .A1(n2755), .A2(n2759), .A3(n2827), .ZN(n2891) );
  NOR3_X1 U35140 ( .A1(n2757), .A2(n4315), .A3(n2756), .ZN(n2761) );
  AND2_X1 U35150 ( .A1(n2759), .A2(n2758), .ZN(n2760) );
  OR2_X1 U35160 ( .A1(n2761), .A2(n4502), .ZN(n2912) );
  INV_X1 U35170 ( .A(n2762), .ZN(n4498) );
  NAND3_X1 U35180 ( .A1(n2796), .A2(n3629), .A3(n2763), .ZN(n3982) );
  OAI22_X1 U35190 ( .A1(n3980), .A2(n4493), .B1(n4498), .B2(n3982), .ZN(n2764)
         );
  AOI21_X1 U35200 ( .B1(REG3_REG_0__SCAN_IN), .B2(n2891), .A(n2764), .ZN(n2765) );
  OAI21_X1 U35210 ( .B1(n3988), .B2(n4004), .A(n2765), .ZN(U3229) );
  NAND2_X1 U35220 ( .A1(n2767), .A2(n2766), .ZN(n2771) );
  NAND2_X2 U35230 ( .A1(n2741), .A2(n2768), .ZN(n2805) );
  NAND2_X1 U35240 ( .A1(n2769), .A2(n3725), .ZN(n2770) );
  NAND2_X1 U35250 ( .A1(n2771), .A2(n2770), .ZN(n2886) );
  NAND2_X1 U35260 ( .A1(n2762), .A2(n2784), .ZN(n2773) );
  NAND2_X1 U35270 ( .A1(n2863), .A2(n3843), .ZN(n2772) );
  AND2_X1 U35280 ( .A1(n2784), .A2(n2863), .ZN(n2775) );
  XNOR2_X1 U35290 ( .A(n2778), .B(n2776), .ZN(n2885) );
  NAND2_X1 U35300 ( .A1(n2886), .A2(n2885), .ZN(n2780) );
  INV_X1 U35310 ( .A(n2776), .ZN(n2777) );
  NAND2_X1 U35320 ( .A1(n2778), .A2(n2777), .ZN(n2779) );
  NAND2_X1 U35330 ( .A1(n2780), .A2(n2779), .ZN(n2791) );
  NAND2_X1 U35340 ( .A1(n2866), .A2(n2784), .ZN(n2782) );
  MUX2_X1 U35350 ( .A(n2136), .B(DATAI_2_), .S(n2682), .Z(n4212) );
  NAND2_X1 U35360 ( .A1(n4212), .A2(n3843), .ZN(n2781) );
  NAND2_X1 U35370 ( .A1(n2782), .A2(n2781), .ZN(n2783) );
  XNOR2_X1 U35380 ( .A(n2783), .B(n3725), .ZN(n2786) );
  AND2_X1 U35390 ( .A1(n2784), .A2(n4212), .ZN(n2785) );
  AOI21_X1 U35400 ( .B1(n2866), .B2(n3830), .A(n2785), .ZN(n2787) );
  NAND2_X1 U35410 ( .A1(n2786), .A2(n2787), .ZN(n2801) );
  INV_X1 U35420 ( .A(n2786), .ZN(n2789) );
  INV_X1 U35430 ( .A(n2787), .ZN(n2788) );
  NAND2_X1 U35440 ( .A1(n2789), .A2(n2788), .ZN(n2790) );
  NAND2_X1 U35450 ( .A1(n2801), .A2(n2790), .ZN(n2795) );
  INV_X1 U35460 ( .A(n2791), .ZN(n2793) );
  NAND2_X1 U35470 ( .A1(n2793), .A2(n2792), .ZN(n2802) );
  INV_X1 U35480 ( .A(n2802), .ZN(n2794) );
  AOI21_X1 U35490 ( .B1(n2791), .B2(n2795), .A(n2794), .ZN(n2800) );
  OAI22_X1 U35500 ( .A1(n2981), .A2(n3982), .B1(n3949), .B2(n4498), .ZN(n2798)
         );
  NOR2_X1 U35510 ( .A1(n3980), .A2(n2948), .ZN(n2797) );
  AOI211_X1 U35520 ( .C1(REG3_REG_2__SCAN_IN), .C2(n2891), .A(n2798), .B(n2797), .ZN(n2799) );
  OAI21_X1 U35530 ( .B1(n2800), .B2(n3988), .A(n2799), .ZN(U3234) );
  NAND2_X1 U35540 ( .A1(n2802), .A2(n2801), .ZN(n2856) );
  NAND2_X1 U35550 ( .A1(n4208), .A2(n2784), .ZN(n2804) );
  MUX2_X1 U35560 ( .A(n4390), .B(DATAI_3_), .S(n2682), .Z(n2977) );
  NAND2_X1 U35570 ( .A1(n2977), .A2(n3843), .ZN(n2803) );
  NAND2_X1 U35580 ( .A1(n2804), .A2(n2803), .ZN(n2806) );
  XNOR2_X1 U35590 ( .A(n2806), .B(n2805), .ZN(n2817) );
  AND2_X1 U35600 ( .A1(n2784), .A2(n2977), .ZN(n2807) );
  AOI21_X1 U35610 ( .B1(n4208), .B2(n3830), .A(n2807), .ZN(n2818) );
  XNOR2_X1 U35620 ( .A(n2817), .B(n2818), .ZN(n2857) );
  NAND2_X1 U35630 ( .A1(n2856), .A2(n2857), .ZN(n2821) );
  NAND2_X1 U35640 ( .A1(n2677), .A2(REG2_REG_4__SCAN_IN), .ZN(n2812) );
  NAND2_X1 U35650 ( .A1(n2133), .A2(REG0_REG_4__SCAN_IN), .ZN(n2811) );
  NAND2_X1 U35660 ( .A1(n2680), .A2(REG1_REG_4__SCAN_IN), .ZN(n2810) );
  NOR2_X1 U35670 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2808) );
  NOR2_X1 U35680 ( .A1(n2829), .A2(n2808), .ZN(n3164) );
  NAND2_X1 U35690 ( .A1(n3488), .A2(n3164), .ZN(n2809) );
  NAND2_X1 U35700 ( .A1(n2983), .A2(n2784), .ZN(n2814) );
  MUX2_X1 U35710 ( .A(n4406), .B(DATAI_4_), .S(n2682), .Z(n2984) );
  NAND2_X1 U35720 ( .A1(n2984), .A2(n3843), .ZN(n2813) );
  NAND2_X1 U35730 ( .A1(n2814), .A2(n2813), .ZN(n2815) );
  XNOR2_X1 U35740 ( .A(n2815), .B(n2805), .ZN(n2896) );
  AND2_X1 U35750 ( .A1(n2784), .A2(n2984), .ZN(n2816) );
  AOI21_X1 U35760 ( .B1(n2983), .B2(n3830), .A(n2816), .ZN(n2894) );
  XNOR2_X1 U35770 ( .A(n2896), .B(n2894), .ZN(n2822) );
  INV_X1 U35780 ( .A(n2817), .ZN(n2819) );
  NAND2_X1 U35790 ( .A1(n2819), .A2(n2818), .ZN(n2823) );
  AND2_X1 U35800 ( .A1(n2822), .A2(n2823), .ZN(n2820) );
  INV_X1 U35810 ( .A(n3988), .ZN(n3966) );
  NAND2_X1 U3582 ( .A1(n2898), .A2(n3966), .ZN(n2837) );
  AOI21_X1 U3583 ( .B1(n2821), .B2(n2823), .A(n2822), .ZN(n2836) );
  NAND2_X1 U3584 ( .A1(n2740), .A2(n2824), .ZN(n2825) );
  OAI21_X1 U3585 ( .B1(n2826), .B2(n2825), .A(STATE_REG_SCAN_IN), .ZN(n2828)
         );
  AOI22_X1 U3586 ( .A1(n2677), .A2(REG2_REG_5__SCAN_IN), .B1(n3489), .B2(
        REG1_REG_5__SCAN_IN), .ZN(n2832) );
  OAI21_X1 U3587 ( .B1(n2829), .B2(REG3_REG_5__SCAN_IN), .A(n2905), .ZN(n2830)
         );
  INV_X1 U3588 ( .A(n2830), .ZN(n2994) );
  AOI22_X1 U3589 ( .A1(n3488), .A2(n2994), .B1(n2133), .B2(REG0_REG_5__SCAN_IN), .ZN(n2831) );
  NAND2_X1 U3590 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n4407) );
  OAI21_X1 U3591 ( .B1(n3982), .B2(n3155), .A(n4407), .ZN(n2834) );
  OAI22_X1 U3592 ( .A1(n3980), .A2(n3154), .B1(n2981), .B2(n3949), .ZN(n2833)
         );
  AOI211_X1 U3593 ( .C1(n3164), .C2(n3985), .A(n2834), .B(n2833), .ZN(n2835)
         );
  OAI21_X1 U3594 ( .B1(n2837), .B2(n2836), .A(n2835), .ZN(U3227) );
  INV_X1 U3595 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n4855) );
  INV_X1 U3596 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3899) );
  INV_X1 U3597 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4661) );
  AND2_X1 U3598 ( .A1(n3452), .A2(n4661), .ZN(n2838) );
  INV_X1 U3599 ( .A(REG2_REG_24__SCAN_IN), .ZN(n2841) );
  NAND2_X1 U3600 ( .A1(n3489), .A2(REG1_REG_24__SCAN_IN), .ZN(n2840) );
  NAND2_X1 U3601 ( .A1(n2133), .A2(REG0_REG_24__SCAN_IN), .ZN(n2839) );
  OAI211_X1 U3602 ( .C1(n2638), .C2(n2841), .A(n2840), .B(n2839), .ZN(n2842)
         );
  INV_X1 U3603 ( .A(n2842), .ZN(n2843) );
  NAND2_X1 U3604 ( .A1(n3862), .A2(U4043), .ZN(n2844) );
  OAI21_X1 U3605 ( .B1(U4043), .B2(n4855), .A(n2844), .ZN(U3574) );
  AOI211_X1 U3606 ( .C1(n2847), .C2(n2846), .A(n4445), .B(n2845), .ZN(n2848)
         );
  INV_X1 U3607 ( .A(n2848), .ZN(n2854) );
  AND2_X1 U3608 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n3214) );
  AOI211_X1 U3609 ( .C1(n2851), .C2(n2850), .A(n2849), .B(n4478), .ZN(n2852)
         );
  AOI211_X1 U3610 ( .C1(n4483), .C2(ADDR_REG_9__SCAN_IN), .A(n3214), .B(n2852), 
        .ZN(n2853) );
  OAI211_X1 U3611 ( .C1(n4490), .C2(n2855), .A(n2854), .B(n2853), .ZN(U3249)
         );
  OAI21_X1 U3612 ( .B1(n2857), .B2(n2856), .A(n2821), .ZN(n2858) );
  NAND2_X1 U3613 ( .A1(n2858), .A2(n3966), .ZN(n2862) );
  INV_X1 U3614 ( .A(n2866), .ZN(n2960) );
  OAI22_X1 U3615 ( .A1(n2960), .A2(n3949), .B1(n3982), .B2(n2989), .ZN(n2860)
         );
  MUX2_X1 U3616 ( .A(n3985), .B(U3149), .S(REG3_REG_3__SCAN_IN), .Z(n2859) );
  AOI211_X1 U3617 ( .C1(n2977), .C2(n2912), .A(n2860), .B(n2859), .ZN(n2861)
         );
  NAND2_X1 U3618 ( .A1(n2862), .A2(n2861), .ZN(U3215) );
  NAND2_X1 U3619 ( .A1(n2762), .A2(n2863), .ZN(n2864) );
  NAND2_X1 U3620 ( .A1(n2866), .A2(n2948), .ZN(n3561) );
  NAND2_X1 U3621 ( .A1(n3558), .A2(n3561), .ZN(n2867) );
  OAI21_X1 U3622 ( .B1(n2868), .B2(n2867), .A(n2950), .ZN(n4214) );
  AOI22_X1 U3623 ( .A1(n4208), .A2(n4327), .B1(n4212), .B2(n4326), .ZN(n2869)
         );
  OAI21_X1 U3624 ( .B1(n4498), .B2(n4330), .A(n2869), .ZN(n2876) );
  NAND2_X1 U3625 ( .A1(n2872), .A2(n2870), .ZN(n2871) );
  NAND2_X1 U3626 ( .A1(n2871), .A2(n3530), .ZN(n2957) );
  NAND3_X1 U3627 ( .A1(n2867), .A2(n2870), .A3(n2872), .ZN(n2873) );
  AOI21_X1 U3628 ( .B1(n2957), .B2(n2873), .A(n4297), .ZN(n2874) );
  AOI21_X1 U3629 ( .B1(n4214), .B2(n4496), .A(n2874), .ZN(n4205) );
  INV_X1 U3630 ( .A(n4205), .ZN(n2875) );
  AOI211_X1 U3631 ( .C1(n4536), .C2(n4214), .A(n2876), .B(n2875), .ZN(n2919)
         );
  NAND2_X1 U3632 ( .A1(n2879), .A2(n2948), .ZN(n2964) );
  INV_X1 U3633 ( .A(n2964), .ZN(n2880) );
  AOI21_X1 U3634 ( .B1(n4212), .B2(n2881), .A(n2880), .ZN(n4213) );
  INV_X2 U3635 ( .A(n4563), .ZN(n4565) );
  INV_X1 U3636 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2882) );
  NOR2_X1 U3637 ( .A1(n4565), .A2(n2882), .ZN(n2883) );
  AOI21_X1 U3638 ( .B1(n4213), .B2(n4346), .A(n2883), .ZN(n2884) );
  OAI21_X1 U3639 ( .B1(n2919), .B2(n4563), .A(n2884), .ZN(U3471) );
  XNOR2_X1 U3640 ( .A(n2886), .B(n2885), .ZN(n2893) );
  OAI22_X1 U3641 ( .A1(n2887), .A2(n3949), .B1(n3982), .B2(n2960), .ZN(n2890)
         );
  NOR2_X1 U3642 ( .A1(n3980), .A2(n2888), .ZN(n2889) );
  AOI211_X1 U3643 ( .C1(REG3_REG_1__SCAN_IN), .C2(n2891), .A(n2890), .B(n2889), 
        .ZN(n2892) );
  OAI21_X1 U3644 ( .B1(n2893), .B2(n3988), .A(n2892), .ZN(U3219) );
  INV_X1 U3645 ( .A(n2894), .ZN(n2895) );
  NAND2_X1 U3646 ( .A1(n2896), .A2(n2895), .ZN(n2897) );
  INV_X1 U3647 ( .A(DATAI_5_), .ZN(n2899) );
  MUX2_X1 U3648 ( .A(n2900), .B(n2899), .S(n2682), .Z(n2997) );
  OAI22_X1 U3649 ( .A1(n3155), .A2(n3837), .B1(n3835), .B2(n2997), .ZN(n2901)
         );
  XNOR2_X1 U3650 ( .A(n2901), .B(n3725), .ZN(n2929) );
  OR2_X1 U3651 ( .A1(n3155), .A2(n3838), .ZN(n2903) );
  NAND2_X1 U3652 ( .A1(n3000), .A2(n3825), .ZN(n2902) );
  NAND2_X1 U3653 ( .A1(n2903), .A2(n2902), .ZN(n2930) );
  XNOR2_X1 U3654 ( .A(n2929), .B(n2930), .ZN(n2927) );
  XNOR2_X1 U3655 ( .A(n2928), .B(n2927), .ZN(n2917) );
  INV_X1 U3656 ( .A(n3982), .ZN(n3970) );
  NAND2_X1 U3657 ( .A1(n2677), .A2(REG2_REG_6__SCAN_IN), .ZN(n2911) );
  AND2_X1 U3658 ( .A1(n2905), .A2(n2904), .ZN(n2906) );
  NOR2_X1 U3659 ( .A1(n2907), .A2(n2906), .ZN(n3094) );
  NAND2_X1 U3660 ( .A1(n3488), .A2(n3094), .ZN(n2910) );
  NAND2_X1 U3661 ( .A1(n3489), .A2(REG1_REG_6__SCAN_IN), .ZN(n2909) );
  NAND2_X1 U3662 ( .A1(n2133), .A2(REG0_REG_6__SCAN_IN), .ZN(n2908) );
  NAND4_X1 U3663 ( .A1(n2911), .A2(n2910), .A3(n2909), .A4(n2908), .ZN(n3992)
         );
  INV_X2 U3664 ( .A(n2912), .ZN(n3980) );
  OAI22_X1 U3665 ( .A1(n3980), .A2(n2997), .B1(n2989), .B2(n3949), .ZN(n2913)
         );
  AOI211_X1 U3666 ( .C1(n3970), .C2(n3992), .A(n2914), .B(n2913), .ZN(n2916)
         );
  NAND2_X1 U3667 ( .A1(n3985), .A2(n2994), .ZN(n2915) );
  OAI211_X1 U3668 ( .C1(n2917), .C2(n3988), .A(n2916), .B(n2915), .ZN(U3224)
         );
  AOI22_X1 U3669 ( .A1(n4244), .A2(n4213), .B1(n4574), .B2(REG1_REG_2__SCAN_IN), .ZN(n2918) );
  OAI21_X1 U3670 ( .B1(n2919), .B2(n4574), .A(n2918), .ZN(U3520) );
  INV_X1 U3671 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n4856) );
  AND2_X1 U3672 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2920) );
  AOI21_X1 U3673 ( .B1(n3466), .B2(REG3_REG_25__SCAN_IN), .A(
        REG3_REG_26__SCAN_IN), .ZN(n2921) );
  INV_X1 U3674 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4089) );
  NAND2_X1 U3675 ( .A1(n3489), .A2(REG1_REG_26__SCAN_IN), .ZN(n2923) );
  NAND2_X1 U3676 ( .A1(n2133), .A2(REG0_REG_26__SCAN_IN), .ZN(n2922) );
  OAI211_X1 U3677 ( .C1(n2638), .C2(n4089), .A(n2923), .B(n2922), .ZN(n2924)
         );
  INV_X1 U3678 ( .A(n2924), .ZN(n2925) );
  NAND2_X1 U3679 ( .A1(n4249), .A2(U4043), .ZN(n2926) );
  OAI21_X1 U3680 ( .B1(U4043), .B2(n4856), .A(n2926), .ZN(U3576) );
  INV_X1 U3681 ( .A(n2929), .ZN(n2931) );
  NAND2_X1 U3682 ( .A1(n3992), .A2(n3825), .ZN(n2933) );
  MUX2_X1 U3683 ( .A(n4388), .B(DATAI_6_), .S(n2682), .Z(n3020) );
  NAND2_X1 U3684 ( .A1(n3020), .A2(n3843), .ZN(n2932) );
  NAND2_X1 U3685 ( .A1(n2933), .A2(n2932), .ZN(n2934) );
  XNOR2_X1 U3686 ( .A(n2934), .B(n2805), .ZN(n2940) );
  INV_X1 U3687 ( .A(n2940), .ZN(n2938) );
  NAND2_X1 U3688 ( .A1(n3992), .A2(n3830), .ZN(n2936) );
  NAND2_X1 U3689 ( .A1(n3825), .A2(n3020), .ZN(n2935) );
  NAND2_X1 U3690 ( .A1(n2936), .A2(n2935), .ZN(n2939) );
  INV_X1 U3691 ( .A(n2939), .ZN(n2937) );
  NAND2_X1 U3692 ( .A1(n2938), .A2(n2937), .ZN(n3051) );
  INV_X1 U3693 ( .A(n3051), .ZN(n2941) );
  AND2_X1 U3694 ( .A1(n2940), .A2(n2939), .ZN(n3048) );
  NOR2_X1 U3695 ( .A1(n2941), .A2(n3048), .ZN(n2942) );
  XNOR2_X1 U3696 ( .A(n3047), .B(n2942), .ZN(n2947) );
  INV_X1 U3697 ( .A(n3020), .ZN(n3005) );
  OAI22_X1 U3698 ( .A1(n3980), .A2(n3005), .B1(n3155), .B2(n3949), .ZN(n2943)
         );
  AOI211_X1 U3699 ( .C1(n3970), .C2(n3058), .A(n2944), .B(n2943), .ZN(n2946)
         );
  NAND2_X1 U3700 ( .A1(n3985), .A2(n3094), .ZN(n2945) );
  OAI211_X1 U3701 ( .C1(n2947), .C2(n3988), .A(n2946), .B(n2945), .ZN(U3236)
         );
  NAND2_X1 U3702 ( .A1(n2960), .A2(n2948), .ZN(n2949) );
  NAND2_X1 U3703 ( .A1(n2950), .A2(n2949), .ZN(n2979) );
  NAND2_X1 U3704 ( .A1(n2981), .A2(n2977), .ZN(n3563) );
  INV_X1 U3705 ( .A(n2977), .ZN(n2980) );
  NAND2_X1 U3706 ( .A1(n4208), .A2(n2980), .ZN(n3560) );
  AND2_X1 U3707 ( .A1(n3563), .A2(n3560), .ZN(n3529) );
  XNOR2_X1 U3708 ( .A(n2979), .B(n3529), .ZN(n4528) );
  NAND4_X1 U3709 ( .A1(n2954), .A2(n2953), .A3(n2952), .A4(n2951), .ZN(n2955)
         );
  OR2_X1 U3710 ( .A1(n2741), .A2(n3627), .ZN(n2975) );
  INV_X1 U3711 ( .A(n2975), .ZN(n2956) );
  NAND2_X1 U3712 ( .A1(n4505), .A2(n2956), .ZN(n3196) );
  NAND2_X1 U3713 ( .A1(n2957), .A2(n3558), .ZN(n2958) );
  OAI21_X1 U3714 ( .B1(n3529), .B2(n2958), .A(n2986), .ZN(n2962) );
  AOI22_X1 U3715 ( .A1(n2983), .A2(n4327), .B1(n4326), .B2(n2977), .ZN(n2959)
         );
  OAI21_X1 U3716 ( .B1(n2960), .B2(n4330), .A(n2959), .ZN(n2961) );
  AOI21_X1 U3717 ( .B1(n2962), .B2(n4495), .A(n2961), .ZN(n2963) );
  OAI21_X1 U3718 ( .B1(n4528), .B2(n3364), .A(n2963), .ZN(n4529) );
  NAND2_X1 U3719 ( .A1(n4529), .A2(n4505), .ZN(n2968) );
  AOI21_X1 U3720 ( .B1(n2977), .B2(n2964), .A(n3151), .ZN(n4531) );
  OAI22_X1 U3721 ( .A1(n4505), .A2(n2965), .B1(REG3_REG_3__SCAN_IN), .B2(n4162), .ZN(n2966) );
  AOI21_X1 U3722 ( .B1(n4531), .B2(n4399), .A(n2966), .ZN(n2967) );
  OAI211_X1 U3723 ( .C1(n4528), .C2(n3196), .A(n2968), .B(n2967), .ZN(U3287)
         );
  MUX2_X1 U3724 ( .A(n2969), .B(REG2_REG_1__SCAN_IN), .S(n4396), .Z(n2970) );
  INV_X1 U3725 ( .A(n2970), .ZN(n2973) );
  INV_X1 U3726 ( .A(n3196), .ZN(n4503) );
  AOI22_X1 U3727 ( .A1(n2971), .A2(n4503), .B1(REG3_REG_1__SCAN_IN), .B2(n4502), .ZN(n2972) );
  OAI211_X1 U3728 ( .C1(n4174), .C2(n2974), .A(n2973), .B(n2972), .ZN(U3289)
         );
  NAND2_X1 U3729 ( .A1(n3364), .A2(n2975), .ZN(n2976) );
  NAND2_X1 U3730 ( .A1(n4208), .A2(n2977), .ZN(n2978) );
  NAND2_X1 U3731 ( .A1(n2981), .A2(n2980), .ZN(n2982) );
  NAND2_X1 U3732 ( .A1(n2983), .A2(n2984), .ZN(n2985) );
  INV_X1 U3733 ( .A(n3155), .ZN(n3993) );
  AND2_X1 U3734 ( .A1(n3993), .A2(n2997), .ZN(n3003) );
  INV_X1 U3735 ( .A(n3003), .ZN(n3566) );
  NAND2_X1 U3736 ( .A1(n3155), .A2(n3000), .ZN(n3576) );
  AND2_X1 U3737 ( .A1(n3566), .A2(n3576), .ZN(n3525) );
  XOR2_X1 U3738 ( .A(n2999), .B(n3525), .Z(n4538) );
  INV_X1 U3739 ( .A(n3564), .ZN(n2987) );
  XOR2_X1 U3740 ( .A(n3525), .B(n3004), .Z(n2991) );
  AOI22_X1 U3741 ( .A1(n3992), .A2(n4327), .B1(n4326), .B2(n3000), .ZN(n2988)
         );
  OAI21_X1 U3742 ( .B1(n2989), .B2(n4330), .A(n2988), .ZN(n2990) );
  AOI21_X1 U3743 ( .B1(n2991), .B2(n4495), .A(n2990), .ZN(n4539) );
  MUX2_X1 U3744 ( .A(n4539), .B(n2992), .S(n4396), .Z(n2996) );
  AND2_X1 U3745 ( .A1(n3011), .A2(n2993), .ZN(n4542) );
  AOI22_X1 U3746 ( .A1(n4542), .A2(n4399), .B1(n2994), .B2(n4502), .ZN(n2995)
         );
  OAI211_X1 U3747 ( .C1(n4182), .C2(n4538), .A(n2996), .B(n2995), .ZN(U3285)
         );
  INV_X1 U3748 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3015) );
  INV_X1 U3749 ( .A(n4536), .ZN(n4557) );
  NAND2_X1 U3750 ( .A1(n3155), .A2(n2997), .ZN(n2998) );
  NAND2_X1 U3751 ( .A1(n2999), .A2(n2998), .ZN(n3002) );
  NAND2_X1 U3752 ( .A1(n3993), .A2(n3000), .ZN(n3001) );
  INV_X1 U3753 ( .A(n3992), .ZN(n3064) );
  NAND2_X1 U3754 ( .A1(n3064), .A2(n3020), .ZN(n3569) );
  NAND2_X1 U3755 ( .A1(n3992), .A2(n3005), .ZN(n3577) );
  AND2_X1 U3756 ( .A1(n3569), .A2(n3577), .ZN(n3516) );
  XNOR2_X1 U3757 ( .A(n3023), .B(n3516), .ZN(n3098) );
  INV_X1 U3758 ( .A(n3098), .ZN(n3010) );
  AOI21_X1 U3759 ( .B1(n3004), .B2(n3576), .A(n3003), .ZN(n3027) );
  XOR2_X1 U3760 ( .A(n3516), .B(n3027), .Z(n3008) );
  INV_X1 U3761 ( .A(n3058), .ZN(n3144) );
  OAI22_X1 U3762 ( .A1(n3144), .A2(n4497), .B1(n4315), .B2(n3005), .ZN(n3006)
         );
  AOI21_X1 U3763 ( .B1(n4321), .B2(n3993), .A(n3006), .ZN(n3007) );
  OAI21_X1 U3764 ( .B1(n3008), .B2(n4297), .A(n3007), .ZN(n3009) );
  AOI21_X1 U3765 ( .B1(n4496), .B2(n3098), .A(n3009), .ZN(n3100) );
  OAI21_X1 U3766 ( .B1(n4557), .B2(n3010), .A(n3100), .ZN(n3016) );
  NAND2_X1 U3767 ( .A1(n3016), .A2(n4565), .ZN(n3014) );
  AND2_X1 U3768 ( .A1(n3011), .A2(n3020), .ZN(n3012) );
  NOR2_X1 U3769 ( .A1(n3106), .A2(n3012), .ZN(n3093) );
  NAND2_X1 U3770 ( .A1(n3093), .A2(n4346), .ZN(n3013) );
  OAI211_X1 U3771 ( .C1(n4565), .C2(n3015), .A(n3014), .B(n3013), .ZN(U3479)
         );
  INV_X1 U3772 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3019) );
  NAND2_X1 U3773 ( .A1(n3016), .A2(n4577), .ZN(n3018) );
  NAND2_X1 U3774 ( .A1(n3093), .A2(n4244), .ZN(n3017) );
  OAI211_X1 U3775 ( .C1(n4577), .C2(n3019), .A(n3018), .B(n3017), .ZN(U3524)
         );
  AND2_X1 U3776 ( .A1(n3992), .A2(n3020), .ZN(n3022) );
  OR2_X1 U3777 ( .A1(n3992), .A2(n3020), .ZN(n3021) );
  OAI21_X1 U3778 ( .B1(n3023), .B2(n3022), .A(n3021), .ZN(n3111) );
  MUX2_X1 U3779 ( .A(n3024), .B(DATAI_7_), .S(n2682), .Z(n3056) );
  NAND2_X1 U3780 ( .A1(n3144), .A2(n3056), .ZN(n3028) );
  NAND2_X1 U3781 ( .A1(n3058), .A2(n3105), .ZN(n3579) );
  NAND2_X1 U3782 ( .A1(n3058), .A2(n3056), .ZN(n3025) );
  INV_X1 U3783 ( .A(DATAI_8_), .ZN(n4649) );
  MUX2_X1 U3784 ( .A(n3026), .B(n4649), .S(n2682), .Z(n3145) );
  INV_X1 U3785 ( .A(n3145), .ZN(n3138) );
  NAND2_X1 U3786 ( .A1(n3211), .A2(n3138), .ZN(n3573) );
  NAND2_X1 U3787 ( .A1(n3083), .A2(n3145), .ZN(n3578) );
  AND2_X1 U3788 ( .A1(n3573), .A2(n3578), .ZN(n3517) );
  XNOR2_X1 U3789 ( .A(n3082), .B(n3517), .ZN(n3038) );
  INV_X1 U3790 ( .A(n3028), .ZN(n3029) );
  XNOR2_X1 U3791 ( .A(n3069), .B(n3517), .ZN(n3045) );
  OAI22_X1 U3792 ( .A1(n3230), .A2(n4497), .B1(n4315), .B2(n3145), .ZN(n3030)
         );
  AOI21_X1 U3793 ( .B1(n4321), .B2(n3058), .A(n3030), .ZN(n3031) );
  OAI21_X1 U3794 ( .B1(n3045), .B2(n4297), .A(n3031), .ZN(n3032) );
  AOI21_X1 U3795 ( .B1(n3038), .B2(n4549), .A(n3032), .ZN(n3037) );
  INV_X1 U3796 ( .A(n3107), .ZN(n3034) );
  INV_X1 U3797 ( .A(n3086), .ZN(n3033) );
  AOI21_X1 U3798 ( .B1(n3138), .B2(n3034), .A(n3033), .ZN(n3042) );
  AOI22_X1 U3799 ( .A1(n3042), .A2(n4244), .B1(n4574), .B2(REG1_REG_8__SCAN_IN), .ZN(n3035) );
  OAI21_X1 U3800 ( .B1(n3037), .B2(n4574), .A(n3035), .ZN(U3526) );
  AOI22_X1 U3801 ( .A1(n3042), .A2(n4346), .B1(n4563), .B2(REG0_REG_8__SCAN_IN), .ZN(n3036) );
  OAI21_X1 U3802 ( .B1(n3037), .B2(n4563), .A(n3036), .ZN(U3483) );
  NAND2_X1 U3803 ( .A1(n4505), .A2(n4495), .ZN(n4204) );
  NAND2_X1 U3804 ( .A1(n3038), .A2(n4192), .ZN(n3044) );
  NAND2_X1 U3805 ( .A1(n4505), .A2(n4327), .ZN(n4207) );
  NAND2_X1 U3806 ( .A1(n4505), .A2(n4326), .ZN(n4068) );
  INV_X1 U3807 ( .A(n4068), .ZN(n4211) );
  NAND2_X1 U3808 ( .A1(n4505), .A2(n4321), .ZN(n4069) );
  INV_X1 U3809 ( .A(n4069), .ZN(n4210) );
  AOI22_X1 U3810 ( .A1(n3138), .A2(n4211), .B1(n4210), .B2(n3058), .ZN(n3040)
         );
  AOI22_X1 U3811 ( .A1(n4396), .A2(REG2_REG_8__SCAN_IN), .B1(n3148), .B2(n4502), .ZN(n3039) );
  OAI211_X1 U3812 ( .C1(n3230), .C2(n4207), .A(n3040), .B(n3039), .ZN(n3041)
         );
  AOI21_X1 U3813 ( .B1(n3042), .B2(n4399), .A(n3041), .ZN(n3043) );
  OAI211_X1 U3814 ( .C1(n3045), .C2(n4204), .A(n3044), .B(n3043), .ZN(U3282)
         );
  INV_X1 U3815 ( .A(n3985), .ZN(n3974) );
  INV_X1 U3816 ( .A(n3046), .ZN(n3109) );
  INV_X1 U3817 ( .A(n3047), .ZN(n3050) );
  INV_X1 U3818 ( .A(n3048), .ZN(n3049) );
  NAND2_X1 U3819 ( .A1(n3050), .A2(n3049), .ZN(n3052) );
  NAND2_X1 U3820 ( .A1(n3052), .A2(n3051), .ZN(n3059) );
  NAND2_X1 U3821 ( .A1(n3058), .A2(n3825), .ZN(n3054) );
  NAND2_X1 U3822 ( .A1(n3056), .A2(n3843), .ZN(n3053) );
  NAND2_X1 U3823 ( .A1(n3054), .A2(n3053), .ZN(n3055) );
  XNOR2_X1 U3824 ( .A(n3055), .B(n3725), .ZN(n3132) );
  AND2_X1 U3825 ( .A1(n3825), .A2(n3056), .ZN(n3057) );
  AOI21_X1 U3826 ( .B1(n3058), .B2(n3830), .A(n3057), .ZN(n3133) );
  XNOR2_X1 U3827 ( .A(n3132), .B(n3133), .ZN(n3060) );
  AOI21_X1 U3828 ( .B1(n3059), .B2(n3060), .A(n3988), .ZN(n3063) );
  INV_X1 U3829 ( .A(n3059), .ZN(n3062) );
  INV_X1 U3830 ( .A(n3060), .ZN(n3061) );
  NAND2_X1 U3831 ( .A1(n3063), .A2(n3137), .ZN(n3068) );
  OAI22_X1 U3832 ( .A1(n3980), .A2(n3105), .B1(n3064), .B2(n3949), .ZN(n3065)
         );
  AOI211_X1 U3833 ( .C1(n3970), .C2(n3083), .A(n3066), .B(n3065), .ZN(n3067)
         );
  OAI211_X1 U3834 ( .C1(n3974), .C2(n3109), .A(n3068), .B(n3067), .ZN(U3210)
         );
  NAND2_X1 U3835 ( .A1(n3069), .A2(n3573), .ZN(n3070) );
  MUX2_X1 U3836 ( .A(n4386), .B(DATAI_9_), .S(n2682), .Z(n3200) );
  INV_X1 U3837 ( .A(n3200), .ZN(n3212) );
  AND2_X1 U3838 ( .A1(n3202), .A2(n3212), .ZN(n3122) );
  INV_X1 U3839 ( .A(n3122), .ZN(n3587) );
  NAND2_X1 U3840 ( .A1(n3230), .A2(n3200), .ZN(n3574) );
  AND2_X1 U3841 ( .A1(n3587), .A2(n3574), .ZN(n3526) );
  INV_X1 U3842 ( .A(n3526), .ZN(n3071) );
  XNOR2_X1 U3843 ( .A(n3123), .B(n3071), .ZN(n3081) );
  NAND2_X1 U3844 ( .A1(n2677), .A2(REG2_REG_10__SCAN_IN), .ZN(n3078) );
  NOR2_X1 U3845 ( .A1(n3072), .A2(REG3_REG_10__SCAN_IN), .ZN(n3073) );
  OR2_X1 U3846 ( .A1(n3074), .A2(n3073), .ZN(n3235) );
  INV_X1 U3847 ( .A(n3235), .ZN(n3125) );
  NAND2_X1 U3848 ( .A1(n3488), .A2(n3125), .ZN(n3077) );
  NAND2_X1 U3849 ( .A1(n3489), .A2(REG1_REG_10__SCAN_IN), .ZN(n3076) );
  NAND2_X1 U3850 ( .A1(n2133), .A2(REG0_REG_10__SCAN_IN), .ZN(n3075) );
  NAND4_X1 U3851 ( .A1(n3078), .A2(n3077), .A3(n3076), .A4(n3075), .ZN(n3991)
         );
  AOI22_X1 U3852 ( .A1(n3991), .A2(n4327), .B1(n4326), .B2(n3200), .ZN(n3079)
         );
  OAI21_X1 U3853 ( .B1(n3211), .B2(n4330), .A(n3079), .ZN(n3080) );
  AOI21_X1 U3854 ( .B1(n3081), .B2(n4495), .A(n3080), .ZN(n4555) );
  NAND2_X1 U3855 ( .A1(n3083), .A2(n3138), .ZN(n3084) );
  NAND2_X1 U3856 ( .A1(n3085), .A2(n3084), .ZN(n3119) );
  XNOR2_X1 U3857 ( .A(n3119), .B(n3526), .ZN(n4550) );
  NAND2_X1 U3858 ( .A1(n3086), .A2(n3200), .ZN(n3087) );
  NAND2_X1 U3859 ( .A1(n3124), .A2(n3087), .ZN(n4552) );
  NOR2_X1 U3860 ( .A1(n4552), .A2(n4174), .ZN(n3091) );
  INV_X1 U3861 ( .A(n3215), .ZN(n3088) );
  OAI22_X1 U3862 ( .A1(n4505), .A2(n3089), .B1(n3088), .B2(n4162), .ZN(n3090)
         );
  AOI211_X1 U3863 ( .C1(n4550), .C2(n4192), .A(n3091), .B(n3090), .ZN(n3092)
         );
  OAI21_X1 U3864 ( .B1(n4396), .B2(n4555), .A(n3092), .ZN(U3281) );
  INV_X1 U3865 ( .A(n3093), .ZN(n3096) );
  AOI22_X1 U3866 ( .A1(n4396), .A2(REG2_REG_6__SCAN_IN), .B1(n3094), .B2(n4502), .ZN(n3095) );
  OAI21_X1 U3867 ( .B1(n3096), .B2(n4174), .A(n3095), .ZN(n3097) );
  AOI21_X1 U3868 ( .B1(n3098), .B2(n4503), .A(n3097), .ZN(n3099) );
  OAI21_X1 U3869 ( .B1(n3100), .B2(n4396), .A(n3099), .ZN(U3284) );
  XOR2_X1 U3870 ( .A(n3570), .B(n3101), .Z(n3104) );
  OAI22_X1 U3871 ( .A1(n3211), .A2(n4497), .B1(n4315), .B2(n3105), .ZN(n3102)
         );
  AOI21_X1 U3872 ( .B1(n4321), .B2(n3992), .A(n3102), .ZN(n3103) );
  OAI21_X1 U3873 ( .B1(n3104), .B2(n4297), .A(n3103), .ZN(n4545) );
  INV_X1 U3874 ( .A(n4545), .ZN(n3116) );
  OAI21_X1 U3875 ( .B1(n3106), .B2(n3105), .A(n4562), .ZN(n3108) );
  NOR2_X1 U3876 ( .A1(n3108), .A2(n3107), .ZN(n4546) );
  OAI22_X1 U3877 ( .A1(n4505), .A2(n2462), .B1(n3109), .B2(n4162), .ZN(n3114)
         );
  INV_X1 U3878 ( .A(n3110), .ZN(n3112) );
  AND2_X1 U3879 ( .A1(n3111), .A2(n3570), .ZN(n4544) );
  NOR3_X1 U3880 ( .A1(n3112), .A2(n4544), .A3(n4182), .ZN(n3113) );
  AOI211_X1 U3881 ( .C1(n3749), .C2(n4546), .A(n3114), .B(n3113), .ZN(n3115)
         );
  OAI21_X1 U3882 ( .B1(n4396), .B2(n3116), .A(n3115), .ZN(U3283) );
  AND2_X1 U3883 ( .A1(n3202), .A2(n3200), .ZN(n3118) );
  NAND2_X1 U3884 ( .A1(n3230), .A2(n3212), .ZN(n3117) );
  MUX2_X1 U3885 ( .A(n3120), .B(DATAI_10_), .S(n2682), .Z(n3224) );
  NAND2_X1 U3886 ( .A1(n3270), .A2(n3224), .ZN(n3584) );
  INV_X1 U3887 ( .A(n3224), .ZN(n3231) );
  NAND2_X1 U3888 ( .A1(n3991), .A2(n3231), .ZN(n3589) );
  AND2_X1 U3889 ( .A1(n3584), .A2(n3589), .ZN(n3524) );
  INV_X1 U3890 ( .A(n3524), .ZN(n3121) );
  XNOR2_X1 U3891 ( .A(n3181), .B(n3121), .ZN(n3172) );
  INV_X1 U3892 ( .A(n3172), .ZN(n3131) );
  XNOR2_X1 U3893 ( .A(n3184), .B(n3524), .ZN(n3171) );
  INV_X1 U3894 ( .A(n4204), .ZN(n3337) );
  OAI21_X1 U3895 ( .B1(n2188), .B2(n3231), .A(n3191), .ZN(n3179) );
  NOR2_X1 U3896 ( .A1(n3179), .A2(n4174), .ZN(n3129) );
  AOI22_X1 U3897 ( .A1(n3224), .A2(n4211), .B1(n4210), .B2(n3202), .ZN(n3127)
         );
  AOI22_X1 U3898 ( .A1(n4396), .A2(REG2_REG_10__SCAN_IN), .B1(n3125), .B2(
        n4502), .ZN(n3126) );
  OAI211_X1 U3899 ( .C1(n3343), .C2(n4207), .A(n3127), .B(n3126), .ZN(n3128)
         );
  AOI211_X1 U3900 ( .C1(n3171), .C2(n3337), .A(n3129), .B(n3128), .ZN(n3130)
         );
  OAI21_X1 U3901 ( .B1(n4182), .B2(n3131), .A(n3130), .ZN(U3280) );
  INV_X1 U3902 ( .A(n3132), .ZN(n3135) );
  INV_X1 U3903 ( .A(n3133), .ZN(n3134) );
  NAND2_X1 U3904 ( .A1(n3135), .A2(n3134), .ZN(n3136) );
  OR2_X1 U3905 ( .A1(n3211), .A2(n3838), .ZN(n3140) );
  NAND2_X1 U3906 ( .A1(n3138), .A2(n3825), .ZN(n3139) );
  NAND2_X1 U3907 ( .A1(n3140), .A2(n3139), .ZN(n3204) );
  OAI22_X1 U3908 ( .A1(n3211), .A2(n3837), .B1(n3835), .B2(n3145), .ZN(n3141)
         );
  XNOR2_X1 U3909 ( .A(n3141), .B(n2805), .ZN(n3203) );
  XOR2_X1 U3910 ( .A(n3204), .B(n3203), .Z(n3142) );
  XNOR2_X1 U3911 ( .A(n3205), .B(n3142), .ZN(n3150) );
  OAI21_X1 U3912 ( .B1(n3982), .B2(n3230), .A(n3143), .ZN(n3147) );
  OAI22_X1 U3913 ( .A1(n3980), .A2(n3145), .B1(n3144), .B2(n3949), .ZN(n3146)
         );
  AOI211_X1 U3914 ( .C1(n3148), .C2(n3985), .A(n3147), .B(n3146), .ZN(n3149)
         );
  OAI21_X1 U3915 ( .B1(n3150), .B2(n3988), .A(n3149), .ZN(U3218) );
  NOR2_X1 U3916 ( .A1(n4533), .A2(n4384), .ZN(n3163) );
  XOR2_X1 U3917 ( .A(n3152), .B(n3153), .Z(n3162) );
  OAI22_X1 U3918 ( .A1(n3155), .A2(n4497), .B1(n3154), .B2(n4315), .ZN(n3160)
         );
  NAND2_X1 U3919 ( .A1(n3156), .A2(n3152), .ZN(n3157) );
  NAND2_X1 U3920 ( .A1(n3158), .A2(n3157), .ZN(n3165) );
  NOR2_X1 U3921 ( .A1(n3165), .A2(n3364), .ZN(n3159) );
  AOI211_X1 U3922 ( .C1(n4321), .C2(n4208), .A(n3160), .B(n3159), .ZN(n3161)
         );
  OAI21_X1 U3923 ( .B1(n4297), .B2(n3162), .A(n3161), .ZN(n4534) );
  AOI211_X1 U3924 ( .C1(n4502), .C2(n3164), .A(n3163), .B(n4534), .ZN(n3167)
         );
  INV_X1 U3925 ( .A(n3165), .ZN(n4537) );
  AOI22_X1 U3926 ( .A1(n4537), .A2(n4503), .B1(REG2_REG_4__SCAN_IN), .B2(n4396), .ZN(n3166) );
  OAI21_X1 U3927 ( .B1(n3167), .B2(n4396), .A(n3166), .ZN(U3286) );
  NAND2_X1 U3928 ( .A1(n3202), .A2(n4321), .ZN(n3169) );
  NAND2_X1 U3929 ( .A1(n3262), .A2(n4327), .ZN(n3168) );
  OAI211_X1 U3930 ( .C1(n4315), .C2(n3231), .A(n3169), .B(n3168), .ZN(n3170)
         );
  AOI21_X1 U3931 ( .B1(n3171), .B2(n4495), .A(n3170), .ZN(n3174) );
  NAND2_X1 U3932 ( .A1(n3172), .A2(n4549), .ZN(n3173) );
  AND2_X1 U3933 ( .A1(n3174), .A2(n3173), .ZN(n3177) );
  MUX2_X1 U3934 ( .A(n3177), .B(n4764), .S(n4574), .Z(n3175) );
  OAI21_X1 U3935 ( .B1(n3179), .B2(n4313), .A(n3175), .ZN(U3528) );
  INV_X1 U3936 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3176) );
  MUX2_X1 U3937 ( .A(n3177), .B(n3176), .S(n4563), .Z(n3178) );
  OAI21_X1 U3938 ( .B1(n3179), .B2(n4378), .A(n3178), .ZN(U3487) );
  NOR2_X1 U3939 ( .A1(n3991), .A2(n3224), .ZN(n3180) );
  MUX2_X1 U3940 ( .A(n4518), .B(DATAI_11_), .S(n2682), .Z(n3260) );
  NAND2_X1 U3941 ( .A1(n3343), .A2(n3260), .ZN(n3591) );
  INV_X1 U3942 ( .A(n3260), .ZN(n3271) );
  NAND2_X1 U3943 ( .A1(n3262), .A2(n3271), .ZN(n3590) );
  NAND2_X1 U3944 ( .A1(n3182), .A2(n3519), .ZN(n3183) );
  NAND2_X1 U3945 ( .A1(n3236), .A2(n3183), .ZN(n3188) );
  INV_X1 U3946 ( .A(n3188), .ZN(n4558) );
  NAND2_X1 U3947 ( .A1(n3185), .A2(n3584), .ZN(n3239) );
  XOR2_X1 U3948 ( .A(n3519), .B(n3239), .Z(n3190) );
  AOI22_X1 U3949 ( .A1(n3362), .A2(n4327), .B1(n4326), .B2(n3260), .ZN(n3186)
         );
  OAI21_X1 U3950 ( .B1(n3270), .B2(n4330), .A(n3186), .ZN(n3187) );
  AOI21_X1 U3951 ( .B1(n3188), .B2(n4496), .A(n3187), .ZN(n3189) );
  OAI21_X1 U3952 ( .B1(n4297), .B2(n3190), .A(n3189), .ZN(n4559) );
  NAND2_X1 U3953 ( .A1(n4559), .A2(n4505), .ZN(n3195) );
  AOI21_X1 U3954 ( .B1(n3260), .B2(n3191), .A(n3243), .ZN(n4561) );
  INV_X1 U3955 ( .A(n3192), .ZN(n3275) );
  OAI22_X1 U3956 ( .A1(n4505), .A2(n4791), .B1(n3275), .B2(n4162), .ZN(n3193)
         );
  AOI21_X1 U3957 ( .B1(n4561), .B2(n4399), .A(n3193), .ZN(n3194) );
  OAI211_X1 U3958 ( .C1(n4558), .C2(n3196), .A(n3195), .B(n3194), .ZN(U3279)
         );
  NAND2_X1 U3959 ( .A1(n3202), .A2(n3825), .ZN(n3198) );
  NAND2_X1 U3960 ( .A1(n3200), .A2(n3843), .ZN(n3197) );
  NAND2_X1 U3961 ( .A1(n3198), .A2(n3197), .ZN(n3199) );
  XNOR2_X1 U3962 ( .A(n3199), .B(n3725), .ZN(n3220) );
  AND2_X1 U3963 ( .A1(n3825), .A2(n3200), .ZN(n3201) );
  AOI21_X1 U3964 ( .B1(n3202), .B2(n3830), .A(n3201), .ZN(n3219) );
  XNOR2_X1 U3965 ( .A(n3220), .B(n3219), .ZN(n3210) );
  INV_X1 U3966 ( .A(n3209), .ZN(n3207) );
  NAND2_X1 U3967 ( .A1(n3207), .A2(n3206), .ZN(n3278) );
  INV_X1 U3968 ( .A(n3278), .ZN(n3208) );
  AOI21_X1 U3969 ( .B1(n3210), .B2(n3209), .A(n3208), .ZN(n3218) );
  OAI22_X1 U3970 ( .A1(n3980), .A2(n3212), .B1(n3211), .B2(n3949), .ZN(n3213)
         );
  AOI211_X1 U3971 ( .C1(n3970), .C2(n3991), .A(n3214), .B(n3213), .ZN(n3217)
         );
  NAND2_X1 U3972 ( .A1(n3985), .A2(n3215), .ZN(n3216) );
  OAI211_X1 U3973 ( .C1(n3218), .C2(n3988), .A(n3217), .B(n3216), .ZN(U3228)
         );
  NAND2_X1 U3974 ( .A1(n3220), .A2(n3219), .ZN(n3226) );
  AND2_X1 U3975 ( .A1(n3278), .A2(n3226), .ZN(n3228) );
  NAND2_X1 U3976 ( .A1(n3991), .A2(n3825), .ZN(n3222) );
  NAND2_X1 U3977 ( .A1(n3224), .A2(n3843), .ZN(n3221) );
  NAND2_X1 U3978 ( .A1(n3222), .A2(n3221), .ZN(n3223) );
  XNOR2_X1 U3979 ( .A(n3223), .B(n2805), .ZN(n3255) );
  AND2_X1 U3980 ( .A1(n3825), .A2(n3224), .ZN(n3225) );
  AOI21_X1 U3981 ( .B1(n3991), .B2(n3830), .A(n3225), .ZN(n3253) );
  XNOR2_X1 U3982 ( .A(n3255), .B(n3253), .ZN(n3227) );
  AND2_X1 U3983 ( .A1(n3227), .A2(n3226), .ZN(n3276) );
  NAND2_X1 U3984 ( .A1(n3278), .A2(n3276), .ZN(n3256) );
  OAI211_X1 U3985 ( .C1(n3228), .C2(n3227), .A(n3966), .B(n3256), .ZN(n3234)
         );
  INV_X1 U3986 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3229) );
  NOR2_X1 U3987 ( .A1(STATE_REG_SCAN_IN), .A2(n3229), .ZN(n4417) );
  OAI22_X1 U3988 ( .A1(n3980), .A2(n3231), .B1(n3230), .B2(n3949), .ZN(n3232)
         );
  AOI211_X1 U3989 ( .C1(n3970), .C2(n3262), .A(n4417), .B(n3232), .ZN(n3233)
         );
  OAI211_X1 U3990 ( .C1(n3974), .C2(n3235), .A(n3234), .B(n3233), .ZN(U3214)
         );
  MUX2_X1 U3991 ( .A(n3237), .B(DATAI_12_), .S(n2682), .Z(n3340) );
  NAND2_X1 U3992 ( .A1(n3362), .A2(n3290), .ZN(n3355) );
  INV_X1 U3993 ( .A(n3355), .ZN(n3238) );
  NOR2_X1 U3994 ( .A1(n3362), .A2(n3290), .ZN(n3356) );
  OR2_X1 U3995 ( .A1(n3238), .A2(n3356), .ZN(n3241) );
  XNOR2_X1 U3996 ( .A(n3318), .B(n3241), .ZN(n3339) );
  INV_X1 U3997 ( .A(n3339), .ZN(n3252) );
  NAND2_X1 U3998 ( .A1(n3239), .A2(n3590), .ZN(n3240) );
  NAND2_X1 U3999 ( .A1(n3240), .A2(n3591), .ZN(n3357) );
  INV_X1 U4000 ( .A(n3241), .ZN(n3527) );
  XNOR2_X1 U4001 ( .A(n3357), .B(n3527), .ZN(n3242) );
  NAND2_X1 U4002 ( .A1(n3242), .A2(n4495), .ZN(n3342) );
  NOR2_X1 U4003 ( .A1(n3342), .A2(n4396), .ZN(n3250) );
  OR2_X1 U4004 ( .A1(n3243), .A2(n3290), .ZN(n3244) );
  NAND2_X1 U4005 ( .A1(n3366), .A2(n3244), .ZN(n3352) );
  NOR2_X1 U4006 ( .A1(n3352), .A2(n4174), .ZN(n3249) );
  NAND2_X1 U4007 ( .A1(n4396), .A2(REG2_REG_12__SCAN_IN), .ZN(n3246) );
  NAND2_X1 U4008 ( .A1(n4502), .A2(n3293), .ZN(n3245) );
  OAI211_X1 U4009 ( .C1(n4207), .C2(n3662), .A(n3246), .B(n3245), .ZN(n3248)
         );
  OAI22_X1 U4010 ( .A1(n3343), .A2(n4069), .B1(n4068), .B2(n3290), .ZN(n3247)
         );
  NOR4_X1 U4011 ( .A1(n3250), .A2(n3249), .A3(n3248), .A4(n3247), .ZN(n3251)
         );
  OAI21_X1 U4012 ( .B1(n3252), .B2(n4182), .A(n3251), .ZN(U3278) );
  INV_X1 U4013 ( .A(n3253), .ZN(n3254) );
  NAND2_X1 U4014 ( .A1(n3255), .A2(n3254), .ZN(n3281) );
  NAND2_X1 U4015 ( .A1(n3256), .A2(n3281), .ZN(n3268) );
  NAND2_X1 U4016 ( .A1(n3262), .A2(n3825), .ZN(n3258) );
  NAND2_X1 U4017 ( .A1(n3260), .A2(n3843), .ZN(n3257) );
  NAND2_X1 U4018 ( .A1(n3258), .A2(n3257), .ZN(n3259) );
  XNOR2_X1 U4019 ( .A(n3259), .B(n3725), .ZN(n3266) );
  INV_X1 U4020 ( .A(n3266), .ZN(n3264) );
  AND2_X1 U4021 ( .A1(n3825), .A2(n3260), .ZN(n3261) );
  AOI21_X1 U4022 ( .B1(n3262), .B2(n3830), .A(n3261), .ZN(n3265) );
  INV_X1 U4023 ( .A(n3265), .ZN(n3263) );
  NAND2_X1 U4024 ( .A1(n3264), .A2(n3263), .ZN(n3280) );
  NAND2_X1 U4025 ( .A1(n3266), .A2(n3265), .ZN(n3279) );
  NAND2_X1 U4026 ( .A1(n3280), .A2(n3279), .ZN(n3267) );
  XNOR2_X1 U4027 ( .A(n3268), .B(n3267), .ZN(n3269) );
  NAND2_X1 U4028 ( .A1(n3269), .A2(n3966), .ZN(n3274) );
  INV_X1 U4029 ( .A(REG3_REG_11__SCAN_IN), .ZN(n4861) );
  NOR2_X1 U4030 ( .A1(STATE_REG_SCAN_IN), .A2(n4861), .ZN(n4425) );
  OAI22_X1 U4031 ( .A1(n3980), .A2(n3271), .B1(n3270), .B2(n3949), .ZN(n3272)
         );
  AOI211_X1 U4032 ( .C1(n3970), .C2(n3362), .A(n4425), .B(n3272), .ZN(n3273)
         );
  OAI211_X1 U4033 ( .C1(n3974), .C2(n3275), .A(n3274), .B(n3273), .ZN(U3233)
         );
  AND2_X1 U4034 ( .A1(n3276), .A2(n3279), .ZN(n3277) );
  NAND2_X1 U4035 ( .A1(n3278), .A2(n3277), .ZN(n3297) );
  INV_X1 U4036 ( .A(n3279), .ZN(n3283) );
  AND2_X1 U4037 ( .A1(n3281), .A2(n3280), .ZN(n3282) );
  NAND2_X1 U4038 ( .A1(n3362), .A2(n3830), .ZN(n3285) );
  NAND2_X1 U4039 ( .A1(n3825), .A2(n3340), .ZN(n3284) );
  NAND2_X1 U4040 ( .A1(n3285), .A2(n3284), .ZN(n3298) );
  NAND2_X1 U4041 ( .A1(n3362), .A2(n3825), .ZN(n3287) );
  NAND2_X1 U4042 ( .A1(n3340), .A2(n3843), .ZN(n3286) );
  NAND2_X1 U40430 ( .A1(n3287), .A2(n3286), .ZN(n3288) );
  XNOR2_X1 U4044 ( .A(n3288), .B(n2805), .ZN(n3299) );
  XOR2_X1 U4045 ( .A(n3298), .B(n3299), .Z(n3289) );
  XNOR2_X1 U4046 ( .A(n2155), .B(n3289), .ZN(n3295) );
  NAND2_X1 U4047 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4436) );
  OAI21_X1 U4048 ( .B1(n3982), .B2(n3662), .A(n4436), .ZN(n3292) );
  OAI22_X1 U4049 ( .A1(n3980), .A2(n3290), .B1(n3343), .B2(n3949), .ZN(n3291)
         );
  AOI211_X1 U4050 ( .C1(n3293), .C2(n3985), .A(n3292), .B(n3291), .ZN(n3294)
         );
  OAI21_X1 U4051 ( .B1(n3295), .B2(n3988), .A(n3294), .ZN(U3221) );
  NAND2_X1 U4052 ( .A1(n3353), .A2(n3825), .ZN(n3302) );
  MUX2_X1 U4053 ( .A(n3300), .B(DATAI_13_), .S(n2682), .Z(n3323) );
  NAND2_X1 U4054 ( .A1(n3323), .A2(n3843), .ZN(n3301) );
  NAND2_X1 U4055 ( .A1(n3302), .A2(n3301), .ZN(n3303) );
  XNOR2_X1 U4056 ( .A(n3303), .B(n2805), .ZN(n3309) );
  INV_X1 U4057 ( .A(n3309), .ZN(n3307) );
  NAND2_X1 U4058 ( .A1(n3353), .A2(n3830), .ZN(n3305) );
  NAND2_X1 U4059 ( .A1(n3825), .A2(n3323), .ZN(n3304) );
  NAND2_X1 U4060 ( .A1(n3305), .A2(n3304), .ZN(n3308) );
  INV_X1 U4061 ( .A(n3308), .ZN(n3306) );
  NOR2_X1 U4062 ( .A1(n2166), .A2(n3384), .ZN(n3310) );
  XNOR2_X1 U4063 ( .A(n3385), .B(n3310), .ZN(n3315) );
  AND2_X1 U4064 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n3405) );
  INV_X1 U4065 ( .A(n3362), .ZN(n3311) );
  OAI22_X1 U4066 ( .A1(n3980), .A2(n3368), .B1(n3311), .B2(n3949), .ZN(n3312)
         );
  AOI211_X1 U4067 ( .C1(n3970), .C2(n3388), .A(n3405), .B(n3312), .ZN(n3314)
         );
  NAND2_X1 U4068 ( .A1(n3985), .A2(n3370), .ZN(n3313) );
  OAI211_X1 U4069 ( .C1(n3315), .C2(n3988), .A(n3314), .B(n3313), .ZN(U3231)
         );
  MUX2_X1 U4070 ( .A(n4514), .B(DATAI_14_), .S(n2682), .Z(n3660) );
  NAND2_X1 U4071 ( .A1(n4331), .A2(n3660), .ZN(n3410) );
  INV_X1 U4072 ( .A(n3660), .ZN(n3393) );
  NAND2_X1 U4073 ( .A1(n3388), .A2(n3393), .ZN(n3411) );
  NAND2_X1 U4074 ( .A1(n3362), .A2(n3340), .ZN(n3317) );
  NOR2_X1 U4075 ( .A1(n3362), .A2(n3340), .ZN(n3316) );
  AOI21_X1 U4076 ( .B1(n3531), .B2(n3319), .A(n3375), .ZN(n3663) );
  NAND2_X1 U4077 ( .A1(n3353), .A2(n3368), .ZN(n3320) );
  NAND2_X1 U4078 ( .A1(n3357), .A2(n3595), .ZN(n3322) );
  NOR2_X1 U4079 ( .A1(n3353), .A2(n3368), .ZN(n3321) );
  AOI21_X1 U4080 ( .B1(n3595), .B2(n3356), .A(n3321), .ZN(n3592) );
  NAND2_X1 U4081 ( .A1(n3322), .A2(n3592), .ZN(n3413) );
  XNOR2_X1 U4082 ( .A(n3413), .B(n3531), .ZN(n3666) );
  INV_X1 U4083 ( .A(n3367), .ZN(n3325) );
  INV_X1 U4084 ( .A(n3652), .ZN(n3324) );
  OAI21_X1 U4085 ( .B1(n3325), .B2(n3393), .A(n3324), .ZN(n3670) );
  NOR2_X1 U4086 ( .A1(n3670), .A2(n4174), .ZN(n3336) );
  NAND2_X1 U4087 ( .A1(n2677), .A2(REG2_REG_15__SCAN_IN), .ZN(n3332) );
  OR2_X1 U4088 ( .A1(n3326), .A2(REG3_REG_15__SCAN_IN), .ZN(n3327) );
  AND2_X1 U4089 ( .A1(n3328), .A2(n3327), .ZN(n3700) );
  NAND2_X1 U4090 ( .A1(n3488), .A2(n3700), .ZN(n3331) );
  NAND2_X1 U4091 ( .A1(n3489), .A2(REG1_REG_15__SCAN_IN), .ZN(n3330) );
  NAND2_X1 U4092 ( .A1(n2133), .A2(REG0_REG_15__SCAN_IN), .ZN(n3329) );
  NAND4_X1 U4093 ( .A1(n3332), .A2(n3331), .A3(n3330), .A4(n3329), .ZN(n4320)
         );
  AOI22_X1 U4094 ( .A1(n3660), .A2(n4211), .B1(n4210), .B2(n3353), .ZN(n3334)
         );
  AOI22_X1 U4095 ( .A1(n4396), .A2(REG2_REG_14__SCAN_IN), .B1(n3396), .B2(
        n4502), .ZN(n3333) );
  OAI211_X1 U4096 ( .C1(n3690), .C2(n4207), .A(n3334), .B(n3333), .ZN(n3335)
         );
  AOI211_X1 U4097 ( .C1(n3666), .C2(n3337), .A(n3336), .B(n3335), .ZN(n3338)
         );
  OAI21_X1 U4098 ( .B1(n3663), .B2(n4182), .A(n3338), .ZN(U3276) );
  NAND2_X1 U4099 ( .A1(n3339), .A2(n4549), .ZN(n3346) );
  AOI22_X1 U4100 ( .A1(n3353), .A2(n4327), .B1(n4326), .B2(n3340), .ZN(n3341)
         );
  OAI211_X1 U4101 ( .C1(n3343), .C2(n4330), .A(n3342), .B(n3341), .ZN(n3344)
         );
  INV_X1 U4102 ( .A(n3344), .ZN(n3345) );
  NAND2_X1 U4103 ( .A1(n3346), .A2(n3345), .ZN(n3349) );
  MUX2_X1 U4104 ( .A(REG0_REG_12__SCAN_IN), .B(n3349), .S(n4565), .Z(n3347) );
  INV_X1 U4105 ( .A(n3347), .ZN(n3348) );
  OAI21_X1 U4106 ( .B1(n3352), .B2(n4378), .A(n3348), .ZN(U3491) );
  MUX2_X1 U4107 ( .A(REG1_REG_12__SCAN_IN), .B(n3349), .S(n4577), .Z(n3350) );
  INV_X1 U4108 ( .A(n3350), .ZN(n3351) );
  OAI21_X1 U4109 ( .B1(n4313), .B2(n3352), .A(n3351), .ZN(U3530) );
  XNOR2_X1 U4110 ( .A(n3353), .B(n3368), .ZN(n3539) );
  XNOR2_X1 U4111 ( .A(n3354), .B(n3539), .ZN(n3365) );
  OAI22_X1 U4112 ( .A1(n4331), .A2(n4497), .B1(n4315), .B2(n3368), .ZN(n3361)
         );
  OAI21_X1 U4113 ( .B1(n3357), .B2(n3356), .A(n3355), .ZN(n3358) );
  XOR2_X1 U4114 ( .A(n3539), .B(n3358), .Z(n3359) );
  NOR2_X1 U4115 ( .A1(n3359), .A2(n4297), .ZN(n3360) );
  AOI211_X1 U4116 ( .C1(n4321), .C2(n3362), .A(n3361), .B(n3360), .ZN(n3363)
         );
  OAI21_X1 U4117 ( .B1(n3365), .B2(n3364), .A(n3363), .ZN(n3635) );
  INV_X1 U4118 ( .A(n3635), .ZN(n3374) );
  INV_X1 U4119 ( .A(n3365), .ZN(n3636) );
  INV_X1 U4120 ( .A(n3366), .ZN(n3369) );
  OAI21_X1 U4121 ( .B1(n3369), .B2(n3368), .A(n3367), .ZN(n3642) );
  AOI22_X1 U4122 ( .A1(n4396), .A2(REG2_REG_13__SCAN_IN), .B1(n3370), .B2(
        n4502), .ZN(n3371) );
  OAI21_X1 U4123 ( .B1(n3642), .B2(n4174), .A(n3371), .ZN(n3372) );
  AOI21_X1 U4124 ( .B1(n3636), .B2(n4503), .A(n3372), .ZN(n3373) );
  OAI21_X1 U4125 ( .B1(n3374), .B2(n4396), .A(n3373), .ZN(U3277) );
  MUX2_X1 U4126 ( .A(n3376), .B(DATAI_15_), .S(n2682), .Z(n4325) );
  NAND2_X1 U4127 ( .A1(n3690), .A2(n4325), .ZN(n3412) );
  NAND2_X1 U4128 ( .A1(n4320), .A2(n3698), .ZN(n3648) );
  NAND2_X1 U4129 ( .A1(n3412), .A2(n3648), .ZN(n3528) );
  XNOR2_X1 U4130 ( .A(n3643), .B(n3528), .ZN(n4336) );
  XNOR2_X1 U4131 ( .A(n3652), .B(n4325), .ZN(n4333) );
  AOI22_X1 U4132 ( .A1(n4325), .A2(n4211), .B1(n4210), .B2(n3388), .ZN(n3378)
         );
  AOI22_X1 U4133 ( .A1(n4396), .A2(REG2_REG_15__SCAN_IN), .B1(n3700), .B2(
        n4502), .ZN(n3377) );
  OAI211_X1 U4134 ( .C1(n3730), .C2(n4207), .A(n3378), .B(n3377), .ZN(n3382)
         );
  AOI21_X1 U4135 ( .B1(n3379), .B2(n3528), .A(n4297), .ZN(n3380) );
  NAND2_X1 U4136 ( .A1(n3380), .A2(n3649), .ZN(n4334) );
  NOR2_X1 U4137 ( .A1(n4334), .A2(n4396), .ZN(n3381) );
  AOI211_X1 U4138 ( .C1(n4399), .C2(n4333), .A(n3382), .B(n3381), .ZN(n3383)
         );
  OAI21_X1 U4139 ( .B1(n4336), .B2(n4182), .A(n3383), .ZN(U3275) );
  NAND2_X1 U4140 ( .A1(n3388), .A2(n3830), .ZN(n3387) );
  NAND2_X1 U4141 ( .A1(n3825), .A2(n3660), .ZN(n3386) );
  NAND2_X1 U4142 ( .A1(n3387), .A2(n3386), .ZN(n3672) );
  NAND2_X1 U4143 ( .A1(n3388), .A2(n3825), .ZN(n3390) );
  NAND2_X1 U4144 ( .A1(n3660), .A2(n3843), .ZN(n3389) );
  NAND2_X1 U4145 ( .A1(n3390), .A2(n3389), .ZN(n3391) );
  XNOR2_X1 U4146 ( .A(n3391), .B(n3725), .ZN(n3675) );
  XOR2_X1 U4147 ( .A(n3672), .B(n3675), .Z(n3392) );
  XNOR2_X1 U4148 ( .A(n3674), .B(n3392), .ZN(n3398) );
  NAND2_X1 U4149 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4451) );
  OAI21_X1 U4150 ( .B1(n3982), .B2(n3690), .A(n4451), .ZN(n3395) );
  OAI22_X1 U4151 ( .A1(n3980), .A2(n3393), .B1(n3662), .B2(n3949), .ZN(n3394)
         );
  AOI211_X1 U4152 ( .C1(n3396), .C2(n3985), .A(n3395), .B(n3394), .ZN(n3397)
         );
  OAI21_X1 U4153 ( .B1(n3398), .B2(n3988), .A(n3397), .ZN(U3212) );
  XNOR2_X1 U4154 ( .A(n3408), .B(REG2_REG_13__SCAN_IN), .ZN(n3400) );
  AOI21_X1 U4155 ( .B1(n3400), .B2(n3401), .A(n4445), .ZN(n3399) );
  OAI21_X1 U4156 ( .B1(n3401), .B2(n3400), .A(n3399), .ZN(n3407) );
  AOI211_X1 U4157 ( .C1(n3403), .C2(n3402), .A(n2313), .B(n4478), .ZN(n3404)
         );
  AOI211_X1 U4158 ( .C1(n4483), .C2(ADDR_REG_13__SCAN_IN), .A(n3405), .B(n3404), .ZN(n3406) );
  OAI211_X1 U4159 ( .C1(n4490), .C2(n3408), .A(n3407), .B(n3406), .ZN(U3253)
         );
  INV_X1 U4160 ( .A(n3409), .ZN(n3626) );
  NAND2_X1 U4161 ( .A1(n2682), .A2(DATAI_31_), .ZN(n4219) );
  INV_X1 U4162 ( .A(n4219), .ZN(n4222) );
  NAND2_X1 U4163 ( .A1(n2682), .A2(DATAI_30_), .ZN(n4229) );
  NAND2_X1 U4164 ( .A1(n3410), .A2(n3412), .ZN(n3594) );
  NAND2_X1 U4165 ( .A1(n3648), .A2(n3411), .ZN(n3582) );
  NAND2_X1 U4166 ( .A1(n3582), .A2(n3412), .ZN(n3585) );
  OAI21_X1 U4167 ( .B1(n3413), .B2(n3594), .A(n3585), .ZN(n3415) );
  INV_X1 U4168 ( .A(n4512), .ZN(n3414) );
  MUX2_X1 U4169 ( .A(n3414), .B(DATAI_16_), .S(n2682), .Z(n3685) );
  NAND2_X1 U4170 ( .A1(n3730), .A2(n3685), .ZN(n3601) );
  NAND2_X1 U4171 ( .A1(n4328), .A2(n4314), .ZN(n3706) );
  AOI21_X1 U4172 ( .B1(n3415), .B2(n3601), .A(n2170), .ZN(n3465) );
  INV_X1 U4173 ( .A(DATAI_19_), .ZN(n3416) );
  NAND2_X1 U4174 ( .A1(n4295), .A2(n3908), .ZN(n3426) );
  AOI22_X1 U4175 ( .A1(n2677), .A2(REG2_REG_18__SCAN_IN), .B1(n3489), .B2(
        REG1_REG_18__SCAN_IN), .ZN(n3424) );
  INV_X1 U4176 ( .A(n3417), .ZN(n3418) );
  AOI21_X1 U4177 ( .B1(n3418), .B2(REG3_REG_17__SCAN_IN), .A(
        REG3_REG_18__SCAN_IN), .ZN(n3420) );
  OR2_X1 U4178 ( .A1(n3420), .A2(n3419), .ZN(n3973) );
  NAND2_X1 U4179 ( .A1(n2133), .A2(REG0_REG_18__SCAN_IN), .ZN(n3421) );
  OAI21_X1 U4180 ( .B1(n3973), .B2(n2679), .A(n3421), .ZN(n3422) );
  INV_X1 U4181 ( .A(n3422), .ZN(n3423) );
  MUX2_X1 U4182 ( .A(n3425), .B(DATAI_18_), .S(n2682), .Z(n3766) );
  NAND2_X1 U4183 ( .A1(n3990), .A2(n3968), .ZN(n3758) );
  AND2_X1 U4184 ( .A1(n3426), .A2(n3758), .ZN(n3448) );
  NAND2_X1 U4185 ( .A1(n3907), .A2(n3766), .ZN(n3757) );
  INV_X1 U4186 ( .A(DATAI_17_), .ZN(n4635) );
  MUX2_X1 U4187 ( .A(n3427), .B(n4635), .S(n2682), .Z(n3741) );
  NAND2_X1 U4188 ( .A1(n4316), .A2(n3742), .ZN(n3737) );
  NAND2_X1 U4189 ( .A1(n3757), .A2(n3737), .ZN(n3428) );
  NAND2_X1 U4190 ( .A1(n3448), .A2(n3428), .ZN(n3430) );
  INV_X1 U4191 ( .A(n3908), .ZN(n3855) );
  NAND2_X1 U4192 ( .A1(n3950), .A2(n3855), .ZN(n3429) );
  NAND2_X1 U4193 ( .A1(n3430), .A2(n3429), .ZN(n4186) );
  INV_X1 U4194 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3948) );
  XNOR2_X1 U4195 ( .A(n3438), .B(n3948), .ZN(n4197) );
  NAND2_X1 U4196 ( .A1(n4197), .A2(n3488), .ZN(n3436) );
  INV_X1 U4197 ( .A(REG2_REG_20__SCAN_IN), .ZN(n3433) );
  NAND2_X1 U4198 ( .A1(n3489), .A2(REG1_REG_20__SCAN_IN), .ZN(n3432) );
  NAND2_X1 U4199 ( .A1(n2133), .A2(REG0_REG_20__SCAN_IN), .ZN(n3431) );
  OAI211_X1 U4200 ( .C1(n2638), .C2(n3433), .A(n3432), .B(n3431), .ZN(n3434)
         );
  INV_X1 U4201 ( .A(n3434), .ZN(n3435) );
  NOR2_X1 U4202 ( .A1(n4288), .A2(n4292), .ZN(n3437) );
  NAND2_X1 U4203 ( .A1(n4288), .A2(n4292), .ZN(n3447) );
  OAI21_X1 U4204 ( .B1(n4186), .B2(n3437), .A(n3447), .ZN(n4130) );
  NAND2_X1 U4205 ( .A1(n2682), .A2(DATAI_22_), .ZN(n3957) );
  NOR2_X1 U4206 ( .A1(n4139), .A2(n3957), .ZN(n4134) );
  INV_X1 U4207 ( .A(REG0_REG_21__SCAN_IN), .ZN(n3444) );
  NAND2_X1 U4208 ( .A1(n3438), .A2(REG3_REG_20__SCAN_IN), .ZN(n3439) );
  INV_X1 U4209 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3919) );
  NAND2_X1 U4210 ( .A1(n3439), .A2(n3919), .ZN(n3441) );
  NAND2_X1 U4211 ( .A1(n3441), .A2(n3440), .ZN(n3918) );
  OR2_X1 U4212 ( .A1(n3918), .A2(n2679), .ZN(n3443) );
  AOI22_X1 U4213 ( .A1(n2677), .A2(REG2_REG_21__SCAN_IN), .B1(n3489), .B2(
        REG1_REG_21__SCAN_IN), .ZN(n3442) );
  OR2_X1 U4214 ( .A1(n4156), .A2(n4283), .ZN(n4133) );
  INV_X1 U4215 ( .A(n4133), .ZN(n3446) );
  NOR2_X1 U4216 ( .A1(n4134), .A2(n3446), .ZN(n3610) );
  AND2_X1 U4217 ( .A1(n4130), .A2(n3610), .ZN(n3874) );
  INV_X1 U4218 ( .A(n3874), .ZN(n3464) );
  NAND2_X1 U4219 ( .A1(n3743), .A2(n3741), .ZN(n3736) );
  NAND2_X1 U4220 ( .A1(n3447), .A2(n3736), .ZN(n3449) );
  INV_X1 U4221 ( .A(n3448), .ZN(n4183) );
  NOR2_X1 U4222 ( .A1(n3449), .A2(n4183), .ZN(n3604) );
  OR2_X1 U4223 ( .A1(n3464), .A2(n3604), .ZN(n3463) );
  NAND2_X1 U4224 ( .A1(n4156), .A2(n4283), .ZN(n3606) );
  NOR2_X1 U4225 ( .A1(n4134), .A2(n3606), .ZN(n3461) );
  AND2_X1 U4226 ( .A1(n4139), .A2(n3957), .ZN(n3547) );
  INV_X1 U4227 ( .A(n3547), .ZN(n3460) );
  NAND2_X1 U4228 ( .A1(n3450), .A2(n3899), .ZN(n3451) );
  AND2_X1 U4229 ( .A1(n3452), .A2(n3451), .ZN(n4146) );
  NAND2_X1 U4230 ( .A1(n4146), .A2(n3488), .ZN(n3458) );
  INV_X1 U4231 ( .A(REG2_REG_23__SCAN_IN), .ZN(n3455) );
  NAND2_X1 U4232 ( .A1(n3489), .A2(REG1_REG_23__SCAN_IN), .ZN(n3454) );
  NAND2_X1 U4233 ( .A1(n2133), .A2(REG0_REG_23__SCAN_IN), .ZN(n3453) );
  OAI211_X1 U4234 ( .C1(n3455), .C2(n2638), .A(n3454), .B(n3453), .ZN(n3456)
         );
  INV_X1 U4235 ( .A(n3456), .ZN(n3457) );
  NAND2_X1 U4236 ( .A1(n2682), .A2(DATAI_23_), .ZN(n4144) );
  NAND2_X1 U4237 ( .A1(n4266), .A2(n4144), .ZN(n3459) );
  NAND2_X1 U4238 ( .A1(n3460), .A2(n3459), .ZN(n3608) );
  NOR2_X1 U4239 ( .A1(n3461), .A2(n3608), .ZN(n3462) );
  OAI21_X1 U4240 ( .B1(n3465), .B2(n3464), .A(n3875), .ZN(n3474) );
  NAND2_X1 U4241 ( .A1(n2682), .A2(DATAI_24_), .ZN(n4120) );
  OR2_X1 U4242 ( .A1(n3862), .A2(n4120), .ZN(n3549) );
  NAND2_X1 U4243 ( .A1(n4158), .A2(n4138), .ZN(n4111) );
  INV_X1 U4244 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3928) );
  XNOR2_X1 U4245 ( .A(n3466), .B(n3928), .ZN(n4106) );
  NAND2_X1 U4246 ( .A1(n4106), .A2(n3488), .ZN(n3472) );
  INV_X1 U4247 ( .A(REG2_REG_25__SCAN_IN), .ZN(n3469) );
  NAND2_X1 U4248 ( .A1(n3489), .A2(REG1_REG_25__SCAN_IN), .ZN(n3468) );
  NAND2_X1 U4249 ( .A1(n2133), .A2(REG0_REG_25__SCAN_IN), .ZN(n3467) );
  OAI211_X1 U4250 ( .C1(n2638), .C2(n3469), .A(n3468), .B(n3467), .ZN(n3470)
         );
  INV_X1 U4251 ( .A(n3470), .ZN(n3471) );
  NAND2_X1 U4252 ( .A1(n2682), .A2(DATAI_25_), .ZN(n4105) );
  NAND2_X1 U4253 ( .A1(n4080), .A2(n4105), .ZN(n3511) );
  NAND2_X1 U4254 ( .A1(n3862), .A2(n4120), .ZN(n4096) );
  AND2_X1 U4255 ( .A1(n3511), .A2(n4096), .ZN(n3877) );
  INV_X1 U4256 ( .A(n3877), .ZN(n3473) );
  AOI21_X1 U4257 ( .B1(n3474), .B2(n3876), .A(n3473), .ZN(n3508) );
  NAND2_X1 U4258 ( .A1(n2682), .A2(DATAI_26_), .ZN(n4088) );
  OR2_X1 U4259 ( .A1(n4249), .A2(n4088), .ZN(n3512) );
  OR2_X1 U4260 ( .A1(n4080), .A2(n4105), .ZN(n4074) );
  AND2_X1 U4261 ( .A1(n3512), .A2(n4074), .ZN(n3879) );
  INV_X1 U4262 ( .A(n4042), .ZN(n3476) );
  INV_X1 U4263 ( .A(n4229), .ZN(n3475) );
  NAND2_X1 U4264 ( .A1(n3476), .A2(n3475), .ZN(n3477) );
  NAND2_X1 U4265 ( .A1(n4221), .A2(n4219), .ZN(n3621) );
  AND2_X1 U4266 ( .A1(n3477), .A2(n3621), .ZN(n3537) );
  NAND2_X1 U4267 ( .A1(n3485), .A2(REG3_REG_27__SCAN_IN), .ZN(n3486) );
  INV_X1 U4268 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3848) );
  NAND2_X1 U4269 ( .A1(n3486), .A2(n3848), .ZN(n3478) );
  NAND2_X1 U4270 ( .A1(n4065), .A2(n3488), .ZN(n3484) );
  INV_X1 U4271 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3481) );
  NAND2_X1 U4272 ( .A1(n3489), .A2(REG1_REG_28__SCAN_IN), .ZN(n3480) );
  NAND2_X1 U4273 ( .A1(n2133), .A2(REG0_REG_28__SCAN_IN), .ZN(n3479) );
  OAI211_X1 U4274 ( .C1(n2638), .C2(n3481), .A(n3480), .B(n3479), .ZN(n3482)
         );
  INV_X1 U4275 ( .A(n3482), .ZN(n3483) );
  NAND2_X1 U4276 ( .A1(n2682), .A2(DATAI_28_), .ZN(n4067) );
  NOR2_X1 U4277 ( .A1(n4247), .A2(n4067), .ZN(n4037) );
  OR2_X1 U4278 ( .A1(n3485), .A2(REG3_REG_27__SCAN_IN), .ZN(n3487) );
  NAND2_X1 U4279 ( .A1(n3892), .A2(n3488), .ZN(n3494) );
  NAND2_X1 U4280 ( .A1(n3489), .A2(REG1_REG_27__SCAN_IN), .ZN(n3491) );
  NAND2_X1 U4281 ( .A1(n2133), .A2(REG0_REG_27__SCAN_IN), .ZN(n3490) );
  OAI211_X1 U4282 ( .C1(n4799), .C2(n2638), .A(n3491), .B(n3490), .ZN(n3492)
         );
  INV_X1 U4283 ( .A(n3492), .ZN(n3493) );
  AND2_X1 U4284 ( .A1(n4241), .A2(n4248), .ZN(n4034) );
  NOR2_X1 U4285 ( .A1(n4037), .A2(n4034), .ZN(n3502) );
  INV_X1 U4286 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3497) );
  NAND2_X1 U4287 ( .A1(n3489), .A2(REG1_REG_29__SCAN_IN), .ZN(n3496) );
  NAND2_X1 U4288 ( .A1(n2133), .A2(REG0_REG_29__SCAN_IN), .ZN(n3495) );
  OAI211_X1 U4289 ( .C1(n2638), .C2(n3497), .A(n3496), .B(n3495), .ZN(n3498)
         );
  INV_X1 U4290 ( .A(n3498), .ZN(n3499) );
  OAI21_X1 U4291 ( .B1(n4033), .B2(n2679), .A(n3499), .ZN(n4238) );
  NAND2_X1 U4292 ( .A1(n2682), .A2(DATAI_29_), .ZN(n4041) );
  OR2_X1 U4293 ( .A1(n4238), .A2(n4041), .ZN(n3515) );
  NAND4_X1 U4294 ( .A1(n3879), .A2(n3537), .A3(n3502), .A4(n3515), .ZN(n3507)
         );
  NAND2_X1 U4295 ( .A1(n4042), .A2(n4229), .ZN(n3535) );
  INV_X1 U4296 ( .A(n3535), .ZN(n3505) );
  INV_X1 U4297 ( .A(n4221), .ZN(n3500) );
  NAND2_X1 U4298 ( .A1(n3500), .A2(n4222), .ZN(n3536) );
  INV_X1 U4299 ( .A(n3536), .ZN(n3504) );
  XNOR2_X1 U4300 ( .A(n4241), .B(n4048), .ZN(n4035) );
  AND2_X1 U4301 ( .A1(n4249), .A2(n4088), .ZN(n3878) );
  NAND2_X1 U4302 ( .A1(n4238), .A2(n4041), .ZN(n3514) );
  NAND2_X1 U4303 ( .A1(n4247), .A2(n4067), .ZN(n4038) );
  NAND2_X1 U4304 ( .A1(n3514), .A2(n4038), .ZN(n3501) );
  NOR2_X1 U4305 ( .A1(n3878), .A2(n3501), .ZN(n3613) );
  OAI211_X1 U4306 ( .C1(n3502), .C2(n3501), .A(n3537), .B(n3515), .ZN(n3617)
         );
  AOI21_X1 U4307 ( .B1(n4035), .B2(n3613), .A(n3617), .ZN(n3503) );
  AOI211_X1 U4308 ( .C1(n4222), .C2(n3505), .A(n3504), .B(n3503), .ZN(n3506)
         );
  OAI21_X1 U4309 ( .B1(n3508), .B2(n3507), .A(n3506), .ZN(n3509) );
  OAI21_X1 U4310 ( .B1(n4222), .B2(n4229), .A(n3509), .ZN(n3625) );
  INV_X1 U4311 ( .A(n4038), .ZN(n3510) );
  INV_X1 U4312 ( .A(n4057), .ZN(n4060) );
  NAND2_X1 U4313 ( .A1(n4074), .A2(n3511), .ZN(n4099) );
  INV_X1 U4314 ( .A(n4099), .ZN(n3546) );
  INV_X1 U4315 ( .A(n3878), .ZN(n3513) );
  NAND2_X1 U4316 ( .A1(n3513), .A2(n3512), .ZN(n4085) );
  NAND2_X1 U4317 ( .A1(n3515), .A2(n3514), .ZN(n4051) );
  NAND2_X1 U4318 ( .A1(n3601), .A2(n3706), .ZN(n3646) );
  INV_X1 U4319 ( .A(n3646), .ZN(n3650) );
  NAND4_X1 U4320 ( .A1(n3518), .A2(n3650), .A3(n3517), .A4(n3516), .ZN(n3523)
         );
  NAND2_X1 U4321 ( .A1(n3757), .A2(n3758), .ZN(n3746) );
  INV_X1 U4322 ( .A(n3746), .ZN(n3521) );
  NAND2_X1 U4323 ( .A1(n3737), .A2(n3736), .ZN(n3708) );
  INV_X1 U4324 ( .A(n3708), .ZN(n3520) );
  NAND4_X1 U4325 ( .A1(n3521), .A2(n3520), .A3(n3519), .A4(n3152), .ZN(n3522)
         );
  NOR2_X1 U4326 ( .A1(n3523), .A2(n3522), .ZN(n3543) );
  NAND4_X1 U4327 ( .A1(n3527), .A2(n3526), .A3(n3525), .A4(n3524), .ZN(n3534)
         );
  INV_X1 U4328 ( .A(n3528), .ZN(n3532) );
  NAND4_X1 U4329 ( .A1(n3532), .A2(n3531), .A3(n3530), .A4(n3529), .ZN(n3533)
         );
  NOR2_X1 U4330 ( .A1(n3534), .A2(n3533), .ZN(n3542) );
  NAND2_X1 U4331 ( .A1(n2688), .A2(n4493), .ZN(n3555) );
  AND2_X1 U4332 ( .A1(n3553), .A2(n3555), .ZN(n4501) );
  NAND2_X1 U4333 ( .A1(n3536), .A2(n3535), .ZN(n3620) );
  NOR2_X1 U4334 ( .A1(n3620), .A2(n3556), .ZN(n3538) );
  NAND4_X1 U4335 ( .A1(n4501), .A2(n3570), .A3(n3538), .A4(n3537), .ZN(n3540)
         );
  NOR2_X1 U4336 ( .A1(n3540), .A2(n3539), .ZN(n3541) );
  NAND3_X1 U4337 ( .A1(n3543), .A2(n3542), .A3(n3541), .ZN(n3544) );
  NOR3_X1 U4338 ( .A1(n4085), .A2(n4051), .A3(n3544), .ZN(n3545) );
  NAND4_X1 U4339 ( .A1(n4060), .A2(n4035), .A3(n3546), .A4(n3545), .ZN(n3552)
         );
  AND2_X1 U4340 ( .A1(n4133), .A2(n3606), .ZN(n4132) );
  NOR2_X1 U4341 ( .A1(n4288), .A2(n4196), .ZN(n3856) );
  NAND2_X1 U4342 ( .A1(n4288), .A2(n4196), .ZN(n3857) );
  INV_X1 U4343 ( .A(n3857), .ZN(n3548) );
  OR2_X1 U4344 ( .A1(n3856), .A2(n3548), .ZN(n4188) );
  INV_X1 U4345 ( .A(n4188), .ZN(n4191) );
  XNOR2_X1 U4346 ( .A(n4266), .B(n4144), .ZN(n4135) );
  NAND2_X1 U4347 ( .A1(n3549), .A2(n4096), .ZN(n4117) );
  XNOR2_X1 U4348 ( .A(n3950), .B(n3855), .ZN(n3762) );
  NOR4_X1 U4349 ( .A1(n4191), .A2(n4135), .A3(n4117), .A4(n3762), .ZN(n3550)
         );
  NAND3_X1 U4350 ( .A1(n4154), .A2(n4132), .A3(n3550), .ZN(n3551) );
  NOR2_X1 U4351 ( .A1(n3552), .A2(n3551), .ZN(n3623) );
  INV_X1 U4352 ( .A(n3553), .ZN(n3557) );
  OAI211_X1 U4353 ( .C1(n3557), .C2(n3556), .A(n3555), .B(n3554), .ZN(n3559)
         );
  NAND3_X1 U4354 ( .A1(n3559), .A2(n3558), .A3(n2870), .ZN(n3562) );
  NAND3_X1 U4355 ( .A1(n3562), .A2(n3561), .A3(n3560), .ZN(n3565) );
  NAND3_X1 U4356 ( .A1(n3565), .A2(n3564), .A3(n3563), .ZN(n3568) );
  NAND4_X1 U4357 ( .A1(n3568), .A2(n3567), .A3(n3577), .A4(n3566), .ZN(n3571)
         );
  NAND3_X1 U4358 ( .A1(n3571), .A2(n3570), .A3(n3569), .ZN(n3572) );
  NAND3_X1 U4359 ( .A1(n3572), .A2(n3579), .A3(n3578), .ZN(n3575) );
  AND3_X1 U4360 ( .A1(n3575), .A2(n3574), .A3(n3573), .ZN(n3583) );
  INV_X1 U4361 ( .A(n3585), .ZN(n3598) );
  INV_X1 U4362 ( .A(n3576), .ZN(n3580) );
  NAND4_X1 U4363 ( .A1(n3580), .A2(n3579), .A3(n3578), .A4(n3577), .ZN(n3581)
         );
  OAI22_X1 U4364 ( .A1(n3583), .A2(n3582), .B1(n3598), .B2(n3581), .ZN(n3588)
         );
  INV_X1 U4365 ( .A(n3584), .ZN(n3586) );
  AOI22_X1 U4366 ( .A1(n3588), .A2(n3587), .B1(n3586), .B2(n3585), .ZN(n3600)
         );
  NAND3_X1 U4367 ( .A1(n3595), .A2(n3590), .A3(n3589), .ZN(n3599) );
  INV_X1 U4368 ( .A(n3591), .ZN(n3596) );
  INV_X1 U4369 ( .A(n3592), .ZN(n3593) );
  AOI211_X1 U4370 ( .C1(n3596), .C2(n3595), .A(n3594), .B(n3593), .ZN(n3597)
         );
  OAI22_X1 U4371 ( .A1(n3600), .A2(n3599), .B1(n3598), .B2(n3597), .ZN(n3603)
         );
  INV_X1 U4372 ( .A(n3601), .ZN(n3602) );
  AOI21_X1 U4373 ( .B1(n3603), .B2(n3706), .A(n3602), .ZN(n3605) );
  INV_X1 U4374 ( .A(n3604), .ZN(n4129) );
  OAI21_X1 U4375 ( .B1(n3605), .B2(n4129), .A(n4130), .ZN(n3607) );
  NAND2_X1 U4376 ( .A1(n3607), .A2(n3606), .ZN(n3609) );
  AOI21_X1 U4377 ( .B1(n3610), .B2(n3609), .A(n3608), .ZN(n3612) );
  INV_X1 U4378 ( .A(n3876), .ZN(n3611) );
  OAI21_X1 U4379 ( .B1(n3612), .B2(n3611), .A(n3877), .ZN(n3616) );
  NOR2_X1 U4380 ( .A1(n4241), .A2(n4248), .ZN(n3615) );
  INV_X1 U4381 ( .A(n3613), .ZN(n3614) );
  AOI211_X1 U4382 ( .C1(n3879), .C2(n3616), .A(n3615), .B(n3614), .ZN(n3618)
         );
  NOR2_X1 U4383 ( .A1(n3618), .A2(n3617), .ZN(n3619) );
  AOI21_X1 U4384 ( .B1(n3621), .B2(n3620), .A(n3619), .ZN(n3622) );
  MUX2_X1 U4385 ( .A(n3623), .B(n3622), .S(n2700), .Z(n3624) );
  AOI21_X1 U4386 ( .B1(n3626), .B2(n3625), .A(n3624), .ZN(n3628) );
  XNOR2_X1 U4387 ( .A(n3628), .B(n3627), .ZN(n3634) );
  NAND2_X1 U4388 ( .A1(n3629), .A2(n4007), .ZN(n3630) );
  OAI211_X1 U4389 ( .C1(n3631), .C2(n3633), .A(n3630), .B(B_REG_SCAN_IN), .ZN(
        n3632) );
  OAI21_X1 U4390 ( .B1(n3634), .B2(n3633), .A(n3632), .ZN(U3239) );
  INV_X1 U4391 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3637) );
  AOI21_X1 U4392 ( .B1(n4536), .B2(n3636), .A(n3635), .ZN(n3639) );
  MUX2_X1 U4393 ( .A(n3637), .B(n3639), .S(n4565), .Z(n3638) );
  OAI21_X1 U4394 ( .B1(n3642), .B2(n4378), .A(n3638), .ZN(U3493) );
  MUX2_X1 U4395 ( .A(n3640), .B(n3639), .S(n4577), .Z(n3641) );
  OAI21_X1 U4396 ( .B1(n4313), .B2(n3642), .A(n3641), .ZN(U3531) );
  AOI21_X1 U4397 ( .B1(n4325), .B2(n4320), .A(n3643), .ZN(n3645) );
  NAND2_X1 U4398 ( .A1(n3647), .A2(n3646), .ZN(n3705) );
  OAI21_X1 U4399 ( .B1(n3647), .B2(n3646), .A(n3705), .ZN(n4324) );
  NAND2_X1 U4400 ( .A1(n3651), .A2(n3650), .ZN(n3707) );
  OAI211_X1 U4401 ( .C1(n3651), .C2(n3650), .A(n3707), .B(n4495), .ZN(n4322)
         );
  INV_X1 U4402 ( .A(n4322), .ZN(n3658) );
  OAI21_X1 U4403 ( .B1(n3653), .B2(n4314), .A(n2158), .ZN(n4317) );
  NOR2_X1 U4404 ( .A1(n4317), .A2(n4174), .ZN(n3657) );
  AOI22_X1 U4405 ( .A1(n3685), .A2(n4211), .B1(n4210), .B2(n4320), .ZN(n3655)
         );
  AOI22_X1 U4406 ( .A1(n4396), .A2(REG2_REG_16__SCAN_IN), .B1(n3693), .B2(
        n4502), .ZN(n3654) );
  OAI211_X1 U4407 ( .C1(n4316), .C2(n4207), .A(n3655), .B(n3654), .ZN(n3656)
         );
  AOI211_X1 U4408 ( .C1(n3658), .C2(n4505), .A(n3657), .B(n3656), .ZN(n3659)
         );
  OAI21_X1 U4409 ( .B1(n4324), .B2(n4182), .A(n3659), .ZN(U3274) );
  INV_X1 U4410 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4756) );
  AOI22_X1 U4411 ( .A1(n4320), .A2(n4327), .B1(n4326), .B2(n3660), .ZN(n3661)
         );
  OAI21_X1 U4412 ( .B1(n3662), .B2(n4330), .A(n3661), .ZN(n3665) );
  NOR2_X1 U4413 ( .A1(n3663), .A2(n4543), .ZN(n3664) );
  AOI211_X1 U4414 ( .C1(n3666), .C2(n4495), .A(n3665), .B(n3664), .ZN(n3668)
         );
  MUX2_X1 U4415 ( .A(n4756), .B(n3668), .S(n4565), .Z(n3667) );
  OAI21_X1 U4416 ( .B1(n3670), .B2(n4378), .A(n3667), .ZN(U3495) );
  MUX2_X1 U4417 ( .A(n4766), .B(n3668), .S(n4577), .Z(n3669) );
  OAI21_X1 U4418 ( .B1(n4313), .B2(n3670), .A(n3669), .ZN(U3532) );
  AND2_X1 U4419 ( .A1(n3825), .A2(n4325), .ZN(n3671) );
  AOI21_X1 U4420 ( .B1(n4320), .B2(n3830), .A(n3671), .ZN(n3719) );
  NAND2_X1 U4421 ( .A1(n3674), .A2(n3675), .ZN(n3673) );
  NAND2_X1 U4422 ( .A1(n3673), .A2(n3672), .ZN(n3679) );
  INV_X1 U4423 ( .A(n3674), .ZN(n3677) );
  INV_X1 U4424 ( .A(n3675), .ZN(n3676) );
  NAND2_X1 U4425 ( .A1(n3677), .A2(n3676), .ZN(n3678) );
  NAND2_X1 U4426 ( .A1(n3679), .A2(n3678), .ZN(n3684) );
  NAND2_X1 U4427 ( .A1(n4320), .A2(n3825), .ZN(n3681) );
  NAND2_X1 U4428 ( .A1(n4325), .A2(n3843), .ZN(n3680) );
  NAND2_X1 U4429 ( .A1(n3681), .A2(n3680), .ZN(n3682) );
  XNOR2_X1 U4430 ( .A(n3682), .B(n2805), .ZN(n3683) );
  NAND2_X1 U4431 ( .A1(n3684), .A2(n3683), .ZN(n3717) );
  AOI21_X1 U4432 ( .B1(n3719), .B2(n3717), .A(n3720), .ZN(n3689) );
  OAI22_X1 U4433 ( .A1(n3730), .A2(n3838), .B1(n3837), .B2(n4314), .ZN(n3721)
         );
  NAND2_X1 U4434 ( .A1(n4328), .A2(n3825), .ZN(n3687) );
  NAND2_X1 U4435 ( .A1(n3685), .A2(n3843), .ZN(n3686) );
  NAND2_X1 U4436 ( .A1(n3687), .A2(n3686), .ZN(n3688) );
  XNOR2_X1 U4437 ( .A(n3688), .B(n2805), .ZN(n3722) );
  XOR2_X1 U4438 ( .A(n3721), .B(n3722), .Z(n3718) );
  XNOR2_X1 U4439 ( .A(n3689), .B(n3718), .ZN(n3695) );
  NAND2_X1 U4440 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4464) );
  OAI21_X1 U4441 ( .B1(n3982), .B2(n4316), .A(n4464), .ZN(n3692) );
  OAI22_X1 U4442 ( .A1(n3980), .A2(n4314), .B1(n3690), .B2(n3949), .ZN(n3691)
         );
  AOI211_X1 U4443 ( .C1(n3693), .C2(n3985), .A(n3692), .B(n3691), .ZN(n3694)
         );
  OAI21_X1 U4444 ( .B1(n3695), .B2(n3988), .A(n3694), .ZN(U3223) );
  INV_X1 U4445 ( .A(n3720), .ZN(n3696) );
  NAND2_X1 U4446 ( .A1(n3696), .A2(n3717), .ZN(n3697) );
  XNOR2_X1 U4447 ( .A(n3697), .B(n3719), .ZN(n3703) );
  AND2_X1 U4448 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4457) );
  OAI22_X1 U4449 ( .A1(n3980), .A2(n3698), .B1(n4331), .B2(n3949), .ZN(n3699)
         );
  AOI211_X1 U4450 ( .C1(n3970), .C2(n4328), .A(n4457), .B(n3699), .ZN(n3702)
         );
  NAND2_X1 U4451 ( .A1(n3985), .A2(n3700), .ZN(n3701) );
  OAI211_X1 U4452 ( .C1(n3703), .C2(n3988), .A(n3702), .B(n3701), .ZN(U3238)
         );
  NAND2_X1 U4453 ( .A1(n3705), .A2(n3704), .ZN(n3745) );
  XOR2_X1 U4454 ( .A(n3708), .B(n3745), .Z(n4311) );
  INV_X1 U4455 ( .A(n4311), .ZN(n3716) );
  XOR2_X1 U4456 ( .A(n3708), .B(n4185), .Z(n3711) );
  OAI22_X1 U4457 ( .A1(n3907), .A2(n4497), .B1(n4315), .B2(n3741), .ZN(n3709)
         );
  AOI21_X1 U4458 ( .B1(n4321), .B2(n4328), .A(n3709), .ZN(n3710) );
  OAI21_X1 U4459 ( .B1(n3711), .B2(n4297), .A(n3710), .ZN(n4310) );
  NAND2_X1 U4460 ( .A1(n2158), .A2(n3742), .ZN(n3712) );
  NAND2_X1 U4461 ( .A1(n2137), .A2(n3712), .ZN(n4379) );
  AOI22_X1 U4462 ( .A1(n4396), .A2(REG2_REG_17__SCAN_IN), .B1(n3732), .B2(
        n4502), .ZN(n3713) );
  OAI21_X1 U4463 ( .B1(n4379), .B2(n4174), .A(n3713), .ZN(n3714) );
  AOI21_X1 U4464 ( .B1(n4310), .B2(n4505), .A(n3714), .ZN(n3715) );
  OAI21_X1 U4465 ( .B1(n3716), .B2(n4182), .A(n3715), .ZN(U3273) );
  OAI211_X1 U4466 ( .C1(n3720), .C2(n3719), .A(n3718), .B(n3717), .ZN(n3724)
         );
  NAND2_X1 U4467 ( .A1(n3724), .A2(n3723), .ZN(n3774) );
  OAI22_X1 U4468 ( .A1(n4316), .A2(n3837), .B1(n3835), .B2(n3741), .ZN(n3726)
         );
  XNOR2_X1 U4469 ( .A(n3726), .B(n3725), .ZN(n3775) );
  OR2_X1 U4470 ( .A1(n4316), .A2(n3838), .ZN(n3728) );
  NAND2_X1 U4471 ( .A1(n3742), .A2(n3825), .ZN(n3727) );
  XNOR2_X1 U4472 ( .A(n3775), .B(n3776), .ZN(n3729) );
  XNOR2_X1 U4473 ( .A(n3774), .B(n3729), .ZN(n3735) );
  AND2_X1 U4474 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4025) );
  OAI22_X1 U4475 ( .A1(n3980), .A2(n3741), .B1(n3730), .B2(n3949), .ZN(n3731)
         );
  AOI211_X1 U4476 ( .C1(n3970), .C2(n3990), .A(n4025), .B(n3731), .ZN(n3734)
         );
  NAND2_X1 U4477 ( .A1(n3985), .A2(n3732), .ZN(n3733) );
  OAI211_X1 U4478 ( .C1(n3735), .C2(n3988), .A(n3734), .B(n3733), .ZN(U3225)
         );
  INV_X1 U4479 ( .A(n3736), .ZN(n4184) );
  OAI21_X1 U4480 ( .B1(n4185), .B2(n4184), .A(n3737), .ZN(n3760) );
  XOR2_X1 U4481 ( .A(n3746), .B(n3760), .Z(n3740) );
  AOI22_X1 U4482 ( .A1(n4295), .A2(n4327), .B1(n3766), .B2(n4326), .ZN(n3738)
         );
  OAI21_X1 U4483 ( .B1(n4316), .B2(n4330), .A(n3738), .ZN(n3739) );
  AOI21_X1 U4484 ( .B1(n3740), .B2(n4495), .A(n3739), .ZN(n4308) );
  NAND2_X1 U4485 ( .A1(n4316), .A2(n3741), .ZN(n3744) );
  OAI21_X1 U4486 ( .B1(n3747), .B2(n3746), .A(n3756), .ZN(n4306) );
  XNOR2_X1 U4487 ( .A(n2137), .B(n3968), .ZN(n3748) );
  NAND2_X1 U4488 ( .A1(n3748), .A2(n4562), .ZN(n4307) );
  INV_X1 U4489 ( .A(n3749), .ZN(n3750) );
  NOR2_X1 U4490 ( .A1(n4307), .A2(n3750), .ZN(n3753) );
  INV_X1 U4491 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3751) );
  OAI22_X1 U4492 ( .A1(n4505), .A2(n3751), .B1(n3973), .B2(n4162), .ZN(n3752)
         );
  AOI211_X1 U4493 ( .C1(n4306), .C2(n4192), .A(n3753), .B(n3752), .ZN(n3754)
         );
  OAI21_X1 U4494 ( .B1(n4396), .B2(n4308), .A(n3754), .ZN(U3272) );
  XNOR2_X1 U4495 ( .A(n3854), .B(n3762), .ZN(n4304) );
  INV_X1 U4496 ( .A(n4304), .ZN(n3773) );
  INV_X1 U4497 ( .A(n3757), .ZN(n3759) );
  OAI21_X1 U4498 ( .B1(n3760), .B2(n3759), .A(n3758), .ZN(n3761) );
  XOR2_X1 U4499 ( .A(n3762), .B(n3761), .Z(n3765) );
  OAI22_X1 U4500 ( .A1(n3907), .A2(n4330), .B1(n4315), .B2(n3908), .ZN(n3763)
         );
  AOI21_X1 U4501 ( .B1(n4327), .B2(n4288), .A(n3763), .ZN(n3764) );
  OAI21_X1 U4502 ( .B1(n3765), .B2(n4297), .A(n3764), .ZN(n4303) );
  OAI21_X1 U4503 ( .B1(n2137), .B2(n3766), .A(n3855), .ZN(n3767) );
  INV_X1 U4504 ( .A(n3767), .ZN(n3769) );
  NAND2_X1 U4505 ( .A1(n3968), .A2(n3908), .ZN(n3768) );
  OR2_X1 U4506 ( .A1(n3769), .A2(n4195), .ZN(n4373) );
  AOI22_X1 U4507 ( .A1(n4396), .A2(REG2_REG_19__SCAN_IN), .B1(n3911), .B2(
        n4502), .ZN(n3770) );
  OAI21_X1 U4508 ( .B1(n4373), .B2(n4174), .A(n3770), .ZN(n3771) );
  AOI21_X1 U4509 ( .B1(n4303), .B2(n4505), .A(n3771), .ZN(n3772) );
  OAI21_X1 U4510 ( .B1(n3773), .B2(n4182), .A(n3772), .ZN(U3271) );
  INV_X1 U4511 ( .A(n3775), .ZN(n3779) );
  INV_X1 U4512 ( .A(n3776), .ZN(n3778) );
  OAI22_X1 U4513 ( .A1(n3907), .A2(n3837), .B1(n3835), .B2(n3968), .ZN(n3780)
         );
  XNOR2_X1 U4514 ( .A(n3780), .B(n2805), .ZN(n3782) );
  OAI22_X1 U4515 ( .A1(n3907), .A2(n3838), .B1(n3837), .B2(n3968), .ZN(n3781)
         );
  NOR2_X1 U4516 ( .A1(n3782), .A2(n3781), .ZN(n3963) );
  OAI22_X1 U4517 ( .A1(n3950), .A2(n3837), .B1(n3835), .B2(n3908), .ZN(n3783)
         );
  XNOR2_X1 U4518 ( .A(n3783), .B(n2805), .ZN(n3785) );
  OAI22_X1 U4519 ( .A1(n3950), .A2(n3838), .B1(n3837), .B2(n3908), .ZN(n3784)
         );
  XNOR2_X1 U4520 ( .A(n3785), .B(n3784), .ZN(n3905) );
  NAND2_X1 U4521 ( .A1(n4288), .A2(n3825), .ZN(n3787) );
  OR2_X1 U4522 ( .A1(n4292), .A2(n3835), .ZN(n3786) );
  NAND2_X1 U4523 ( .A1(n3787), .A2(n3786), .ZN(n3788) );
  XNOR2_X1 U4524 ( .A(n3788), .B(n3725), .ZN(n3791) );
  NOR2_X1 U4525 ( .A1(n3837), .A2(n4292), .ZN(n3789) );
  AOI21_X1 U4526 ( .B1(n4288), .B2(n3830), .A(n3789), .ZN(n3790) );
  OR2_X1 U4527 ( .A1(n3791), .A2(n3790), .ZN(n3944) );
  NAND2_X1 U4528 ( .A1(n3791), .A2(n3790), .ZN(n3946) );
  NAND2_X1 U4529 ( .A1(n4156), .A2(n3825), .ZN(n3793) );
  OR2_X1 U4530 ( .A1(n3835), .A2(n4283), .ZN(n3792) );
  NAND2_X1 U4531 ( .A1(n3793), .A2(n3792), .ZN(n3794) );
  XNOR2_X1 U4532 ( .A(n3794), .B(n2805), .ZN(n3915) );
  NAND2_X1 U4533 ( .A1(n4156), .A2(n3830), .ZN(n3796) );
  OR2_X1 U4534 ( .A1(n3837), .A2(n4283), .ZN(n3795) );
  NAND2_X1 U4535 ( .A1(n3796), .A2(n3795), .ZN(n3914) );
  NOR2_X1 U4536 ( .A1(n3915), .A2(n3914), .ZN(n3799) );
  INV_X1 U4537 ( .A(n3915), .ZN(n3798) );
  INV_X1 U4538 ( .A(n3914), .ZN(n3797) );
  AOI22_X1 U4539 ( .A1(n4139), .A2(n3825), .B1(n3843), .B2(n4161), .ZN(n3800)
         );
  XNOR2_X1 U4540 ( .A(n3800), .B(n2805), .ZN(n3805) );
  AOI22_X1 U4541 ( .A1(n4139), .A2(n3830), .B1(n3825), .B2(n4161), .ZN(n3806)
         );
  XNOR2_X1 U4542 ( .A(n3805), .B(n3806), .ZN(n3956) );
  NAND2_X1 U4543 ( .A1(n4266), .A2(n3825), .ZN(n3802) );
  OR2_X1 U4544 ( .A1(n3835), .A2(n4144), .ZN(n3801) );
  NAND2_X1 U4545 ( .A1(n3802), .A2(n3801), .ZN(n3803) );
  XNOR2_X1 U4546 ( .A(n3803), .B(n3725), .ZN(n3811) );
  NOR2_X1 U4547 ( .A1(n3837), .A2(n4144), .ZN(n3804) );
  AOI21_X1 U4548 ( .B1(n4266), .B2(n3830), .A(n3804), .ZN(n3810) );
  XNOR2_X1 U4549 ( .A(n3811), .B(n3810), .ZN(n3895) );
  INV_X1 U4550 ( .A(n3805), .ZN(n3808) );
  INV_X1 U4551 ( .A(n3806), .ZN(n3807) );
  NOR2_X1 U4552 ( .A1(n3808), .A2(n3807), .ZN(n3896) );
  NAND2_X1 U4553 ( .A1(n3862), .A2(n3830), .ZN(n3813) );
  OR2_X1 U4554 ( .A1(n3837), .A2(n4120), .ZN(n3812) );
  NAND2_X1 U4555 ( .A1(n3813), .A2(n3812), .ZN(n3817) );
  INV_X1 U4556 ( .A(n3817), .ZN(n3814) );
  NAND2_X1 U4557 ( .A1(n3898), .A2(n2309), .ZN(n3815) );
  OAI22_X1 U4558 ( .A1(n4142), .A2(n3837), .B1(n3835), .B2(n4120), .ZN(n3816)
         );
  XOR2_X1 U4559 ( .A(n2805), .B(n3816), .Z(n3935) );
  INV_X1 U4560 ( .A(n3898), .ZN(n3818) );
  NAND2_X1 U4561 ( .A1(n4080), .A2(n3825), .ZN(n3820) );
  OR2_X1 U4562 ( .A1(n3835), .A2(n4105), .ZN(n3819) );
  NAND2_X1 U4563 ( .A1(n3820), .A2(n3819), .ZN(n3821) );
  XNOR2_X1 U4564 ( .A(n3821), .B(n3725), .ZN(n3824) );
  NOR2_X1 U4565 ( .A1(n3837), .A2(n4105), .ZN(n3822) );
  AOI21_X1 U4566 ( .B1(n4080), .B2(n3830), .A(n3822), .ZN(n3823) );
  NOR2_X1 U4567 ( .A1(n3824), .A2(n3823), .ZN(n3925) );
  NAND2_X1 U4568 ( .A1(n4249), .A2(n3825), .ZN(n3827) );
  OR2_X1 U4569 ( .A1(n3835), .A2(n4088), .ZN(n3826) );
  NAND2_X1 U4570 ( .A1(n3827), .A2(n3826), .ZN(n3828) );
  XNOR2_X1 U4571 ( .A(n3828), .B(n3725), .ZN(n3834) );
  INV_X1 U4572 ( .A(n3834), .ZN(n3832) );
  NOR2_X1 U4573 ( .A1(n3837), .A2(n4088), .ZN(n3829) );
  AOI21_X1 U4574 ( .B1(n4249), .B2(n3830), .A(n3829), .ZN(n3833) );
  INV_X1 U4575 ( .A(n3833), .ZN(n3831) );
  NAND2_X1 U4576 ( .A1(n3832), .A2(n3831), .ZN(n3976) );
  AND2_X1 U4577 ( .A1(n3834), .A2(n3833), .ZN(n3975) );
  OAI22_X1 U4578 ( .A1(n4241), .A2(n3837), .B1(n4048), .B2(n3835), .ZN(n3836)
         );
  XNOR2_X1 U4579 ( .A(n3836), .B(n3725), .ZN(n3839) );
  OAI22_X1 U4580 ( .A1(n4241), .A2(n3838), .B1(n4048), .B2(n3837), .ZN(n3840)
         );
  XNOR2_X1 U4581 ( .A(n3839), .B(n3840), .ZN(n3887) );
  INV_X1 U4582 ( .A(n3839), .ZN(n3841) );
  INV_X1 U4583 ( .A(n4067), .ZN(n4237) );
  AOI22_X1 U4584 ( .A1(n4247), .A2(n3830), .B1(n3825), .B2(n4237), .ZN(n3842)
         );
  XNOR2_X1 U4585 ( .A(n3842), .B(n2805), .ZN(n3845) );
  AOI22_X1 U4586 ( .A1(n4247), .A2(n3825), .B1(n3843), .B2(n4237), .ZN(n3844)
         );
  XNOR2_X1 U4587 ( .A(n3845), .B(n3844), .ZN(n3846) );
  XNOR2_X1 U4588 ( .A(n3847), .B(n3846), .ZN(n3852) );
  OAI22_X1 U4589 ( .A1(n4241), .A2(n3949), .B1(n3980), .B2(n4067), .ZN(n3850)
         );
  INV_X1 U4590 ( .A(n4238), .ZN(n4578) );
  OAI22_X1 U4591 ( .A1(n4578), .A2(n3982), .B1(STATE_REG_SCAN_IN), .B2(n3848), 
        .ZN(n3849) );
  AOI211_X1 U4592 ( .C1(n4065), .C2(n3985), .A(n3850), .B(n3849), .ZN(n3851)
         );
  OAI21_X1 U4593 ( .B1(n3852), .B2(n3988), .A(n3851), .ZN(U3217) );
  INV_X1 U4594 ( .A(n4156), .ZN(n4293) );
  NOR2_X1 U4595 ( .A1(n4293), .A2(n4283), .ZN(n3859) );
  NOR2_X1 U4596 ( .A1(n4266), .A2(n4138), .ZN(n3861) );
  NOR2_X1 U4597 ( .A1(n4142), .A2(n4120), .ZN(n3863) );
  INV_X1 U4598 ( .A(n4105), .ZN(n3865) );
  NOR2_X1 U4599 ( .A1(n4080), .A2(n3865), .ZN(n4081) );
  INV_X1 U4600 ( .A(n4249), .ZN(n3929) );
  AND2_X1 U4601 ( .A1(n3929), .A2(n4088), .ZN(n3868) );
  OR2_X1 U4602 ( .A1(n4081), .A2(n3868), .ZN(n3864) );
  NOR2_X1 U4603 ( .A1(n4095), .A2(n3864), .ZN(n3870) );
  NAND2_X1 U4604 ( .A1(n4080), .A2(n3865), .ZN(n4082) );
  OR2_X1 U4605 ( .A1(n3929), .A2(n4088), .ZN(n3866) );
  AND2_X1 U4606 ( .A1(n4082), .A2(n3866), .ZN(n3867) );
  NOR2_X1 U4607 ( .A1(n3868), .A2(n3867), .ZN(n3869) );
  XNOR2_X1 U4608 ( .A(n4050), .B(n4035), .ZN(n4256) );
  OR2_X1 U4609 ( .A1(n4086), .A2(n4048), .ZN(n3871) );
  AND2_X1 U4610 ( .A1(n3871), .A2(n4062), .ZN(n4253) );
  INV_X1 U4611 ( .A(n4247), .ZN(n3889) );
  AOI22_X1 U4612 ( .A1(n3892), .A2(n4502), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4396), .ZN(n3873) );
  AOI22_X1 U4613 ( .A1(n4249), .A2(n4210), .B1(n4248), .B2(n4211), .ZN(n3872)
         );
  OAI211_X1 U4614 ( .C1(n3889), .C2(n4207), .A(n3873), .B(n3872), .ZN(n3882)
         );
  NAND2_X1 U4615 ( .A1(n4097), .A2(n3877), .ZN(n4075) );
  AOI21_X1 U4616 ( .B1(n4075), .B2(n3879), .A(n3878), .ZN(n4036) );
  XNOR2_X1 U4617 ( .A(n4036), .B(n4035), .ZN(n3880) );
  NAND2_X1 U4618 ( .A1(n3880), .A2(n4495), .ZN(n4254) );
  NOR2_X1 U4619 ( .A1(n4254), .A2(n4396), .ZN(n3881) );
  AOI211_X1 U4620 ( .C1(n4399), .C2(n4253), .A(n3882), .B(n3881), .ZN(n3883)
         );
  OAI21_X1 U4621 ( .B1(n4256), .B2(n4182), .A(n3883), .ZN(U3263) );
  NAND3_X1 U4622 ( .A1(n3884), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3886) );
  INV_X1 U4623 ( .A(DATAI_31_), .ZN(n3885) );
  OAI22_X1 U4624 ( .A1(n2517), .A2(n3886), .B1(STATE_REG_SCAN_IN), .B2(n3885), 
        .ZN(U3321) );
  XNOR2_X1 U4625 ( .A(n3888), .B(n3887), .ZN(n3894) );
  INV_X1 U4626 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4864) );
  OAI22_X1 U4627 ( .A1(n3929), .A2(n3949), .B1(STATE_REG_SCAN_IN), .B2(n4864), 
        .ZN(n3891) );
  OAI22_X1 U4628 ( .A1(n3889), .A2(n3982), .B1(n3980), .B2(n4048), .ZN(n3890)
         );
  AOI211_X1 U4629 ( .C1(n3892), .C2(n3985), .A(n3891), .B(n3890), .ZN(n3893)
         );
  OAI21_X1 U4630 ( .B1(n3894), .B2(n3988), .A(n3893), .ZN(U3211) );
  OAI21_X1 U4631 ( .B1(n2144), .B2(n3896), .A(n3895), .ZN(n3897) );
  NAND3_X1 U4632 ( .A1(n3898), .A2(n3966), .A3(n3897), .ZN(n3903) );
  INV_X1 U4633 ( .A(n4139), .ZN(n4284) );
  OAI22_X1 U4634 ( .A1(n3980), .A2(n4144), .B1(n4284), .B2(n3949), .ZN(n3901)
         );
  OAI22_X1 U4635 ( .A1(n4142), .A2(n3982), .B1(STATE_REG_SCAN_IN), .B2(n3899), 
        .ZN(n3900) );
  AOI211_X1 U4636 ( .C1(n4146), .C2(n3985), .A(n3901), .B(n3900), .ZN(n3902)
         );
  NAND2_X1 U4637 ( .A1(n3903), .A2(n3902), .ZN(U3213) );
  XOR2_X1 U4638 ( .A(n3905), .B(n3904), .Z(n3913) );
  INV_X1 U4639 ( .A(n4288), .ZN(n3920) );
  OAI21_X1 U4640 ( .B1(n3982), .B2(n3920), .A(n3906), .ZN(n3910) );
  OAI22_X1 U4641 ( .A1(n3980), .A2(n3908), .B1(n3907), .B2(n3949), .ZN(n3909)
         );
  AOI211_X1 U4642 ( .C1(n3911), .C2(n3985), .A(n3910), .B(n3909), .ZN(n3912)
         );
  OAI21_X1 U4643 ( .B1(n3913), .B2(n3988), .A(n3912), .ZN(U3216) );
  XNOR2_X1 U4644 ( .A(n3915), .B(n3914), .ZN(n3916) );
  XNOR2_X1 U4645 ( .A(n3917), .B(n3916), .ZN(n3924) );
  INV_X1 U4646 ( .A(n3918), .ZN(n4175) );
  OAI22_X1 U4647 ( .A1(n3982), .A2(n4284), .B1(STATE_REG_SCAN_IN), .B2(n3919), 
        .ZN(n3922) );
  OAI22_X1 U4648 ( .A1(n3980), .A2(n4283), .B1(n3920), .B2(n3949), .ZN(n3921)
         );
  AOI211_X1 U4649 ( .C1(n4175), .C2(n3985), .A(n3922), .B(n3921), .ZN(n3923)
         );
  OAI21_X1 U4650 ( .B1(n3924), .B2(n3988), .A(n3923), .ZN(U3220) );
  NOR2_X1 U4651 ( .A1(n3925), .A2(n2157), .ZN(n3926) );
  XNOR2_X1 U4652 ( .A(n3927), .B(n3926), .ZN(n3933) );
  OAI22_X1 U4653 ( .A1(n4142), .A2(n3949), .B1(n3980), .B2(n4105), .ZN(n3931)
         );
  OAI22_X1 U4654 ( .A1(n3929), .A2(n3982), .B1(STATE_REG_SCAN_IN), .B2(n3928), 
        .ZN(n3930) );
  AOI211_X1 U4655 ( .C1(n4106), .C2(n3985), .A(n3931), .B(n3930), .ZN(n3932)
         );
  OAI21_X1 U4656 ( .B1(n3933), .B2(n3988), .A(n3932), .ZN(U3222) );
  NAND2_X1 U4657 ( .A1(n3815), .A2(n3934), .ZN(n3936) );
  XNOR2_X1 U4658 ( .A(n3936), .B(n3935), .ZN(n3941) );
  INV_X1 U4659 ( .A(n3937), .ZN(n4122) );
  OAI22_X1 U4660 ( .A1(n4158), .A2(n3949), .B1(STATE_REG_SCAN_IN), .B2(n4661), 
        .ZN(n3939) );
  INV_X1 U4661 ( .A(n4080), .ZN(n4269) );
  OAI22_X1 U4662 ( .A1(n4269), .A2(n3982), .B1(n3980), .B2(n4120), .ZN(n3938)
         );
  AOI211_X1 U4663 ( .C1(n4122), .C2(n3985), .A(n3939), .B(n3938), .ZN(n3940)
         );
  OAI21_X1 U4664 ( .B1(n3941), .B2(n3988), .A(n3940), .ZN(U3226) );
  INV_X1 U4665 ( .A(n3942), .ZN(n3947) );
  AOI21_X1 U4666 ( .B1(n3946), .B2(n3944), .A(n3943), .ZN(n3945) );
  AOI21_X1 U4667 ( .B1(n3947), .B2(n3946), .A(n3945), .ZN(n3954) );
  OAI22_X1 U4668 ( .A1(n3982), .A2(n4293), .B1(STATE_REG_SCAN_IN), .B2(n3948), 
        .ZN(n3952) );
  OAI22_X1 U4669 ( .A1(n3980), .A2(n4292), .B1(n3950), .B2(n3949), .ZN(n3951)
         );
  AOI211_X1 U4670 ( .C1(n4197), .C2(n3985), .A(n3952), .B(n3951), .ZN(n3953)
         );
  OAI21_X1 U4671 ( .B1(n3954), .B2(n3988), .A(n3953), .ZN(U3230) );
  AOI21_X1 U4672 ( .B1(n3956), .B2(n3955), .A(n2144), .ZN(n3962) );
  INV_X1 U4673 ( .A(n4163), .ZN(n3960) );
  OAI22_X1 U4674 ( .A1(n4158), .A2(n3982), .B1(STATE_REG_SCAN_IN), .B2(n4862), 
        .ZN(n3959) );
  OAI22_X1 U4675 ( .A1(n3980), .A2(n3957), .B1(n4293), .B2(n3949), .ZN(n3958)
         );
  AOI211_X1 U4676 ( .C1(n3960), .C2(n3985), .A(n3959), .B(n3958), .ZN(n3961)
         );
  OAI21_X1 U4677 ( .B1(n3962), .B2(n3988), .A(n3961), .ZN(U3232) );
  NOR2_X1 U4678 ( .A1(n3963), .A2(n2165), .ZN(n3964) );
  XNOR2_X1 U4679 ( .A(n3965), .B(n3964), .ZN(n3967) );
  NAND2_X1 U4680 ( .A1(n3967), .A2(n3966), .ZN(n3972) );
  AND2_X1 U4681 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4482) );
  OAI22_X1 U4682 ( .A1(n3980), .A2(n3968), .B1(n4316), .B2(n3949), .ZN(n3969)
         );
  AOI211_X1 U4683 ( .C1(n3970), .C2(n4295), .A(n4482), .B(n3969), .ZN(n3971)
         );
  OAI211_X1 U4684 ( .C1(n3974), .C2(n3973), .A(n3972), .B(n3971), .ZN(U3235)
         );
  INV_X1 U4685 ( .A(n3975), .ZN(n3977) );
  NAND2_X1 U4686 ( .A1(n3977), .A2(n3976), .ZN(n3978) );
  XNOR2_X1 U4687 ( .A(n3979), .B(n3978), .ZN(n3989) );
  INV_X1 U4688 ( .A(n4090), .ZN(n3986) );
  OAI22_X1 U4689 ( .A1(n4269), .A2(n3949), .B1(n3980), .B2(n4088), .ZN(n3984)
         );
  INV_X1 U4690 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3981) );
  OAI22_X1 U4691 ( .A1(n4241), .A2(n3982), .B1(STATE_REG_SCAN_IN), .B2(n3981), 
        .ZN(n3983) );
  AOI211_X1 U4692 ( .C1(n3986), .C2(n3985), .A(n3984), .B(n3983), .ZN(n3987)
         );
  OAI21_X1 U4693 ( .B1(n3989), .B2(n3988), .A(n3987), .ZN(U3237) );
  MUX2_X1 U4694 ( .A(n4247), .B(DATAO_REG_28__SCAN_IN), .S(n3994), .Z(U3578)
         );
  INV_X1 U4695 ( .A(n4241), .ZN(n4047) );
  MUX2_X1 U4696 ( .A(n4047), .B(DATAO_REG_27__SCAN_IN), .S(n3994), .Z(U3577)
         );
  MUX2_X1 U4697 ( .A(n4080), .B(DATAO_REG_25__SCAN_IN), .S(n3994), .Z(U3575)
         );
  MUX2_X1 U4698 ( .A(n4266), .B(DATAO_REG_23__SCAN_IN), .S(n3994), .Z(U3573)
         );
  MUX2_X1 U4699 ( .A(n4156), .B(DATAO_REG_21__SCAN_IN), .S(n3994), .Z(U3571)
         );
  MUX2_X1 U4700 ( .A(DATAO_REG_20__SCAN_IN), .B(n4288), .S(U4043), .Z(U3570)
         );
  MUX2_X1 U4701 ( .A(DATAO_REG_18__SCAN_IN), .B(n3990), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4702 ( .A(n4320), .B(DATAO_REG_15__SCAN_IN), .S(n3994), .Z(U3565)
         );
  MUX2_X1 U4703 ( .A(n3991), .B(DATAO_REG_10__SCAN_IN), .S(n3994), .Z(U3560)
         );
  MUX2_X1 U4704 ( .A(n3992), .B(DATAO_REG_6__SCAN_IN), .S(n3994), .Z(U3556) );
  MUX2_X1 U4705 ( .A(DATAO_REG_5__SCAN_IN), .B(n3993), .S(U4043), .Z(U3555) );
  MUX2_X1 U4706 ( .A(n2983), .B(DATAO_REG_4__SCAN_IN), .S(n3994), .Z(U3554) );
  MUX2_X1 U4707 ( .A(n2762), .B(DATAO_REG_1__SCAN_IN), .S(n3994), .Z(U3551) );
  OAI211_X1 U4708 ( .C1(n4006), .C2(n3995), .A(n4488), .B(n4015), .ZN(n4002)
         );
  OAI211_X1 U4709 ( .C1(n3998), .C2(n3997), .A(n4474), .B(n3996), .ZN(n4001)
         );
  AOI22_X1 U4710 ( .A1(n4483), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4000) );
  NAND2_X1 U4711 ( .A1(n4450), .A2(n4392), .ZN(n3999) );
  NAND4_X1 U4712 ( .A1(n4002), .A2(n4001), .A3(n4000), .A4(n3999), .ZN(U3241)
         );
  NAND3_X1 U4713 ( .A1(n4004), .A2(n4382), .A3(n4003), .ZN(n4009) );
  AOI22_X1 U4714 ( .A1(n4007), .A2(n4006), .B1(n4005), .B2(n4669), .ZN(n4008)
         );
  NAND3_X1 U4715 ( .A1(n4009), .A2(U4043), .A3(n4008), .ZN(n4413) );
  AOI22_X1 U4716 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4483), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4020) );
  XOR2_X1 U4717 ( .A(n4011), .B(n4010), .Z(n4012) );
  AOI22_X1 U4718 ( .A1(n2136), .A2(n4450), .B1(n4474), .B2(n4012), .ZN(n4019)
         );
  MUX2_X1 U4719 ( .A(n4206), .B(REG2_REG_2__SCAN_IN), .S(n2136), .Z(n4013) );
  NAND3_X1 U4720 ( .A1(n4015), .A2(n4014), .A3(n4013), .ZN(n4016) );
  NAND3_X1 U4721 ( .A1(n4488), .A2(n4017), .A3(n4016), .ZN(n4018) );
  NAND4_X1 U4722 ( .A1(n4413), .A2(n4020), .A3(n4019), .A4(n4018), .ZN(U3242)
         );
  OAI21_X1 U4723 ( .B1(n4023), .B2(n4022), .A(n4021), .ZN(n4024) );
  AOI22_X1 U4724 ( .A1(n4385), .A2(n4450), .B1(n4474), .B2(n4024), .ZN(n4032)
         );
  AOI21_X1 U4725 ( .B1(n4483), .B2(ADDR_REG_17__SCAN_IN), .A(n4025), .ZN(n4031) );
  OAI21_X1 U4726 ( .B1(n4028), .B2(n4027), .A(n4026), .ZN(n4029) );
  NAND2_X1 U4727 ( .A1(n4488), .A2(n4029), .ZN(n4030) );
  NAND3_X1 U4728 ( .A1(n4032), .A2(n4031), .A3(n4030), .ZN(U3257) );
  INV_X1 U4729 ( .A(n4033), .ZN(n4046) );
  AOI21_X1 U4730 ( .B1(n4036), .B2(n4035), .A(n4034), .ZN(n4058) );
  INV_X1 U4731 ( .A(n4058), .ZN(n4039) );
  AOI21_X1 U4732 ( .B1(n4039), .B2(n4038), .A(n4037), .ZN(n4040) );
  XOR2_X1 U4733 ( .A(n4051), .B(n4040), .Z(n4045) );
  AOI21_X1 U4734 ( .B1(B_REG_SCAN_IN), .B2(n4383), .A(n4497), .ZN(n4220) );
  INV_X1 U4735 ( .A(n4041), .ZN(n4053) );
  AOI22_X1 U4736 ( .A1(n4042), .A2(n4220), .B1(n4326), .B2(n4053), .ZN(n4044)
         );
  NAND2_X1 U4737 ( .A1(n4247), .A2(n4321), .ZN(n4043) );
  OAI211_X1 U4738 ( .C1(n4045), .C2(n4297), .A(n4044), .B(n4043), .ZN(n4233)
         );
  AOI21_X1 U4739 ( .B1(n4046), .B2(n4502), .A(n4233), .ZN(n4056) );
  NOR2_X1 U4740 ( .A1(n4047), .A2(n4248), .ZN(n4049) );
  OAI22_X1 U4741 ( .A1(n4050), .A2(n4049), .B1(n4241), .B2(n4048), .ZN(n4061)
         );
  AOI22_X1 U4742 ( .A1(n4061), .A2(n4057), .B1(n4237), .B2(n4247), .ZN(n4052)
         );
  XNOR2_X1 U4743 ( .A(n4052), .B(n4051), .ZN(n4232) );
  NAND2_X1 U4744 ( .A1(n4232), .A2(n4192), .ZN(n4055) );
  AOI21_X1 U4745 ( .B1(n4053), .B2(n4064), .A(n4226), .ZN(n4234) );
  AOI22_X1 U4746 ( .A1(n4234), .A2(n4399), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4396), .ZN(n4054) );
  OAI211_X1 U4747 ( .C1(n4396), .C2(n4056), .A(n4055), .B(n4054), .ZN(U3354)
         );
  XNOR2_X1 U4748 ( .A(n4058), .B(n4057), .ZN(n4059) );
  NAND2_X1 U4749 ( .A1(n4059), .A2(n4495), .ZN(n4240) );
  XNOR2_X1 U4750 ( .A(n4061), .B(n4060), .ZN(n4243) );
  NAND2_X1 U4751 ( .A1(n4243), .A2(n4192), .ZN(n4073) );
  NAND2_X1 U4752 ( .A1(n4062), .A2(n4237), .ZN(n4063) );
  AOI22_X1 U4753 ( .A1(n4065), .A2(n4502), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4396), .ZN(n4066) );
  OAI21_X1 U4754 ( .B1(n4578), .B2(n4207), .A(n4066), .ZN(n4071) );
  OAI22_X1 U4755 ( .A1(n4241), .A2(n4069), .B1(n4068), .B2(n4067), .ZN(n4070)
         );
  AOI211_X1 U4756 ( .C1(n4347), .C2(n4399), .A(n4071), .B(n4070), .ZN(n4072)
         );
  OAI211_X1 U4757 ( .C1(n4396), .C2(n4240), .A(n4073), .B(n4072), .ZN(U3262)
         );
  OAI22_X1 U4758 ( .A1(n4241), .A2(n4497), .B1(n4315), .B2(n4088), .ZN(n4079)
         );
  NAND2_X1 U4759 ( .A1(n4075), .A2(n4074), .ZN(n4076) );
  XNOR2_X1 U4760 ( .A(n4076), .B(n4085), .ZN(n4077) );
  NOR2_X1 U4761 ( .A1(n4077), .A2(n4297), .ZN(n4078) );
  AOI211_X1 U4762 ( .C1(n4321), .C2(n4080), .A(n4079), .B(n4078), .ZN(n4257)
         );
  OR2_X1 U4763 ( .A1(n4095), .A2(n4081), .ZN(n4083) );
  NAND2_X1 U4764 ( .A1(n4083), .A2(n4082), .ZN(n4084) );
  XOR2_X1 U4765 ( .A(n4085), .B(n4084), .Z(n4259) );
  NAND2_X1 U4766 ( .A1(n4259), .A2(n4192), .ZN(n4094) );
  INV_X1 U4767 ( .A(n4086), .ZN(n4087) );
  OAI21_X1 U4768 ( .B1(n4103), .B2(n4088), .A(n4087), .ZN(n4354) );
  INV_X1 U4769 ( .A(n4354), .ZN(n4092) );
  OAI22_X1 U4770 ( .A1(n4090), .A2(n4162), .B1(n4089), .B2(n4505), .ZN(n4091)
         );
  AOI21_X1 U4771 ( .B1(n4092), .B2(n4399), .A(n4091), .ZN(n4093) );
  OAI211_X1 U4772 ( .C1(n4396), .C2(n4257), .A(n4094), .B(n4093), .ZN(U3264)
         );
  XNOR2_X1 U4773 ( .A(n4095), .B(n4099), .ZN(n4263) );
  INV_X1 U4774 ( .A(n4263), .ZN(n4110) );
  NAND2_X1 U4775 ( .A1(n4097), .A2(n4096), .ZN(n4098) );
  XOR2_X1 U4776 ( .A(n4099), .B(n4098), .Z(n4102) );
  OAI22_X1 U4777 ( .A1(n4142), .A2(n4330), .B1(n4105), .B2(n4315), .ZN(n4100)
         );
  AOI21_X1 U4778 ( .B1(n4327), .B2(n4249), .A(n4100), .ZN(n4101) );
  OAI21_X1 U4779 ( .B1(n4102), .B2(n4297), .A(n4101), .ZN(n4262) );
  INV_X1 U4780 ( .A(n4103), .ZN(n4104) );
  OAI21_X1 U4781 ( .B1(n4118), .B2(n4105), .A(n4104), .ZN(n4358) );
  AOI22_X1 U4782 ( .A1(n4106), .A2(n4502), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4396), .ZN(n4107) );
  OAI21_X1 U4783 ( .B1(n4358), .B2(n4174), .A(n4107), .ZN(n4108) );
  AOI21_X1 U4784 ( .B1(n4262), .B2(n4505), .A(n4108), .ZN(n4109) );
  OAI21_X1 U4785 ( .B1(n4110), .B2(n4182), .A(n4109), .ZN(U3265) );
  NAND2_X1 U4786 ( .A1(n4112), .A2(n4111), .ZN(n4114) );
  INV_X1 U4787 ( .A(n4117), .ZN(n4113) );
  XNOR2_X1 U4788 ( .A(n4114), .B(n4113), .ZN(n4115) );
  NAND2_X1 U4789 ( .A1(n4115), .A2(n4495), .ZN(n4268) );
  XOR2_X1 U4790 ( .A(n4117), .B(n4116), .Z(n4271) );
  NAND2_X1 U4791 ( .A1(n4271), .A2(n4192), .ZN(n4128) );
  INV_X1 U4792 ( .A(n4143), .ZN(n4121) );
  INV_X1 U4793 ( .A(n4118), .ZN(n4119) );
  OAI21_X1 U4794 ( .B1(n4121), .B2(n4120), .A(n4119), .ZN(n4361) );
  INV_X1 U4795 ( .A(n4361), .ZN(n4126) );
  AOI22_X1 U4796 ( .A1(n4122), .A2(n4502), .B1(REG2_REG_24__SCAN_IN), .B2(
        n4396), .ZN(n4124) );
  AOI22_X1 U4797 ( .A1(n4210), .A2(n4266), .B1(n4211), .B2(n4265), .ZN(n4123)
         );
  OAI211_X1 U4798 ( .C1(n4269), .C2(n4207), .A(n4124), .B(n4123), .ZN(n4125)
         );
  AOI21_X1 U4799 ( .B1(n4126), .B2(n4399), .A(n4125), .ZN(n4127) );
  OAI211_X1 U4800 ( .C1(n4396), .C2(n4268), .A(n4128), .B(n4127), .ZN(U3266)
         );
  XNOR2_X1 U4801 ( .A(n2153), .B(n4135), .ZN(n4275) );
  INV_X1 U4802 ( .A(n4275), .ZN(n4150) );
  OR2_X1 U4803 ( .A1(n4185), .A2(n4129), .ZN(n4131) );
  OAI21_X1 U4804 ( .B1(n4171), .B2(n4170), .A(n4133), .ZN(n4155) );
  AOI21_X1 U4805 ( .B1(n4155), .B2(n4154), .A(n4134), .ZN(n4136) );
  XNOR2_X1 U4806 ( .A(n4136), .B(n4135), .ZN(n4137) );
  NAND2_X1 U4807 ( .A1(n4137), .A2(n4495), .ZN(n4141) );
  AOI22_X1 U4808 ( .A1(n4139), .A2(n4321), .B1(n4326), .B2(n4138), .ZN(n4140)
         );
  OAI211_X1 U4809 ( .C1(n4142), .C2(n4497), .A(n4141), .B(n4140), .ZN(n4274)
         );
  INV_X1 U4810 ( .A(n4279), .ZN(n4145) );
  OAI21_X1 U4811 ( .B1(n4145), .B2(n4144), .A(n4143), .ZN(n4365) );
  AOI22_X1 U4812 ( .A1(n4396), .A2(REG2_REG_23__SCAN_IN), .B1(n4146), .B2(
        n4502), .ZN(n4147) );
  OAI21_X1 U4813 ( .B1(n4365), .B2(n4174), .A(n4147), .ZN(n4148) );
  AOI21_X1 U4814 ( .B1(n4274), .B2(n4505), .A(n4148), .ZN(n4149) );
  OAI21_X1 U4815 ( .B1(n4150), .B2(n4182), .A(n4149), .ZN(U3267) );
  AOI21_X1 U4816 ( .B1(n4154), .B2(n4152), .A(n4151), .ZN(n4153) );
  INV_X1 U4817 ( .A(n4153), .ZN(n4282) );
  XNOR2_X1 U4818 ( .A(n4155), .B(n4154), .ZN(n4160) );
  AOI22_X1 U4819 ( .A1(n4156), .A2(n4321), .B1(n4161), .B2(n4326), .ZN(n4157)
         );
  OAI21_X1 U4820 ( .B1(n4158), .B2(n4497), .A(n4157), .ZN(n4159) );
  AOI21_X1 U4821 ( .B1(n4160), .B2(n4495), .A(n4159), .ZN(n4281) );
  INV_X1 U4822 ( .A(n4281), .ZN(n4167) );
  NAND2_X1 U4823 ( .A1(n4173), .A2(n4161), .ZN(n4278) );
  AND3_X1 U4824 ( .A1(n4279), .A2(n4399), .A3(n4278), .ZN(n4166) );
  INV_X1 U4825 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4164) );
  OAI22_X1 U4826 ( .A1(n4505), .A2(n4164), .B1(n4163), .B2(n4162), .ZN(n4165)
         );
  AOI211_X1 U4827 ( .C1(n4167), .C2(n4505), .A(n4166), .B(n4165), .ZN(n4168)
         );
  OAI21_X1 U4828 ( .B1(n4282), .B2(n4182), .A(n4168), .ZN(U3268) );
  XNOR2_X1 U4829 ( .A(n4169), .B(n4170), .ZN(n4291) );
  XNOR2_X1 U4830 ( .A(n4171), .B(n4170), .ZN(n4172) );
  NAND2_X1 U4831 ( .A1(n4172), .A2(n4495), .ZN(n4289) );
  INV_X1 U4832 ( .A(n4289), .ZN(n4180) );
  OAI21_X1 U4833 ( .B1(n4193), .B2(n4283), .A(n4173), .ZN(n4285) );
  NOR2_X1 U4834 ( .A1(n4285), .A2(n4174), .ZN(n4179) );
  AOI22_X1 U4835 ( .A1(n2187), .A2(n4211), .B1(n4210), .B2(n4288), .ZN(n4177)
         );
  AOI22_X1 U4836 ( .A1(n4396), .A2(REG2_REG_21__SCAN_IN), .B1(n4175), .B2(
        n4502), .ZN(n4176) );
  OAI211_X1 U4837 ( .C1(n4284), .C2(n4207), .A(n4177), .B(n4176), .ZN(n4178)
         );
  AOI211_X1 U4838 ( .C1(n4180), .C2(n4505), .A(n4179), .B(n4178), .ZN(n4181)
         );
  OAI21_X1 U4839 ( .B1(n4291), .B2(n4182), .A(n4181), .ZN(U3269) );
  NOR3_X1 U4840 ( .A1(n4185), .A2(n4184), .A3(n4183), .ZN(n4187) );
  NOR2_X1 U4841 ( .A1(n4187), .A2(n4186), .ZN(n4189) );
  XNOR2_X1 U4842 ( .A(n4189), .B(n4188), .ZN(n4298) );
  XNOR2_X1 U4843 ( .A(n4190), .B(n4191), .ZN(n4300) );
  NAND2_X1 U4844 ( .A1(n4300), .A2(n4192), .ZN(n4203) );
  INV_X1 U4845 ( .A(n4193), .ZN(n4194) );
  OAI21_X1 U4846 ( .B1(n4195), .B2(n4292), .A(n4194), .ZN(n4370) );
  INV_X1 U4847 ( .A(n4370), .ZN(n4201) );
  AOI22_X1 U4848 ( .A1(n4196), .A2(n4211), .B1(n4210), .B2(n4295), .ZN(n4199)
         );
  AOI22_X1 U4849 ( .A1(n4396), .A2(REG2_REG_20__SCAN_IN), .B1(n4197), .B2(
        n4502), .ZN(n4198) );
  OAI211_X1 U4850 ( .C1(n4293), .C2(n4207), .A(n4199), .B(n4198), .ZN(n4200)
         );
  AOI21_X1 U4851 ( .B1(n4201), .B2(n4399), .A(n4200), .ZN(n4202) );
  OAI211_X1 U4852 ( .C1(n4298), .C2(n4204), .A(n4203), .B(n4202), .ZN(U3270)
         );
  MUX2_X1 U4853 ( .A(n4206), .B(n4205), .S(n4505), .Z(n4218) );
  INV_X1 U4854 ( .A(n4207), .ZN(n4209) );
  AOI22_X1 U4855 ( .A1(n4209), .A2(n4208), .B1(REG3_REG_2__SCAN_IN), .B2(n4502), .ZN(n4217) );
  AOI22_X1 U4856 ( .A1(n4212), .A2(n4211), .B1(n4210), .B2(n2762), .ZN(n4216)
         );
  AOI22_X1 U4857 ( .A1(n4214), .A2(n4503), .B1(n4399), .B2(n4213), .ZN(n4215)
         );
  NAND4_X1 U4858 ( .A1(n4218), .A2(n4217), .A3(n4216), .A4(n4215), .ZN(U3288)
         );
  NAND2_X1 U4859 ( .A1(n4226), .A2(n4229), .ZN(n4225) );
  XNOR2_X1 U4860 ( .A(n4225), .B(n4219), .ZN(n4393) );
  INV_X1 U4861 ( .A(n4393), .ZN(n4339) );
  INV_X1 U4862 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4223) );
  AND2_X1 U4863 ( .A1(n4221), .A2(n4220), .ZN(n4227) );
  AOI21_X1 U4864 ( .B1(n4222), .B2(n4326), .A(n4227), .ZN(n4395) );
  MUX2_X1 U4865 ( .A(n4223), .B(n4395), .S(n4577), .Z(n4224) );
  OAI21_X1 U4866 ( .B1(n4339), .B2(n4313), .A(n4224), .ZN(U3549) );
  INV_X1 U4867 ( .A(n4227), .ZN(n4228) );
  OAI21_X1 U4868 ( .B1(n4229), .B2(n4315), .A(n4228), .ZN(n4398) );
  INV_X1 U4869 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4779) );
  NOR2_X1 U4870 ( .A1(n4577), .A2(n4779), .ZN(n4230) );
  AOI21_X1 U4871 ( .B1(n4577), .B2(n4398), .A(n4230), .ZN(n4231) );
  OAI21_X1 U4872 ( .B1(n4397), .B2(n4313), .A(n4231), .ZN(U3548) );
  NAND2_X1 U4873 ( .A1(n4232), .A2(n4549), .ZN(n4236) );
  NAND2_X1 U4874 ( .A1(n4236), .A2(n4235), .ZN(n4343) );
  MUX2_X1 U4875 ( .A(REG1_REG_29__SCAN_IN), .B(n4343), .S(n4577), .Z(U3547) );
  INV_X1 U4876 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4772) );
  AOI22_X1 U4877 ( .A1(n4238), .A2(n4327), .B1(n4237), .B2(n4326), .ZN(n4239)
         );
  OAI211_X1 U4878 ( .C1(n4241), .C2(n4330), .A(n4240), .B(n4239), .ZN(n4242)
         );
  AOI21_X1 U4879 ( .B1(n4243), .B2(n4549), .A(n4242), .ZN(n4344) );
  NAND2_X1 U4880 ( .A1(n4347), .A2(n4244), .ZN(n4245) );
  NAND2_X1 U4881 ( .A1(n4246), .A2(n4245), .ZN(U3546) );
  NAND2_X1 U4882 ( .A1(n4247), .A2(n4327), .ZN(n4251) );
  AOI22_X1 U4883 ( .A1(n4249), .A2(n4321), .B1(n4248), .B2(n4326), .ZN(n4250)
         );
  NAND2_X1 U4884 ( .A1(n4251), .A2(n4250), .ZN(n4252) );
  AOI21_X1 U4885 ( .B1(n4253), .B2(n4562), .A(n4252), .ZN(n4255) );
  OAI211_X1 U4886 ( .C1(n4256), .C2(n4543), .A(n4255), .B(n4254), .ZN(n4350)
         );
  MUX2_X1 U4887 ( .A(REG1_REG_27__SCAN_IN), .B(n4350), .S(n4577), .Z(U3545) );
  INV_X1 U4888 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4260) );
  INV_X1 U4889 ( .A(n4257), .ZN(n4258) );
  AOI21_X1 U4890 ( .B1(n4259), .B2(n4549), .A(n4258), .ZN(n4351) );
  MUX2_X1 U4891 ( .A(n4260), .B(n4351), .S(n4577), .Z(n4261) );
  OAI21_X1 U4892 ( .B1(n4313), .B2(n4354), .A(n4261), .ZN(U3544) );
  INV_X1 U4893 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4773) );
  AOI21_X1 U4894 ( .B1(n4263), .B2(n4549), .A(n4262), .ZN(n4355) );
  MUX2_X1 U4895 ( .A(n4773), .B(n4355), .S(n4577), .Z(n4264) );
  OAI21_X1 U4896 ( .B1(n4313), .B2(n4358), .A(n4264), .ZN(U3543) );
  INV_X1 U4897 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4272) );
  AOI22_X1 U4898 ( .A1(n4266), .A2(n4321), .B1(n4326), .B2(n4265), .ZN(n4267)
         );
  OAI211_X1 U4899 ( .C1(n4269), .C2(n4497), .A(n4268), .B(n4267), .ZN(n4270)
         );
  AOI21_X1 U4900 ( .B1(n4271), .B2(n4549), .A(n4270), .ZN(n4359) );
  MUX2_X1 U4901 ( .A(n4272), .B(n4359), .S(n4577), .Z(n4273) );
  OAI21_X1 U4902 ( .B1(n4313), .B2(n4361), .A(n4273), .ZN(U3542) );
  INV_X1 U4903 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4276) );
  AOI21_X1 U4904 ( .B1(n4275), .B2(n4549), .A(n4274), .ZN(n4362) );
  MUX2_X1 U4905 ( .A(n4276), .B(n4362), .S(n4577), .Z(n4277) );
  OAI21_X1 U4906 ( .B1(n4313), .B2(n4365), .A(n4277), .ZN(U3541) );
  NAND3_X1 U4907 ( .A1(n4279), .A2(n4562), .A3(n4278), .ZN(n4280) );
  OAI211_X1 U4908 ( .C1(n4282), .C2(n4543), .A(n4281), .B(n4280), .ZN(n4366)
         );
  MUX2_X1 U4909 ( .A(REG1_REG_22__SCAN_IN), .B(n4366), .S(n4577), .Z(U3540) );
  OAI22_X1 U4910 ( .A1(n4284), .A2(n4497), .B1(n4315), .B2(n4283), .ZN(n4287)
         );
  NOR2_X1 U4911 ( .A1(n4285), .A2(n4551), .ZN(n4286) );
  AOI211_X1 U4912 ( .C1(n4321), .C2(n4288), .A(n4287), .B(n4286), .ZN(n4290)
         );
  OAI211_X1 U4913 ( .C1(n4291), .C2(n4543), .A(n4290), .B(n4289), .ZN(n4367)
         );
  MUX2_X1 U4914 ( .A(REG1_REG_21__SCAN_IN), .B(n4367), .S(n4577), .Z(U3539) );
  INV_X1 U4915 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4301) );
  OAI22_X1 U4916 ( .A1(n4293), .A2(n4497), .B1(n4315), .B2(n4292), .ZN(n4294)
         );
  AOI21_X1 U4917 ( .B1(n4321), .B2(n4295), .A(n4294), .ZN(n4296) );
  OAI21_X1 U4918 ( .B1(n4298), .B2(n4297), .A(n4296), .ZN(n4299) );
  AOI21_X1 U4919 ( .B1(n4300), .B2(n4549), .A(n4299), .ZN(n4368) );
  MUX2_X1 U4920 ( .A(n4301), .B(n4368), .S(n4577), .Z(n4302) );
  OAI21_X1 U4921 ( .B1(n4313), .B2(n4370), .A(n4302), .ZN(U3538) );
  INV_X1 U4922 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4770) );
  AOI21_X1 U4923 ( .B1(n4304), .B2(n4549), .A(n4303), .ZN(n4371) );
  MUX2_X1 U4924 ( .A(n4770), .B(n4371), .S(n4577), .Z(n4305) );
  OAI21_X1 U4925 ( .B1(n4313), .B2(n4373), .A(n4305), .ZN(U3537) );
  INV_X1 U4926 ( .A(n4306), .ZN(n4309) );
  OAI211_X1 U4927 ( .C1(n4309), .C2(n4543), .A(n4308), .B(n4307), .ZN(n4374)
         );
  MUX2_X1 U4928 ( .A(REG1_REG_18__SCAN_IN), .B(n4374), .S(n4577), .Z(U3536) );
  INV_X1 U4929 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4767) );
  AOI21_X1 U4930 ( .B1(n4311), .B2(n4549), .A(n4310), .ZN(n4375) );
  MUX2_X1 U4931 ( .A(n4767), .B(n4375), .S(n4577), .Z(n4312) );
  OAI21_X1 U4932 ( .B1(n4313), .B2(n4379), .A(n4312), .ZN(U3535) );
  OAI22_X1 U4933 ( .A1(n4316), .A2(n4497), .B1(n4315), .B2(n4314), .ZN(n4319)
         );
  NOR2_X1 U4934 ( .A1(n4317), .A2(n4551), .ZN(n4318) );
  AOI211_X1 U4935 ( .C1(n4321), .C2(n4320), .A(n4319), .B(n4318), .ZN(n4323)
         );
  OAI211_X1 U4936 ( .C1(n4324), .C2(n4543), .A(n4323), .B(n4322), .ZN(n4380)
         );
  MUX2_X1 U4937 ( .A(REG1_REG_16__SCAN_IN), .B(n4380), .S(n4577), .Z(U3534) );
  AOI22_X1 U4938 ( .A1(n4328), .A2(n4327), .B1(n4326), .B2(n4325), .ZN(n4329)
         );
  OAI21_X1 U4939 ( .B1(n4331), .B2(n4330), .A(n4329), .ZN(n4332) );
  AOI21_X1 U4940 ( .B1(n4333), .B2(n4562), .A(n4332), .ZN(n4335) );
  OAI211_X1 U4941 ( .C1(n4336), .C2(n4543), .A(n4335), .B(n4334), .ZN(n4381)
         );
  MUX2_X1 U4942 ( .A(REG1_REG_15__SCAN_IN), .B(n4381), .S(n4577), .Z(U3533) );
  INV_X1 U4943 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4337) );
  MUX2_X1 U4944 ( .A(n4337), .B(n4395), .S(n4565), .Z(n4338) );
  OAI21_X1 U4945 ( .B1(n4339), .B2(n4378), .A(n4338), .ZN(U3517) );
  INV_X1 U4946 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4340) );
  NOR2_X1 U4947 ( .A1(n4565), .A2(n4340), .ZN(n4341) );
  AOI21_X1 U4948 ( .B1(n4565), .B2(n4398), .A(n4341), .ZN(n4342) );
  OAI21_X1 U4949 ( .B1(n4397), .B2(n4378), .A(n4342), .ZN(U3516) );
  MUX2_X1 U4950 ( .A(REG0_REG_29__SCAN_IN), .B(n4343), .S(n4565), .Z(U3515) );
  INV_X1 U4951 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4345) );
  NAND2_X1 U4952 ( .A1(n4347), .A2(n4346), .ZN(n4348) );
  NAND2_X1 U4953 ( .A1(n4349), .A2(n4348), .ZN(U3514) );
  MUX2_X1 U4954 ( .A(REG0_REG_27__SCAN_IN), .B(n4350), .S(n4565), .Z(U3513) );
  INV_X1 U4955 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4352) );
  MUX2_X1 U4956 ( .A(n4352), .B(n4351), .S(n4565), .Z(n4353) );
  OAI21_X1 U4957 ( .B1(n4354), .B2(n4378), .A(n4353), .ZN(U3512) );
  INV_X1 U4958 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4356) );
  MUX2_X1 U4959 ( .A(n4356), .B(n4355), .S(n4565), .Z(n4357) );
  OAI21_X1 U4960 ( .B1(n4358), .B2(n4378), .A(n4357), .ZN(U3511) );
  INV_X1 U4961 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4752) );
  MUX2_X1 U4962 ( .A(n4752), .B(n4359), .S(n4565), .Z(n4360) );
  OAI21_X1 U4963 ( .B1(n4361), .B2(n4378), .A(n4360), .ZN(U3510) );
  INV_X1 U4964 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4363) );
  MUX2_X1 U4965 ( .A(n4363), .B(n4362), .S(n4565), .Z(n4364) );
  OAI21_X1 U4966 ( .B1(n4365), .B2(n4378), .A(n4364), .ZN(U3509) );
  MUX2_X1 U4967 ( .A(REG0_REG_22__SCAN_IN), .B(n4366), .S(n4565), .Z(U3508) );
  MUX2_X1 U4968 ( .A(REG0_REG_21__SCAN_IN), .B(n4367), .S(n4565), .Z(U3507) );
  INV_X1 U4969 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4749) );
  MUX2_X1 U4970 ( .A(n4749), .B(n4368), .S(n4565), .Z(n4369) );
  OAI21_X1 U4971 ( .B1(n4370), .B2(n4378), .A(n4369), .ZN(U3506) );
  INV_X1 U4972 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4750) );
  MUX2_X1 U4973 ( .A(n4750), .B(n4371), .S(n4565), .Z(n4372) );
  OAI21_X1 U4974 ( .B1(n4373), .B2(n4378), .A(n4372), .ZN(U3505) );
  MUX2_X1 U4975 ( .A(REG0_REG_18__SCAN_IN), .B(n4374), .S(n4565), .Z(U3503) );
  INV_X1 U4976 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4376) );
  MUX2_X1 U4977 ( .A(n4376), .B(n4375), .S(n4565), .Z(n4377) );
  OAI21_X1 U4978 ( .B1(n4379), .B2(n4378), .A(n4377), .ZN(U3501) );
  MUX2_X1 U4979 ( .A(REG0_REG_16__SCAN_IN), .B(n4380), .S(n4565), .Z(U3499) );
  MUX2_X1 U4980 ( .A(REG0_REG_15__SCAN_IN), .B(n4381), .S(n4565), .Z(U3497) );
  MUX2_X1 U4981 ( .A(n4382), .B(DATAI_28_), .S(U3149), .Z(U3324) );
  MUX2_X1 U4982 ( .A(n4383), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U4983 ( .A(n4384), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4984 ( .A(n4385), .B(DATAI_17_), .S(U3149), .Z(U3335) );
  MUX2_X1 U4985 ( .A(n4386), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U4986 ( .A(DATAI_8_), .B(n4387), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U4987 ( .A(n4388), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U4988 ( .A(n4389), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U4989 ( .A(n4390), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4990 ( .A(n2136), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4991 ( .A(n4392), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI22_X1 U4992 ( .A1(n4393), .A2(n4399), .B1(n4396), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n4394) );
  OAI21_X1 U4993 ( .B1(n4396), .B2(n4395), .A(n4394), .ZN(U3260) );
  INV_X1 U4994 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4809) );
  INV_X1 U4995 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4400) );
  XNOR2_X1 U4996 ( .A(n4401), .B(n4400), .ZN(n4402) );
  NAND2_X1 U4997 ( .A1(n4474), .A2(n4402), .ZN(n4412) );
  INV_X1 U4998 ( .A(REG2_REG_4__SCAN_IN), .ZN(n4403) );
  XNOR2_X1 U4999 ( .A(n4404), .B(n4403), .ZN(n4405) );
  NAND2_X1 U5000 ( .A1(n4488), .A2(n4405), .ZN(n4411) );
  NAND2_X1 U5001 ( .A1(n4450), .A2(n4406), .ZN(n4410) );
  INV_X1 U5002 ( .A(n4407), .ZN(n4408) );
  AOI21_X1 U5003 ( .B1(n4483), .B2(ADDR_REG_4__SCAN_IN), .A(n4408), .ZN(n4409)
         );
  AND4_X1 U5004 ( .A1(n4412), .A2(n4411), .A3(n4410), .A4(n4409), .ZN(n4414)
         );
  NAND2_X1 U5005 ( .A1(n4414), .A2(n4413), .ZN(U3244) );
  AOI211_X1 U5006 ( .C1(n4764), .C2(n4416), .A(n4415), .B(n4478), .ZN(n4418)
         );
  AOI211_X1 U5007 ( .C1(n4483), .C2(ADDR_REG_10__SCAN_IN), .A(n4418), .B(n4417), .ZN(n4422) );
  OAI211_X1 U5008 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4420), .A(n4488), .B(n4419), .ZN(n4421) );
  OAI211_X1 U5009 ( .C1(n4490), .C2(n4520), .A(n4422), .B(n4421), .ZN(U3250)
         );
  AOI211_X1 U5010 ( .C1(n2167), .C2(n4424), .A(n4423), .B(n4478), .ZN(n4426)
         );
  AOI211_X1 U5011 ( .C1(n4483), .C2(ADDR_REG_11__SCAN_IN), .A(n4426), .B(n4425), .ZN(n4431) );
  OAI211_X1 U5012 ( .C1(n4429), .C2(n4428), .A(n4488), .B(n4427), .ZN(n4430)
         );
  OAI211_X1 U5013 ( .C1(n4490), .C2(n4432), .A(n4431), .B(n4430), .ZN(U3251)
         );
  AOI211_X1 U5014 ( .C1(n4435), .C2(n4434), .A(n4433), .B(n4478), .ZN(n4438)
         );
  INV_X1 U5015 ( .A(n4436), .ZN(n4437) );
  AOI211_X1 U5016 ( .C1(n4483), .C2(ADDR_REG_12__SCAN_IN), .A(n4438), .B(n4437), .ZN(n4442) );
  OAI211_X1 U5017 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4440), .A(n4488), .B(n4439), .ZN(n4441) );
  OAI211_X1 U5018 ( .C1(n4490), .C2(n4517), .A(n4442), .B(n4441), .ZN(U3252)
         );
  INV_X1 U5019 ( .A(ADDR_REG_14__SCAN_IN), .ZN(n4814) );
  AOI211_X1 U5020 ( .C1(n4766), .C2(n4444), .A(n4443), .B(n4478), .ZN(n4449)
         );
  AOI211_X1 U5021 ( .C1(n4794), .C2(n4447), .A(n4446), .B(n4445), .ZN(n4448)
         );
  AOI211_X1 U5022 ( .C1(n4450), .C2(n4514), .A(n4449), .B(n4448), .ZN(n4452)
         );
  OAI211_X1 U5023 ( .C1(n4465), .C2(n4814), .A(n4452), .B(n4451), .ZN(U3254)
         );
  AOI211_X1 U5024 ( .C1(n4455), .C2(n4454), .A(n4453), .B(n4478), .ZN(n4456)
         );
  AOI211_X1 U5025 ( .C1(n4483), .C2(ADDR_REG_15__SCAN_IN), .A(n4457), .B(n4456), .ZN(n4463) );
  AOI21_X1 U5026 ( .B1(n4460), .B2(n4459), .A(n4458), .ZN(n4461) );
  NAND2_X1 U5027 ( .A1(n4488), .A2(n4461), .ZN(n4462) );
  OAI211_X1 U5028 ( .C1(n4490), .C2(n4513), .A(n4463), .B(n4462), .ZN(U3255)
         );
  INV_X1 U5029 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n4811) );
  OAI21_X1 U5030 ( .B1(n4465), .B2(n4811), .A(n4464), .ZN(n4466) );
  INV_X1 U5031 ( .A(n4466), .ZN(n4477) );
  OAI21_X1 U5032 ( .B1(n4469), .B2(n4468), .A(n4467), .ZN(n4475) );
  OAI21_X1 U5033 ( .B1(n4472), .B2(n4471), .A(n4470), .ZN(n4473) );
  AOI22_X1 U5034 ( .A1(n4488), .A2(n4475), .B1(n4474), .B2(n4473), .ZN(n4476)
         );
  OAI211_X1 U5035 ( .C1(n4512), .C2(n4490), .A(n4477), .B(n4476), .ZN(U3256)
         );
  AOI21_X1 U5036 ( .B1(n4486), .B2(n4485), .A(n4484), .ZN(n4487) );
  NAND2_X1 U5037 ( .A1(n4488), .A2(n4487), .ZN(n4489) );
  INV_X1 U5038 ( .A(n4491), .ZN(n4492) );
  NOR2_X1 U5039 ( .A1(n4493), .A2(n4492), .ZN(n4523) );
  INV_X1 U5040 ( .A(n4494), .ZN(n4500) );
  NOR2_X1 U5041 ( .A1(n4496), .A2(n4495), .ZN(n4499) );
  OAI22_X1 U5042 ( .A1(n4501), .A2(n4499), .B1(n4498), .B2(n4497), .ZN(n4522)
         );
  AOI21_X1 U5043 ( .B1(n4523), .B2(n4500), .A(n4522), .ZN(n4506) );
  INV_X1 U5044 ( .A(n4501), .ZN(n4524) );
  AOI22_X1 U5045 ( .A1(n4524), .A2(n4503), .B1(REG3_REG_0__SCAN_IN), .B2(n4502), .ZN(n4504) );
  OAI221_X1 U5046 ( .B1(n4396), .B2(n4506), .C1(n4505), .C2(n4780), .A(n4504), 
        .ZN(U3290) );
  INV_X1 U5047 ( .A(D_REG_31__SCAN_IN), .ZN(n4733) );
  NOR2_X1 U5048 ( .A1(n4508), .A2(n4733), .ZN(U3291) );
  INV_X1 U5049 ( .A(D_REG_30__SCAN_IN), .ZN(n4732) );
  NOR2_X1 U5050 ( .A1(n4508), .A2(n4732), .ZN(U3292) );
  INV_X1 U5051 ( .A(D_REG_29__SCAN_IN), .ZN(n4730) );
  NOR2_X1 U5052 ( .A1(n4508), .A2(n4730), .ZN(U3293) );
  INV_X1 U5053 ( .A(D_REG_28__SCAN_IN), .ZN(n4729) );
  NOR2_X1 U5054 ( .A1(n4508), .A2(n4729), .ZN(U3294) );
  NOR2_X1 U5055 ( .A1(n4508), .A2(n4722), .ZN(U3295) );
  AND2_X1 U5056 ( .A1(D_REG_26__SCAN_IN), .A2(n4507), .ZN(U3296) );
  INV_X1 U5057 ( .A(D_REG_25__SCAN_IN), .ZN(n4723) );
  NOR2_X1 U5058 ( .A1(n4508), .A2(n4723), .ZN(U3297) );
  INV_X1 U5059 ( .A(D_REG_24__SCAN_IN), .ZN(n4720) );
  NOR2_X1 U5060 ( .A1(n4508), .A2(n4720), .ZN(U3298) );
  AND2_X1 U5061 ( .A1(D_REG_23__SCAN_IN), .A2(n4507), .ZN(U3299) );
  NOR2_X1 U5062 ( .A1(n4508), .A2(n4719), .ZN(U3300) );
  INV_X1 U5063 ( .A(D_REG_21__SCAN_IN), .ZN(n4716) );
  NOR2_X1 U5064 ( .A1(n4508), .A2(n4716), .ZN(U3301) );
  AND2_X1 U5065 ( .A1(D_REG_20__SCAN_IN), .A2(n4507), .ZN(U3302) );
  AND2_X1 U5066 ( .A1(D_REG_19__SCAN_IN), .A2(n4507), .ZN(U3303) );
  NOR2_X1 U5067 ( .A1(n4508), .A2(n4717), .ZN(U3304) );
  AND2_X1 U5068 ( .A1(D_REG_17__SCAN_IN), .A2(n4507), .ZN(U3305) );
  AND2_X1 U5069 ( .A1(D_REG_16__SCAN_IN), .A2(n4507), .ZN(U3306) );
  AND2_X1 U5070 ( .A1(D_REG_15__SCAN_IN), .A2(n4507), .ZN(U3307) );
  INV_X1 U5071 ( .A(D_REG_14__SCAN_IN), .ZN(n4713) );
  NOR2_X1 U5072 ( .A1(n4508), .A2(n4713), .ZN(U3308) );
  AND2_X1 U5073 ( .A1(D_REG_13__SCAN_IN), .A2(n4507), .ZN(U3309) );
  AND2_X1 U5074 ( .A1(D_REG_12__SCAN_IN), .A2(n4507), .ZN(U3310) );
  INV_X1 U5075 ( .A(D_REG_11__SCAN_IN), .ZN(n4714) );
  NOR2_X1 U5076 ( .A1(n4508), .A2(n4714), .ZN(U3311) );
  INV_X1 U5077 ( .A(D_REG_10__SCAN_IN), .ZN(n4699) );
  NOR2_X1 U5078 ( .A1(n4508), .A2(n4699), .ZN(U3312) );
  AND2_X1 U5079 ( .A1(D_REG_9__SCAN_IN), .A2(n4507), .ZN(U3313) );
  AND2_X1 U5080 ( .A1(D_REG_8__SCAN_IN), .A2(n4507), .ZN(U3314) );
  INV_X1 U5081 ( .A(D_REG_7__SCAN_IN), .ZN(n4698) );
  NOR2_X1 U5082 ( .A1(n4508), .A2(n4698), .ZN(U3315) );
  INV_X1 U5083 ( .A(D_REG_6__SCAN_IN), .ZN(n4704) );
  NOR2_X1 U5084 ( .A1(n4508), .A2(n4704), .ZN(U3316) );
  AND2_X1 U5085 ( .A1(D_REG_5__SCAN_IN), .A2(n4507), .ZN(U3317) );
  INV_X1 U5086 ( .A(D_REG_4__SCAN_IN), .ZN(n4705) );
  NOR2_X1 U5087 ( .A1(n4508), .A2(n4705), .ZN(U3318) );
  NOR2_X1 U5088 ( .A1(n4508), .A2(n4702), .ZN(U3319) );
  INV_X1 U5089 ( .A(D_REG_2__SCAN_IN), .ZN(n4701) );
  NOR2_X1 U5090 ( .A1(n4508), .A2(n4701), .ZN(U3320) );
  OAI21_X1 U5091 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4509), .ZN(
        n4510) );
  INV_X1 U5092 ( .A(n4510), .ZN(U3329) );
  INV_X1 U5093 ( .A(DATAI_18_), .ZN(n4636) );
  AOI22_X1 U5094 ( .A1(STATE_REG_SCAN_IN), .A2(n4511), .B1(n4636), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U5095 ( .A(DATAI_16_), .ZN(n4638) );
  AOI22_X1 U5096 ( .A1(STATE_REG_SCAN_IN), .A2(n4512), .B1(n4638), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5097 ( .A(DATAI_15_), .ZN(n4639) );
  AOI22_X1 U5098 ( .A1(STATE_REG_SCAN_IN), .A2(n4513), .B1(n4639), .B2(U3149), 
        .ZN(U3337) );
  OAI22_X1 U5099 ( .A1(U3149), .A2(n4514), .B1(DATAI_14_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4515) );
  INV_X1 U5100 ( .A(n4515), .ZN(U3338) );
  INV_X1 U5101 ( .A(DATAI_12_), .ZN(n4516) );
  AOI22_X1 U5102 ( .A1(STATE_REG_SCAN_IN), .A2(n4517), .B1(n4516), .B2(U3149), 
        .ZN(U3340) );
  OAI22_X1 U5103 ( .A1(U3149), .A2(n4518), .B1(DATAI_11_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4519) );
  INV_X1 U5104 ( .A(n4519), .ZN(U3341) );
  INV_X1 U5105 ( .A(DATAI_10_), .ZN(n4647) );
  AOI22_X1 U5106 ( .A1(STATE_REG_SCAN_IN), .A2(n4520), .B1(n4647), .B2(U3149), 
        .ZN(U3342) );
  OAI22_X1 U5107 ( .A1(U3149), .A2(n4603), .B1(DATAI_0_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4521) );
  INV_X1 U5108 ( .A(n4521), .ZN(U3352) );
  AOI211_X1 U5109 ( .C1(n4536), .C2(n4524), .A(n4523), .B(n4522), .ZN(n4566)
         );
  INV_X1 U5110 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4525) );
  AOI22_X1 U5111 ( .A1(n4565), .A2(n4566), .B1(n4525), .B2(n4563), .ZN(U3467)
         );
  INV_X1 U5112 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4526) );
  AOI22_X1 U5113 ( .A1(n4565), .A2(n4527), .B1(n4526), .B2(n4563), .ZN(U3469)
         );
  NOR2_X1 U5114 ( .A1(n4528), .A2(n4557), .ZN(n4530) );
  AOI211_X1 U5115 ( .C1(n4562), .C2(n4531), .A(n4530), .B(n4529), .ZN(n4568)
         );
  INV_X1 U5116 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4532) );
  AOI22_X1 U5117 ( .A1(n4565), .A2(n4568), .B1(n4532), .B2(n4563), .ZN(U3473)
         );
  INV_X1 U5118 ( .A(n4533), .ZN(n4535) );
  AOI211_X1 U5119 ( .C1(n4537), .C2(n4536), .A(n4535), .B(n4534), .ZN(n4569)
         );
  INV_X1 U5120 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4736) );
  AOI22_X1 U5121 ( .A1(n4565), .A2(n4569), .B1(n4736), .B2(n4563), .ZN(U3475)
         );
  NOR2_X1 U5122 ( .A1(n4538), .A2(n4543), .ZN(n4541) );
  INV_X1 U5123 ( .A(n4539), .ZN(n4540) );
  AOI211_X1 U5124 ( .C1(n4562), .C2(n4542), .A(n4541), .B(n4540), .ZN(n4570)
         );
  INV_X1 U5125 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4735) );
  AOI22_X1 U5126 ( .A1(n4565), .A2(n4570), .B1(n4735), .B2(n4563), .ZN(U3477)
         );
  NOR2_X1 U5127 ( .A1(n4544), .A2(n4543), .ZN(n4547) );
  AOI211_X1 U5128 ( .C1(n4547), .C2(n3110), .A(n4546), .B(n4545), .ZN(n4572)
         );
  INV_X1 U5129 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4548) );
  AOI22_X1 U5130 ( .A1(n4565), .A2(n4572), .B1(n4548), .B2(n4563), .ZN(U3481)
         );
  NAND2_X1 U5131 ( .A1(n4550), .A2(n4549), .ZN(n4554) );
  OR2_X1 U5132 ( .A1(n4552), .A2(n4551), .ZN(n4553) );
  AND3_X1 U5133 ( .A1(n4555), .A2(n4554), .A3(n4553), .ZN(n4573) );
  INV_X1 U5134 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4556) );
  AOI22_X1 U5135 ( .A1(n4565), .A2(n4573), .B1(n4556), .B2(n4563), .ZN(U3485)
         );
  NOR2_X1 U5136 ( .A1(n4558), .A2(n4557), .ZN(n4560) );
  AOI211_X1 U5137 ( .C1(n4562), .C2(n4561), .A(n4560), .B(n4559), .ZN(n4576)
         );
  INV_X1 U5138 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4564) );
  AOI22_X1 U5139 ( .A1(n4565), .A2(n4576), .B1(n4564), .B2(n4563), .ZN(U3489)
         );
  AOI22_X1 U5140 ( .A1(n4577), .A2(n4566), .B1(n2742), .B2(n4574), .ZN(U3518)
         );
  INV_X1 U5141 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4567) );
  AOI22_X1 U5142 ( .A1(n4577), .A2(n4568), .B1(n4567), .B2(n4574), .ZN(U3521)
         );
  AOI22_X1 U5143 ( .A1(n4577), .A2(n4569), .B1(n4400), .B2(n4574), .ZN(U3522)
         );
  AOI22_X1 U5144 ( .A1(n4577), .A2(n4570), .B1(n2365), .B2(n4574), .ZN(U3523)
         );
  AOI22_X1 U5145 ( .A1(n4577), .A2(n4572), .B1(n4571), .B2(n4574), .ZN(U3525)
         );
  AOI22_X1 U5146 ( .A1(n4577), .A2(n4573), .B1(n2383), .B2(n4574), .ZN(U3527)
         );
  AOI22_X1 U5147 ( .A1(n4577), .A2(n4576), .B1(n4575), .B2(n4574), .ZN(U3529)
         );
  NAND2_X1 U5148 ( .A1(n4578), .A2(U4043), .ZN(n4579) );
  OAI21_X1 U5149 ( .B1(U4043), .B2(DATAO_REG_29__SCAN_IN), .A(n4579), .ZN(
        n4881) );
  NOR4_X1 U5150 ( .A1(REG0_REG_28__SCAN_IN), .A2(REG1_REG_28__SCAN_IN), .A3(
        REG1_REG_25__SCAN_IN), .A4(REG0_REG_24__SCAN_IN), .ZN(n4584) );
  NOR4_X1 U5151 ( .A1(REG1_REG_30__SCAN_IN), .A2(ADDR_REG_13__SCAN_IN), .A3(
        ADDR_REG_5__SCAN_IN), .A4(DATAO_REG_31__SCAN_IN), .ZN(n4583) );
  NOR4_X1 U5152 ( .A1(REG0_REG_12__SCAN_IN), .A2(REG2_REG_7__SCAN_IN), .A3(
        REG0_REG_5__SCAN_IN), .A4(REG1_REG_2__SCAN_IN), .ZN(n4582) );
  NOR4_X1 U5153 ( .A1(REG0_REG_16__SCAN_IN), .A2(DATAI_10_), .A3(DATAI_8_), 
        .A4(REG0_REG_8__SCAN_IN), .ZN(n4581) );
  NAND4_X1 U5154 ( .A1(n4584), .A2(n4583), .A3(n4582), .A4(n4581), .ZN(n4627)
         );
  NOR4_X1 U5155 ( .A1(DATAO_REG_9__SCAN_IN), .A2(DATAO_REG_11__SCAN_IN), .A3(
        DATAO_REG_3__SCAN_IN), .A4(DATAO_REG_12__SCAN_IN), .ZN(n4589) );
  NOR4_X1 U5156 ( .A1(REG3_REG_3__SCAN_IN), .A2(DATAI_9_), .A3(DATAI_3_), .A4(
        DATAO_REG_8__SCAN_IN), .ZN(n4588) );
  NOR4_X1 U5157 ( .A1(D_REG_21__SCAN_IN), .A2(DATAO_REG_24__SCAN_IN), .A3(
        DATAO_REG_19__SCAN_IN), .A4(DATAO_REG_7__SCAN_IN), .ZN(n4587) );
  INV_X1 U5158 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4585) );
  AND4_X1 U5159 ( .A1(n4585), .A2(REG3_REG_8__SCAN_IN), .A3(
        REG3_REG_10__SCAN_IN), .A4(REG3_REG_4__SCAN_IN), .ZN(n4586) );
  NAND4_X1 U5160 ( .A1(n4589), .A2(n4588), .A3(n4587), .A4(n4586), .ZN(n4626)
         );
  NOR4_X1 U5161 ( .A1(DATAI_21_), .A2(DATAI_17_), .A3(REG2_REG_6__SCAN_IN), 
        .A4(ADDR_REG_0__SCAN_IN), .ZN(n4599) );
  NOR4_X1 U5162 ( .A1(REG1_REG_17__SCAN_IN), .A2(REG2_REG_12__SCAN_IN), .A3(
        ADDR_REG_16__SCAN_IN), .A4(ADDR_REG_12__SCAN_IN), .ZN(n4598) );
  NOR4_X1 U5163 ( .A1(REG2_REG_22__SCAN_IN), .A2(REG2_REG_4__SCAN_IN), .A3(
        REG1_REG_18__SCAN_IN), .A4(n4814), .ZN(n4590) );
  NAND3_X1 U5164 ( .A1(DATAO_REG_13__SCAN_IN), .A2(DATAO_REG_2__SCAN_IN), .A3(
        n4590), .ZN(n4591) );
  NOR3_X1 U5165 ( .A1(DATAI_27_), .A2(DATAI_25_), .A3(n4591), .ZN(n4597) );
  NAND4_X1 U5166 ( .A1(DATAI_30_), .A2(DATAO_REG_0__SCAN_IN), .A3(
        DATAO_REG_26__SCAN_IN), .A4(DATAO_REG_30__SCAN_IN), .ZN(n4595) );
  NAND4_X1 U5167 ( .A1(DATAO_REG_16__SCAN_IN), .A2(DATAO_REG_17__SCAN_IN), 
        .A3(DATAO_REG_14__SCAN_IN), .A4(DATAO_REG_22__SCAN_IN), .ZN(n4594) );
  NAND4_X1 U5168 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_30__SCAN_IN), .A4(REG0_REG_20__SCAN_IN), .ZN(n4593) );
  NAND4_X1 U5169 ( .A1(D_REG_0__SCAN_IN), .A2(REG0_REG_22__SCAN_IN), .A3(
        REG0_REG_19__SCAN_IN), .A4(DATAI_16_), .ZN(n4592) );
  NOR4_X1 U5170 ( .A1(n4595), .A2(n4594), .A3(n4593), .A4(n4592), .ZN(n4596)
         );
  NAND4_X1 U5171 ( .A1(n4599), .A2(n4598), .A3(n4597), .A4(n4596), .ZN(n4625)
         );
  NAND4_X1 U5172 ( .A1(n4600), .A2(REG2_REG_21__SCAN_IN), .A3(
        REG2_REG_3__SCAN_IN), .A4(REG2_REG_30__SCAN_IN), .ZN(n4617) );
  NOR4_X1 U5173 ( .A1(n4602), .A2(n4601), .A3(n2437), .A4(IR_REG_17__SCAN_IN), 
        .ZN(n4612) );
  INV_X1 U5174 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4865) );
  NAND4_X1 U5175 ( .A1(REG3_REG_11__SCAN_IN), .A2(n4862), .A3(n4865), .A4(
        n4658), .ZN(n4610) );
  NAND4_X1 U5176 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .A3(
        IR_REG_7__SCAN_IN), .A4(n4685), .ZN(n4609) );
  NAND4_X1 U5177 ( .A1(DATAI_15_), .A2(REG2_REG_5__SCAN_IN), .A3(
        REG1_REG_5__SCAN_IN), .A4(ADDR_REG_8__SCAN_IN), .ZN(n4607) );
  NAND4_X1 U5178 ( .A1(REG2_REG_27__SCAN_IN), .A2(REG2_REG_10__SCAN_IN), .A3(
        REG2_REG_8__SCAN_IN), .A4(DATAI_18_), .ZN(n4606) );
  NAND4_X1 U5179 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .A3(
        IR_REG_2__SCAN_IN), .A4(n4603), .ZN(n4605) );
  NAND4_X1 U5180 ( .A1(REG2_REG_29__SCAN_IN), .A2(REG3_REG_23__SCAN_IN), .A3(
        n4661), .A4(n4864), .ZN(n4604) );
  OR4_X1 U5181 ( .A1(n4607), .A2(n4606), .A3(n4605), .A4(n4604), .ZN(n4608) );
  NOR4_X1 U5182 ( .A1(IR_REG_28__SCAN_IN), .A2(n4610), .A3(n4609), .A4(n4608), 
        .ZN(n4611) );
  NAND3_X1 U5183 ( .A1(n4612), .A2(IR_REG_18__SCAN_IN), .A3(n4611), .ZN(n4616)
         );
  NAND4_X1 U5184 ( .A1(n4613), .A2(IR_REG_24__SCAN_IN), .A3(IR_REG_23__SCAN_IN), .A4(STATE_REG_SCAN_IN), .ZN(n4615) );
  NAND4_X1 U5185 ( .A1(REG3_REG_0__SCAN_IN), .A2(REG1_REG_19__SCAN_IN), .A3(
        REG2_REG_28__SCAN_IN), .A4(ADDR_REG_19__SCAN_IN), .ZN(n4614) );
  NOR4_X1 U5186 ( .A1(n4617), .A2(n4616), .A3(n4615), .A4(n4614), .ZN(n4623)
         );
  NAND4_X1 U5187 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_29__SCAN_IN), .A4(DATAI_6_), .ZN(n4621) );
  NAND4_X1 U5188 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_25__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n4620) );
  NAND4_X1 U5189 ( .A1(REG2_REG_14__SCAN_IN), .A2(REG2_REG_11__SCAN_IN), .A3(
        REG0_REG_4__SCAN_IN), .A4(REG2_REG_0__SCAN_IN), .ZN(n4619) );
  NAND4_X1 U5190 ( .A1(REG0_REG_14__SCAN_IN), .A2(REG1_REG_14__SCAN_IN), .A3(
        REG1_REG_10__SCAN_IN), .A4(DATAI_2_), .ZN(n4618) );
  NOR4_X1 U5191 ( .A1(n4621), .A2(n4620), .A3(n4619), .A4(n4618), .ZN(n4622)
         );
  NAND2_X1 U5192 ( .A1(n4623), .A2(n4622), .ZN(n4624) );
  NOR4_X1 U5193 ( .A1(n4627), .A2(n4626), .A3(n4625), .A4(n4624), .ZN(n4879)
         );
  INV_X1 U5194 ( .A(DATAI_27_), .ZN(n4630) );
  AOI22_X1 U5195 ( .A1(n4630), .A2(keyinput117), .B1(keyinput112), .B2(n4629), 
        .ZN(n4628) );
  OAI221_X1 U5196 ( .B1(n4630), .B2(keyinput117), .C1(n4629), .C2(keyinput112), 
        .A(n4628), .ZN(n4643) );
  INV_X1 U5197 ( .A(DATAI_25_), .ZN(n4633) );
  AOI22_X1 U5198 ( .A1(n4633), .A2(keyinput64), .B1(keyinput54), .B2(n4632), 
        .ZN(n4631) );
  OAI221_X1 U5199 ( .B1(n4633), .B2(keyinput64), .C1(n4632), .C2(keyinput54), 
        .A(n4631), .ZN(n4642) );
  AOI22_X1 U5200 ( .A1(n4636), .A2(keyinput61), .B1(n4635), .B2(keyinput98), 
        .ZN(n4634) );
  OAI221_X1 U5201 ( .B1(n4636), .B2(keyinput61), .C1(n4635), .C2(keyinput98), 
        .A(n4634), .ZN(n4641) );
  AOI22_X1 U5202 ( .A1(n4639), .A2(keyinput2), .B1(n4638), .B2(keyinput113), 
        .ZN(n4637) );
  OAI221_X1 U5203 ( .B1(n4639), .B2(keyinput2), .C1(n4638), .C2(keyinput113), 
        .A(n4637), .ZN(n4640) );
  NOR4_X1 U5204 ( .A1(n4643), .A2(n4642), .A3(n4641), .A4(n4640), .ZN(n4683)
         );
  AOI22_X1 U5205 ( .A1(U3149), .A2(keyinput59), .B1(keyinput101), .B2(n4585), 
        .ZN(n4644) );
  OAI221_X1 U5206 ( .B1(U3149), .B2(keyinput59), .C1(n4585), .C2(keyinput101), 
        .A(n4644), .ZN(n4656) );
  INV_X1 U5207 ( .A(DATAI_9_), .ZN(n4646) );
  AOI22_X1 U5208 ( .A1(n4647), .A2(keyinput84), .B1(keyinput85), .B2(n4646), 
        .ZN(n4645) );
  OAI221_X1 U5209 ( .B1(n4647), .B2(keyinput84), .C1(n4646), .C2(keyinput85), 
        .A(n4645), .ZN(n4655) );
  INV_X1 U5210 ( .A(DATAI_6_), .ZN(n4650) );
  AOI22_X1 U5211 ( .A1(n4650), .A2(keyinput51), .B1(n4649), .B2(keyinput92), 
        .ZN(n4648) );
  OAI221_X1 U5212 ( .B1(n4650), .B2(keyinput51), .C1(n4649), .C2(keyinput92), 
        .A(n4648), .ZN(n4654) );
  XNOR2_X1 U5213 ( .A(DATAI_2_), .B(keyinput119), .ZN(n4652) );
  XNOR2_X1 U5214 ( .A(keyinput21), .B(DATAI_3_), .ZN(n4651) );
  NAND2_X1 U5215 ( .A1(n4652), .A2(n4651), .ZN(n4653) );
  NOR4_X1 U5216 ( .A1(n4656), .A2(n4655), .A3(n4654), .A4(n4653), .ZN(n4682)
         );
  AOI22_X1 U5217 ( .A1(n4658), .A2(keyinput43), .B1(n3899), .B2(keyinput90), 
        .ZN(n4657) );
  OAI221_X1 U5218 ( .B1(n4658), .B2(keyinput43), .C1(n3899), .C2(keyinput90), 
        .A(n4657), .ZN(n4668) );
  AOI22_X1 U5219 ( .A1(n4661), .A2(keyinput6), .B1(keyinput17), .B2(n4660), 
        .ZN(n4659) );
  OAI221_X1 U5220 ( .B1(n4661), .B2(keyinput6), .C1(n4660), .C2(keyinput17), 
        .A(n4659), .ZN(n4667) );
  XNOR2_X1 U5221 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput33), .ZN(n4665) );
  XNOR2_X1 U5222 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput75), .ZN(n4664) );
  XNOR2_X1 U5223 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput37), .ZN(n4663) );
  XNOR2_X1 U5224 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput46), .ZN(n4662) );
  NAND4_X1 U5225 ( .A1(n4665), .A2(n4664), .A3(n4663), .A4(n4662), .ZN(n4666)
         );
  NOR3_X1 U5226 ( .A1(n4668), .A2(n4667), .A3(n4666), .ZN(n4681) );
  XOR2_X1 U5227 ( .A(n4669), .B(keyinput29), .Z(n4673) );
  XNOR2_X1 U5228 ( .A(IR_REG_8__SCAN_IN), .B(keyinput30), .ZN(n4672) );
  XNOR2_X1 U5229 ( .A(IR_REG_7__SCAN_IN), .B(keyinput80), .ZN(n4671) );
  XNOR2_X1 U5230 ( .A(IR_REG_9__SCAN_IN), .B(keyinput95), .ZN(n4670) );
  NAND4_X1 U5231 ( .A1(n4673), .A2(n4672), .A3(n4671), .A4(n4670), .ZN(n4679)
         );
  XNOR2_X1 U5232 ( .A(IR_REG_3__SCAN_IN), .B(keyinput56), .ZN(n4677) );
  XNOR2_X1 U5233 ( .A(IR_REG_2__SCAN_IN), .B(keyinput87), .ZN(n4676) );
  XNOR2_X1 U5234 ( .A(IR_REG_6__SCAN_IN), .B(keyinput23), .ZN(n4675) );
  XNOR2_X1 U5235 ( .A(IR_REG_5__SCAN_IN), .B(keyinput109), .ZN(n4674) );
  NAND4_X1 U5236 ( .A1(n4677), .A2(n4676), .A3(n4675), .A4(n4674), .ZN(n4678)
         );
  NOR2_X1 U5237 ( .A1(n4679), .A2(n4678), .ZN(n4680) );
  NAND4_X1 U5238 ( .A1(n4683), .A2(n4682), .A3(n4681), .A4(n4680), .ZN(n4877)
         );
  AOI22_X1 U5239 ( .A1(n4686), .A2(keyinput31), .B1(keyinput99), .B2(n4685), 
        .ZN(n4684) );
  OAI221_X1 U5240 ( .B1(n4686), .B2(keyinput31), .C1(n4685), .C2(keyinput99), 
        .A(n4684), .ZN(n4696) );
  XNOR2_X1 U5241 ( .A(IR_REG_17__SCAN_IN), .B(keyinput8), .ZN(n4690) );
  XNOR2_X1 U5242 ( .A(IR_REG_13__SCAN_IN), .B(keyinput50), .ZN(n4689) );
  XNOR2_X1 U5243 ( .A(IR_REG_22__SCAN_IN), .B(keyinput42), .ZN(n4688) );
  XNOR2_X1 U5244 ( .A(IR_REG_21__SCAN_IN), .B(keyinput67), .ZN(n4687) );
  NAND4_X1 U5245 ( .A1(n4690), .A2(n4689), .A3(n4688), .A4(n4687), .ZN(n4695)
         );
  XNOR2_X1 U5246 ( .A(n4691), .B(keyinput106), .ZN(n4694) );
  XNOR2_X1 U5247 ( .A(n4692), .B(keyinput79), .ZN(n4693) );
  NOR4_X1 U5248 ( .A1(n4696), .A2(n4695), .A3(n4694), .A4(n4693), .ZN(n4747)
         );
  AOI22_X1 U5249 ( .A1(n4699), .A2(keyinput16), .B1(keyinput10), .B2(n4698), 
        .ZN(n4697) );
  OAI221_X1 U5250 ( .B1(n4699), .B2(keyinput16), .C1(n4698), .C2(keyinput10), 
        .A(n4697), .ZN(n4711) );
  AOI22_X1 U5251 ( .A1(n4702), .A2(keyinput11), .B1(keyinput41), .B2(n4701), 
        .ZN(n4700) );
  OAI221_X1 U5252 ( .B1(n4702), .B2(keyinput11), .C1(n4701), .C2(keyinput41), 
        .A(n4700), .ZN(n4710) );
  AOI22_X1 U5253 ( .A1(n4705), .A2(keyinput121), .B1(n4704), .B2(keyinput14), 
        .ZN(n4703) );
  OAI221_X1 U5254 ( .B1(n4705), .B2(keyinput121), .C1(n4704), .C2(keyinput14), 
        .A(n4703), .ZN(n4709) );
  XNOR2_X1 U5255 ( .A(D_REG_0__SCAN_IN), .B(keyinput39), .ZN(n4707) );
  XNOR2_X1 U5256 ( .A(IR_REG_28__SCAN_IN), .B(keyinput100), .ZN(n4706) );
  NAND2_X1 U5257 ( .A1(n4707), .A2(n4706), .ZN(n4708) );
  NOR4_X1 U5258 ( .A1(n4711), .A2(n4710), .A3(n4709), .A4(n4708), .ZN(n4746)
         );
  AOI22_X1 U5259 ( .A1(n4714), .A2(keyinput76), .B1(n4713), .B2(keyinput65), 
        .ZN(n4712) );
  OAI221_X1 U5260 ( .B1(n4714), .B2(keyinput76), .C1(n4713), .C2(keyinput65), 
        .A(n4712), .ZN(n4727) );
  AOI22_X1 U5261 ( .A1(n4717), .A2(keyinput110), .B1(keyinput1), .B2(n4716), 
        .ZN(n4715) );
  OAI221_X1 U5262 ( .B1(n4717), .B2(keyinput110), .C1(n4716), .C2(keyinput1), 
        .A(n4715), .ZN(n4726) );
  AOI22_X1 U5263 ( .A1(n4720), .A2(keyinput52), .B1(n4719), .B2(keyinput25), 
        .ZN(n4718) );
  OAI221_X1 U5264 ( .B1(n4720), .B2(keyinput52), .C1(n4719), .C2(keyinput25), 
        .A(n4718), .ZN(n4725) );
  AOI22_X1 U5265 ( .A1(n4723), .A2(keyinput94), .B1(n4722), .B2(keyinput63), 
        .ZN(n4721) );
  OAI221_X1 U5266 ( .B1(n4723), .B2(keyinput94), .C1(n4722), .C2(keyinput63), 
        .A(n4721), .ZN(n4724) );
  NOR4_X1 U5267 ( .A1(n4727), .A2(n4726), .A3(n4725), .A4(n4724), .ZN(n4745)
         );
  AOI22_X1 U5268 ( .A1(n4730), .A2(keyinput83), .B1(n4729), .B2(keyinput115), 
        .ZN(n4728) );
  OAI221_X1 U5269 ( .B1(n4730), .B2(keyinput83), .C1(n4729), .C2(keyinput115), 
        .A(n4728), .ZN(n4743) );
  AOI22_X1 U5270 ( .A1(n4733), .A2(keyinput44), .B1(keyinput0), .B2(n4732), 
        .ZN(n4731) );
  OAI221_X1 U5271 ( .B1(n4733), .B2(keyinput44), .C1(n4732), .C2(keyinput0), 
        .A(n4731), .ZN(n4742) );
  AOI22_X1 U5272 ( .A1(n4736), .A2(keyinput125), .B1(n4735), .B2(keyinput82), 
        .ZN(n4734) );
  OAI221_X1 U5273 ( .B1(n4736), .B2(keyinput125), .C1(n4735), .C2(keyinput82), 
        .A(n4734), .ZN(n4741) );
  INV_X1 U5274 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4739) );
  INV_X1 U5275 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4738) );
  AOI22_X1 U5276 ( .A1(n4739), .A2(keyinput62), .B1(keyinput38), .B2(n4738), 
        .ZN(n4737) );
  OAI221_X1 U5277 ( .B1(n4739), .B2(keyinput62), .C1(n4738), .C2(keyinput38), 
        .A(n4737), .ZN(n4740) );
  NOR4_X1 U5278 ( .A1(n4743), .A2(n4742), .A3(n4741), .A4(n4740), .ZN(n4744)
         );
  NAND4_X1 U5279 ( .A1(n4747), .A2(n4746), .A3(n4745), .A4(n4744), .ZN(n4876)
         );
  AOI22_X1 U5280 ( .A1(n4750), .A2(keyinput49), .B1(n4749), .B2(keyinput72), 
        .ZN(n4748) );
  OAI221_X1 U5281 ( .B1(n4750), .B2(keyinput49), .C1(n4749), .C2(keyinput72), 
        .A(n4748), .ZN(n4762) );
  AOI22_X1 U5282 ( .A1(n4753), .A2(keyinput116), .B1(keyinput47), .B2(n4752), 
        .ZN(n4751) );
  OAI221_X1 U5283 ( .B1(n4753), .B2(keyinput116), .C1(n4752), .C2(keyinput47), 
        .A(n4751), .ZN(n4761) );
  INV_X1 U5284 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4755) );
  AOI22_X1 U5285 ( .A1(n4756), .A2(keyinput91), .B1(n4755), .B2(keyinput22), 
        .ZN(n4754) );
  OAI221_X1 U5286 ( .B1(n4756), .B2(keyinput91), .C1(n4755), .C2(keyinput22), 
        .A(n4754), .ZN(n4760) );
  XNOR2_X1 U5287 ( .A(REG1_REG_2__SCAN_IN), .B(keyinput88), .ZN(n4758) );
  XNOR2_X1 U5288 ( .A(REG0_REG_28__SCAN_IN), .B(keyinput45), .ZN(n4757) );
  NAND2_X1 U5289 ( .A1(n4758), .A2(n4757), .ZN(n4759) );
  NOR4_X1 U5290 ( .A1(n4762), .A2(n4761), .A3(n4760), .A4(n4759), .ZN(n4807)
         );
  AOI22_X1 U5291 ( .A1(n2365), .A2(keyinput71), .B1(n4764), .B2(keyinput20), 
        .ZN(n4763) );
  OAI221_X1 U5292 ( .B1(n2365), .B2(keyinput71), .C1(n4764), .C2(keyinput20), 
        .A(n4763), .ZN(n4777) );
  AOI22_X1 U5293 ( .A1(n4767), .A2(keyinput127), .B1(keyinput55), .B2(n4766), 
        .ZN(n4765) );
  OAI221_X1 U5294 ( .B1(n4767), .B2(keyinput127), .C1(n4766), .C2(keyinput55), 
        .A(n4765), .ZN(n4776) );
  AOI22_X1 U5295 ( .A1(n4770), .A2(keyinput111), .B1(keyinput12), .B2(n4769), 
        .ZN(n4768) );
  OAI221_X1 U5296 ( .B1(n4770), .B2(keyinput111), .C1(n4769), .C2(keyinput12), 
        .A(n4768), .ZN(n4775) );
  AOI22_X1 U5297 ( .A1(n4773), .A2(keyinput108), .B1(n4772), .B2(keyinput34), 
        .ZN(n4771) );
  OAI221_X1 U5298 ( .B1(n4773), .B2(keyinput108), .C1(n4772), .C2(keyinput34), 
        .A(n4771), .ZN(n4774) );
  NOR4_X1 U5299 ( .A1(n4777), .A2(n4776), .A3(n4775), .A4(n4774), .ZN(n4806)
         );
  AOI22_X1 U5300 ( .A1(n4780), .A2(keyinput19), .B1(keyinput48), .B2(n4779), 
        .ZN(n4778) );
  OAI221_X1 U5301 ( .B1(n4780), .B2(keyinput19), .C1(n4779), .C2(keyinput48), 
        .A(n4778), .ZN(n4789) );
  AOI22_X1 U5302 ( .A1(n4403), .A2(keyinput120), .B1(keyinput114), .B2(n2965), 
        .ZN(n4781) );
  OAI221_X1 U5303 ( .B1(n4403), .B2(keyinput120), .C1(n2965), .C2(keyinput114), 
        .A(n4781), .ZN(n4788) );
  INV_X1 U5304 ( .A(REG2_REG_6__SCAN_IN), .ZN(n4783) );
  AOI22_X1 U5305 ( .A1(n4783), .A2(keyinput126), .B1(keyinput89), .B2(n2992), 
        .ZN(n4782) );
  OAI221_X1 U5306 ( .B1(n4783), .B2(keyinput126), .C1(n2992), .C2(keyinput89), 
        .A(n4782), .ZN(n4787) );
  INV_X1 U5307 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4785) );
  AOI22_X1 U5308 ( .A1(n4785), .A2(keyinput96), .B1(keyinput53), .B2(n2462), 
        .ZN(n4784) );
  OAI221_X1 U5309 ( .B1(n4785), .B2(keyinput96), .C1(n2462), .C2(keyinput53), 
        .A(n4784), .ZN(n4786) );
  NOR4_X1 U5310 ( .A1(n4789), .A2(n4788), .A3(n4787), .A4(n4786), .ZN(n4805)
         );
  INV_X1 U5311 ( .A(REG2_REG_10__SCAN_IN), .ZN(n4792) );
  AOI22_X1 U5312 ( .A1(n4792), .A2(keyinput32), .B1(n4791), .B2(keyinput26), 
        .ZN(n4790) );
  OAI221_X1 U5313 ( .B1(n4792), .B2(keyinput32), .C1(n4791), .C2(keyinput26), 
        .A(n4790), .ZN(n4803) );
  INV_X1 U5314 ( .A(REG2_REG_12__SCAN_IN), .ZN(n4795) );
  AOI22_X1 U5315 ( .A1(n4795), .A2(keyinput97), .B1(n4794), .B2(keyinput77), 
        .ZN(n4793) );
  OAI221_X1 U5316 ( .B1(n4795), .B2(keyinput97), .C1(n4794), .C2(keyinput77), 
        .A(n4793), .ZN(n4802) );
  INV_X1 U5317 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4797) );
  AOI22_X1 U5318 ( .A1(n4164), .A2(keyinput66), .B1(keyinput93), .B2(n4797), 
        .ZN(n4796) );
  OAI221_X1 U5319 ( .B1(n4164), .B2(keyinput66), .C1(n4797), .C2(keyinput93), 
        .A(n4796), .ZN(n4801) );
  INV_X1 U5320 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4799) );
  AOI22_X1 U5321 ( .A1(n3481), .A2(keyinput58), .B1(keyinput13), .B2(n4799), 
        .ZN(n4798) );
  OAI221_X1 U5322 ( .B1(n3481), .B2(keyinput58), .C1(n4799), .C2(keyinput13), 
        .A(n4798), .ZN(n4800) );
  NOR4_X1 U5323 ( .A1(n4803), .A2(n4802), .A3(n4801), .A4(n4800), .ZN(n4804)
         );
  NAND4_X1 U5324 ( .A1(n4807), .A2(n4806), .A3(n4805), .A4(n4804), .ZN(n4875)
         );
  AOI22_X1 U5325 ( .A1(n3497), .A2(keyinput60), .B1(keyinput7), .B2(n4809), 
        .ZN(n4808) );
  OAI221_X1 U5326 ( .B1(n3497), .B2(keyinput60), .C1(n4809), .C2(keyinput7), 
        .A(n4808), .ZN(n4821) );
  AOI22_X1 U5327 ( .A1(n4812), .A2(keyinput35), .B1(keyinput123), .B2(n4811), 
        .ZN(n4810) );
  OAI221_X1 U5328 ( .B1(n4812), .B2(keyinput35), .C1(n4811), .C2(keyinput123), 
        .A(n4810), .ZN(n4820) );
  INV_X1 U5329 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n4815) );
  AOI22_X1 U5330 ( .A1(n4815), .A2(keyinput18), .B1(n4814), .B2(keyinput78), 
        .ZN(n4813) );
  OAI221_X1 U5331 ( .B1(n4815), .B2(keyinput18), .C1(n4814), .C2(keyinput78), 
        .A(n4813), .ZN(n4819) );
  INV_X1 U5332 ( .A(ADDR_REG_12__SCAN_IN), .ZN(n4817) );
  AOI22_X1 U5333 ( .A1(n2725), .A2(keyinput103), .B1(n4817), .B2(keyinput81), 
        .ZN(n4816) );
  OAI221_X1 U5334 ( .B1(n2725), .B2(keyinput103), .C1(n4817), .C2(keyinput81), 
        .A(n4816), .ZN(n4818) );
  NOR4_X1 U5335 ( .A1(n4821), .A2(n4820), .A3(n4819), .A4(n4818), .ZN(n4873)
         );
  INV_X1 U5336 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n4824) );
  AOI22_X1 U5337 ( .A1(n4824), .A2(keyinput36), .B1(n4823), .B2(keyinput102), 
        .ZN(n4822) );
  OAI221_X1 U5338 ( .B1(n4824), .B2(keyinput36), .C1(n4823), .C2(keyinput102), 
        .A(n4822), .ZN(n4837) );
  AOI22_X1 U5339 ( .A1(n4827), .A2(keyinput118), .B1(n4826), .B2(keyinput15), 
        .ZN(n4825) );
  OAI221_X1 U5340 ( .B1(n4827), .B2(keyinput118), .C1(n4826), .C2(keyinput15), 
        .A(n4825), .ZN(n4836) );
  AOI22_X1 U5341 ( .A1(n4830), .A2(keyinput86), .B1(n4829), .B2(keyinput74), 
        .ZN(n4828) );
  OAI221_X1 U5342 ( .B1(n4830), .B2(keyinput86), .C1(n4829), .C2(keyinput74), 
        .A(n4828), .ZN(n4835) );
  AOI22_X1 U5343 ( .A1(n4833), .A2(keyinput70), .B1(n4832), .B2(keyinput104), 
        .ZN(n4831) );
  OAI221_X1 U5344 ( .B1(n4833), .B2(keyinput70), .C1(n4832), .C2(keyinput104), 
        .A(n4831), .ZN(n4834) );
  NOR4_X1 U5345 ( .A1(n4837), .A2(n4836), .A3(n4835), .A4(n4834), .ZN(n4872)
         );
  AOI22_X1 U5346 ( .A1(n4840), .A2(keyinput3), .B1(n4839), .B2(keyinput68), 
        .ZN(n4838) );
  OAI221_X1 U5347 ( .B1(n4840), .B2(keyinput3), .C1(n4839), .C2(keyinput68), 
        .A(n4838), .ZN(n4853) );
  AOI22_X1 U5348 ( .A1(n4843), .A2(keyinput105), .B1(keyinput28), .B2(n4842), 
        .ZN(n4841) );
  OAI221_X1 U5349 ( .B1(n4843), .B2(keyinput105), .C1(n4842), .C2(keyinput28), 
        .A(n4841), .ZN(n4852) );
  AOI22_X1 U5350 ( .A1(n4846), .A2(keyinput4), .B1(keyinput5), .B2(n4845), 
        .ZN(n4844) );
  OAI221_X1 U5351 ( .B1(n4846), .B2(keyinput4), .C1(n4845), .C2(keyinput5), 
        .A(n4844), .ZN(n4851) );
  AOI22_X1 U5352 ( .A1(n4849), .A2(keyinput24), .B1(keyinput124), .B2(n4848), 
        .ZN(n4847) );
  OAI221_X1 U5353 ( .B1(n4849), .B2(keyinput24), .C1(n4848), .C2(keyinput124), 
        .A(n4847), .ZN(n4850) );
  NOR4_X1 U5354 ( .A1(n4853), .A2(n4852), .A3(n4851), .A4(n4850), .ZN(n4871)
         );
  AOI22_X1 U5355 ( .A1(n4856), .A2(keyinput27), .B1(n4855), .B2(keyinput40), 
        .ZN(n4854) );
  OAI221_X1 U5356 ( .B1(n4856), .B2(keyinput27), .C1(n4855), .C2(keyinput40), 
        .A(n4854), .ZN(n4869) );
  AOI22_X1 U5357 ( .A1(n4859), .A2(keyinput57), .B1(keyinput73), .B2(n4858), 
        .ZN(n4857) );
  OAI221_X1 U5358 ( .B1(n4859), .B2(keyinput57), .C1(n4858), .C2(keyinput73), 
        .A(n4857), .ZN(n4868) );
  AOI22_X1 U5359 ( .A1(n4862), .A2(keyinput9), .B1(keyinput122), .B2(n4861), 
        .ZN(n4860) );
  OAI221_X1 U5360 ( .B1(n4862), .B2(keyinput9), .C1(n4861), .C2(keyinput122), 
        .A(n4860), .ZN(n4867) );
  AOI22_X1 U5361 ( .A1(n4865), .A2(keyinput69), .B1(n4864), .B2(keyinput107), 
        .ZN(n4863) );
  OAI221_X1 U5362 ( .B1(n4865), .B2(keyinput69), .C1(n4864), .C2(keyinput107), 
        .A(n4863), .ZN(n4866) );
  NOR4_X1 U5363 ( .A1(n4869), .A2(n4868), .A3(n4867), .A4(n4866), .ZN(n4870)
         );
  NAND4_X1 U5364 ( .A1(n4873), .A2(n4872), .A3(n4871), .A4(n4870), .ZN(n4874)
         );
  NOR4_X1 U5365 ( .A1(n4877), .A2(n4876), .A3(n4875), .A4(n4874), .ZN(n4878)
         );
  XOR2_X1 U5366 ( .A(n4879), .B(n4878), .Z(n4880) );
  XNOR2_X1 U5367 ( .A(n4881), .B(n4880), .ZN(U3579) );
  OR2_X1 U2383 ( .A1(n4416), .A2(n2207), .ZN(n2205) );
  CLKBUF_X3 U2398 ( .A(n2681), .Z(n2133) );
  CLKBUF_X1 U2403 ( .A(n4391), .Z(n2136) );
endmodule

