

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, keyinput58, 
        keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, keyinput52, 
        keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, keyinput46, 
        keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, keyinput40, 
        keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, keyinput34, 
        keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, keyinput28, 
        keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, keyinput22, 
        keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, keyinput16, 
        keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, 
        keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, 
        keyinput3, keyinput2, keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086;

  AND2_X1 U4770 ( .A1(n8298), .A2(n8190), .ZN(n8189) );
  NAND2_X1 U4771 ( .A1(n5535), .A2(n4349), .ZN(n9406) );
  OR2_X1 U4772 ( .A1(n5476), .A2(n9109), .ZN(n6284) );
  INV_X1 U4773 ( .A(n5676), .ZN(n8113) );
  AND2_X1 U4774 ( .A1(n6852), .A2(n6851), .ZN(n6853) );
  INV_X2 U4775 ( .A(n5649), .ZN(n5670) );
  INV_X2 U4776 ( .A(n6196), .ZN(n5446) );
  NAND4_X2 U4777 ( .A1(n5653), .A2(n5650), .A3(n5651), .A4(n5652), .ZN(n8383)
         );
  AND2_X1 U4778 ( .A1(n8890), .A2(n7914), .ZN(n5671) );
  NAND2_X1 U4779 ( .A1(n6329), .A2(n6348), .ZN(n5287) );
  NAND2_X1 U4780 ( .A1(n5464), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5466) );
  INV_X1 U4782 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4505) );
  INV_X1 U4783 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5465) );
  INV_X1 U4784 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5456) );
  INV_X1 U4785 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5190) );
  CLKBUF_X1 U4786 ( .A(n9175), .Z(n4264) );
  OAI21_X1 U4787 ( .B1(n6558), .B2(n6624), .A(n9471), .ZN(n9175) );
  INV_X1 U4788 ( .A(n5960), .ZN(n4265) );
  AND2_X1 U4789 ( .A1(n5783), .A2(n5566), .ZN(n5959) );
  INV_X1 U4790 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5506) );
  INV_X2 U4791 ( .A(n9058), .ZN(n4497) );
  INV_X1 U4792 ( .A(n5671), .ZN(n4267) );
  INV_X2 U4793 ( .A(n7121), .ZN(n7593) );
  INV_X1 U4794 ( .A(n6329), .ZN(n5256) );
  NAND2_X1 U4795 ( .A1(n5991), .A2(n5992), .ZN(n5665) );
  OR2_X1 U4796 ( .A1(n8883), .A2(n8884), .ZN(n5590) );
  NOR2_X1 U4797 ( .A1(n5510), .A2(n7906), .ZN(n5511) );
  BUF_X1 U4798 ( .A(n5035), .Z(n5447) );
  AND2_X1 U4799 ( .A1(n6479), .A2(n7551), .ZN(n6632) );
  INV_X1 U4800 ( .A(n7605), .ZN(n6479) );
  OAI21_X1 U4801 ( .B1(n9406), .B2(n4791), .A(n4789), .ZN(n4795) );
  OAI21_X1 U4802 ( .B1(n7632), .B2(n5968), .A(n8032), .ZN(n7705) );
  BUF_X1 U4803 ( .A(n5665), .Z(n6324) );
  NAND2_X1 U4804 ( .A1(n7846), .A2(n5511), .ZN(n6521) );
  AOI21_X1 U4805 ( .B1(P1_REG1_REG_0__SCAN_IN), .B2(n6484), .A(n6527), .ZN(
        n6529) );
  INV_X1 U4806 ( .A(n9268), .ZN(n6623) );
  INV_X2 U4807 ( .A(n5287), .ZN(n6191) );
  BUF_X4 U4808 ( .A(n5120), .Z(n4266) );
  NAND2_X1 U4809 ( .A1(n4799), .A2(n4996), .ZN(n5120) );
  NAND2_X1 U4810 ( .A1(n6850), .A2(n6849), .ZN(n6854) );
  NAND2_X2 U4811 ( .A1(n4489), .A2(n5696), .ZN(n7165) );
  NAND2_X2 U4813 ( .A1(n7705), .A2(n7798), .ZN(n5969) );
  OAI21_X2 U4815 ( .B1(n7959), .B2(n5941), .A(n5940), .ZN(n8552) );
  AND2_X4 U4816 ( .A1(n6532), .A2(n6485), .ZN(n9058) );
  AOI21_X2 U4817 ( .B1(n8562), .B2(n8350), .A(n5942), .ZN(n8543) );
  AOI21_X2 U4818 ( .B1(n8546), .B2(n8812), .A(n8552), .ZN(n5942) );
  AOI21_X4 U4819 ( .B1(n6391), .B2(n6394), .A(n4854), .ZN(n6850) );
  INV_X4 U4820 ( .A(n4267), .ZN(n4268) );
  XNOR2_X2 U4821 ( .A(n5507), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6481) );
  XNOR2_X2 U4822 ( .A(n5570), .B(n5588), .ZN(n5991) );
  XNOR2_X2 U4823 ( .A(n4993), .B(n4992), .ZN(n4997) );
  AOI22_X2 U4825 ( .A1(n6955), .A2(n6954), .B1(n6958), .B2(n6953), .ZN(n6957)
         );
  AND2_X2 U4826 ( .A1(n6623), .A2(n7551), .ZN(n6480) );
  XNOR2_X2 U4827 ( .A(n5131), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6409) );
  XNOR2_X1 U4828 ( .A(n8197), .B(n8198), .ZN(n8346) );
  AND2_X1 U4829 ( .A1(n4476), .A2(n4333), .ZN(n8565) );
  OR2_X1 U4830 ( .A1(n8592), .A2(n8081), .ZN(n8586) );
  NAND2_X1 U4831 ( .A1(n8322), .A2(n8185), .ZN(n8186) );
  NAND2_X1 U4832 ( .A1(n8324), .A2(n8323), .ZN(n8322) );
  XNOR2_X1 U4833 ( .A(n7666), .B(n4296), .ZN(n7595) );
  NOR2_X1 U4834 ( .A1(n9215), .A2(n7092), .ZN(n5522) );
  NAND2_X1 U4835 ( .A1(n7997), .A2(n8003), .ZN(n8131) );
  AND2_X1 U4836 ( .A1(n5154), .A2(n5153), .ZN(n7092) );
  NAND2_X1 U4837 ( .A1(n6046), .A2(n5962), .ZN(n8719) );
  INV_X1 U4838 ( .A(n8381), .ZN(n6958) );
  INV_X2 U4839 ( .A(n8988), .ZN(n6689) );
  INV_X2 U4840 ( .A(n9761), .ZN(n7051) );
  INV_X1 U4841 ( .A(n5649), .ZN(n4269) );
  XNOR2_X1 U4842 ( .A(n5590), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5592) );
  CLKBUF_X2 U4843 ( .A(n5992), .Z(n8474) );
  MUX2_X1 U4844 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4983), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n4984) );
  NAND2_X1 U4845 ( .A1(n5455), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5059) );
  INV_X8 U4846 ( .A(n6345), .ZN(n6348) );
  OAI21_X1 U4847 ( .B1(n9163), .B2(n9162), .A(n9161), .ZN(n9166) );
  AOI21_X1 U4848 ( .B1(n4490), .B2(n8719), .A(n4352), .ZN(n8804) );
  AND2_X1 U4849 ( .A1(n4626), .A2(n4871), .ZN(n4428) );
  NAND2_X1 U4850 ( .A1(n8346), .A2(n8553), .ZN(n8201) );
  NAND2_X1 U4851 ( .A1(n8196), .A2(n8195), .ZN(n8197) );
  NOR2_X1 U4852 ( .A1(n8127), .A2(n8165), .ZN(n4724) );
  AND2_X1 U4853 ( .A1(n9325), .A2(n4389), .ZN(n9275) );
  NAND2_X1 U4854 ( .A1(n4364), .A2(n6144), .ZN(n9363) );
  NAND2_X1 U4855 ( .A1(n8188), .A2(n8187), .ZN(n8298) );
  NAND2_X1 U4856 ( .A1(n5335), .A2(n6293), .ZN(n9389) );
  NOR2_X1 U4857 ( .A1(n4607), .A2(n4604), .ZN(n4603) );
  OAI21_X1 U4858 ( .B1(n9206), .B2(n7861), .A(n7727), .ZN(n7783) );
  NAND2_X1 U4859 ( .A1(n7729), .A2(n7728), .ZN(n7727) );
  XNOR2_X1 U4860 ( .A(n8408), .B(n8409), .ZN(n8386) );
  AND2_X1 U4861 ( .A1(n4710), .A2(n4709), .ZN(n8408) );
  NAND2_X1 U4862 ( .A1(n7623), .A2(n7622), .ZN(n7621) );
  AOI21_X1 U4863 ( .B1(n4792), .B2(n4790), .A(n4346), .ZN(n4789) );
  INV_X1 U4864 ( .A(n4792), .ZN(n4791) );
  INV_X1 U4865 ( .A(n8074), .ZN(n4604) );
  NAND2_X1 U4866 ( .A1(n8733), .A2(n8052), .ZN(n8702) );
  XNOR2_X1 U4867 ( .A(n7815), .B(n7816), .ZN(n7685) );
  AOI21_X1 U4868 ( .B1(n4637), .B2(n4635), .A(n4634), .ZN(n4633) );
  AND2_X1 U4869 ( .A1(n4696), .A2(n4695), .ZN(n7815) );
  AND2_X1 U4870 ( .A1(n4638), .A2(n9452), .ZN(n4637) );
  NAND2_X1 U4871 ( .A1(n6284), .A2(n6287), .ZN(n9468) );
  NAND2_X1 U4872 ( .A1(n5062), .A2(n5061), .ZN(n9540) );
  NAND2_X1 U4873 ( .A1(n8307), .A2(n7775), .ZN(n7848) );
  NAND2_X1 U4874 ( .A1(n8309), .A2(n8308), .ZN(n8307) );
  XNOR2_X1 U4875 ( .A(n7437), .B(n7438), .ZN(n7339) );
  AND2_X1 U4876 ( .A1(n4712), .A2(n4711), .ZN(n7437) );
  NAND2_X1 U4877 ( .A1(n7125), .A2(n7126), .ZN(n7206) );
  NAND2_X1 U4878 ( .A1(n5292), .A2(n5291), .ZN(n7861) );
  AND2_X1 U4879 ( .A1(n7042), .A2(n7044), .ZN(n4382) );
  NOR2_X2 U4880 ( .A1(n7264), .A2(n7484), .ZN(n7430) );
  NAND2_X1 U4881 ( .A1(n5284), .A2(n4858), .ZN(n5286) );
  NAND2_X1 U4882 ( .A1(n5223), .A2(n5222), .ZN(n7564) );
  NAND2_X1 U4883 ( .A1(n6788), .A2(n6787), .ZN(n8365) );
  NAND2_X1 U4884 ( .A1(n4650), .A2(n6263), .ZN(n7016) );
  INV_X1 U4885 ( .A(n6857), .ZN(n8202) );
  XNOR2_X2 U4886 ( .A(n6857), .B(n6941), .ZN(n6856) );
  INV_X2 U4887 ( .A(n9142), .ZN(n4270) );
  CLKBUF_X1 U4888 ( .A(n5104), .Z(n6559) );
  NAND4_X1 U4889 ( .A1(n5703), .A2(n5702), .A3(n5701), .A4(n5700), .ZN(n8379)
         );
  NAND4_X1 U4890 ( .A1(n5675), .A2(n5674), .A3(n5673), .A4(n5672), .ZN(n8381)
         );
  AND3_X1 U4891 ( .A1(n5695), .A2(n5694), .A3(n5693), .ZN(n7228) );
  NAND2_X1 U4892 ( .A1(n4800), .A2(n4796), .ZN(n5104) );
  NAND2_X1 U4893 ( .A1(n5658), .A2(n5657), .ZN(n6941) );
  CLKBUF_X3 U4894 ( .A(n5668), .Z(n7108) );
  NAND2_X2 U4895 ( .A1(n5592), .A2(n7914), .ZN(n5649) );
  AND2_X1 U4896 ( .A1(n8890), .A2(n5593), .ZN(n5668) );
  INV_X1 U4897 ( .A(n5592), .ZN(n8890) );
  NAND2_X2 U4898 ( .A1(n4799), .A2(n9628), .ZN(n5141) );
  INV_X2 U4899 ( .A(n6324), .ZN(n5897) );
  XNOR2_X1 U4900 ( .A(n6007), .B(n4365), .ZN(n6016) );
  INV_X1 U4901 ( .A(n5593), .ZN(n7914) );
  NAND2_X1 U4902 ( .A1(n5880), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U4903 ( .A1(n4853), .A2(n6009), .ZN(n7902) );
  XNOR2_X1 U4904 ( .A(n5591), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5593) );
  INV_X1 U4905 ( .A(n4996), .ZN(n9628) );
  NAND2_X1 U4906 ( .A1(n4804), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5591) );
  XNOR2_X1 U4907 ( .A(n5489), .B(P1_IR_REG_24__SCAN_IN), .ZN(n7846) );
  NAND2_X1 U4908 ( .A1(n4685), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5489) );
  NAND2_X1 U4909 ( .A1(n5488), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5507) );
  INV_X1 U4910 ( .A(n5455), .ZN(n5463) );
  AND2_X1 U4911 ( .A1(n4684), .A2(n4332), .ZN(n4683) );
  NOR2_X1 U4912 ( .A1(n5565), .A2(n5564), .ZN(n5566) );
  NAND2_X2 U4913 ( .A1(n4452), .A2(n4450), .ZN(n4901) );
  NAND3_X1 U4914 ( .A1(n8505), .A2(n4879), .A3(n4453), .ZN(n4452) );
  INV_X1 U4915 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8505) );
  INV_X1 U4916 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5239) );
  NOR3_X1 U4917 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n5568) );
  INV_X1 U4918 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4879) );
  INV_X4 U4919 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U4920 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4757) );
  INV_X1 U4921 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5168) );
  INV_X1 U4922 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4714) );
  NOR2_X1 U4923 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5559) );
  INV_X1 U4924 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5854) );
  INV_X1 U4925 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5849) );
  INV_X4 U4926 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U4927 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5881) );
  INV_X1 U4928 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4992) );
  INV_X2 U4929 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n10035) );
  NOR2_X1 U4930 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5560) );
  NOR2_X1 U4931 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5558) );
  NAND2_X1 U4932 ( .A1(n4271), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U4933 ( .A1(n5959), .A2(n4847), .ZN(n4271) );
  NAND2_X1 U4934 ( .A1(n8910), .A2(n8911), .ZN(n4678) );
  NAND2_X1 U4935 ( .A1(n4677), .A2(n4676), .ZN(n4675) );
  NAND2_X1 U4936 ( .A1(n8297), .A2(n8189), .ZN(n4272) );
  NAND2_X2 U4937 ( .A1(n8246), .A2(n8326), .ZN(n8297) );
  OAI22_X1 U4938 ( .A1(n6866), .A2(n6865), .B1(n8383), .B2(n6856), .ZN(n6955)
         );
  NOR2_X2 U4939 ( .A1(n7062), .A2(n7063), .ZN(n7286) );
  AOI21_X2 U4940 ( .B1(n8257), .B2(n4824), .A(n4822), .ZN(n8324) );
  OR2_X2 U4941 ( .A1(n8226), .A2(n8227), .ZN(n8228) );
  NAND2_X2 U4942 ( .A1(n8201), .A2(n8200), .ZN(n8226) );
  OAI222_X1 U4943 ( .A1(n8901), .A2(n7903), .B1(P2_U3151), .B2(n7902), .C1(
        n7901), .C2(n8893), .ZN(P2_U3271) );
  OAI222_X1 U4944 ( .A1(n8901), .A2(n7905), .B1(P2_U3151), .B2(n6016), .C1(
        n7900), .C2(n8893), .ZN(P2_U3270) );
  NOR2_X2 U4945 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5677) );
  XNOR2_X1 U4946 ( .A(n6856), .B(n8383), .ZN(n6866) );
  NOR2_X2 U4947 ( .A1(n9529), .A2(n9432), .ZN(n9414) );
  XNOR2_X2 U4948 ( .A(n8186), .B(n8187), .ZN(n8246) );
  OAI21_X2 U4949 ( .B1(n8358), .B2(n4835), .A(n4832), .ZN(n8290) );
  OAI21_X2 U4950 ( .B1(n8237), .B2(n8236), .A(n8235), .ZN(n8234) );
  NOR2_X2 U4951 ( .A1(n7949), .A2(n7950), .ZN(n8237) );
  NAND2_X1 U4952 ( .A1(n9628), .A2(n4997), .ZN(n5035) );
  NAND2_X1 U4953 ( .A1(n4716), .A2(n5406), .ZN(n5423) );
  NAND2_X1 U4954 ( .A1(n5405), .A2(n5404), .ZN(n4716) );
  NAND2_X1 U4955 ( .A1(n5189), .A2(n4459), .ZN(n4460) );
  AND2_X1 U4956 ( .A1(n4931), .A2(n4279), .ZN(n4459) );
  AND2_X1 U4957 ( .A1(n8035), .A2(n8037), .ZN(n7798) );
  NAND2_X1 U4958 ( .A1(n4624), .A2(n4307), .ZN(n4623) );
  NOR2_X1 U4959 ( .A1(n8536), .A2(n8086), .ZN(n4625) );
  INV_X1 U4960 ( .A(n9014), .ZN(n4676) );
  INV_X1 U4961 ( .A(n5322), .ZN(n6190) );
  INV_X1 U4962 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4985) );
  NAND2_X1 U4963 ( .A1(n4521), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4986) );
  INV_X1 U4964 ( .A(n7016), .ZN(n4539) );
  NOR2_X1 U4965 ( .A1(n4446), .A2(n8110), .ZN(n4441) );
  INV_X1 U4966 ( .A(n8129), .ZN(n4446) );
  OR2_X1 U4967 ( .A1(n9518), .A2(n6075), .ZN(n6215) );
  INV_X1 U4968 ( .A(n4445), .ZN(n4438) );
  OR2_X1 U4969 ( .A1(n6040), .A2(n8370), .ZN(n8118) );
  NAND2_X1 U4970 ( .A1(n4745), .A2(n4343), .ZN(n4455) );
  AND2_X1 U4971 ( .A1(n4275), .A2(n4353), .ZN(n4457) );
  AND2_X1 U4972 ( .A1(n4274), .A2(n4305), .ZN(n4471) );
  OR2_X1 U4973 ( .A1(n9860), .A2(n8310), .ZN(n8034) );
  OR2_X1 U4974 ( .A1(n8380), .A2(n7228), .ZN(n7997) );
  OR2_X1 U4975 ( .A1(n8822), .A2(n8251), .ZN(n8129) );
  INV_X1 U4976 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4451) );
  NOR2_X1 U4977 ( .A1(n6207), .A2(n4570), .ZN(n4569) );
  NAND2_X1 U4978 ( .A1(n6164), .A2(n6168), .ZN(n4570) );
  NOR2_X1 U4979 ( .A1(n6229), .A2(n4568), .ZN(n4567) );
  NAND2_X1 U4980 ( .A1(n6165), .A2(n6310), .ZN(n4568) );
  OAI21_X1 U4981 ( .B1(n4266), .B2(n5087), .A(n4802), .ZN(n4801) );
  NAND2_X1 U4982 ( .A1(n9349), .A2(n4873), .ZN(n4629) );
  INV_X1 U4983 ( .A(n6273), .ZN(n4647) );
  NOR2_X1 U4984 ( .A1(n6059), .A2(n4765), .ZN(n4764) );
  INV_X1 U4985 ( .A(n5543), .ZN(n4765) );
  NAND2_X1 U4986 ( .A1(n4395), .A2(n9137), .ZN(n4788) );
  OR2_X1 U4987 ( .A1(n9616), .A2(n9098), .ZN(n6283) );
  OR2_X1 U4988 ( .A1(n7861), .A2(n7863), .ZN(n6276) );
  NAND2_X1 U4989 ( .A1(n9792), .A2(n7644), .ZN(n4756) );
  NAND2_X1 U4990 ( .A1(n5423), .A2(n5422), .ZN(n5442) );
  NAND2_X1 U4991 ( .A1(n5389), .A2(n5388), .ZN(n5405) );
  INV_X1 U4992 ( .A(n4738), .ZN(n4737) );
  AOI21_X1 U4993 ( .B1(n4738), .B2(n4736), .A(n4735), .ZN(n4734) );
  OAI211_X1 U4994 ( .C1(n4455), .C2(n4295), .A(n4368), .B(n4742), .ZN(n5016)
         );
  AOI21_X1 U4995 ( .B1(n4744), .B2(n4745), .A(n4743), .ZN(n4742) );
  NAND2_X1 U4996 ( .A1(n4370), .A2(n4369), .ZN(n4368) );
  INV_X1 U4997 ( .A(n4958), .ZN(n4743) );
  NAND2_X1 U4998 ( .A1(n4778), .A2(n4514), .ZN(n5455) );
  NAND2_X1 U4999 ( .A1(n5206), .A2(n4918), .ZN(n5189) );
  OAI21_X1 U5000 ( .B1(n4820), .B2(n4816), .A(n4815), .ZN(n4814) );
  NOR2_X1 U5001 ( .A1(n4819), .A2(n4817), .ZN(n4816) );
  NAND2_X1 U5002 ( .A1(n4820), .A2(n8204), .ZN(n4815) );
  INV_X1 U5003 ( .A(n8204), .ZN(n4817) );
  INV_X1 U5004 ( .A(n8255), .ZN(n4828) );
  OAI21_X1 U5005 ( .B1(n8126), .B2(n8125), .A(n8168), .ZN(n4626) );
  INV_X1 U5006 ( .A(n8167), .ZN(n8168) );
  OAI21_X1 U5007 ( .B1(n8166), .B2(n6945), .A(n8165), .ZN(n8167) );
  CLKBUF_X1 U5008 ( .A(n5649), .Z(n7111) );
  INV_X1 U5009 ( .A(n8499), .ZN(n4694) );
  OR2_X1 U5010 ( .A1(n5932), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5934) );
  NAND2_X1 U5011 ( .A1(n5796), .A2(n5795), .ZN(n7716) );
  OAI21_X1 U5012 ( .B1(n8005), .B2(n4612), .A(n8010), .ZN(n4611) );
  OAI21_X1 U5013 ( .B1(n7165), .B2(n5708), .A(n5709), .ZN(n7253) );
  OR2_X1 U5014 ( .A1(n8812), .A2(n8350), .ZN(n8540) );
  XNOR2_X1 U5015 ( .A(n8806), .B(n8554), .ZN(n8544) );
  AND2_X1 U5016 ( .A1(n5575), .A2(n5574), .ZN(n8095) );
  NAND2_X1 U5017 ( .A1(n5987), .A2(n5986), .ZN(n7957) );
  INV_X1 U5018 ( .A(n5656), .ZN(n5898) );
  OR2_X1 U5019 ( .A1(n6945), .A2(n8172), .ZN(n9842) );
  INV_X1 U5020 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4627) );
  NAND2_X1 U5021 ( .A1(n6257), .A2(n9268), .ZN(n6260) );
  AND3_X1 U5022 ( .A1(n5056), .A2(n5055), .A3(n5054), .ZN(n9110) );
  AND4_X1 U5023 ( .A1(n5314), .A2(n5313), .A3(n5312), .A4(n5311), .ZN(n8914)
         );
  NOR2_X1 U5024 ( .A1(n7918), .A2(n4390), .ZN(n4389) );
  INV_X1 U5025 ( .A(n4392), .ZN(n4390) );
  NAND2_X1 U5026 ( .A1(n9321), .A2(n6153), .ZN(n9304) );
  AND2_X1 U5027 ( .A1(n5480), .A2(n9196), .ZN(n9320) );
  NAND2_X1 U5028 ( .A1(n4632), .A2(n4637), .ZN(n9451) );
  NAND2_X1 U5029 ( .A1(n9461), .A2(n6284), .ZN(n4632) );
  NAND2_X1 U5030 ( .A1(n9268), .A2(n6481), .ZN(n6627) );
  NAND2_X1 U5031 ( .A1(n4775), .A2(n4773), .ZN(n4772) );
  INV_X1 U5032 ( .A(n5530), .ZN(n4773) );
  XNOR2_X1 U5033 ( .A(n6189), .B(n6188), .ZN(n8882) );
  OAI21_X1 U5034 ( .B1(n6185), .B2(n6184), .A(n6183), .ZN(n6189) );
  OR2_X1 U5035 ( .A1(n9621), .A2(n5457), .ZN(n5026) );
  AND2_X1 U5036 ( .A1(n4939), .A2(n4937), .ZN(n4725) );
  INV_X1 U5037 ( .A(n5267), .ZN(n4939) );
  NAND2_X1 U5038 ( .A1(n6003), .A2(n6002), .ZN(n8528) );
  INV_X1 U5039 ( .A(n6001), .ZN(n6002) );
  OAI21_X1 U5040 ( .B1(n8535), .B2(n7612), .A(n6000), .ZN(n6001) );
  NAND2_X1 U5041 ( .A1(n5030), .A2(n5029), .ZN(n9529) );
  NAND2_X1 U5042 ( .A1(n5413), .A2(n5412), .ZN(n9010) );
  NOR2_X1 U5043 ( .A1(n6081), .A2(n6310), .ZN(n4538) );
  NAND2_X1 U5044 ( .A1(n4432), .A2(n4431), .ZN(n8065) );
  AOI21_X1 U5045 ( .B1(n4433), .B2(n4436), .A(n5875), .ZN(n4431) );
  NOR2_X1 U5046 ( .A1(n4435), .A2(n4434), .ZN(n4433) );
  NAND2_X1 U5047 ( .A1(n4520), .A2(n9452), .ZN(n6138) );
  AOI21_X1 U5048 ( .B1(n6128), .B2(n4519), .A(n4516), .ZN(n4518) );
  AND2_X1 U5049 ( .A1(n8571), .A2(n4440), .ZN(n4439) );
  AOI21_X1 U5050 ( .B1(n4441), .B2(n8080), .A(n4326), .ZN(n4440) );
  NOR2_X1 U5051 ( .A1(n8088), .A2(n8159), .ZN(n4445) );
  AOI211_X1 U5052 ( .C1(n8079), .C2(n8078), .A(n8081), .B(n8077), .ZN(n8083)
         );
  NAND2_X1 U5053 ( .A1(n4419), .A2(n8072), .ZN(n8078) );
  NAND2_X1 U5054 ( .A1(n4454), .A2(n6168), .ZN(n4575) );
  NAND2_X1 U5055 ( .A1(n6219), .A2(n6154), .ZN(n4454) );
  AOI21_X1 U5056 ( .B1(n4541), .B2(n6145), .A(n4540), .ZN(n6149) );
  INV_X1 U5057 ( .A(n9364), .ZN(n4540) );
  NAND2_X1 U5058 ( .A1(n4543), .A2(n4542), .ZN(n4541) );
  INV_X1 U5059 ( .A(n4575), .ZN(n4580) );
  NOR2_X1 U5060 ( .A1(n6156), .A2(n6168), .ZN(n4577) );
  INV_X1 U5061 ( .A(n6151), .ZN(n4582) );
  NAND2_X1 U5062 ( .A1(n6154), .A2(n4313), .ZN(n4579) );
  OR2_X1 U5063 ( .A1(n5973), .A2(n5972), .ZN(n5975) );
  AOI21_X1 U5064 ( .B1(n6226), .B2(n9389), .A(n6295), .ZN(n6227) );
  NOR2_X1 U5065 ( .A1(n9513), .A2(n4397), .ZN(n4396) );
  INV_X1 U5066 ( .A(n4398), .ZN(n4397) );
  NOR2_X1 U5067 ( .A1(n9518), .A2(n9520), .ZN(n4398) );
  INV_X1 U5068 ( .A(n5070), .ZN(n4753) );
  NAND2_X1 U5069 ( .A1(n5300), .A2(SI_14_), .ZN(n4755) );
  NOR2_X1 U5070 ( .A1(n5300), .A2(SI_14_), .ZN(n4754) );
  AOI21_X1 U5071 ( .B1(n7935), .B2(n8357), .A(n8289), .ZN(n4836) );
  INV_X1 U5072 ( .A(n7935), .ZN(n4834) );
  AND2_X1 U5073 ( .A1(n5735), .A2(n6891), .ZN(n5752) );
  OAI21_X1 U5074 ( .B1(n8098), .B2(n4416), .A(n4413), .ZN(n8109) );
  NOR2_X1 U5075 ( .A1(n8094), .A2(n8093), .ZN(n8098) );
  NAND2_X1 U5076 ( .A1(n8099), .A2(n4417), .ZN(n4416) );
  NOR2_X1 U5077 ( .A1(n4415), .A2(n4414), .ZN(n4413) );
  INV_X1 U5078 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6891) );
  NAND2_X1 U5079 ( .A1(n4411), .A2(n4410), .ZN(n7153) );
  NAND2_X1 U5080 ( .A1(n7041), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4410) );
  NAND2_X1 U5081 ( .A1(n4407), .A2(n4406), .ZN(n8466) );
  NAND2_X1 U5082 ( .A1(n8443), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4406) );
  NAND2_X1 U5083 ( .A1(n8445), .A2(n8444), .ZN(n4407) );
  NOR2_X1 U5084 ( .A1(n5801), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5800) );
  AND2_X1 U5085 ( .A1(n4472), .A2(n4305), .ZN(n4468) );
  OR2_X1 U5086 ( .A1(n5777), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U5087 ( .A1(n4449), .A2(n8374), .ZN(n8024) );
  INV_X1 U5088 ( .A(n9856), .ZN(n4449) );
  OR2_X1 U5089 ( .A1(n8377), .A2(n7360), .ZN(n8010) );
  AND3_X1 U5090 ( .A1(n5682), .A2(n5681), .A3(n5680), .ZN(n6860) );
  OR2_X1 U5091 ( .A1(n8353), .A2(n8553), .ZN(n8537) );
  INV_X1 U5092 ( .A(n8769), .ZN(n8179) );
  OR2_X1 U5093 ( .A1(n8848), .A2(n8667), .ZN(n8069) );
  OR2_X1 U5094 ( .A1(n8699), .A2(n8682), .ZN(n8060) );
  OR2_X1 U5095 ( .A1(n8858), .A2(n8668), .ZN(n8650) );
  OR2_X1 U5096 ( .A1(n8871), .A2(n8725), .ZN(n4488) );
  INV_X1 U5097 ( .A(n8042), .ZN(n4619) );
  AND2_X1 U5098 ( .A1(n4847), .A2(n5568), .ZN(n4845) );
  NAND2_X1 U5099 ( .A1(n5882), .A2(n5881), .ZN(n5895) );
  AND2_X1 U5100 ( .A1(n4496), .A2(n4495), .ZN(n6688) );
  NAND2_X1 U5101 ( .A1(n9216), .A2(n7593), .ZN(n4495) );
  NAND2_X1 U5102 ( .A1(n4497), .A2(n9747), .ZN(n4496) );
  NAND2_X1 U5103 ( .A1(n4672), .A2(n7302), .ZN(n4671) );
  INV_X1 U5104 ( .A(n7219), .ZN(n4672) );
  NAND2_X1 U5105 ( .A1(n7481), .A2(n7480), .ZN(n4673) );
  AND2_X1 U5106 ( .A1(n4571), .A2(n9562), .ZN(n4561) );
  NAND2_X1 U5107 ( .A1(n4571), .A2(n4563), .ZN(n4562) );
  INV_X1 U5108 ( .A(n6300), .ZN(n6314) );
  NAND3_X1 U5109 ( .A1(n4799), .A2(n9628), .A3(P1_REG3_REG_1__SCAN_IN), .ZN(
        n4798) );
  NAND2_X1 U5110 ( .A1(n4394), .A2(n9569), .ZN(n4393) );
  NAND2_X1 U5111 ( .A1(n9468), .A2(n6284), .ZN(n4638) );
  OAI21_X1 U5112 ( .B1(n4648), .B2(n4647), .A(n6276), .ZN(n4646) );
  NOR2_X1 U5113 ( .A1(n7622), .A2(n4649), .ZN(n4648) );
  INV_X1 U5114 ( .A(n6114), .ZN(n4649) );
  OAI21_X1 U5115 ( .B1(n6175), .B2(n6174), .A(n6173), .ZN(n6185) );
  INV_X1 U5116 ( .A(n5072), .ZN(n4631) );
  NOR2_X1 U5117 ( .A1(n4372), .A2(n4977), .ZN(n4630) );
  AND2_X1 U5118 ( .A1(n5388), .A2(n5373), .ZN(n5386) );
  AND2_X1 U5119 ( .A1(n5368), .A2(n5357), .ZN(n5366) );
  AOI21_X1 U5120 ( .B1(n5286), .B2(n4302), .A(n4754), .ZN(n5069) );
  OR2_X1 U5121 ( .A1(n4729), .A2(n4926), .ZN(n4280) );
  AOI21_X1 U5122 ( .B1(n4731), .B2(n4922), .A(n4730), .ZN(n4729) );
  XNOR2_X1 U5123 ( .A(n4919), .B(SI_8_), .ZN(n4731) );
  OAI21_X1 U5124 ( .B1(n6348), .B2(n4903), .A(n4902), .ZN(n4906) );
  NAND2_X1 U5125 ( .A1(n6348), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n4902) );
  OAI21_X1 U5126 ( .B1(n4901), .B2(n4886), .A(n4885), .ZN(n4888) );
  NAND2_X1 U5127 ( .A1(n4840), .A2(n4839), .ZN(n4843) );
  INV_X1 U5128 ( .A(n8216), .ZN(n4842) );
  AND2_X1 U5129 ( .A1(n8279), .A2(n8280), .ZN(n7935) );
  INV_X1 U5130 ( .A(n8263), .ZN(n4823) );
  AOI21_X1 U5131 ( .B1(n4827), .B2(n4826), .A(n4289), .ZN(n4825) );
  INV_X1 U5132 ( .A(n4358), .ZN(n4826) );
  INV_X1 U5133 ( .A(n8176), .ZN(n4831) );
  OR2_X1 U5134 ( .A1(n7774), .A2(n7773), .ZN(n7775) );
  XNOR2_X1 U5135 ( .A(n6857), .B(n6860), .ZN(n6952) );
  INV_X1 U5136 ( .A(n4843), .ZN(n7567) );
  XNOR2_X1 U5137 ( .A(n5896), .B(P2_IR_REG_19__SCAN_IN), .ZN(n5989) );
  NAND2_X1 U5138 ( .A1(n5895), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5896) );
  INV_X1 U5139 ( .A(n4848), .ZN(n4846) );
  AND2_X1 U5140 ( .A1(n7114), .A2(n5953), .ZN(n8370) );
  XNOR2_X1 U5141 ( .A(n6603), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n6721) );
  AOI21_X1 U5142 ( .B1(n6658), .B2(P2_REG1_REG_3__SCAN_IN), .A(n4404), .ZN(
        n6595) );
  NOR2_X1 U5143 ( .A1(n4405), .A2(n6668), .ZN(n4404) );
  INV_X1 U5144 ( .A(n6594), .ZN(n4405) );
  OR2_X1 U5145 ( .A1(n6595), .A2(n6596), .ZN(n4403) );
  NAND2_X1 U5146 ( .A1(n4403), .A2(n4402), .ZN(n4401) );
  NAND2_X1 U5147 ( .A1(n6749), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4402) );
  OR2_X1 U5148 ( .A1(n6889), .A2(n6890), .ZN(n4411) );
  XNOR2_X1 U5149 ( .A(n7153), .B(n7044), .ZN(n7039) );
  INV_X1 U5150 ( .A(n7138), .ZN(n4383) );
  NAND2_X1 U5151 ( .A1(n7446), .A2(n7447), .ZN(n7448) );
  NAND2_X1 U5152 ( .A1(n7448), .A2(n7449), .ZN(n7686) );
  OR2_X1 U5153 ( .A1(n7821), .A2(n7820), .ZN(n4710) );
  OR2_X1 U5154 ( .A1(n8413), .A2(n8414), .ZN(n8440) );
  INV_X1 U5155 ( .A(n4691), .ZN(n4690) );
  OAI21_X1 U5156 ( .B1(n4694), .B2(n8494), .A(n4692), .ZN(n4691) );
  NAND2_X1 U5157 ( .A1(n4694), .A2(n4693), .ZN(n4692) );
  NAND2_X1 U5158 ( .A1(n5584), .A2(n5583), .ZN(n5932) );
  NAND2_X1 U5159 ( .A1(n5969), .A2(n4620), .ZN(n7713) );
  INV_X1 U5160 ( .A(n5760), .ZN(n4474) );
  INV_X1 U5161 ( .A(n4473), .ZN(n4472) );
  OAI21_X1 U5162 ( .B1(n5759), .B2(n4274), .A(n4475), .ZN(n4473) );
  OR2_X1 U5163 ( .A1(n8374), .A2(n9856), .ZN(n4475) );
  AND2_X1 U5164 ( .A1(n8034), .A2(n8032), .ZN(n8143) );
  NAND2_X1 U5165 ( .A1(n6971), .A2(n8131), .ZN(n4489) );
  NAND2_X1 U5166 ( .A1(n5948), .A2(n5947), .ZN(n6040) );
  NAND2_X1 U5167 ( .A1(n8586), .A2(n5985), .ZN(n4601) );
  NAND2_X1 U5168 ( .A1(n4477), .A2(n4285), .ZN(n4476) );
  NAND2_X1 U5169 ( .A1(n4329), .A2(n4608), .ZN(n4607) );
  NAND2_X1 U5170 ( .A1(n4278), .A2(n8071), .ZN(n4608) );
  NAND2_X1 U5171 ( .A1(n8649), .A2(n4609), .ZN(n4605) );
  AND2_X1 U5172 ( .A1(n8071), .A2(n5974), .ZN(n4609) );
  CLKBUF_X1 U5173 ( .A(n5989), .Z(n8495) );
  OR2_X1 U5174 ( .A1(n8779), .A2(n8683), .ZN(n8651) );
  NAND2_X1 U5175 ( .A1(n6858), .A2(n8051), .ZN(n9665) );
  OAI21_X1 U5176 ( .B1(n8704), .B2(n4479), .A(n4478), .ZN(n8681) );
  INV_X1 U5177 ( .A(n4480), .ZN(n4479) );
  AOI21_X1 U5178 ( .B1(n4480), .B2(n4482), .A(n8679), .ZN(n4478) );
  AOI21_X1 U5179 ( .B1(n4483), .B2(n5847), .A(n4481), .ZN(n4480) );
  INV_X1 U5180 ( .A(n8726), .ZN(n9663) );
  NAND2_X1 U5181 ( .A1(n8716), .A2(n8717), .ZN(n8704) );
  AND2_X1 U5182 ( .A1(n5747), .A2(n5746), .ZN(n9843) );
  AND3_X1 U5183 ( .A1(n5719), .A2(n5718), .A3(n5717), .ZN(n9832) );
  INV_X1 U5184 ( .A(n6016), .ZN(n6017) );
  XNOR2_X1 U5185 ( .A(n7902), .B(P2_B_REG_SCAN_IN), .ZN(n6015) );
  INV_X1 U5186 ( .A(n5587), .ZN(n5589) );
  INV_X1 U5187 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5588) );
  INV_X1 U5188 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5557) );
  AND2_X1 U5189 ( .A1(n5156), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5214) );
  OR2_X1 U5190 ( .A1(n7589), .A2(n7588), .ZN(n4874) );
  NAND2_X1 U5191 ( .A1(n6686), .A2(n6685), .ZN(n9041) );
  OR2_X1 U5192 ( .A1(n9148), .A2(n4344), .ZN(n4679) );
  INV_X1 U5193 ( .A(n7123), .ZN(n4506) );
  NAND2_X1 U5194 ( .A1(n9041), .A2(n9042), .ZN(n6700) );
  NAND2_X1 U5195 ( .A1(n4513), .A2(n4511), .ZN(n9125) );
  AOI21_X1 U5196 ( .B1(n4277), .B2(n4344), .A(n4512), .ZN(n4511) );
  INV_X1 U5197 ( .A(n9050), .ZN(n4512) );
  OR2_X1 U5198 ( .A1(n5033), .A2(n9996), .ZN(n5344) );
  NAND2_X1 U5199 ( .A1(n8997), .A2(n9761), .ZN(n6531) );
  NOR2_X1 U5200 ( .A1(n4660), .A2(n4664), .ZN(n4659) );
  INV_X1 U5201 ( .A(n9107), .ZN(n4664) );
  INV_X1 U5202 ( .A(n9096), .ZN(n4660) );
  INV_X1 U5203 ( .A(n9106), .ZN(n4662) );
  AND2_X1 U5204 ( .A1(n6481), .A2(n6479), .ZN(n6549) );
  INV_X1 U5205 ( .A(n9180), .ZN(n4507) );
  NAND2_X1 U5206 ( .A1(n4508), .A2(n8917), .ZN(n8920) );
  NAND2_X1 U5207 ( .A1(n4675), .A2(n4678), .ZN(n4508) );
  NOR2_X1 U5208 ( .A1(n4561), .A2(n4555), .ZN(n4554) );
  INV_X1 U5209 ( .A(n4569), .ZN(n4555) );
  NOR2_X1 U5210 ( .A1(n4561), .A2(n4557), .ZN(n4556) );
  INV_X1 U5211 ( .A(n4567), .ZN(n4557) );
  AOI21_X1 U5212 ( .B1(n6160), .B2(n4554), .A(n4550), .ZN(n4549) );
  NAND2_X1 U5213 ( .A1(n4552), .A2(n4551), .ZN(n4550) );
  NAND2_X1 U5214 ( .A1(n4556), .A2(n6166), .ZN(n4551) );
  NAND2_X1 U5215 ( .A1(n4553), .A2(n4562), .ZN(n4552) );
  NOR2_X1 U5216 ( .A1(n6304), .A2(n6303), .ZN(n6307) );
  NAND2_X1 U5217 ( .A1(n6303), .A2(n6168), .ZN(n4534) );
  OR2_X1 U5218 ( .A1(n6161), .A2(n6160), .ZN(n4559) );
  INV_X1 U5219 ( .A(n6166), .ZN(n4464) );
  NOR2_X1 U5220 ( .A1(n4560), .A2(n6301), .ZN(n4466) );
  INV_X1 U5221 ( .A(n4563), .ZN(n4560) );
  AND2_X1 U5222 ( .A1(n6301), .A2(n6310), .ZN(n6197) );
  AND2_X1 U5223 ( .A1(n5011), .A2(n5010), .ZN(n9079) );
  INV_X1 U5224 ( .A(n5141), .ZN(n5051) );
  AND3_X1 U5225 ( .A1(n5040), .A2(n5039), .A3(n5038), .ZN(n9152) );
  AND4_X1 U5226 ( .A1(n5333), .A2(n5332), .A3(n5331), .A4(n5330), .ZN(n9109)
         );
  AND4_X1 U5227 ( .A1(n5298), .A2(n5297), .A3(n5296), .A4(n5295), .ZN(n7863)
         );
  AND4_X1 U5228 ( .A1(n5265), .A2(n5264), .A3(n5263), .A4(n5262), .ZN(n7669)
         );
  AND4_X1 U5229 ( .A1(n5231), .A2(n5230), .A3(n5229), .A4(n5228), .ZN(n7554)
         );
  AOI21_X1 U5230 ( .B1(n9649), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9644), .ZN(
        n9684) );
  NOR2_X1 U5231 ( .A1(n9641), .A2(n4599), .ZN(n9679) );
  AND2_X1 U5232 ( .A1(n9649), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4599) );
  NAND2_X1 U5233 ( .A1(n9244), .A2(n4380), .ZN(n9262) );
  OR2_X1 U5234 ( .A1(n9245), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n4380) );
  INV_X1 U5235 ( .A(n9319), .ZN(n5385) );
  INV_X1 U5236 ( .A(n4629), .ZN(n9334) );
  NOR2_X1 U5237 ( .A1(n9394), .A2(n4793), .ZN(n4792) );
  INV_X1 U5238 ( .A(n4864), .ZN(n4793) );
  OR2_X1 U5239 ( .A1(n9529), .A2(n9200), .ZN(n5536) );
  OR2_X1 U5240 ( .A1(n9419), .A2(n9152), .ZN(n4864) );
  INV_X1 U5241 ( .A(n6247), .ZN(n9394) );
  NAND2_X1 U5242 ( .A1(n4376), .A2(n4375), .ZN(n5316) );
  INV_X1 U5243 ( .A(n7891), .ZN(n4375) );
  INV_X1 U5244 ( .A(n7890), .ZN(n4376) );
  NAND2_X1 U5245 ( .A1(n4640), .A2(n4639), .ZN(n9464) );
  INV_X1 U5246 ( .A(n9468), .ZN(n4639) );
  INV_X1 U5247 ( .A(n9461), .ZN(n4640) );
  NAND2_X1 U5248 ( .A1(n5266), .A2(n4648), .ZN(n4644) );
  OR2_X1 U5249 ( .A1(n7680), .A2(n7669), .ZN(n6114) );
  NAND2_X1 U5250 ( .A1(n6115), .A2(n6273), .ZN(n7622) );
  NAND2_X1 U5251 ( .A1(n7640), .A2(n5528), .ZN(n7623) );
  OR2_X1 U5252 ( .A1(n7680), .A2(n9208), .ZN(n5528) );
  NAND2_X1 U5253 ( .A1(n7017), .A2(n9775), .ZN(n4371) );
  NAND2_X1 U5254 ( .A1(n6918), .A2(n5520), .ZN(n4650) );
  NAND2_X1 U5255 ( .A1(n5445), .A2(n5444), .ZN(n7918) );
  NAND2_X1 U5256 ( .A1(n4760), .A2(n4758), .ZN(n9282) );
  AOI21_X1 U5257 ( .B1(n4761), .B2(n4763), .A(n4759), .ZN(n4758) );
  INV_X1 U5258 ( .A(n9283), .ZN(n4759) );
  AND2_X1 U5259 ( .A1(n5384), .A2(n6216), .ZN(n9339) );
  NAND2_X1 U5260 ( .A1(n4328), .A2(n4788), .ZN(n4783) );
  AND2_X1 U5261 ( .A1(n4788), .A2(n5539), .ZN(n4784) );
  AND2_X1 U5262 ( .A1(n6147), .A2(n9333), .ZN(n9351) );
  NAND2_X1 U5263 ( .A1(n5479), .A2(n9079), .ZN(n5539) );
  AND2_X1 U5264 ( .A1(n9513), .A2(n9198), .ZN(n5538) );
  OR2_X1 U5265 ( .A1(n9434), .A2(n9201), .ZN(n5534) );
  OR2_X1 U5266 ( .A1(n9616), .A2(n9204), .ZN(n5531) );
  AND2_X1 U5267 ( .A1(n5243), .A2(n5242), .ZN(n9792) );
  INV_X1 U5268 ( .A(n9798), .ZN(n9541) );
  XNOR2_X1 U5269 ( .A(n6185), .B(n6184), .ZN(n8889) );
  NAND2_X1 U5270 ( .A1(n4994), .A2(n4651), .ZN(n4996) );
  AOI21_X1 U5271 ( .B1(n4995), .B2(n4315), .A(n4652), .ZN(n4651) );
  NOR2_X1 U5272 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n4652) );
  XNOR2_X1 U5273 ( .A(n5425), .B(n5439), .ZN(n8894) );
  XNOR2_X1 U5274 ( .A(n5423), .B(n5422), .ZN(n8897) );
  XNOR2_X1 U5275 ( .A(n5405), .B(n5404), .ZN(n7907) );
  INV_X1 U5276 ( .A(n4778), .ZN(n5025) );
  XNOR2_X1 U5277 ( .A(n5387), .B(n5386), .ZN(n7899) );
  XNOR2_X1 U5278 ( .A(n5367), .B(n5366), .ZN(n7845) );
  NOR2_X1 U5279 ( .A1(n5001), .A2(n4741), .ZN(n4740) );
  INV_X1 U5280 ( .A(n4961), .ZN(n4741) );
  AOI21_X1 U5281 ( .B1(n4740), .B2(n4962), .A(n4739), .ZN(n4738) );
  INV_X1 U5282 ( .A(n4967), .ZN(n4739) );
  NAND2_X1 U5283 ( .A1(n4960), .A2(n4959), .ZN(n5340) );
  AND3_X1 U5284 ( .A1(n5457), .A2(n5456), .A3(n4505), .ZN(n5462) );
  NAND2_X1 U5285 ( .A1(n4747), .A2(n4953), .ZN(n5024) );
  NAND2_X1 U5286 ( .A1(n4951), .A2(n4748), .ZN(n4747) );
  NAND2_X1 U5287 ( .A1(n4951), .A2(n4950), .ZN(n5043) );
  INV_X1 U5288 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5457) );
  NAND2_X1 U5289 ( .A1(n4456), .A2(n4946), .ZN(n5058) );
  NAND2_X1 U5290 ( .A1(n5286), .A2(n4945), .ZN(n5299) );
  NAND2_X1 U5291 ( .A1(n4461), .A2(n4460), .ZN(n5253) );
  NAND2_X1 U5292 ( .A1(n4728), .A2(n4280), .ZN(n5233) );
  NAND2_X1 U5293 ( .A1(n5189), .A2(n4279), .ZN(n4728) );
  XNOR2_X1 U5294 ( .A(n4412), .B(n5219), .ZN(n6384) );
  OAI21_X1 U5295 ( .B1(n5189), .B2(n4731), .A(n4922), .ZN(n4412) );
  AND4_X1 U5296 ( .A1(n5794), .A2(n5793), .A3(n5792), .A4(n5791), .ZN(n7795)
         );
  NOR2_X1 U5297 ( .A1(n4282), .A2(n8356), .ZN(n4811) );
  NAND2_X1 U5298 ( .A1(n8206), .A2(n8204), .ZN(n4818) );
  NAND2_X1 U5299 ( .A1(n4814), .A2(n4322), .ZN(n4813) );
  NAND2_X1 U5300 ( .A1(n5811), .A2(n5810), .ZN(n9654) );
  INV_X1 U5301 ( .A(n8380), .ZN(n7241) );
  AND2_X1 U5302 ( .A1(n5609), .A2(n5608), .ZN(n8350) );
  NAND2_X1 U5303 ( .A1(n6773), .A2(n9656), .ZN(n8352) );
  OR2_X1 U5304 ( .A1(n7443), .A2(n7442), .ZN(n4696) );
  NOR2_X1 U5305 ( .A1(n8463), .A2(n8462), .ZN(n8465) );
  AND2_X1 U5306 ( .A1(n8461), .A2(n8441), .ZN(n8462) );
  AND2_X1 U5307 ( .A1(n6589), .A2(n8474), .ZN(n8516) );
  NAND2_X1 U5308 ( .A1(n5799), .A2(n5798), .ZN(n9871) );
  NAND2_X1 U5309 ( .A1(n5776), .A2(n5775), .ZN(n9860) );
  INV_X1 U5310 ( .A(n8785), .ZN(n8789) );
  INV_X1 U5311 ( .A(n6040), .ZN(n8529) );
  NOR2_X1 U5312 ( .A1(n8535), .A2(n9852), .ZN(n6004) );
  INV_X1 U5313 ( .A(n8095), .ZN(n8806) );
  NAND2_X1 U5314 ( .A1(n5630), .A2(n5629), .ZN(n5984) );
  NOR2_X1 U5315 ( .A1(n4273), .A2(n4532), .ZN(n4525) );
  AND2_X1 U5316 ( .A1(n4593), .A2(n4592), .ZN(n6453) );
  NAND2_X1 U5317 ( .A1(n6451), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4592) );
  XNOR2_X1 U5318 ( .A(n9259), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n4591) );
  OAI21_X1 U5319 ( .B1(n4591), .B2(n9730), .A(n4589), .ZN(n4588) );
  NAND2_X1 U5320 ( .A1(n9267), .A2(n9733), .ZN(n4589) );
  NAND2_X1 U5321 ( .A1(n5275), .A2(n5274), .ZN(n7629) );
  NAND2_X1 U5322 ( .A1(n6480), .A2(n6479), .ZN(n6989) );
  AOI21_X1 U5323 ( .B1(n8882), .B2(n6191), .A(n4866), .ZN(n9558) );
  NAND2_X1 U5324 ( .A1(n4387), .A2(n9521), .ZN(n9482) );
  XNOR2_X1 U5325 ( .A(n9274), .B(n9558), .ZN(n4387) );
  OR2_X1 U5326 ( .A1(n9293), .A2(n9299), .ZN(n6068) );
  NAND2_X1 U5327 ( .A1(n4504), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n4503) );
  NAND2_X1 U5328 ( .A1(n5059), .A2(n4286), .ZN(n4501) );
  OR2_X1 U5329 ( .A1(n5059), .A2(n4505), .ZN(n4502) );
  NAND2_X1 U5330 ( .A1(n7016), .A2(n4536), .ZN(n4535) );
  NAND2_X1 U5331 ( .A1(n4539), .A2(n4538), .ZN(n4537) );
  AND2_X1 U5332 ( .A1(n6084), .A2(n6310), .ZN(n4536) );
  NAND2_X1 U5333 ( .A1(n4448), .A2(n4447), .ZN(n8017) );
  NAND2_X1 U5334 ( .A1(n8021), .A2(n8110), .ZN(n4447) );
  NAND2_X1 U5335 ( .A1(n8058), .A2(n8063), .ZN(n4435) );
  NOR2_X1 U5336 ( .A1(n4436), .A2(n8049), .ZN(n4434) );
  NAND2_X1 U5337 ( .A1(n4517), .A2(n6131), .ZN(n4516) );
  NAND2_X1 U5338 ( .A1(n6127), .A2(n6168), .ZN(n4517) );
  AOI21_X1 U5339 ( .B1(n4515), .B2(n4310), .A(n6310), .ZN(n4519) );
  INV_X1 U5340 ( .A(n6127), .ZN(n4515) );
  OAI21_X1 U5341 ( .B1(n4422), .B2(n8062), .A(n8066), .ZN(n4421) );
  AOI21_X1 U5342 ( .B1(n8061), .B2(n8060), .A(n8151), .ZN(n4422) );
  NOR2_X1 U5343 ( .A1(n4427), .A2(n4426), .ZN(n4425) );
  NAND2_X1 U5344 ( .A1(n8066), .A2(n8067), .ZN(n4426) );
  NOR2_X1 U5345 ( .A1(n8068), .A2(n8130), .ZN(n4427) );
  OAI21_X1 U5346 ( .B1(n4423), .B2(n8051), .A(n4420), .ZN(n4419) );
  NOR2_X1 U5347 ( .A1(n4425), .A2(n4424), .ZN(n4423) );
  AOI21_X1 U5348 ( .B1(n4421), .B2(n8051), .A(n8073), .ZN(n4420) );
  NAND2_X1 U5349 ( .A1(n8069), .A2(n8621), .ZN(n4424) );
  NAND2_X1 U5350 ( .A1(n6142), .A2(n6143), .ZN(n4545) );
  NAND2_X1 U5351 ( .A1(n6141), .A2(n6168), .ZN(n4544) );
  NAND2_X1 U5352 ( .A1(n6140), .A2(n6310), .ZN(n4546) );
  INV_X1 U5353 ( .A(n6146), .ZN(n4542) );
  NOR2_X1 U5354 ( .A1(n6209), .A2(n6208), .ZN(n6222) );
  INV_X1 U5355 ( .A(n8104), .ZN(n4415) );
  MUX2_X1 U5356 ( .A(n8163), .B(n8162), .S(n8110), .Z(n8104) );
  NOR2_X1 U5357 ( .A1(n4418), .A2(n4288), .ZN(n4414) );
  NAND2_X1 U5358 ( .A1(n8096), .A2(n8097), .ZN(n4417) );
  AOI211_X1 U5359 ( .C1(n8083), .C2(n4284), .A(n4437), .B(n4442), .ZN(n8094)
         );
  NAND2_X1 U5360 ( .A1(n4444), .A2(n4443), .ZN(n4442) );
  NOR2_X1 U5361 ( .A1(n4439), .A2(n4438), .ZN(n4437) );
  NOR2_X1 U5362 ( .A1(n4848), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n4847) );
  INV_X1 U5363 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4453) );
  AND2_X1 U5364 ( .A1(n6165), .A2(n6158), .ZN(n6223) );
  OR2_X1 U5365 ( .A1(n6152), .A2(n4309), .ZN(n4574) );
  INV_X1 U5366 ( .A(n4573), .ZN(n4572) );
  NOR2_X1 U5367 ( .A1(n6155), .A2(n4582), .ZN(n4581) );
  AOI21_X1 U5368 ( .B1(n4580), .B2(n4578), .A(n4577), .ZN(n4576) );
  INV_X1 U5369 ( .A(n6268), .ZN(n6112) );
  AND2_X1 U5370 ( .A1(n4463), .A2(n4462), .ZN(n6208) );
  AND2_X1 U5371 ( .A1(n9194), .A2(n4356), .ZN(n4462) );
  AOI21_X1 U5372 ( .B1(n5442), .B2(n5441), .A(n4875), .ZN(n6169) );
  INV_X1 U5373 ( .A(n4740), .ZN(n4736) );
  INV_X1 U5374 ( .A(n5349), .ZN(n4735) );
  INV_X1 U5375 ( .A(n4457), .ZN(n4370) );
  INV_X1 U5376 ( .A(n4455), .ZN(n4369) );
  INV_X1 U5377 ( .A(n4953), .ZN(n4746) );
  INV_X1 U5378 ( .A(n4748), .ZN(n4744) );
  NAND2_X1 U5379 ( .A1(n4955), .A2(n4954), .ZN(n4958) );
  INV_X1 U5380 ( .A(SI_19_), .ZN(n4954) );
  INV_X1 U5381 ( .A(n5057), .ZN(n4458) );
  INV_X1 U5382 ( .A(n8121), .ZN(n8123) );
  NAND2_X1 U5383 ( .A1(n5567), .A2(n4849), .ZN(n4848) );
  INV_X1 U5384 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4849) );
  NAND2_X1 U5385 ( .A1(n4708), .A2(n6668), .ZN(n4707) );
  NAND2_X1 U5386 ( .A1(n4707), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4706) );
  INV_X1 U5387 ( .A(n6756), .ZN(n4702) );
  AND2_X1 U5388 ( .A1(n4699), .A2(n4340), .ZN(n4698) );
  OAI22_X1 U5389 ( .A1(n4698), .A2(n6813), .B1(n4697), .B2(n6756), .ZN(n6893)
         );
  NAND2_X1 U5390 ( .A1(n4276), .A2(n4703), .ZN(n4697) );
  NAND2_X1 U5391 ( .A1(n7341), .A2(n7342), .ZN(n7444) );
  NAND2_X1 U5392 ( .A1(n7686), .A2(n4357), .ZN(n7822) );
  NAND2_X1 U5393 ( .A1(n8464), .A2(n8493), .ZN(n4693) );
  NAND2_X1 U5394 ( .A1(n4281), .A2(n4316), .ZN(n4624) );
  AND2_X1 U5395 ( .A1(n5613), .A2(n5580), .ZN(n5612) );
  NOR2_X1 U5396 ( .A1(n5903), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5613) );
  NOR2_X1 U5397 ( .A1(n5841), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5840) );
  INV_X1 U5398 ( .A(n6932), .ZN(n7983) );
  CLKBUF_X1 U5399 ( .A(n6855), .Z(n7977) );
  NAND2_X1 U5400 ( .A1(n8383), .A2(n6941), .ZN(n7979) );
  INV_X1 U5401 ( .A(n5978), .ZN(n7973) );
  NAND2_X1 U5402 ( .A1(n8179), .A2(n8643), .ZN(n5978) );
  INV_X1 U5403 ( .A(n8678), .ZN(n4481) );
  INV_X1 U5404 ( .A(n4483), .ZN(n4482) );
  NAND2_X1 U5405 ( .A1(n4487), .A2(n4486), .ZN(n4485) );
  INV_X1 U5406 ( .A(n8704), .ZN(n4487) );
  NOR2_X1 U5407 ( .A1(n8690), .A2(n4484), .ZN(n4483) );
  INV_X1 U5408 ( .A(n4488), .ZN(n4484) );
  OR2_X1 U5409 ( .A1(n6945), .A2(n7499), .ZN(n6848) );
  INV_X1 U5410 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6032) );
  INV_X1 U5411 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5878) );
  INV_X1 U5412 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5808) );
  INV_X1 U5413 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5561) );
  INV_X1 U5414 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5848) );
  INV_X1 U5415 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5785) );
  INV_X1 U5416 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5556) );
  NOR2_X1 U5417 ( .A1(n5727), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5744) );
  OR2_X1 U5418 ( .A1(n5691), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5727) );
  OR2_X1 U5419 ( .A1(n8959), .A2(n9077), .ZN(n9022) );
  AND2_X1 U5420 ( .A1(n5138), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5156) );
  INV_X1 U5421 ( .A(n9058), .ZN(n8997) );
  INV_X1 U5422 ( .A(n4561), .ZN(n4553) );
  AOI21_X1 U5423 ( .B1(n6230), .B2(n6301), .A(n6229), .ZN(n4366) );
  OR2_X1 U5424 ( .A1(n6228), .A2(n6227), .ZN(n4367) );
  AND2_X1 U5425 ( .A1(n9558), .A2(n9271), .ZN(n6300) );
  NAND2_X1 U5426 ( .A1(n6164), .A2(n6163), .ZN(n6166) );
  NAND2_X1 U5427 ( .A1(n6207), .A2(n6168), .ZN(n4565) );
  NAND2_X1 U5428 ( .A1(n6229), .A2(n6310), .ZN(n4564) );
  AOI21_X1 U5429 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9714), .A(n9709), .ZN(
        n9221) );
  AND2_X1 U5430 ( .A1(n5414), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5448) );
  NOR2_X1 U5431 ( .A1(n7918), .A2(n9065), .ZN(n6207) );
  NOR2_X1 U5432 ( .A1(n9289), .A2(n4393), .ZN(n4392) );
  AND2_X1 U5433 ( .A1(n5376), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5396) );
  AND2_X1 U5434 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n5361), .ZN(n5376) );
  INV_X1 U5435 ( .A(n9424), .ZN(n4634) );
  INV_X1 U5436 ( .A(n6284), .ZN(n4635) );
  NAND2_X1 U5437 ( .A1(n7175), .A2(n4656), .ZN(n4655) );
  NOR2_X1 U5438 ( .A1(n6239), .A2(n4657), .ZN(n4656) );
  NAND2_X1 U5439 ( .A1(n5251), .A2(n6240), .ZN(n4377) );
  AND2_X1 U5440 ( .A1(n6112), .A2(n6110), .ZN(n5527) );
  NAND2_X1 U5441 ( .A1(n9217), .A2(n9775), .ZN(n6263) );
  NAND2_X1 U5442 ( .A1(n7055), .A2(n9216), .ZN(n6265) );
  INV_X1 U5443 ( .A(n6206), .ZN(n6164) );
  NAND2_X1 U5444 ( .A1(n9289), .A2(n9057), .ZN(n6165) );
  INV_X1 U5445 ( .A(n6208), .ZN(n6154) );
  AND2_X1 U5446 ( .A1(n9414), .A2(n4291), .ZN(n9356) );
  NAND2_X1 U5447 ( .A1(n9414), .A2(n4396), .ZN(n9369) );
  INV_X1 U5448 ( .A(n5536), .ZN(n4790) );
  NAND2_X1 U5449 ( .A1(n9414), .A2(n9401), .ZN(n9396) );
  NAND2_X1 U5450 ( .A1(n9431), .A2(n9605), .ZN(n9432) );
  NAND2_X1 U5451 ( .A1(n7641), .A2(n7643), .ZN(n7640) );
  NAND2_X1 U5452 ( .A1(n5518), .A2(n7051), .ZN(n5519) );
  NAND2_X1 U5453 ( .A1(n6263), .A2(n5520), .ZN(n6921) );
  XNOR2_X1 U5454 ( .A(n6169), .B(n6170), .ZN(n6175) );
  AND2_X1 U5455 ( .A1(n5437), .A2(n5411), .ZN(n5422) );
  AND2_X1 U5456 ( .A1(n5406), .A2(n5394), .ZN(n5404) );
  INV_X1 U5457 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4979) );
  INV_X1 U5458 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5487) );
  XNOR2_X1 U5459 ( .A(n5509), .B(P1_IR_REG_23__SCAN_IN), .ZN(n6305) );
  INV_X1 U5460 ( .A(SI_20_), .ZN(n5013) );
  NOR2_X1 U5461 ( .A1(n5041), .A2(n4749), .ZN(n4748) );
  INV_X1 U5462 ( .A(n4950), .ZN(n4749) );
  NAND2_X1 U5463 ( .A1(n4947), .A2(n10038), .ZN(n4950) );
  NAND2_X1 U5464 ( .A1(n4456), .A2(n4343), .ZN(n4951) );
  NAND2_X1 U5465 ( .A1(n4295), .A2(n4457), .ZN(n4456) );
  OAI21_X1 U5466 ( .B1(n4754), .B2(n4752), .A(n4753), .ZN(n4751) );
  INV_X1 U5467 ( .A(SI_15_), .ZN(n4752) );
  NAND2_X1 U5468 ( .A1(n4941), .A2(SI_13_), .ZN(n4945) );
  INV_X1 U5469 ( .A(n8227), .ZN(n4819) );
  NOR2_X1 U5470 ( .A1(n5964), .A2(n6886), .ZN(n6855) );
  AOI21_X1 U5471 ( .B1(n4836), .B2(n4834), .A(n4833), .ZN(n4832) );
  INV_X1 U5472 ( .A(n4836), .ZN(n4835) );
  INV_X1 U5473 ( .A(n8288), .ZN(n4833) );
  XNOR2_X1 U5474 ( .A(n6857), .B(n7228), .ZN(n7059) );
  NAND2_X1 U5475 ( .A1(n5752), .A2(n5577), .ZN(n5777) );
  AND2_X1 U5476 ( .A1(n6050), .A2(n6049), .ZN(n6786) );
  INV_X1 U5477 ( .A(n8341), .ZN(n8361) );
  NAND2_X1 U5478 ( .A1(n8107), .A2(n8110), .ZN(n4430) );
  NOR2_X1 U5479 ( .A1(n8106), .A2(n8122), .ZN(n8107) );
  NAND2_X1 U5480 ( .A1(n8111), .A2(n8051), .ZN(n8112) );
  AND2_X1 U5481 ( .A1(n5637), .A2(n5636), .ZN(n8326) );
  AOI22_X1 U5482 ( .A1(n6592), .A2(n6591), .B1(n6593), .B2(n6590), .ZN(n4400)
         );
  OAI22_X1 U5483 ( .A1(n4400), .A2(n6645), .B1(n6593), .B2(n6466), .ZN(n6716)
         );
  NAND2_X1 U5484 ( .A1(n4707), .A2(n6609), .ZN(n6662) );
  CLKBUF_X1 U5485 ( .A(n5690), .Z(n5691) );
  NAND2_X1 U5486 ( .A1(n6606), .A2(n6605), .ZN(n6609) );
  NAND2_X1 U5487 ( .A1(n4705), .A2(n6609), .ZN(n6660) );
  INV_X1 U5488 ( .A(n4706), .ZN(n4705) );
  NAND2_X1 U5489 ( .A1(n4702), .A2(n4276), .ZN(n4701) );
  NAND2_X1 U5490 ( .A1(n4700), .A2(n4704), .ZN(n4699) );
  INV_X1 U5491 ( .A(n6830), .ZN(n4700) );
  NAND2_X1 U5492 ( .A1(n6755), .A2(n6754), .ZN(n6830) );
  NAND2_X1 U5493 ( .A1(n4702), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6832) );
  INV_X1 U5494 ( .A(n4401), .ZN(n6791) );
  OR2_X1 U5495 ( .A1(n5748), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5761) );
  NAND2_X1 U5496 ( .A1(n7155), .A2(n7156), .ZN(n7157) );
  NAND2_X1 U5497 ( .A1(n7157), .A2(n7158), .ZN(n7341) );
  XNOR2_X1 U5498 ( .A(n7444), .B(n7438), .ZN(n7343) );
  NAND2_X1 U5499 ( .A1(n7340), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4711) );
  XNOR2_X1 U5500 ( .A(n7822), .B(n7816), .ZN(n7688) );
  NAND2_X1 U5501 ( .A1(n7684), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4695) );
  NAND2_X1 U5502 ( .A1(n8385), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4709) );
  NAND2_X1 U5503 ( .A1(n8417), .A2(n8418), .ZN(n8445) );
  XNOR2_X1 U5504 ( .A(n8466), .B(n8470), .ZN(n8446) );
  NAND2_X1 U5505 ( .A1(n8440), .A2(n8439), .ZN(n8461) );
  OR2_X1 U5506 ( .A1(n5603), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8522) );
  XNOR2_X1 U5507 ( .A(n5954), .B(n8099), .ZN(n5963) );
  NAND2_X1 U5508 ( .A1(n8806), .A2(n5943), .ZN(n5944) );
  OR2_X1 U5509 ( .A1(n5631), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U5510 ( .A1(n5612), .A2(n5581), .ZN(n5624) );
  OR2_X1 U5511 ( .A1(n5624), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5631) );
  OR2_X1 U5512 ( .A1(n5886), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5903) );
  AND4_X1 U5513 ( .A1(n5874), .A2(n5873), .A3(n5872), .A4(n5871), .ZN(n8668)
         );
  NAND2_X1 U5514 ( .A1(n5800), .A2(n5578), .ZN(n5829) );
  AND4_X1 U5515 ( .A1(n5782), .A2(n5781), .A3(n5780), .A4(n5779), .ZN(n8310)
         );
  NAND2_X1 U5516 ( .A1(n4467), .A2(n4469), .ZN(n7706) );
  AOI21_X1 U5517 ( .B1(n4472), .B2(n4471), .A(n4470), .ZN(n4469) );
  INV_X1 U5518 ( .A(n7797), .ZN(n4470) );
  INV_X1 U5519 ( .A(n7798), .ZN(n8145) );
  AND2_X1 U5520 ( .A1(n8024), .A2(n8022), .ZN(n8142) );
  NAND2_X1 U5521 ( .A1(n7411), .A2(n5760), .ZN(n7608) );
  AND2_X1 U5522 ( .A1(n8016), .A2(n8021), .ZN(n8141) );
  NAND2_X1 U5523 ( .A1(n7467), .A2(n5759), .ZN(n7411) );
  AND4_X1 U5524 ( .A1(n5758), .A2(n5757), .A3(n5756), .A4(n5755), .ZN(n8313)
         );
  AND3_X1 U5525 ( .A1(n5731), .A2(n5730), .A3(n5729), .ZN(n7360) );
  OR2_X1 U5526 ( .A1(n5721), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5736) );
  OR2_X1 U5527 ( .A1(n6880), .A2(n5990), .ZN(n7612) );
  AND2_X1 U5528 ( .A1(n6045), .A2(n6033), .ZN(n6877) );
  AND2_X1 U5529 ( .A1(n6035), .A2(n8110), .ZN(n6874) );
  INV_X1 U5530 ( .A(n8544), .ZN(n4494) );
  OR2_X1 U5531 ( .A1(n8604), .A2(n5638), .ZN(n8576) );
  OR2_X1 U5532 ( .A1(n8607), .A2(n8611), .ZN(n8604) );
  AND2_X1 U5533 ( .A1(n5983), .A2(n8585), .ZN(n8596) );
  NAND2_X1 U5534 ( .A1(n4859), .A2(n8156), .ZN(n8606) );
  INV_X1 U5535 ( .A(n5979), .ZN(n8621) );
  NAND2_X1 U5536 ( .A1(n5978), .A2(n7972), .ZN(n8625) );
  AND2_X1 U5537 ( .A1(n5611), .A2(n5610), .ZN(n7943) );
  OR2_X1 U5538 ( .A1(n8575), .A2(n8639), .ZN(n8640) );
  AND2_X1 U5539 ( .A1(n8621), .A2(n8622), .ZN(n8639) );
  AOI21_X1 U5540 ( .B1(n8676), .B2(n5974), .A(n4278), .ZN(n4606) );
  AND2_X1 U5541 ( .A1(n8069), .A2(n8066), .ZN(n8653) );
  AND2_X1 U5542 ( .A1(n8651), .A2(n8067), .ZN(n8664) );
  AND4_X1 U5543 ( .A1(n5865), .A2(n5864), .A3(n5863), .A4(n5862), .ZN(n8682)
         );
  NAND2_X1 U5544 ( .A1(n4485), .A2(n4488), .ZN(n8691) );
  NAND2_X1 U5545 ( .A1(n4485), .A2(n4483), .ZN(n8693) );
  INV_X1 U5546 ( .A(n8149), .ZN(n8690) );
  AND2_X1 U5547 ( .A1(n6766), .A2(n8051), .ZN(n8726) );
  INV_X1 U5548 ( .A(n4618), .ZN(n4617) );
  AOI21_X1 U5549 ( .B1(n4621), .B2(n4618), .A(n8047), .ZN(n4616) );
  NOR2_X1 U5550 ( .A1(n8046), .A2(n4619), .ZN(n4618) );
  NAND2_X1 U5551 ( .A1(n5828), .A2(n5827), .ZN(n8793) );
  AND3_X1 U5552 ( .A1(n5707), .A2(n5706), .A3(n5705), .ZN(n9827) );
  OR2_X1 U5553 ( .A1(n6852), .A2(n8110), .ZN(n6783) );
  INV_X1 U5554 ( .A(n9842), .ZN(n9872) );
  NAND2_X1 U5555 ( .A1(n6777), .A2(n6393), .ZN(n6784) );
  XNOR2_X1 U5556 ( .A(n6031), .B(n6032), .ZN(n6776) );
  NAND2_X1 U5557 ( .A1(n8884), .A2(n4714), .ZN(n4713) );
  NAND2_X1 U5558 ( .A1(n5678), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n4715) );
  INV_X1 U5559 ( .A(n6305), .ZN(n6328) );
  INV_X1 U5560 ( .A(n5448), .ZN(n5430) );
  NAND2_X1 U5561 ( .A1(n4682), .A2(n4681), .ZN(n4680) );
  OAI211_X1 U5562 ( .C1(n7595), .C2(n4327), .A(n4498), .B(n7758), .ZN(n7760)
         );
  INV_X1 U5563 ( .A(n7594), .ZN(n4499) );
  NAND2_X1 U5564 ( .A1(n9094), .A2(n9096), .ZN(n9095) );
  INV_X1 U5565 ( .A(n4673), .ZN(n4668) );
  NAND2_X1 U5566 ( .A1(n7302), .A2(n4673), .ZN(n4669) );
  AND2_X1 U5567 ( .A1(n7482), .A2(n4671), .ZN(n4670) );
  AND2_X1 U5568 ( .A1(n6366), .A2(n6549), .ZN(n9129) );
  INV_X1 U5569 ( .A(n8969), .ZN(n9135) );
  INV_X1 U5570 ( .A(n9129), .ZN(n9167) );
  NAND2_X1 U5571 ( .A1(n7218), .A2(n7219), .ZN(n7303) );
  NAND2_X1 U5572 ( .A1(n4675), .A2(n4509), .ZN(n4510) );
  AND2_X1 U5573 ( .A1(n4678), .A2(n8918), .ZN(n4509) );
  AND4_X1 U5574 ( .A1(n5383), .A2(n5382), .A3(n5381), .A4(n5380), .ZN(n9170)
         );
  AOI21_X1 U5575 ( .B1(n9357), .B2(n5051), .A(n5000), .ZN(n9137) );
  NOR2_X1 U5576 ( .A1(n5068), .A2(n5067), .ZN(n9154) );
  AND4_X1 U5577 ( .A1(n5085), .A2(n5084), .A3(n5083), .A4(n5082), .ZN(n9098)
         );
  AND4_X1 U5578 ( .A1(n5218), .A2(n5217), .A3(n5216), .A4(n5215), .ZN(n7298)
         );
  AND4_X1 U5579 ( .A1(n5188), .A2(n5187), .A3(n5186), .A4(n5185), .ZN(n7211)
         );
  AND4_X1 U5580 ( .A1(n5164), .A2(n5163), .A3(n5162), .A4(n5161), .ZN(n7196)
         );
  AND4_X2 U5581 ( .A1(n5111), .A2(n5110), .A3(n5109), .A4(n5108), .ZN(n7017)
         );
  INV_X1 U5582 ( .A(n4797), .ZN(n4796) );
  OAI21_X1 U5583 ( .B1(n5035), .B2(n6326), .A(n4798), .ZN(n4797) );
  OR2_X1 U5584 ( .A1(n6426), .A2(n6425), .ZN(n4595) );
  OR2_X1 U5585 ( .A1(n6413), .A2(n6412), .ZN(n4593) );
  AOI21_X1 U5586 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n6739), .A(n6730), .ZN(
        n6731) );
  NOR2_X1 U5587 ( .A1(n9679), .A2(n9680), .ZN(n9678) );
  NOR2_X1 U5588 ( .A1(n9706), .A2(n4596), .ZN(n9234) );
  AND2_X1 U5589 ( .A1(n9714), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4596) );
  AOI21_X1 U5590 ( .B1(n9262), .B2(n9261), .A(n4379), .ZN(n9736) );
  AND2_X1 U5591 ( .A1(n9260), .A2(n9542), .ZN(n4379) );
  NAND2_X1 U5592 ( .A1(n4583), .A2(n9255), .ZN(n9732) );
  NAND2_X1 U5593 ( .A1(n9254), .A2(n9253), .ZN(n4583) );
  NAND2_X1 U5594 ( .A1(n9631), .A2(n6549), .ZN(n9169) );
  NOR2_X1 U5595 ( .A1(n6061), .A2(n5421), .ZN(n9279) );
  AOI21_X1 U5596 ( .B1(n6062), .B2(n6156), .A(n6251), .ZN(n6061) );
  NAND2_X1 U5597 ( .A1(n9304), .A2(n9303), .ZN(n6062) );
  INV_X1 U5598 ( .A(n4393), .ZN(n4391) );
  NAND2_X1 U5599 ( .A1(n9325), .A2(n9569), .ZN(n9312) );
  NAND2_X1 U5600 ( .A1(n7907), .A2(n6191), .ZN(n4463) );
  INV_X1 U5601 ( .A(n5360), .ZN(n5361) );
  OR2_X1 U5602 ( .A1(n9434), .A2(n9110), .ZN(n9407) );
  INV_X1 U5603 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9101) );
  NAND2_X1 U5604 ( .A1(n5309), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5327) );
  AOI21_X1 U5605 ( .B1(n4645), .B2(n4647), .A(n4642), .ZN(n4641) );
  INV_X1 U5606 ( .A(n6272), .ZN(n4642) );
  AND2_X1 U5607 ( .A1(n5293), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5309) );
  INV_X1 U5608 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5277) );
  NOR2_X1 U5609 ( .A1(n5278), .A2(n5277), .ZN(n5293) );
  INV_X1 U5610 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5259) );
  OR2_X1 U5611 ( .A1(n5260), .A2(n5259), .ZN(n5278) );
  INV_X1 U5612 ( .A(n4655), .ZN(n7420) );
  INV_X1 U5613 ( .A(n4377), .ZN(n7419) );
  INV_X1 U5614 ( .A(n5527), .ZN(n7427) );
  OR2_X1 U5615 ( .A1(n7564), .A2(n9210), .ZN(n5526) );
  NOR2_X1 U5616 ( .A1(n5224), .A2(n4989), .ZN(n5245) );
  AND2_X1 U5617 ( .A1(n6093), .A2(n7325), .ZN(n7324) );
  NOR2_X1 U5618 ( .A1(n7077), .A2(n7131), .ZN(n7191) );
  NAND2_X1 U5619 ( .A1(n7020), .A2(n7092), .ZN(n7077) );
  AND2_X1 U5620 ( .A1(n7071), .A2(n6262), .ZN(n6983) );
  NAND2_X1 U5621 ( .A1(n7014), .A2(n7015), .ZN(n7013) );
  AND2_X1 U5622 ( .A1(n7022), .A2(n7055), .ZN(n7020) );
  AOI21_X1 U5623 ( .B1(n6378), .B2(n5515), .A(n6380), .ZN(n6520) );
  AOI21_X1 U5624 ( .B1(n4764), .B2(n4762), .A(n4323), .ZN(n4761) );
  INV_X1 U5625 ( .A(n5542), .ZN(n4762) );
  INV_X1 U5626 ( .A(n4764), .ZN(n4763) );
  NAND2_X1 U5627 ( .A1(n6164), .A2(n6165), .ZN(n9283) );
  NAND2_X1 U5628 ( .A1(n5375), .A2(n5374), .ZN(n9500) );
  AND2_X1 U5629 ( .A1(n4784), .A2(n5540), .ZN(n4782) );
  OAI21_X1 U5630 ( .B1(n4783), .B2(n4781), .A(n4351), .ZN(n4780) );
  INV_X1 U5631 ( .A(n5540), .ZN(n4781) );
  AND2_X1 U5632 ( .A1(n6625), .A2(n7551), .ZN(n9521) );
  AND2_X1 U5633 ( .A1(n6136), .A2(n6293), .ZN(n9409) );
  AND2_X1 U5634 ( .A1(n9407), .A2(n6135), .ZN(n9423) );
  OAI21_X1 U5635 ( .B1(n7783), .B2(n4769), .A(n4768), .ZN(n4767) );
  NAND2_X1 U5636 ( .A1(n9468), .A2(n4775), .ZN(n4769) );
  NOR2_X1 U5637 ( .A1(n4283), .A2(n5532), .ZN(n4768) );
  AND2_X1 U5638 ( .A1(n6120), .A2(n6278), .ZN(n7784) );
  OR2_X1 U5639 ( .A1(n7629), .A2(n9207), .ZN(n5529) );
  NAND2_X1 U5640 ( .A1(n5197), .A2(n5196), .ZN(n7484) );
  NAND2_X1 U5641 ( .A1(n7269), .A2(n7268), .ZN(n7267) );
  INV_X1 U5642 ( .A(n6983), .ZN(n6987) );
  NAND2_X1 U5643 ( .A1(n6988), .A2(n6987), .ZN(n6986) );
  XNOR2_X1 U5644 ( .A(n6175), .B(SI_29_), .ZN(n5946) );
  XNOR2_X1 U5645 ( .A(n5492), .B(n4522), .ZN(n5510) );
  NAND2_X1 U5646 ( .A1(n4778), .A2(n4777), .ZN(n5491) );
  AND2_X1 U5647 ( .A1(n5458), .A2(n5459), .ZN(n4684) );
  OAI21_X1 U5648 ( .B1(n5340), .B2(n4962), .A(n4961), .ZN(n5002) );
  NAND2_X1 U5649 ( .A1(n5027), .A2(n5026), .ZN(n4504) );
  NAND2_X1 U5650 ( .A1(n5025), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5321) );
  INV_X1 U5651 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9928) );
  INV_X1 U5652 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5193) );
  XNOR2_X1 U5653 ( .A(n5189), .B(n4731), .ZN(n6372) );
  INV_X1 U5654 ( .A(n4913), .ZN(n4722) );
  NAND2_X1 U5655 ( .A1(n5174), .A2(n4868), .ZN(n5176) );
  NAND2_X1 U5656 ( .A1(n5165), .A2(n4870), .ZN(n5167) );
  CLKBUF_X1 U5657 ( .A(n5072), .Z(n5073) );
  NOR2_X2 U5658 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5112) );
  OAI21_X1 U5659 ( .B1(n5089), .B2(n4718), .A(n4884), .ZN(n5114) );
  AND2_X1 U5660 ( .A1(n4889), .A2(n4890), .ZN(n5113) );
  NAND2_X1 U5661 ( .A1(n4717), .A2(n4884), .ZN(n4719) );
  INV_X1 U5662 ( .A(n4718), .ZN(n4717) );
  XNOR2_X1 U5663 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput27), .ZN(n10026) );
  NAND2_X1 U5664 ( .A1(n4843), .A2(n4841), .ZN(n8215) );
  AND2_X1 U5665 ( .A1(n5647), .A2(n5646), .ZN(n8251) );
  AOI21_X1 U5666 ( .B1(n4841), .B2(n7365), .A(n4320), .ZN(n4838) );
  NAND2_X1 U5667 ( .A1(n4821), .A2(n4825), .ZN(n8264) );
  NAND2_X1 U5668 ( .A1(n8257), .A2(n4827), .ZN(n4821) );
  INV_X1 U5669 ( .A(n8724), .ZN(n8242) );
  AND2_X1 U5670 ( .A1(n5939), .A2(n5938), .ZN(n8553) );
  AND2_X1 U5671 ( .A1(n5928), .A2(n5927), .ZN(n8303) );
  AND3_X1 U5672 ( .A1(n5908), .A2(n5907), .A3(n5906), .ZN(n8667) );
  NAND2_X1 U5673 ( .A1(n4830), .A2(n4358), .ZN(n4829) );
  INV_X1 U5674 ( .A(n8257), .ZN(n4830) );
  AND4_X1 U5675 ( .A1(n5834), .A2(n5833), .A3(n5832), .A4(n5831), .ZN(n9662)
         );
  AND2_X1 U5676 ( .A1(n4827), .A2(n8263), .ZN(n4824) );
  OAI21_X1 U5677 ( .B1(n4825), .B2(n4823), .A(n4324), .ZN(n4822) );
  OR2_X1 U5678 ( .A1(n8358), .A2(n8357), .ZN(n8359) );
  XNOR2_X1 U5679 ( .A(n5955), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8172) );
  AND2_X1 U5680 ( .A1(n7114), .A2(n7113), .ZN(n8521) );
  INV_X1 U5681 ( .A(n8350), .ZN(n8546) );
  INV_X1 U5682 ( .A(n8303), .ZN(n8580) );
  INV_X1 U5683 ( .A(n8251), .ZN(n8598) );
  INV_X1 U5684 ( .A(n8326), .ZN(n8614) );
  INV_X1 U5685 ( .A(n8667), .ZN(n8642) );
  INV_X1 U5686 ( .A(n8682), .ZN(n8706) );
  INV_X1 U5687 ( .A(n9662), .ZN(n8705) );
  INV_X1 U5688 ( .A(n8310), .ZN(n8373) );
  INV_X1 U5689 ( .A(n8313), .ZN(n8375) );
  NAND2_X1 U5690 ( .A1(n5670), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5686) );
  OR2_X1 U5691 ( .A1(n6777), .A2(n6322), .ZN(n8382) );
  INV_X1 U5692 ( .A(n4403), .ZN(n6748) );
  XNOR2_X1 U5693 ( .A(n4401), .B(n6754), .ZN(n6793) );
  INV_X1 U5694 ( .A(n4411), .ZN(n7038) );
  INV_X1 U5695 ( .A(n4710), .ZN(n8384) );
  XNOR2_X1 U5696 ( .A(n8461), .B(n8441), .ZN(n8442) );
  INV_X1 U5697 ( .A(n8464), .ZN(n4381) );
  OR2_X1 U5698 ( .A1(n4690), .A2(n4362), .ZN(n4689) );
  NOR2_X1 U5699 ( .A1(n4690), .A2(n4361), .ZN(n4687) );
  INV_X1 U5700 ( .A(n8518), .ZN(n4409) );
  NAND2_X1 U5701 ( .A1(n5619), .A2(n5618), .ZN(n8769) );
  NAND2_X1 U5702 ( .A1(n5885), .A2(n5884), .ZN(n8779) );
  NAND2_X1 U5703 ( .A1(n5858), .A2(n5857), .ZN(n8699) );
  NAND2_X1 U5704 ( .A1(n7713), .A2(n8042), .ZN(n9653) );
  OAI21_X1 U5705 ( .B1(n7467), .B2(n4274), .A(n4472), .ZN(n7633) );
  NAND2_X1 U5706 ( .A1(n5763), .A2(n5762), .ZN(n9856) );
  NAND2_X1 U5707 ( .A1(n4614), .A2(n8009), .ZN(n7374) );
  NAND2_X1 U5708 ( .A1(n4615), .A2(n8005), .ZN(n4614) );
  INV_X1 U5709 ( .A(n7255), .ZN(n4615) );
  NAND2_X1 U5710 ( .A1(n6772), .A2(n8880), .ZN(n9656) );
  NAND2_X1 U5711 ( .A1(n8672), .A2(n9667), .ZN(n8713) );
  INV_X1 U5712 ( .A(n8561), .ZN(n8710) );
  INV_X1 U5713 ( .A(n9656), .ZN(n8731) );
  NAND2_X1 U5714 ( .A1(n8116), .A2(n8115), .ZN(n8797) );
  NAND2_X1 U5715 ( .A1(n8101), .A2(n8100), .ZN(n8120) );
  NAND2_X1 U5716 ( .A1(n5601), .A2(n5600), .ZN(n8812) );
  NAND2_X1 U5717 ( .A1(n5931), .A2(n5930), .ZN(n8353) );
  NAND2_X1 U5718 ( .A1(n5921), .A2(n5920), .ZN(n8816) );
  NAND2_X1 U5719 ( .A1(n5640), .A2(n5639), .ZN(n8822) );
  NAND2_X1 U5720 ( .A1(n8321), .A2(n8320), .ZN(n5912) );
  INV_X1 U5721 ( .A(n4607), .ZN(n4602) );
  INV_X1 U5722 ( .A(n7943), .ZN(n8842) );
  NAND2_X1 U5723 ( .A1(n5900), .A2(n5899), .ZN(n8848) );
  NAND2_X1 U5724 ( .A1(n5868), .A2(n5867), .ZN(n8858) );
  NAND2_X1 U5725 ( .A1(n5839), .A2(n5838), .ZN(n8871) );
  INV_X1 U5726 ( .A(n8863), .ZN(n8870) );
  INV_X1 U5727 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4805) );
  MUX2_X1 U5728 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6012), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6013) );
  INV_X1 U5729 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4365) );
  NAND2_X1 U5730 ( .A1(n6009), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6007) );
  INV_X1 U5731 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n9968) );
  INV_X1 U5732 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7498) );
  INV_X1 U5733 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7405) );
  CLKBUF_X1 U5734 ( .A(n7404), .Z(n8502) );
  INV_X1 U5735 ( .A(n8388), .ZN(n8385) );
  INV_X1 U5736 ( .A(n7687), .ZN(n7684) );
  INV_X1 U5737 ( .A(n7152), .ZN(n7340) );
  INV_X1 U5738 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6388) );
  AND2_X1 U5739 ( .A1(n6328), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6321) );
  NAND2_X1 U5740 ( .A1(n7303), .A2(n7302), .ZN(n7483) );
  INV_X1 U5741 ( .A(n4678), .ZN(n4674) );
  NAND2_X1 U5742 ( .A1(n4677), .A2(n4678), .ZN(n9013) );
  INV_X1 U5743 ( .A(n9031), .ZN(n9032) );
  NOR2_X1 U5744 ( .A1(n7595), .A2(n7594), .ZN(n7668) );
  OR2_X1 U5745 ( .A1(n5322), .A2(n5129), .ZN(n5135) );
  NAND2_X1 U5746 ( .A1(n4679), .A2(n8934), .ZN(n9049) );
  NAND2_X1 U5747 ( .A1(n5342), .A2(n5341), .ZN(n9518) );
  INV_X1 U5748 ( .A(n7629), .ZN(n9799) );
  AND2_X1 U5749 ( .A1(n6701), .A2(n6698), .ZN(n6699) );
  INV_X1 U5750 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9996) );
  INV_X1 U5751 ( .A(n7861), .ZN(n5478) );
  INV_X1 U5752 ( .A(n4385), .ZN(n5117) );
  OAI21_X1 U5753 ( .B1(n5287), .B2(n6362), .A(n4386), .ZN(n4385) );
  AOI21_X1 U5754 ( .B1(n6526), .B2(P1_STATE_REG_SCAN_IN), .A(n7743), .ZN(n9157) );
  AOI21_X1 U5755 ( .B1(n4663), .B2(n9107), .A(n4662), .ZN(n4661) );
  INV_X1 U5756 ( .A(n8926), .ZN(n4663) );
  NOR2_X2 U5757 ( .A1(n6558), .A2(n6551), .ZN(n9165) );
  NAND2_X1 U5758 ( .A1(n8920), .A2(n4510), .ZN(n9181) );
  NAND2_X1 U5759 ( .A1(n6161), .A2(n4556), .ZN(n4548) );
  INV_X1 U5760 ( .A(n4533), .ZN(n4529) );
  NOR2_X1 U5761 ( .A1(n6310), .A2(n6312), .ZN(n4531) );
  OAI21_X1 U5762 ( .B1(n6309), .B2(n7551), .A(n6308), .ZN(n6318) );
  OR2_X1 U5763 ( .A1(n4534), .A2(n4533), .ZN(n4528) );
  NOR2_X1 U5764 ( .A1(n6198), .A2(n6197), .ZN(n6201) );
  AND3_X1 U5765 ( .A1(n5022), .A2(n5021), .A3(n5020), .ZN(n9078) );
  INV_X1 U5766 ( .A(n7196), .ZN(n9214) );
  NAND4_X1 U5767 ( .A1(n5145), .A2(n5144), .A3(n5143), .A4(n5142), .ZN(n9215)
         );
  INV_X1 U5768 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4881) );
  NAND4_X2 U5769 ( .A1(n5101), .A2(n5100), .A3(n5099), .A4(n5098), .ZN(n9219)
         );
  OR2_X1 U5770 ( .A1(n5141), .A2(n5097), .ZN(n5098) );
  AOI21_X1 U5771 ( .B1(n6408), .B2(P1_REG1_REG_1__SCAN_IN), .A(n6402), .ZN(
        n6510) );
  AOI21_X1 U5772 ( .B1(n6433), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6439), .ZN(
        n6496) );
  INV_X1 U5773 ( .A(n4595), .ZN(n6424) );
  AND2_X1 U5774 ( .A1(n4595), .A2(n4594), .ZN(n6413) );
  NAND2_X1 U5775 ( .A1(n6427), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4594) );
  INV_X1 U5776 ( .A(n4593), .ZN(n6450) );
  AOI21_X1 U5777 ( .B1(n6427), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6421), .ZN(
        n6406) );
  AOI21_X1 U5778 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n6568), .A(n6564), .ZN(
        n6566) );
  NOR2_X1 U5779 ( .A1(n6567), .A2(n4350), .ZN(n6571) );
  NOR2_X1 U5780 ( .A1(n6570), .A2(n6571), .ZN(n6738) );
  AOI21_X1 U5781 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6739), .A(n6738), .ZN(
        n6740) );
  NAND2_X1 U5782 ( .A1(n6740), .A2(n6741), .ZN(n7386) );
  NOR2_X1 U5783 ( .A1(n9678), .A2(n4598), .ZN(n7388) );
  AND2_X1 U5784 ( .A1(n9677), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4598) );
  NAND2_X1 U5785 ( .A1(n7388), .A2(n7389), .ZN(n9229) );
  AOI21_X1 U5786 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n9702), .A(n9694), .ZN(
        n9711) );
  NOR2_X1 U5787 ( .A1(n9697), .A2(n4597), .ZN(n9708) );
  NOR2_X1 U5788 ( .A1(n9232), .A2(n9231), .ZN(n4597) );
  NOR2_X1 U5789 ( .A1(n9708), .A2(n9707), .ZN(n9706) );
  XNOR2_X1 U5790 ( .A(n9234), .B(n9717), .ZN(n9722) );
  NOR2_X1 U5791 ( .A1(n9243), .A2(n4584), .ZN(n9254) );
  AND2_X1 U5792 ( .A1(n9245), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4584) );
  OR2_X1 U5793 ( .A1(n9732), .A2(n9731), .ZN(n9741) );
  OAI21_X1 U5794 ( .B1(n9746), .B2(n4879), .A(n9269), .ZN(n4586) );
  NAND2_X1 U5795 ( .A1(n4463), .A2(n4356), .ZN(n9315) );
  OR2_X1 U5796 ( .A1(n9324), .A2(n9323), .ZN(n9499) );
  INV_X1 U5797 ( .A(n5480), .ZN(n9346) );
  NAND2_X1 U5798 ( .A1(n4794), .A2(n4864), .ZN(n9393) );
  NAND2_X1 U5799 ( .A1(n9406), .A2(n5536), .ZN(n4794) );
  NAND2_X1 U5800 ( .A1(n9464), .A2(n6284), .ZN(n9453) );
  NAND2_X1 U5801 ( .A1(n4644), .A2(n6273), .ZN(n7723) );
  NAND2_X1 U5802 ( .A1(n5266), .A2(n6114), .ZN(n7617) );
  AND2_X1 U5803 ( .A1(n7655), .A2(n6990), .ZN(n9460) );
  OR2_X1 U5804 ( .A1(n6556), .A2(n6555), .ZN(n9471) );
  INV_X1 U5805 ( .A(n9765), .ZN(n9450) );
  OR2_X1 U5806 ( .A1(n9749), .A2(n6623), .ZN(n9765) );
  NAND2_X1 U5808 ( .A1(n5258), .A2(n5257), .ZN(n7680) );
  AND2_X1 U5809 ( .A1(n6182), .A2(n6181), .ZN(n9562) );
  OR2_X1 U5810 ( .A1(n5483), .A2(n5482), .ZN(n5484) );
  AND2_X1 U5811 ( .A1(n5427), .A2(n5426), .ZN(n9568) );
  NAND2_X1 U5812 ( .A1(n4779), .A2(n4783), .ZN(n9338) );
  NAND2_X1 U5813 ( .A1(n4787), .A2(n4784), .ZN(n4779) );
  INV_X1 U5814 ( .A(n5538), .ZN(n4785) );
  NAND2_X1 U5815 ( .A1(n4787), .A2(n5539), .ZN(n4786) );
  OAI21_X1 U5816 ( .B1(n7783), .B2(n4774), .A(n4770), .ZN(n9469) );
  NAND2_X1 U5817 ( .A1(n5081), .A2(n5080), .ZN(n9616) );
  AND2_X1 U5818 ( .A1(n4776), .A2(n4306), .ZN(n7885) );
  NAND2_X1 U5819 ( .A1(n7783), .A2(n5530), .ZN(n4776) );
  NAND2_X1 U5820 ( .A1(n5308), .A2(n5307), .ZN(n9019) );
  NOR2_X1 U5821 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n4803) );
  INV_X1 U5822 ( .A(n5510), .ZN(n7908) );
  NAND2_X1 U5823 ( .A1(n4733), .A2(n4738), .ZN(n5350) );
  INV_X1 U5824 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7748) );
  XNOR2_X1 U5825 ( .A(n5461), .B(n5459), .ZN(n7605) );
  INV_X1 U5826 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8212) );
  AND2_X1 U5827 ( .A1(n5059), .A2(n5026), .ZN(n5044) );
  INV_X1 U5828 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7205) );
  NAND2_X1 U5829 ( .A1(n4726), .A2(n4937), .ZN(n5268) );
  NAND2_X1 U5830 ( .A1(n5233), .A2(n4931), .ZN(n5237) );
  AND2_X1 U5831 ( .A1(n5254), .A2(n5241), .ZN(n9649) );
  NAND2_X1 U5832 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4600) );
  INV_X1 U5833 ( .A(n8382), .ZN(P2_U3893) );
  NAND2_X1 U5834 ( .A1(n4813), .A2(n8336), .ZN(n4812) );
  INV_X1 U5835 ( .A(n4696), .ZN(n7683) );
  XNOR2_X1 U5836 ( .A(n8465), .B(n4381), .ZN(n8492) );
  OAI21_X1 U5837 ( .B1(n4686), .B2(n4688), .A(n4408), .ZN(P2_U3201) );
  AOI21_X1 U5838 ( .B1(n8517), .B2(n8516), .A(n4409), .ZN(n4408) );
  AND2_X1 U5839 ( .A1(n8465), .A2(n4687), .ZN(n4686) );
  OAI21_X1 U5840 ( .B1(n8465), .B2(n4689), .A(n6759), .ZN(n4688) );
  OAI21_X1 U5841 ( .B1(n8804), .B2(n9670), .A(n4491), .ZN(P2_U3205) );
  INV_X1 U5842 ( .A(n4492), .ZN(n4491) );
  OAI21_X1 U5843 ( .B1(n8809), .B2(n8713), .A(n4493), .ZN(n4492) );
  AND2_X1 U5844 ( .A1(n8551), .A2(n4355), .ZN(n4493) );
  OAI21_X1 U5845 ( .B1(n8529), .B2(n8785), .A(n4851), .ZN(n6042) );
  NAND2_X1 U5846 ( .A1(n8748), .A2(n8747), .ZN(n8750) );
  NAND2_X1 U5847 ( .A1(n8746), .A2(n8745), .ZN(n8747) );
  OAI21_X1 U5848 ( .B1(n8529), .B2(n8863), .A(n6055), .ZN(n6056) );
  INV_X1 U5849 ( .A(n4586), .ZN(n4585) );
  NAND2_X1 U5850 ( .A1(n4588), .A2(n9268), .ZN(n4587) );
  AOI21_X1 U5851 ( .B1(n4591), .B2(n9682), .A(n9266), .ZN(n4590) );
  AND2_X1 U5852 ( .A1(n9482), .A2(n9485), .ZN(n9555) );
  OAI21_X1 U5853 ( .B1(n6319), .B2(n9812), .A(n4373), .ZN(P1_U3549) );
  NOR2_X1 U5854 ( .A1(n4348), .A2(n4374), .ZN(n4373) );
  NOR2_X1 U5855 ( .A1(n9811), .A2(n6320), .ZN(n4374) );
  NAND2_X1 U5856 ( .A1(n4388), .A2(n4294), .ZN(n9557) );
  AOI21_X1 U5857 ( .B1(n9010), .B2(n6071), .A(n6070), .ZN(n6072) );
  NOR2_X1 U5858 ( .A1(n9795), .A2(n6069), .ZN(n6070) );
  NAND2_X1 U5859 ( .A1(n4528), .A2(n4363), .ZN(n4273) );
  CLKBUF_X3 U5860 ( .A(n6857), .Z(n8205) );
  NAND2_X1 U5861 ( .A1(n6521), .A2(n6632), .ZN(n7121) );
  OR2_X1 U5862 ( .A1(n5770), .A2(n4474), .ZN(n4274) );
  INV_X1 U5863 ( .A(n6481), .ZN(n4682) );
  AND2_X1 U5864 ( .A1(n4750), .A2(n4751), .ZN(n4275) );
  AND2_X1 U5865 ( .A1(n4704), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4276) );
  AND2_X1 U5866 ( .A1(n8934), .A2(n4852), .ZN(n4277) );
  NOR2_X1 U5867 ( .A1(n5977), .A2(n5976), .ZN(n4278) );
  INV_X1 U5868 ( .A(n8044), .ZN(n4622) );
  AND2_X1 U5869 ( .A1(n4732), .A2(n4922), .ZN(n4279) );
  NOR2_X1 U5870 ( .A1(n8383), .A2(n6941), .ZN(n7980) );
  AND2_X1 U5871 ( .A1(n5988), .A2(n8539), .ZN(n4281) );
  INV_X1 U5872 ( .A(n9010), .ZN(n4394) );
  NAND3_X1 U5873 ( .A1(n4574), .A2(n4572), .A3(n4465), .ZN(n6162) );
  INV_X1 U5874 ( .A(n7365), .ZN(n4839) );
  AND2_X1 U5875 ( .A1(n4814), .A2(n4818), .ZN(n4282) );
  AND2_X1 U5876 ( .A1(n9468), .A2(n4771), .ZN(n4283) );
  AND2_X1 U5877 ( .A1(n4445), .A2(n4312), .ZN(n4284) );
  NOR2_X1 U5878 ( .A1(n8576), .A2(n5648), .ZN(n4285) );
  NAND2_X1 U5879 ( .A1(n9414), .A2(n4398), .ZN(n4399) );
  AND2_X1 U5880 ( .A1(n5027), .A2(n4318), .ZN(n4286) );
  NOR2_X1 U5881 ( .A1(n6318), .A2(n4531), .ZN(n4287) );
  OR2_X1 U5882 ( .A1(n8096), .A2(n8097), .ZN(n4288) );
  INV_X1 U5883 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4980) );
  AND2_X1 U5884 ( .A1(n4831), .A2(n8631), .ZN(n4289) );
  AND4_X1 U5885 ( .A1(n5487), .A2(n4505), .A3(n4979), .A4(n5506), .ZN(n4290)
         );
  NOR2_X1 U5886 ( .A1(n5023), .A2(n4746), .ZN(n4745) );
  INV_X1 U5887 ( .A(n6303), .ZN(n6311) );
  AND2_X1 U5888 ( .A1(n6200), .A2(n6199), .ZN(n6303) );
  AND2_X1 U5889 ( .A1(n4396), .A2(n4395), .ZN(n4291) );
  NAND2_X1 U5890 ( .A1(n4559), .A2(n4569), .ZN(n4292) );
  INV_X1 U5891 ( .A(n8683), .ZN(n8655) );
  AND4_X1 U5892 ( .A1(n5891), .A2(n5890), .A3(n5889), .A4(n5888), .ZN(n8683)
         );
  NOR2_X1 U5893 ( .A1(n4675), .A2(n4674), .ZN(n4293) );
  OR2_X1 U5894 ( .A1(n9804), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n4294) );
  INV_X1 U5895 ( .A(n6532), .ZN(n6687) );
  INV_X2 U5896 ( .A(n6687), .ZN(n8978) );
  NAND3_X2 U5897 ( .A1(n6627), .A2(n6521), .A3(n6482), .ZN(n6532) );
  OR2_X1 U5898 ( .A1(n5069), .A2(SI_15_), .ZN(n4295) );
  INV_X1 U5899 ( .A(n9362), .ZN(n4787) );
  XOR2_X1 U5900 ( .A(n7592), .B(n8978), .Z(n4296) );
  INV_X1 U5901 ( .A(n4266), .ZN(n5137) );
  NAND2_X1 U5902 ( .A1(n4988), .A2(n4987), .ZN(n5475) );
  AND2_X1 U5903 ( .A1(n5359), .A2(n5358), .ZN(n5480) );
  NAND2_X1 U5904 ( .A1(n5677), .A2(n4714), .ZN(n5679) );
  NAND2_X1 U5905 ( .A1(n4265), .A2(n4846), .ZN(n4297) );
  OR2_X1 U5906 ( .A1(n7136), .A2(n4382), .ZN(n4298) );
  NAND2_X1 U5907 ( .A1(n5980), .A2(n8074), .ZN(n8156) );
  AND2_X1 U5908 ( .A1(n8128), .A2(n8110), .ZN(n4299) );
  OR2_X1 U5909 ( .A1(n8919), .A2(n9098), .ZN(n4300) );
  OR2_X1 U5910 ( .A1(n7124), .A2(n7123), .ZN(n4301) );
  AND2_X1 U5911 ( .A1(n4945), .A2(n4755), .ZN(n4302) );
  INV_X1 U5912 ( .A(n7911), .ZN(n6018) );
  NAND2_X1 U5913 ( .A1(n6014), .A2(n6013), .ZN(n7911) );
  AND4_X1 U5914 ( .A1(n4845), .A2(n5566), .A3(n5783), .A4(n4627), .ZN(n6010)
         );
  NAND2_X1 U5915 ( .A1(n5018), .A2(n5017), .ZN(n9520) );
  INV_X1 U5916 ( .A(n6690), .ZN(n9216) );
  AND4_X1 U5917 ( .A1(n5125), .A2(n5124), .A3(n5123), .A4(n5122), .ZN(n6690)
         );
  NOR2_X1 U5918 ( .A1(n8177), .A2(n4828), .ZN(n4827) );
  NAND2_X1 U5919 ( .A1(n4658), .A2(n4661), .ZN(n9148) );
  NAND2_X1 U5920 ( .A1(n9095), .A2(n8926), .ZN(n9105) );
  NAND2_X1 U5921 ( .A1(n4829), .A2(n8255), .ZN(n8178) );
  INV_X1 U5922 ( .A(n6236), .ZN(n4657) );
  INV_X1 U5923 ( .A(n6485), .ZN(n8988) );
  NAND3_X2 U5924 ( .A1(n6989), .A2(n4680), .A3(n6521), .ZN(n6485) );
  INV_X1 U5925 ( .A(n8557), .ZN(n4443) );
  OR2_X1 U5926 ( .A1(n9027), .A2(n9026), .ZN(n4303) );
  AND2_X1 U5927 ( .A1(n9325), .A2(n4391), .ZN(n4304) );
  OR2_X1 U5928 ( .A1(n9860), .A2(n8373), .ZN(n4305) );
  INV_X1 U5929 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9621) );
  NAND2_X1 U5930 ( .A1(n8915), .A2(n8914), .ZN(n4306) );
  OR2_X1 U5931 ( .A1(n8806), .A2(n8554), .ZN(n4307) );
  NAND2_X1 U5932 ( .A1(n4265), .A2(n5567), .ZN(n5956) );
  NAND2_X1 U5933 ( .A1(n5959), .A2(n4845), .ZN(n6011) );
  NAND2_X1 U5934 ( .A1(n4757), .A2(n5112), .ZN(n5150) );
  AND4_X1 U5935 ( .A1(n5769), .A2(n5768), .A3(n5767), .A4(n5766), .ZN(n7773)
         );
  INV_X1 U5936 ( .A(n7773), .ZN(n8374) );
  INV_X1 U5937 ( .A(n9513), .ZN(n5479) );
  NAND2_X1 U5938 ( .A1(n5004), .A2(n5003), .ZN(n9513) );
  INV_X1 U5939 ( .A(n8138), .ZN(n7465) );
  INV_X1 U5940 ( .A(n5477), .ZN(n9775) );
  AND2_X1 U5941 ( .A1(n5475), .A2(n9197), .ZN(n4308) );
  AND2_X1 U5942 ( .A1(n4575), .A2(n4579), .ZN(n4309) );
  OR2_X1 U5943 ( .A1(n6130), .A2(n6122), .ZN(n4310) );
  AND2_X1 U5944 ( .A1(n4679), .A2(n4277), .ZN(n4311) );
  OR2_X1 U5945 ( .A1(n4441), .A2(n4299), .ZN(n4312) );
  INV_X1 U5946 ( .A(n5847), .ZN(n4486) );
  AND2_X1 U5947 ( .A1(n6221), .A2(n6310), .ZN(n4313) );
  AND2_X1 U5948 ( .A1(n4794), .A2(n4792), .ZN(n4314) );
  AND2_X1 U5949 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n4315) );
  NAND2_X1 U5950 ( .A1(n8537), .A2(n8540), .ZN(n4316) );
  INV_X1 U5951 ( .A(n4606), .ZN(n8620) );
  AND2_X1 U5952 ( .A1(n4701), .A2(n4698), .ZN(n4317) );
  INV_X1 U5953 ( .A(n9568), .ZN(n9289) );
  AND2_X1 U5954 ( .A1(n5026), .A2(n4505), .ZN(n4318) );
  AND2_X1 U5955 ( .A1(n7288), .A2(n7287), .ZN(n4319) );
  INV_X1 U5956 ( .A(n4775), .ZN(n4774) );
  AND2_X1 U5957 ( .A1(n5531), .A2(n4306), .ZN(n4775) );
  NOR2_X1 U5958 ( .A1(n7570), .A2(n8376), .ZN(n4320) );
  INV_X1 U5959 ( .A(n4771), .ZN(n4770) );
  NAND2_X1 U5960 ( .A1(n4772), .A2(n4300), .ZN(n4771) );
  OR2_X1 U5961 ( .A1(n5025), .A2(n4862), .ZN(n4321) );
  NAND2_X1 U5962 ( .A1(n5911), .A2(n5910), .ZN(n8575) );
  INV_X1 U5963 ( .A(n8575), .ZN(n4477) );
  INV_X1 U5964 ( .A(n6831), .ZN(n4704) );
  OR2_X1 U5965 ( .A1(n8120), .A2(n8102), .ZN(n8105) );
  NAND2_X1 U5966 ( .A1(n4820), .A2(n4819), .ZN(n4322) );
  NOR2_X1 U5967 ( .A1(n9010), .A2(n9193), .ZN(n4323) );
  INV_X1 U5968 ( .A(n8206), .ZN(n4820) );
  XOR2_X1 U5969 ( .A(n8205), .B(n8544), .Z(n8206) );
  NAND2_X1 U5970 ( .A1(n8182), .A2(n8181), .ZN(n4324) );
  AOI21_X1 U5971 ( .B1(n6202), .B2(n6201), .A(n6303), .ZN(n6203) );
  INV_X1 U5972 ( .A(n6203), .ZN(n4530) );
  AND2_X1 U5973 ( .A1(n9871), .A2(n8371), .ZN(n4325) );
  AND2_X1 U5974 ( .A1(n8650), .A2(n8059), .ZN(n8679) );
  AND2_X1 U5975 ( .A1(n8082), .A2(n4299), .ZN(n4326) );
  INV_X1 U5976 ( .A(n4621), .ZN(n4620) );
  NAND2_X1 U5977 ( .A1(n4622), .A2(n8037), .ZN(n4621) );
  NAND2_X1 U5978 ( .A1(n4500), .A2(n4499), .ZN(n4327) );
  OR2_X1 U5979 ( .A1(n4308), .A2(n5538), .ZN(n4328) );
  NAND2_X1 U5980 ( .A1(n6156), .A2(n6153), .ZN(n6219) );
  OR2_X1 U5981 ( .A1(n7973), .A2(n8070), .ZN(n4329) );
  AND2_X1 U5982 ( .A1(n8118), .A2(n8103), .ZN(n8099) );
  INV_X1 U5983 ( .A(n8099), .ZN(n4418) );
  AND2_X1 U5984 ( .A1(n4786), .A2(n4785), .ZN(n4330) );
  AND3_X1 U5985 ( .A1(n4514), .A2(n5456), .A3(n5465), .ZN(n4331) );
  NOR2_X1 U5986 ( .A1(n4842), .A2(n4844), .ZN(n4841) );
  INV_X1 U5987 ( .A(n4926), .ZN(n4732) );
  AND2_X1 U5988 ( .A1(n5506), .A2(n5487), .ZN(n4332) );
  NAND2_X1 U5989 ( .A1(n5919), .A2(n5918), .ZN(n4333) );
  AND2_X1 U5990 ( .A1(n5588), .A2(n4805), .ZN(n4334) );
  OR2_X1 U5991 ( .A1(n7060), .A2(n7241), .ZN(n4335) );
  AND2_X1 U5992 ( .A1(n4367), .A2(n4366), .ZN(n4336) );
  AND2_X1 U5993 ( .A1(n4281), .A2(n4625), .ZN(n4337) );
  AND2_X1 U5994 ( .A1(n5385), .A2(n5384), .ZN(n4338) );
  AND2_X1 U5995 ( .A1(n5454), .A2(n6297), .ZN(n6167) );
  INV_X1 U5996 ( .A(n6167), .ZN(n4566) );
  OR2_X1 U5997 ( .A1(n9500), .A2(n9170), .ZN(n6221) );
  AND2_X1 U5998 ( .A1(n4302), .A2(n4753), .ZN(n4339) );
  INV_X1 U5999 ( .A(n8081), .ZN(n5983) );
  AND2_X1 U6000 ( .A1(n5982), .A2(n8614), .ZN(n8081) );
  OR2_X1 U6001 ( .A1(n6808), .A2(n6807), .ZN(n4340) );
  NAND2_X1 U6002 ( .A1(n4558), .A2(n4567), .ZN(n4341) );
  INV_X1 U6003 ( .A(n7759), .ZN(n4500) );
  INV_X1 U6004 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4514) );
  INV_X1 U6005 ( .A(n6813), .ZN(n4703) );
  INV_X1 U6006 ( .A(n7154), .ZN(n7044) );
  INV_X1 U6007 ( .A(n5475), .ZN(n4395) );
  INV_X1 U6008 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4522) );
  XNOR2_X1 U6009 ( .A(n5716), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6802) );
  AND2_X1 U6010 ( .A1(n8359), .A2(n7935), .ZN(n4342) );
  AND2_X1 U6011 ( .A1(n4458), .A2(n4946), .ZN(n4343) );
  NAND2_X1 U6012 ( .A1(n5049), .A2(n5048), .ZN(n9434) );
  INV_X1 U6013 ( .A(n9434), .ZN(n9605) );
  NOR2_X1 U6014 ( .A1(n9150), .A2(n9149), .ZN(n4344) );
  NOR2_X1 U6015 ( .A1(n7668), .A2(n7667), .ZN(n4345) );
  AND2_X1 U6016 ( .A1(n9401), .A2(n9078), .ZN(n4346) );
  AND2_X1 U6017 ( .A1(n5969), .A2(n8037), .ZN(n4347) );
  NOR2_X1 U6018 ( .A1(n4394), .A2(n9537), .ZN(n4348) );
  NOR2_X1 U6019 ( .A1(n9475), .A2(n9540), .ZN(n9431) );
  AND4_X1 U6020 ( .A1(n5203), .A2(n5202), .A3(n5201), .A4(n5200), .ZN(n7485)
         );
  OR2_X1 U6021 ( .A1(n9110), .A2(n9605), .ZN(n4349) );
  AND2_X1 U6022 ( .A1(n6568), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4350) );
  NAND2_X1 U6023 ( .A1(n9346), .A2(n9196), .ZN(n4351) );
  INV_X1 U6024 ( .A(n9792), .ZN(n7600) );
  AND4_X1 U6025 ( .A1(n5806), .A2(n5805), .A3(n5804), .A4(n5803), .ZN(n9664)
         );
  NAND2_X1 U6026 ( .A1(n8548), .A2(n8547), .ZN(n4352) );
  OR2_X1 U6027 ( .A1(n5318), .A2(SI_16_), .ZN(n4353) );
  AND2_X1 U6028 ( .A1(n4605), .A2(n4602), .ZN(n4354) );
  OR2_X1 U6029 ( .A1(n9668), .A2(n8549), .ZN(n4355) );
  NAND2_X1 U6030 ( .A1(n6190), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n4356) );
  OR2_X1 U6031 ( .A1(n7687), .A2(n10012), .ZN(n4357) );
  OR2_X1 U6032 ( .A1(n7942), .A2(n8642), .ZN(n4358) );
  NOR2_X1 U6033 ( .A1(n7625), .A2(n7629), .ZN(n7626) );
  INV_X1 U6034 ( .A(n8356), .ZN(n8336) );
  INV_X1 U6035 ( .A(n6168), .ZN(n6310) );
  NAND2_X2 U6036 ( .A1(n8172), .A2(n6945), .ZN(n8110) );
  INV_X1 U6037 ( .A(n6557), .ZN(n4681) );
  AND2_X1 U6038 ( .A1(n9804), .A2(n9485), .ZN(n4359) );
  INV_X1 U6039 ( .A(n5989), .ZN(n7404) );
  AND2_X1 U6040 ( .A1(n4701), .A2(n4699), .ZN(n4360) );
  AND2_X1 U6041 ( .A1(n4694), .A2(n8493), .ZN(n4361) );
  NOR2_X1 U6042 ( .A1(n4694), .A2(n8464), .ZN(n4362) );
  NAND2_X1 U6043 ( .A1(n4850), .A2(n6317), .ZN(n4363) );
  AND2_X1 U6044 ( .A1(n5958), .A2(n4297), .ZN(n6945) );
  NAND3_X2 U6045 ( .A1(n4502), .A2(n4501), .A3(n4503), .ZN(n9268) );
  INV_X1 U6046 ( .A(n4997), .ZN(n4799) );
  AND2_X1 U6047 ( .A1(n5589), .A2(n4334), .ZN(n8883) );
  INV_X1 U6048 ( .A(n8165), .ZN(n7499) );
  XNOR2_X1 U6049 ( .A(n5961), .B(P2_IR_REG_20__SCAN_IN), .ZN(n8165) );
  NAND2_X1 U6050 ( .A1(n6623), .A2(n6205), .ZN(n4532) );
  INV_X1 U6051 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4806) );
  OAI21_X1 U6052 ( .B1(n7927), .B2(n8371), .A(n7926), .ZN(n4809) );
  OAI22_X1 U6053 ( .A1(n7363), .A2(n7362), .B1(n7361), .B2(n8378), .ZN(n7364)
         );
  AOI21_X2 U6054 ( .B1(n7772), .B2(n7771), .A(n7770), .ZN(n8309) );
  NAND2_X1 U6055 ( .A1(n9378), .A2(n9377), .ZN(n4364) );
  NAND2_X1 U6056 ( .A1(n9389), .A2(n9394), .ZN(n5336) );
  OAI211_X1 U6057 ( .C1(n4868), .C2(n4722), .A(n4720), .B(n4865), .ZN(n5206)
         );
  NAND2_X1 U6058 ( .A1(n5325), .A2(n5324), .ZN(n5476) );
  NAND2_X1 U6059 ( .A1(n4726), .A2(n4725), .ZN(n5269) );
  AOI21_X2 U6060 ( .B1(n6015), .B2(n6016), .A(n7911), .ZN(n6391) );
  OAI21_X1 U6061 ( .B1(n5340), .B2(n4737), .A(n4734), .ZN(n5352) );
  NAND2_X1 U6062 ( .A1(n6256), .A2(n6258), .ZN(n6257) );
  NAND2_X1 U6063 ( .A1(n6920), .A2(n4371), .ZN(n7014) );
  NAND2_X1 U6064 ( .A1(n4766), .A2(n5543), .ZN(n6060) );
  NAND2_X1 U6065 ( .A1(n7426), .A2(n4756), .ZN(n7641) );
  NAND4_X1 U6066 ( .A1(n4974), .A2(n4975), .A3(n4976), .A4(n5190), .ZN(n4372)
         );
  INV_X1 U6067 ( .A(n4767), .ZN(n9441) );
  NAND2_X1 U6068 ( .A1(n4601), .A2(n8129), .ZN(n8570) );
  INV_X1 U6069 ( .A(n8009), .ZN(n4610) );
  NAND2_X1 U6070 ( .A1(n4429), .A2(n4428), .ZN(n4723) );
  INV_X1 U6071 ( .A(n4613), .ZN(n4612) );
  AOI21_X1 U6072 ( .B1(n7255), .B2(n4613), .A(n4611), .ZN(n7466) );
  NAND2_X1 U6073 ( .A1(n5315), .A2(n6278), .ZN(n7890) );
  NAND2_X1 U6074 ( .A1(n5232), .A2(n6107), .ZN(n6239) );
  NAND3_X1 U6075 ( .A1(n4655), .A2(n5527), .A3(n4377), .ZN(n7421) );
  NAND2_X1 U6076 ( .A1(n5176), .A2(n4913), .ZN(n5204) );
  NAND2_X1 U6077 ( .A1(n9350), .A2(n9351), .ZN(n9349) );
  NAND2_X1 U6078 ( .A1(n4629), .A2(n4338), .ZN(n9321) );
  NOR2_X1 U6079 ( .A1(n4882), .A2(SI_1_), .ZN(n4718) );
  XNOR2_X1 U6080 ( .A(n4654), .B(n4566), .ZN(n4653) );
  NAND2_X2 U6081 ( .A1(n6854), .A2(n6853), .ZN(n6857) );
  NOR2_X2 U6082 ( .A1(n4378), .A2(n5690), .ZN(n5783) );
  NAND4_X1 U6083 ( .A1(n5559), .A2(n5558), .A3(n5560), .A4(n5557), .ZN(n4378)
         );
  NAND2_X1 U6084 ( .A1(n7927), .A2(n8371), .ZN(n4808) );
  NAND2_X1 U6085 ( .A1(n7803), .A2(n7802), .ZN(n7927) );
  NAND2_X1 U6086 ( .A1(n7061), .A2(n4335), .ZN(n7062) );
  NAND2_X1 U6087 ( .A1(n4809), .A2(n4808), .ZN(n7949) );
  NAND2_X2 U6088 ( .A1(n8335), .A2(n7941), .ZN(n8257) );
  OAI211_X1 U6089 ( .C1(n4590), .C2(n9268), .A(n4587), .B(n4585), .ZN(P1_U3262) );
  AND2_X2 U6090 ( .A1(n5316), .A2(n6283), .ZN(n9461) );
  NAND2_X1 U6091 ( .A1(n4628), .A2(n6073), .ZN(n9350) );
  OAI21_X1 U6092 ( .B1(n4280), .B2(n5234), .A(n4932), .ZN(n4727) );
  OAI21_X1 U6093 ( .B1(n9279), .B2(n9283), .A(n6165), .ZN(n4654) );
  INV_X1 U6094 ( .A(n4646), .ZN(n4645) );
  NAND2_X1 U6095 ( .A1(n4643), .A2(n4641), .ZN(n7785) );
  INV_X1 U6096 ( .A(n4384), .ZN(n7139) );
  NAND2_X1 U6097 ( .A1(n4384), .A2(n4383), .ZN(n4712) );
  OR2_X1 U6098 ( .A1(n7135), .A2(n7136), .ZN(n4384) );
  INV_X1 U6099 ( .A(n5219), .ZN(n4730) );
  NOR2_X1 U6100 ( .A1(n7922), .A2(n5484), .ZN(n5551) );
  NOR2_X1 U6101 ( .A1(n7439), .A2(n7440), .ZN(n7443) );
  NOR2_X1 U6102 ( .A1(n8410), .A2(n8411), .ZN(n8413) );
  NOR2_X1 U6103 ( .A1(n7817), .A2(n7818), .ZN(n7821) );
  NAND2_X4 U6104 ( .A1(n6366), .A2(n6489), .ZN(n6329) );
  NAND2_X1 U6105 ( .A1(n5256), .A2(n6409), .ZN(n4386) );
  NOR2_X2 U6106 ( .A1(n5477), .A2(n7008), .ZN(n7022) );
  NAND2_X1 U6107 ( .A1(n9482), .A2(n4359), .ZN(n4388) );
  NAND2_X1 U6108 ( .A1(n9325), .A2(n4392), .ZN(n9285) );
  INV_X1 U6109 ( .A(n4399), .ZN(n9368) );
  XNOR2_X1 U6110 ( .A(n4400), .B(n6645), .ZN(n6646) );
  XNOR2_X2 U6111 ( .A(n5654), .B(P2_IR_REG_1__SCAN_IN), .ZN(n6651) );
  INV_X1 U6112 ( .A(n8109), .ZN(n8106) );
  NAND3_X1 U6113 ( .A1(n4430), .A2(n4724), .A3(n8112), .ZN(n4429) );
  NAND2_X1 U6114 ( .A1(n8050), .A2(n4433), .ZN(n4432) );
  NAND2_X1 U6115 ( .A1(n8054), .A2(n8703), .ZN(n4436) );
  INV_X1 U6116 ( .A(n8090), .ZN(n4444) );
  NAND3_X1 U6117 ( .A1(n8016), .A2(n8051), .A3(n8024), .ZN(n4448) );
  INV_X2 U6118 ( .A(n4901), .ZN(n6345) );
  NAND3_X1 U6119 ( .A1(n4451), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4450) );
  NAND2_X1 U6120 ( .A1(n4295), .A2(n4275), .ZN(n5317) );
  NAND3_X1 U6121 ( .A1(n4461), .A2(n4460), .A3(n4933), .ZN(n4726) );
  INV_X1 U6122 ( .A(n4727), .ZN(n4461) );
  INV_X1 U6123 ( .A(n9315), .ZN(n9569) );
  NAND2_X1 U6124 ( .A1(n4572), .A2(n4574), .ZN(n6159) );
  NAND2_X1 U6125 ( .A1(n6162), .A2(n4464), .ZN(n4558) );
  INV_X1 U6126 ( .A(n6157), .ZN(n4465) );
  NAND3_X1 U6127 ( .A1(n4341), .A2(n4466), .A3(n4292), .ZN(n6202) );
  NAND2_X1 U6128 ( .A1(n4468), .A2(n7467), .ZN(n4467) );
  OAI21_X2 U6129 ( .B1(n8565), .B2(n5929), .A(n8085), .ZN(n7959) );
  OAI21_X2 U6130 ( .B1(n7716), .B2(n4325), .A(n5807), .ZN(n9660) );
  XNOR2_X1 U6131 ( .A(n8543), .B(n4494), .ZN(n4490) );
  NAND2_X1 U6132 ( .A1(n7667), .A2(n4500), .ZN(n4498) );
  XNOR2_X1 U6133 ( .A(n7124), .B(n4506), .ZN(n7125) );
  NAND2_X2 U6134 ( .A1(n7206), .A2(n4301), .ZN(n7218) );
  NAND3_X1 U6135 ( .A1(n8920), .A2(n4510), .A3(n4507), .ZN(n9178) );
  NAND2_X1 U6136 ( .A1(n9148), .A2(n4277), .ZN(n4513) );
  AND2_X2 U6137 ( .A1(n4630), .A2(n4631), .ZN(n4778) );
  OAI21_X1 U6138 ( .B1(n6129), .B2(n6168), .A(n4518), .ZN(n4520) );
  NAND3_X1 U6139 ( .A1(n4778), .A2(n4777), .A3(n4522), .ZN(n4521) );
  NOR2_X2 U6140 ( .A1(n4862), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4777) );
  NAND2_X1 U6141 ( .A1(n4526), .A2(n4523), .ZN(P1_U3242) );
  OAI22_X1 U6142 ( .A1(n4530), .A2(n4524), .B1(n4273), .B2(n4287), .ZN(n4523)
         );
  NAND2_X1 U6143 ( .A1(n6204), .A2(n4525), .ZN(n4524) );
  OR2_X1 U6144 ( .A1(n4527), .A2(n4530), .ZN(n4526) );
  NAND2_X1 U6145 ( .A1(n6204), .A2(n4529), .ZN(n4527) );
  OAI21_X1 U6146 ( .B1(n6314), .B2(n9268), .A(n6313), .ZN(n4533) );
  NAND3_X1 U6147 ( .A1(n4537), .A2(n6983), .A3(n4535), .ZN(n6086) );
  NAND3_X1 U6148 ( .A1(n4546), .A2(n4545), .A3(n4544), .ZN(n4543) );
  NAND2_X1 U6149 ( .A1(n6161), .A2(n4554), .ZN(n4547) );
  NAND3_X1 U6150 ( .A1(n4549), .A2(n4548), .A3(n4547), .ZN(n6192) );
  NAND3_X1 U6151 ( .A1(n4566), .A2(n4565), .A3(n4564), .ZN(n4563) );
  NAND2_X1 U6152 ( .A1(n9562), .A2(n6310), .ZN(n4571) );
  OAI21_X1 U6153 ( .B1(n4579), .B2(n4581), .A(n4576), .ZN(n4573) );
  NAND3_X1 U6154 ( .A1(n6154), .A2(n6151), .A3(n6221), .ZN(n4578) );
  MUX2_X1 U6155 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n5087), .S(n6401), .Z(n6334)
         );
  XNOR2_X2 U6156 ( .A(n4600), .B(n5088), .ZN(n6401) );
  NAND2_X1 U6157 ( .A1(n4605), .A2(n4603), .ZN(n5981) );
  NAND4_X1 U6158 ( .A1(n5685), .A2(n5686), .A3(n5688), .A4(n5687), .ZN(n8380)
         );
  NOR2_X1 U6159 ( .A1(n8137), .A2(n4610), .ZN(n4613) );
  NAND2_X1 U6160 ( .A1(n7466), .A2(n7465), .ZN(n7406) );
  OAI21_X1 U6161 ( .B1(n5969), .B2(n4617), .A(n4616), .ZN(n8732) );
  AOI21_X1 U6162 ( .B1(n5987), .B2(n4337), .A(n4623), .ZN(n8119) );
  AOI21_X1 U6163 ( .B1(n7406), .B2(n8025), .A(n5967), .ZN(n7607) );
  AOI21_X1 U6164 ( .B1(n8119), .B2(n8118), .A(n8117), .ZN(n8121) );
  NAND2_X1 U6165 ( .A1(n5971), .A2(n8060), .ZN(n8677) );
  NAND2_X1 U6166 ( .A1(n6970), .A2(n6969), .ZN(n6968) );
  NAND2_X1 U6167 ( .A1(n6968), .A2(n7997), .ZN(n7167) );
  XNOR2_X1 U6168 ( .A(n4723), .B(n7404), .ZN(n8175) );
  NAND2_X1 U6169 ( .A1(n9363), .A2(n9364), .ZN(n4628) );
  NAND3_X1 U6170 ( .A1(n4777), .A2(n4778), .A3(n4872), .ZN(n4982) );
  NAND3_X1 U6171 ( .A1(n4290), .A2(n4978), .A3(n4331), .ZN(n4862) );
  OAI21_X1 U6172 ( .B1(n9461), .B2(n4636), .A(n4633), .ZN(n5334) );
  INV_X1 U6173 ( .A(n4637), .ZN(n4636) );
  NAND2_X1 U6174 ( .A1(n5266), .A2(n4645), .ZN(n4643) );
  OAI21_X1 U6175 ( .B1(n7016), .B2(n7015), .A(n6084), .ZN(n6982) );
  NAND2_X1 U6176 ( .A1(n6265), .A2(n6084), .ZN(n7015) );
  OAI21_X2 U6178 ( .B1(n4653), .B2(n9412), .A(n5474), .ZN(n7922) );
  NAND2_X1 U6179 ( .A1(n9094), .A2(n4659), .ZN(n4658) );
  NOR2_X1 U6180 ( .A1(n6677), .A2(n6678), .ZN(n6545) );
  NAND3_X1 U6181 ( .A1(n6546), .A2(n4666), .A3(n4665), .ZN(n6686) );
  NAND2_X1 U6182 ( .A1(n4667), .A2(n6677), .ZN(n4665) );
  NAND2_X1 U6183 ( .A1(n4667), .A2(n6678), .ZN(n4666) );
  INV_X1 U6184 ( .A(n6547), .ZN(n4667) );
  AND2_X1 U6185 ( .A1(n6544), .A2(n6685), .ZN(n6546) );
  AOI21_X2 U6186 ( .B1(n7591), .B2(n7590), .A(n4874), .ZN(n7666) );
  OAI22_X2 U6187 ( .A1(n7218), .A2(n4669), .B1(n4668), .B2(n4670), .ZN(n7591)
         );
  NAND2_X1 U6188 ( .A1(n8913), .A2(n8912), .ZN(n4677) );
  NAND2_X1 U6189 ( .A1(n5463), .A2(n4684), .ZN(n5488) );
  NAND2_X1 U6190 ( .A1(n5463), .A2(n4683), .ZN(n4685) );
  NAND2_X1 U6191 ( .A1(n5463), .A2(n5458), .ZN(n5460) );
  NAND2_X1 U6192 ( .A1(n4706), .A2(n6609), .ZN(n6607) );
  INV_X1 U6193 ( .A(n6606), .ZN(n4708) );
  INV_X1 U6194 ( .A(n4712), .ZN(n7338) );
  AND3_X2 U6195 ( .A1(n5679), .A2(n4715), .A3(n4713), .ZN(n6603) );
  XNOR2_X1 U6196 ( .A(n5090), .B(n4719), .ZN(n6351) );
  NAND2_X1 U6197 ( .A1(n5167), .A2(n4908), .ZN(n5174) );
  NAND2_X1 U6198 ( .A1(n5167), .A2(n4721), .ZN(n4720) );
  AND2_X1 U6199 ( .A1(n4913), .A2(n4908), .ZN(n4721) );
  NAND2_X1 U6200 ( .A1(n5340), .A2(n4740), .ZN(n4733) );
  NAND2_X1 U6201 ( .A1(n5286), .A2(n4339), .ZN(n4750) );
  NAND3_X1 U6202 ( .A1(n4757), .A2(n5112), .A3(n4973), .ZN(n5072) );
  NAND2_X1 U6203 ( .A1(n9308), .A2(n4761), .ZN(n4760) );
  NAND2_X1 U6204 ( .A1(n9308), .A2(n5542), .ZN(n4766) );
  OAI21_X1 U6205 ( .B1(n9308), .B2(n4763), .A(n4761), .ZN(n9284) );
  AOI21_X2 U6206 ( .B1(n4787), .B2(n4782), .A(n4780), .ZN(n9318) );
  INV_X1 U6207 ( .A(n4795), .ZN(n9376) );
  NAND3_X1 U6209 ( .A1(n4997), .A2(n4996), .A3(P1_REG0_REG_1__SCAN_IN), .ZN(
        n4802) );
  INV_X1 U6210 ( .A(n4801), .ZN(n4800) );
  NAND2_X1 U6211 ( .A1(n4981), .A2(n4980), .ZN(n4995) );
  NAND2_X1 U6212 ( .A1(n4981), .A2(n4803), .ZN(n4994) );
  NAND2_X1 U6213 ( .A1(n5589), .A2(n5588), .ZN(n4804) );
  INV_X2 U6214 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4807) );
  NOR2_X2 U6215 ( .A1(n7286), .A2(n4319), .ZN(n7363) );
  NAND2_X1 U6216 ( .A1(n6957), .A2(n6956), .ZN(n7061) );
  OAI211_X1 U6217 ( .C1(n8226), .C2(n4812), .A(n4810), .B(n8210), .ZN(P2_U3160) );
  NAND2_X1 U6218 ( .A1(n8226), .A2(n4811), .ZN(n4810) );
  INV_X1 U6219 ( .A(n7364), .ZN(n4840) );
  NAND2_X1 U6220 ( .A1(n4837), .A2(n4838), .ZN(n7772) );
  NAND2_X1 U6221 ( .A1(n7364), .A2(n4841), .ZN(n4837) );
  NOR2_X1 U6222 ( .A1(n7567), .A2(n4844), .ZN(n8214) );
  AND2_X1 U6223 ( .A1(n7568), .A2(n8377), .ZN(n4844) );
  NAND2_X1 U6224 ( .A1(n9133), .A2(n4303), .ZN(n9033) );
  NAND2_X1 U6225 ( .A1(n6321), .A2(n6521), .ZN(n6556) );
  XNOR2_X1 U6226 ( .A(n6533), .B(n6687), .ZN(n6536) );
  XNOR2_X1 U6227 ( .A(n6536), .B(n6535), .ZN(n6677) );
  XNOR2_X1 U6228 ( .A(n5340), .B(n5339), .ZN(n5617) );
  CLKBUF_X1 U6229 ( .A(n8649), .Z(n8676) );
  NAND2_X1 U6230 ( .A1(n6008), .A2(n6006), .ZN(n6009) );
  NAND2_X1 U6231 ( .A1(n5671), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5660) );
  NAND2_X1 U6232 ( .A1(n8889), .A2(n8113), .ZN(n8101) );
  NAND2_X2 U6233 ( .A1(n5665), .A2(n6348), .ZN(n5656) );
  AOI21_X1 U6234 ( .B1(n6391), .B2(n6020), .A(n6019), .ZN(n8881) );
  NAND2_X1 U6235 ( .A1(n5965), .A2(n7979), .ZN(n6932) );
  AOI22_X2 U6236 ( .A1(n9441), .A2(n5533), .B1(n9154), .B2(n9445), .ZN(n9422)
         );
  AOI22_X2 U6237 ( .A1(n9318), .A2(n5541), .B1(n9170), .B2(n9330), .ZN(n9308)
         );
  OR4_X1 U6238 ( .A1(n6556), .A2(n6366), .A3(n6627), .A4(n6315), .ZN(n4850) );
  AND2_X2 U6239 ( .A1(n5550), .A2(n6520), .ZN(n9811) );
  INV_X1 U6240 ( .A(n9619), .ZN(n9795) );
  AND2_X1 U6241 ( .A1(n5550), .A2(n6621), .ZN(n9804) );
  INV_X1 U6242 ( .A(n8110), .ZN(n8051) );
  AND2_X1 U6243 ( .A1(n6053), .A2(n6052), .ZN(n9875) );
  OR2_X1 U6244 ( .A1(n9890), .A2(n6041), .ZN(n4851) );
  AND2_X2 U6245 ( .A1(n6877), .A2(n6039), .ZN(n9890) );
  INV_X1 U6246 ( .A(n9890), .ZN(n8746) );
  OR2_X1 U6247 ( .A1(n8940), .A2(n8939), .ZN(n4852) );
  NAND2_X1 U6248 ( .A1(n6622), .A2(n9471), .ZN(n9457) );
  INV_X1 U6249 ( .A(n9474), .ZN(n9405) );
  OR2_X1 U6250 ( .A1(n6008), .A2(n6006), .ZN(n4853) );
  AND2_X1 U6251 ( .A1(n7911), .A2(n7902), .ZN(n4854) );
  AND2_X1 U6252 ( .A1(n5849), .A2(n5848), .ZN(n4855) );
  AND3_X1 U6253 ( .A1(n9062), .A2(n9165), .A3(n9061), .ZN(n4856) );
  OR2_X1 U6254 ( .A1(n9214), .A2(n7131), .ZN(n4857) );
  AND2_X1 U6255 ( .A1(n4945), .A2(n4944), .ZN(n4858) );
  INV_X1 U6256 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4973) );
  NAND2_X1 U6257 ( .A1(n8610), .A2(n8608), .ZN(n4859) );
  NOR2_X1 U6258 ( .A1(n8967), .A2(n9024), .ZN(n4860) );
  OR2_X1 U6259 ( .A1(n6994), .A2(n9215), .ZN(n4861) );
  OR2_X1 U6260 ( .A1(n9212), .A2(n7308), .ZN(n4863) );
  AND2_X1 U6261 ( .A1(n4918), .A2(n4917), .ZN(n4865) );
  AND2_X1 U6262 ( .A1(n6190), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n4866) );
  NAND2_X1 U6263 ( .A1(n9795), .A2(n9801), .ZN(n9613) );
  INV_X1 U6264 ( .A(n9613), .ZN(n5547) );
  INV_X1 U6265 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4886) );
  AND2_X1 U6266 ( .A1(n4895), .A2(n4894), .ZN(n4867) );
  AND2_X1 U6267 ( .A1(n4913), .A2(n4912), .ZN(n4868) );
  AND2_X1 U6268 ( .A1(n4900), .A2(n4899), .ZN(n4869) );
  INV_X1 U6269 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n4903) );
  AND2_X1 U6270 ( .A1(n4907), .A2(n4908), .ZN(n4870) );
  INV_X1 U6271 ( .A(n9604), .ZN(n6071) );
  NAND2_X1 U6272 ( .A1(n9811), .A2(n9801), .ZN(n9548) );
  AND2_X1 U6273 ( .A1(n5598), .A2(n5597), .ZN(n8554) );
  NAND2_X1 U6274 ( .A1(n8797), .A2(n8521), .ZN(n4871) );
  NOR2_X1 U6275 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n4872) );
  AND2_X1 U6276 ( .A1(n9339), .A2(n9333), .ZN(n4873) );
  NOR2_X1 U6277 ( .A1(n5440), .A2(n5439), .ZN(n4875) );
  INV_X1 U6278 ( .A(n7484), .ZN(n5524) );
  OR2_X1 U6279 ( .A1(n8822), .A2(n8598), .ZN(n4876) );
  AND2_X1 U6280 ( .A1(n7852), .A2(n7794), .ZN(n4877) );
  AND2_X1 U6281 ( .A1(n5734), .A2(n5733), .ZN(n4878) );
  INV_X1 U6282 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U6283 ( .A1(n8108), .A2(n8103), .ZN(n8117) );
  OR2_X1 U6284 ( .A1(n7849), .A2(n8373), .ZN(n7794) );
  INV_X1 U6285 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5567) );
  INV_X1 U6286 ( .A(n8554), .ZN(n5943) );
  INV_X1 U6287 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5569) );
  OAI22_X1 U6288 ( .A1(n9058), .A2(n9775), .B1(n7017), .B2(n7121), .ZN(n6537)
         );
  INV_X1 U6289 ( .A(n9320), .ZN(n5384) );
  INV_X1 U6290 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5075) );
  NAND2_X1 U6291 ( .A1(n4901), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4885) );
  OR2_X1 U6292 ( .A1(n7801), .A2(n7800), .ZN(n7802) );
  INV_X1 U6293 ( .A(n5641), .ZN(n5582) );
  OR2_X1 U6294 ( .A1(n5789), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U6295 ( .A1(n8606), .A2(n5913), .ZN(n8593) );
  NAND2_X1 U6296 ( .A1(n7988), .A2(n7987), .ZN(n8133) );
  OAI22_X1 U6297 ( .A1(n5676), .A2(n6351), .B1(n6651), .B2(n5665), .ZN(n5655)
         );
  INV_X1 U6298 ( .A(n9022), .ZN(n9023) );
  AND2_X1 U6299 ( .A1(n5396), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5414) );
  INV_X1 U6300 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9967) );
  INV_X1 U6301 ( .A(SI_17_), .ZN(n10038) );
  NOR2_X1 U6302 ( .A1(n5736), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5735) );
  INV_X1 U6303 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5577) );
  NAND2_X1 U6304 ( .A1(n5582), .A2(n10054), .ZN(n5922) );
  AND2_X1 U6305 ( .A1(n5840), .A2(n8282), .ZN(n5859) );
  INV_X1 U6306 ( .A(n7445), .ZN(n7438) );
  INV_X1 U6307 ( .A(n8133), .ZN(n7984) );
  INV_X1 U6308 ( .A(n5655), .ZN(n5658) );
  NAND2_X1 U6309 ( .A1(n6531), .A2(n6530), .ZN(n6533) );
  OR2_X1 U6310 ( .A1(n8925), .A2(n8924), .ZN(n8926) );
  OAI22_X1 U6311 ( .A1(n9057), .A2(n9169), .B1(n5472), .B2(n6302), .ZN(n5473)
         );
  NOR2_X1 U6312 ( .A1(n5328), .A2(n9967), .ZN(n5063) );
  OR3_X1 U6313 ( .A1(n5327), .A2(n5326), .A3(n9101), .ZN(n5328) );
  AND2_X1 U6314 ( .A1(n7918), .A2(n9541), .ZN(n5482) );
  AND2_X1 U6315 ( .A1(n5476), .A2(n9203), .ZN(n5532) );
  AOI21_X1 U6316 ( .B1(n7003), .B2(n6233), .A(n5105), .ZN(n6918) );
  AOI21_X1 U6317 ( .B1(n6378), .B2(n5494), .A(n6382), .ZN(n6619) );
  AND2_X1 U6318 ( .A1(n5462), .A2(n5465), .ZN(n5458) );
  OR3_X1 U6319 ( .A1(n5238), .A2(P1_IR_REG_10__SCAN_IN), .A3(
        P1_IR_REG_11__SCAN_IN), .ZN(n5271) );
  AND2_X1 U6320 ( .A1(n7769), .A2(n8313), .ZN(n7770) );
  NAND2_X1 U6321 ( .A1(n6797), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6896) );
  NOR2_X1 U6322 ( .A1(n7028), .A2(n4298), .ZN(n7135) );
  INV_X1 U6323 ( .A(n8470), .ZN(n8441) );
  NAND2_X1 U6324 ( .A1(n5859), .A2(n5579), .ZN(n5886) );
  OR2_X1 U6325 ( .A1(n5829), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5841) );
  OR2_X1 U6326 ( .A1(n7239), .A2(n8172), .ZN(n9852) );
  INV_X1 U6327 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6006) );
  AND2_X1 U6328 ( .A1(n5345), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5006) );
  OR2_X1 U6329 ( .A1(n6548), .A2(n6556), .ZN(n6558) );
  NOR2_X1 U6330 ( .A1(n5344), .A2(n5343), .ZN(n5345) );
  OR2_X1 U6331 ( .A1(n5141), .A2(n9930), .ZN(n5108) );
  INV_X1 U6332 ( .A(n9616), .ZN(n8919) );
  INV_X1 U6333 ( .A(n9019), .ZN(n8915) );
  NAND2_X1 U6334 ( .A1(n7626), .A2(n5478), .ZN(n7789) );
  INV_X1 U6335 ( .A(n9521), .ZN(n9443) );
  AND2_X1 U6336 ( .A1(n5467), .A2(n6312), .ZN(n9412) );
  AND2_X1 U6337 ( .A1(n5351), .A2(n4972), .ZN(n5349) );
  INV_X1 U6338 ( .A(n8363), .ZN(n8339) );
  NAND2_X1 U6339 ( .A1(n6017), .A2(n6030), .ZN(n6777) );
  INV_X1 U6340 ( .A(n8503), .ZN(n8486) );
  NOR2_X1 U6341 ( .A1(n8382), .A2(n8169), .ZN(n8509) );
  INV_X1 U6342 ( .A(n9665), .ZN(n8723) );
  INV_X1 U6343 ( .A(n9670), .ZN(n8672) );
  NAND2_X1 U6344 ( .A1(n8804), .A2(n9890), .ZN(n8748) );
  AND2_X1 U6345 ( .A1(n6038), .A2(n6037), .ZN(n6039) );
  AND2_X1 U6346 ( .A1(n8129), .A2(n8128), .ZN(n8588) );
  NAND2_X1 U6347 ( .A1(n7612), .A2(n9852), .ZN(n9835) );
  OR2_X1 U6348 ( .A1(n6771), .A2(n6047), .ZN(n6053) );
  AND2_X1 U6349 ( .A1(n5836), .A2(n5826), .ZN(n8388) );
  NAND2_X1 U6350 ( .A1(n6260), .A2(n6259), .ZN(n6309) );
  AND4_X1 U6351 ( .A1(n5420), .A2(n5419), .A3(n5418), .A4(n5417), .ZN(n9168)
         );
  AND4_X1 U6352 ( .A1(n5283), .A2(n5282), .A3(n5281), .A4(n5280), .ZN(n7755)
         );
  INV_X1 U6353 ( .A(n9739), .ZN(n9726) );
  INV_X1 U6354 ( .A(n9718), .ZN(n9733) );
  INV_X1 U6355 ( .A(n9460), .ZN(n9754) );
  INV_X1 U6356 ( .A(n9412), .ZN(n9463) );
  INV_X1 U6357 ( .A(n9444), .ZN(n9762) );
  INV_X1 U6358 ( .A(n9548), .ZN(n9551) );
  NOR2_X1 U6359 ( .A1(n6481), .A2(n6479), .ZN(n6625) );
  NAND2_X1 U6360 ( .A1(n8894), .A2(n6191), .ZN(n5427) );
  NAND2_X1 U6361 ( .A1(n7647), .A2(n7657), .ZN(n9801) );
  NOR2_X1 U6362 ( .A1(n5514), .A2(n6618), .ZN(n5550) );
  AND2_X1 U6363 ( .A1(n5493), .A2(n7908), .ZN(n6378) );
  AND2_X1 U6364 ( .A1(n5305), .A2(n5304), .ZN(n9714) );
  INV_X1 U6365 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7507) );
  NAND2_X1 U6366 ( .A1(n6859), .A2(n6766), .ZN(n8363) );
  AND2_X1 U6367 ( .A1(n6770), .A2(n6769), .ZN(n8356) );
  INV_X1 U6368 ( .A(n8352), .ZN(n8368) );
  INV_X1 U6369 ( .A(n8553), .ZN(n8566) );
  INV_X1 U6370 ( .A(n8509), .ZN(n8481) );
  OR2_X1 U6371 ( .A1(n6611), .A2(n8474), .ZN(n8519) );
  INV_X1 U6372 ( .A(n9670), .ZN(n9668) );
  AND2_X1 U6373 ( .A1(n6882), .A2(n9656), .ZN(n9670) );
  INV_X1 U6374 ( .A(n6042), .ZN(n6043) );
  NAND2_X1 U6375 ( .A1(n9890), .A2(n9835), .ZN(n8796) );
  NOR2_X1 U6376 ( .A1(n8528), .A2(n6004), .ZN(n6058) );
  NAND2_X1 U6377 ( .A1(n9873), .A2(n9835), .ZN(n8878) );
  INV_X2 U6378 ( .A(n9875), .ZN(n9873) );
  INV_X1 U6379 ( .A(n6784), .ZN(n8880) );
  AND2_X1 U6380 ( .A1(n6776), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6393) );
  INV_X1 U6381 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7203) );
  XNOR2_X1 U6382 ( .A(n9033), .B(n9032), .ZN(n9040) );
  NAND2_X1 U6383 ( .A1(n9063), .A2(n4856), .ZN(n9073) );
  INV_X1 U6384 ( .A(n5476), .ZN(n9477) );
  INV_X1 U6385 ( .A(n9520), .ZN(n9401) );
  INV_X1 U6386 ( .A(n9165), .ZN(n9189) );
  AND4_X1 U6387 ( .A1(n5453), .A2(n5452), .A3(n5451), .A4(n5450), .ZN(n9065)
         );
  INV_X1 U6388 ( .A(n9079), .ZN(n9198) );
  INV_X1 U6389 ( .A(P1_U3973), .ZN(n9218) );
  NAND2_X1 U6390 ( .A1(n6369), .A2(n6333), .ZN(n9730) );
  NAND2_X1 U6391 ( .A1(n6338), .A2(n6337), .ZN(n9746) );
  OR2_X1 U6392 ( .A1(n9749), .A2(n6989), .ZN(n7655) );
  INV_X1 U6393 ( .A(n9474), .ZN(n9749) );
  OR2_X1 U6394 ( .A1(n9405), .A2(n6624), .ZN(n9444) );
  NAND2_X1 U6395 ( .A1(n9811), .A2(n9541), .ZN(n9537) );
  INV_X1 U6396 ( .A(n9811), .ZN(n9812) );
  NAND2_X1 U6397 ( .A1(n9795), .A2(n9541), .ZN(n9604) );
  INV_X1 U6398 ( .A(n9804), .ZN(n9619) );
  NOR2_X1 U6399 ( .A1(n6378), .A2(n6556), .ZN(n9771) );
  INV_X1 U6400 ( .A(n9771), .ZN(n9772) );
  INV_X1 U6401 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7904) );
  AND2_X2 U6402 ( .A1(n6484), .A2(n6321), .ZN(P1_U3973) );
  INV_X1 U6403 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U6404 ( .A1(n4901), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4880) );
  OAI21_X1 U6405 ( .B1(n4901), .B2(n4881), .A(n4880), .ZN(n4882) );
  NAND2_X1 U6406 ( .A1(n4882), .A2(SI_1_), .ZN(n4884) );
  MUX2_X1 U6407 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(P2_DATAO_REG_0__SCAN_IN), 
        .S(n4901), .Z(n4883) );
  NAND2_X1 U6408 ( .A1(n4883), .A2(SI_0_), .ZN(n5089) );
  INV_X1 U6409 ( .A(n4888), .ZN(n4887) );
  INV_X1 U6410 ( .A(SI_2_), .ZN(n9924) );
  NAND2_X1 U6411 ( .A1(n4887), .A2(n9924), .ZN(n4889) );
  NAND2_X1 U6412 ( .A1(n4888), .A2(SI_2_), .ZN(n4890) );
  NAND2_X1 U6413 ( .A1(n5114), .A2(n5113), .ZN(n5116) );
  NAND2_X1 U6414 ( .A1(n5116), .A2(n4890), .ZN(n5126) );
  MUX2_X1 U6415 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n4901), .Z(n4891) );
  NAND2_X1 U6416 ( .A1(n4891), .A2(SI_3_), .ZN(n4895) );
  INV_X1 U6417 ( .A(n4891), .ZN(n4893) );
  INV_X1 U6418 ( .A(SI_3_), .ZN(n4892) );
  NAND2_X1 U6419 ( .A1(n4893), .A2(n4892), .ZN(n4894) );
  NAND2_X1 U6420 ( .A1(n5126), .A2(n4867), .ZN(n5128) );
  NAND2_X1 U6421 ( .A1(n5128), .A2(n4895), .ZN(n5146) );
  MUX2_X1 U6422 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n4901), .Z(n4896) );
  NAND2_X1 U6423 ( .A1(n4896), .A2(SI_4_), .ZN(n4900) );
  INV_X1 U6424 ( .A(n4896), .ZN(n4898) );
  INV_X1 U6425 ( .A(SI_4_), .ZN(n4897) );
  NAND2_X1 U6426 ( .A1(n4898), .A2(n4897), .ZN(n4899) );
  NAND2_X1 U6427 ( .A1(n5146), .A2(n4869), .ZN(n5148) );
  NAND2_X1 U6428 ( .A1(n5148), .A2(n4900), .ZN(n5165) );
  INV_X1 U6429 ( .A(n4906), .ZN(n4905) );
  INV_X1 U6430 ( .A(SI_5_), .ZN(n4904) );
  NAND2_X1 U6431 ( .A1(n4905), .A2(n4904), .ZN(n4907) );
  NAND2_X1 U6432 ( .A1(n4906), .A2(SI_5_), .ZN(n4908) );
  MUX2_X1 U6433 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6348), .Z(n4909) );
  NAND2_X1 U6434 ( .A1(n4909), .A2(SI_6_), .ZN(n4913) );
  INV_X1 U6435 ( .A(n4909), .ZN(n4911) );
  INV_X1 U6436 ( .A(SI_6_), .ZN(n4910) );
  NAND2_X1 U6437 ( .A1(n4911), .A2(n4910), .ZN(n4912) );
  MUX2_X1 U6438 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6348), .Z(n4914) );
  NAND2_X1 U6439 ( .A1(n4914), .A2(SI_7_), .ZN(n4918) );
  INV_X1 U6440 ( .A(n4914), .ZN(n4916) );
  INV_X1 U6441 ( .A(SI_7_), .ZN(n4915) );
  NAND2_X1 U6442 ( .A1(n4916), .A2(n4915), .ZN(n4917) );
  MUX2_X1 U6443 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n6348), .Z(n4919) );
  INV_X1 U6444 ( .A(n4919), .ZN(n4921) );
  INV_X1 U6445 ( .A(SI_8_), .ZN(n4920) );
  NAND2_X1 U6446 ( .A1(n4921), .A2(n4920), .ZN(n4922) );
  INV_X1 U6447 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n4923) );
  MUX2_X1 U6448 ( .A(n6388), .B(n4923), .S(n6348), .Z(n4924) );
  XNOR2_X1 U6449 ( .A(n4924), .B(SI_9_), .ZN(n5219) );
  INV_X1 U6450 ( .A(n4924), .ZN(n4925) );
  NOR2_X1 U6451 ( .A1(n4925), .A2(SI_9_), .ZN(n4926) );
  MUX2_X1 U6452 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6348), .Z(n4927) );
  NAND2_X1 U6453 ( .A1(n4927), .A2(SI_10_), .ZN(n4932) );
  INV_X1 U6454 ( .A(n4927), .ZN(n4929) );
  INV_X1 U6455 ( .A(SI_10_), .ZN(n4928) );
  NAND2_X1 U6456 ( .A1(n4929), .A2(n4928), .ZN(n4930) );
  NAND2_X1 U6457 ( .A1(n4932), .A2(n4930), .ZN(n5234) );
  INV_X1 U6458 ( .A(n5234), .ZN(n4931) );
  MUX2_X1 U6459 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6348), .Z(n4934) );
  XNOR2_X1 U6460 ( .A(n4934), .B(SI_11_), .ZN(n5252) );
  INV_X1 U6461 ( .A(n5252), .ZN(n4933) );
  INV_X1 U6462 ( .A(n4934), .ZN(n4936) );
  INV_X1 U6463 ( .A(SI_11_), .ZN(n4935) );
  NAND2_X1 U6464 ( .A1(n4936), .A2(n4935), .ZN(n4937) );
  MUX2_X1 U6465 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6348), .Z(n4938) );
  NAND2_X1 U6466 ( .A1(n4938), .A2(SI_12_), .ZN(n4940) );
  OAI21_X1 U6467 ( .B1(n4938), .B2(SI_12_), .A(n4940), .ZN(n5267) );
  NAND2_X1 U6468 ( .A1(n5269), .A2(n4940), .ZN(n5284) );
  MUX2_X1 U6469 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6348), .Z(n4941) );
  INV_X1 U6470 ( .A(n4941), .ZN(n4943) );
  INV_X1 U6471 ( .A(SI_13_), .ZN(n4942) );
  NAND2_X1 U6472 ( .A1(n4943), .A2(n4942), .ZN(n4944) );
  MUX2_X1 U6473 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6348), .Z(n5300) );
  MUX2_X1 U6474 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6348), .Z(n5070) );
  MUX2_X1 U6475 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n6348), .Z(n5318) );
  NAND2_X1 U6476 ( .A1(n5318), .A2(SI_16_), .ZN(n4946) );
  MUX2_X1 U6477 ( .A(n7203), .B(n7205), .S(n6348), .Z(n4947) );
  INV_X1 U6478 ( .A(n4947), .ZN(n4948) );
  NAND2_X1 U6479 ( .A1(n4948), .A2(SI_17_), .ZN(n4949) );
  NAND2_X1 U6480 ( .A1(n4950), .A2(n4949), .ZN(n5057) );
  MUX2_X1 U6481 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6348), .Z(n4952) );
  XNOR2_X1 U6482 ( .A(n4952), .B(SI_18_), .ZN(n5041) );
  NAND2_X1 U6483 ( .A1(n4952), .A2(SI_18_), .ZN(n4953) );
  MUX2_X1 U6484 ( .A(n7405), .B(n8212), .S(n6348), .Z(n4955) );
  INV_X1 U6485 ( .A(n4955), .ZN(n4956) );
  NAND2_X1 U6486 ( .A1(n4956), .A2(SI_19_), .ZN(n4957) );
  NAND2_X1 U6487 ( .A1(n4958), .A2(n4957), .ZN(n5023) );
  INV_X1 U6488 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7549) );
  MUX2_X1 U6489 ( .A(n7498), .B(n7549), .S(n6348), .Z(n5012) );
  OAI21_X1 U6490 ( .B1(n5016), .B2(n5013), .A(n5012), .ZN(n4960) );
  NAND2_X1 U6491 ( .A1(n5016), .A2(n5013), .ZN(n4959) );
  MUX2_X1 U6492 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n6348), .Z(n5337) );
  NOR2_X1 U6493 ( .A1(n5337), .A2(SI_21_), .ZN(n4962) );
  NAND2_X1 U6494 ( .A1(n5337), .A2(SI_21_), .ZN(n4961) );
  MUX2_X1 U6495 ( .A(n9968), .B(n7748), .S(n6348), .Z(n4964) );
  INV_X1 U6496 ( .A(SI_22_), .ZN(n4963) );
  NAND2_X1 U6497 ( .A1(n4964), .A2(n4963), .ZN(n4967) );
  INV_X1 U6498 ( .A(n4964), .ZN(n4965) );
  NAND2_X1 U6499 ( .A1(n4965), .A2(SI_22_), .ZN(n4966) );
  NAND2_X1 U6500 ( .A1(n4967), .A2(n4966), .ZN(n5001) );
  INV_X1 U6501 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7753) );
  INV_X1 U6502 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n4968) );
  MUX2_X1 U6503 ( .A(n7753), .B(n4968), .S(n6348), .Z(n4970) );
  INV_X1 U6504 ( .A(SI_23_), .ZN(n4969) );
  NAND2_X1 U6505 ( .A1(n4970), .A2(n4969), .ZN(n5351) );
  INV_X1 U6506 ( .A(n4970), .ZN(n4971) );
  NAND2_X1 U6507 ( .A1(n4971), .A2(SI_23_), .ZN(n4972) );
  XNOR2_X1 U6508 ( .A(n5350), .B(n5349), .ZN(n7750) );
  NOR2_X1 U6509 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n4976) );
  NOR2_X1 U6510 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n4975) );
  NOR2_X1 U6511 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4974) );
  NAND4_X1 U6512 ( .A1(n5168), .A2(n10035), .A3(n5239), .A4(n5075), .ZN(n4977)
         );
  NOR2_X1 U6513 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n4978) );
  INV_X1 U6514 ( .A(n4982), .ZN(n4981) );
  NAND2_X1 U6515 ( .A1(n4982), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4983) );
  NAND2_X2 U6516 ( .A1(n4995), .A2(n4984), .ZN(n6366) );
  XNOR2_X2 U6517 ( .A(n4986), .B(n4985), .ZN(n6489) );
  NAND2_X1 U6518 ( .A1(n7750), .A2(n6191), .ZN(n4988) );
  NAND2_X4 U6519 ( .A1(n6329), .A2(n6345), .ZN(n5322) );
  NAND2_X1 U6520 ( .A1(n6190), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n4987) );
  AND2_X1 U6521 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5138) );
  NAND2_X1 U6522 ( .A1(n5214), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U6523 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n4989) );
  NAND2_X1 U6524 ( .A1(n5245), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5260) );
  INV_X1 U6525 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5326) );
  AND2_X1 U6526 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n4990) );
  NAND2_X1 U6527 ( .A1(n5063), .A2(n4990), .ZN(n5033) );
  INV_X1 U6528 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5343) );
  OR2_X1 U6529 ( .A1(n5006), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n4991) );
  NAND2_X1 U6530 ( .A1(n5006), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5360) );
  AND2_X1 U6531 ( .A1(n4991), .A2(n5360), .ZN(n9357) );
  INV_X1 U6532 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9583) );
  NAND2_X1 U6533 ( .A1(n5137), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n4999) );
  NAND2_X1 U6534 ( .A1(n6193), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n4998) );
  OAI211_X1 U6535 ( .C1(n6196), .C2(n9583), .A(n4999), .B(n4998), .ZN(n5000)
         );
  OR2_X1 U6536 ( .A1(n5475), .A2(n9137), .ZN(n6147) );
  NAND2_X1 U6537 ( .A1(n5475), .A2(n9137), .ZN(n9333) );
  XNOR2_X1 U6538 ( .A(n5002), .B(n5001), .ZN(n7746) );
  NAND2_X1 U6539 ( .A1(n7746), .A2(n6191), .ZN(n5004) );
  NAND2_X1 U6540 ( .A1(n6190), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5003) );
  NOR2_X1 U6541 ( .A1(n5345), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5005) );
  NOR2_X1 U6542 ( .A1(n5006), .A2(n5005), .ZN(n9371) );
  NAND2_X1 U6543 ( .A1(n9371), .A2(n5051), .ZN(n5011) );
  INV_X1 U6544 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9587) );
  NAND2_X1 U6545 ( .A1(n5137), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5008) );
  NAND2_X1 U6546 ( .A1(n6193), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5007) );
  OAI211_X1 U6547 ( .C1(n6196), .C2(n9587), .A(n5008), .B(n5007), .ZN(n5009)
         );
  INV_X1 U6548 ( .A(n5009), .ZN(n5010) );
  XNOR2_X1 U6549 ( .A(n9513), .B(n9198), .ZN(n9364) );
  INV_X1 U6550 ( .A(n5012), .ZN(n5014) );
  XNOR2_X1 U6551 ( .A(n5014), .B(n5013), .ZN(n5015) );
  XNOR2_X1 U6552 ( .A(n5016), .B(n5015), .ZN(n7497) );
  NAND2_X1 U6553 ( .A1(n7497), .A2(n6191), .ZN(n5018) );
  NAND2_X1 U6554 ( .A1(n6190), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5017) );
  NAND2_X1 U6555 ( .A1(n5033), .A2(n9996), .ZN(n5019) );
  AND2_X1 U6556 ( .A1(n5344), .A2(n5019), .ZN(n9398) );
  NAND2_X1 U6557 ( .A1(n9398), .A2(n5051), .ZN(n5022) );
  AOI22_X1 U6558 ( .A1(n5446), .A2(P1_REG0_REG_20__SCAN_IN), .B1(n6193), .B2(
        P1_REG1_REG_20__SCAN_IN), .ZN(n5021) );
  NAND2_X1 U6559 ( .A1(n5137), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5020) );
  OR2_X1 U6560 ( .A1(n9520), .A2(n9078), .ZN(n6078) );
  NAND2_X1 U6561 ( .A1(n9520), .A2(n9078), .ZN(n6077) );
  NAND2_X1 U6562 ( .A1(n6078), .A2(n6077), .ZN(n6247) );
  XNOR2_X1 U6563 ( .A(n5024), .B(n5023), .ZN(n7403) );
  NAND2_X1 U6564 ( .A1(n7403), .A2(n6191), .ZN(n5030) );
  OR2_X1 U6565 ( .A1(n9621), .A2(n5456), .ZN(n5027) );
  OAI22_X1 U6566 ( .A1(n5322), .A2(n8212), .B1(n9268), .B2(n6329), .ZN(n5028)
         );
  INV_X1 U6567 ( .A(n5028), .ZN(n5029) );
  NAND2_X1 U6568 ( .A1(n5063), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5032) );
  INV_X1 U6569 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5031) );
  NAND2_X1 U6570 ( .A1(n5032), .A2(n5031), .ZN(n5034) );
  NAND2_X1 U6571 ( .A1(n5034), .A2(n5033), .ZN(n9415) );
  OR2_X1 U6572 ( .A1(n9415), .A2(n5141), .ZN(n5040) );
  INV_X1 U6573 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9530) );
  OR2_X1 U6574 ( .A1(n5447), .A2(n9530), .ZN(n5037) );
  INV_X1 U6575 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9596) );
  OR2_X1 U6576 ( .A1(n6196), .A2(n9596), .ZN(n5036) );
  AND2_X1 U6577 ( .A1(n5037), .A2(n5036), .ZN(n5039) );
  NAND2_X1 U6578 ( .A1(n5137), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5038) );
  OR2_X1 U6579 ( .A1(n9529), .A2(n9152), .ZN(n6136) );
  NAND2_X1 U6580 ( .A1(n9529), .A2(n9152), .ZN(n6293) );
  INV_X1 U6581 ( .A(n5041), .ZN(n5042) );
  XNOR2_X1 U6582 ( .A(n5043), .B(n5042), .ZN(n7296) );
  NAND2_X1 U6583 ( .A1(n7296), .A2(n6191), .ZN(n5049) );
  INV_X1 U6584 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7297) );
  NAND2_X1 U6585 ( .A1(n5044), .A2(n5456), .ZN(n5046) );
  OR2_X1 U6586 ( .A1(n5044), .A2(n5456), .ZN(n5045) );
  NAND2_X1 U6587 ( .A1(n5046), .A2(n5045), .ZN(n9738) );
  OAI22_X1 U6588 ( .A1(n5322), .A2(n7297), .B1(n6329), .B2(n9738), .ZN(n5047)
         );
  INV_X1 U6589 ( .A(n5047), .ZN(n5048) );
  INV_X1 U6590 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5050) );
  XNOR2_X1 U6591 ( .A(n5063), .B(n5050), .ZN(n9435) );
  NAND2_X1 U6592 ( .A1(n9435), .A2(n5051), .ZN(n5056) );
  INV_X1 U6593 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9534) );
  OR2_X1 U6594 ( .A1(n5447), .A2(n9534), .ZN(n5053) );
  INV_X1 U6595 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10055) );
  OR2_X1 U6596 ( .A1(n4266), .A2(n10055), .ZN(n5052) );
  AND2_X1 U6597 ( .A1(n5053), .A2(n5052), .ZN(n5055) );
  NAND2_X1 U6598 ( .A1(n5446), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5054) );
  NAND2_X1 U6599 ( .A1(n9434), .A2(n9110), .ZN(n6135) );
  XNOR2_X1 U6600 ( .A(n5058), .B(n5057), .ZN(n7202) );
  NAND2_X1 U6601 ( .A1(n7202), .A2(n6191), .ZN(n5062) );
  XNOR2_X1 U6602 ( .A(n5059), .B(n5457), .ZN(n9260) );
  OAI22_X1 U6603 ( .A1(n5322), .A2(n7205), .B1(n6329), .B2(n9260), .ZN(n5060)
         );
  INV_X1 U6604 ( .A(n5060), .ZN(n5061) );
  AND2_X1 U6605 ( .A1(n5328), .A2(n9967), .ZN(n5064) );
  OR2_X1 U6606 ( .A1(n5064), .A2(n5063), .ZN(n9446) );
  NAND2_X1 U6607 ( .A1(n5137), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5065) );
  OAI21_X1 U6608 ( .B1(n9446), .B2(n5141), .A(n5065), .ZN(n5068) );
  INV_X1 U6609 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9607) );
  INV_X1 U6610 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9542) );
  OR2_X1 U6611 ( .A1(n5447), .A2(n9542), .ZN(n5066) );
  OAI21_X1 U6612 ( .B1(n6196), .B2(n9607), .A(n5066), .ZN(n5067) );
  INV_X1 U6613 ( .A(n9154), .ZN(n9202) );
  XNOR2_X1 U6614 ( .A(n9540), .B(n9202), .ZN(n9452) );
  XNOR2_X1 U6615 ( .A(n5070), .B(SI_15_), .ZN(n5071) );
  XNOR2_X1 U6616 ( .A(n5069), .B(n5071), .ZN(n6845) );
  NAND2_X1 U6617 ( .A1(n6845), .A2(n6191), .ZN(n5081) );
  INV_X1 U6618 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9925) );
  NAND4_X1 U6619 ( .A1(n5168), .A2(n10035), .A3(n5190), .A4(n5193), .ZN(n5074)
         );
  NOR2_X1 U6620 ( .A1(n5073), .A2(n5074), .ZN(n5220) );
  NAND2_X1 U6621 ( .A1(n5220), .A2(n5075), .ZN(n5238) );
  NOR2_X1 U6622 ( .A1(n5271), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5288) );
  NAND2_X1 U6623 ( .A1(n5288), .A2(n9928), .ZN(n5076) );
  NAND2_X1 U6624 ( .A1(n5076), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5303) );
  INV_X1 U6625 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5302) );
  NAND2_X1 U6626 ( .A1(n5303), .A2(n5302), .ZN(n5305) );
  NAND2_X1 U6627 ( .A1(n5305), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5078) );
  INV_X1 U6628 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5077) );
  XNOR2_X1 U6629 ( .A(n5078), .B(n5077), .ZN(n9717) );
  OAI22_X1 U6630 ( .A1(n5322), .A2(n9925), .B1(n9717), .B2(n6329), .ZN(n5079)
         );
  INV_X1 U6631 ( .A(n5079), .ZN(n5080) );
  NAND2_X1 U6632 ( .A1(n5446), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5085) );
  INV_X1 U6633 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10024) );
  OR2_X1 U6634 ( .A1(n5447), .A2(n10024), .ZN(n5084) );
  XNOR2_X1 U6635 ( .A(n5327), .B(n5326), .ZN(n9185) );
  OR2_X1 U6636 ( .A1(n5141), .A2(n9185), .ZN(n5083) );
  INV_X1 U6637 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7887) );
  OR2_X1 U6638 ( .A1(n4266), .A2(n7887), .ZN(n5082) );
  NAND2_X1 U6639 ( .A1(n9616), .A2(n9098), .ZN(n6279) );
  NAND2_X1 U6640 ( .A1(n6283), .A2(n6279), .ZN(n7891) );
  INV_X1 U6641 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6339) );
  INV_X1 U6642 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5086) );
  INV_X1 U6643 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5087) );
  INV_X1 U6644 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5088) );
  INV_X1 U6645 ( .A(n5089), .ZN(n5090) );
  INV_X1 U6646 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6360) );
  NOR2_X1 U6647 ( .A1(n6348), .A2(n6360), .ZN(n5091) );
  AOI21_X1 U6648 ( .B1(n6351), .B2(n6348), .A(n5091), .ZN(n5092) );
  OR2_X1 U6649 ( .A1(n6366), .A2(n5092), .ZN(n5095) );
  INV_X1 U6650 ( .A(n6489), .ZN(n9635) );
  NAND2_X1 U6651 ( .A1(n6345), .A2(n6360), .ZN(n5093) );
  OAI211_X1 U6652 ( .C1(n6351), .C2(n6345), .A(n9635), .B(n5093), .ZN(n5094)
         );
  OAI211_X2 U6653 ( .C1(n6329), .C2(n6401), .A(n5095), .B(n5094), .ZN(n9761)
         );
  XNOR2_X2 U6654 ( .A(n5104), .B(n9761), .ZN(n7003) );
  NAND2_X1 U6655 ( .A1(n5137), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5101) );
  INV_X1 U6656 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6327) );
  OR2_X1 U6657 ( .A1(n5447), .A2(n6327), .ZN(n5100) );
  INV_X1 U6658 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5096) );
  OR2_X1 U6659 ( .A1(n6196), .A2(n5096), .ZN(n5099) );
  INV_X1 U6660 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5097) );
  INV_X1 U6661 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6486) );
  NAND2_X1 U6662 ( .A1(n6348), .A2(SI_0_), .ZN(n5103) );
  INV_X1 U6663 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5102) );
  XNOR2_X1 U6664 ( .A(n5103), .B(n5102), .ZN(n9639) );
  MUX2_X1 U6665 ( .A(n6486), .B(n9639), .S(n6329), .Z(n6487) );
  NOR2_X1 U6666 ( .A1(n9219), .A2(n6487), .ZN(n6233) );
  NOR2_X1 U6667 ( .A1(n6559), .A2(n7051), .ZN(n5105) );
  NAND2_X1 U6668 ( .A1(n6193), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5111) );
  INV_X1 U6669 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5106) );
  OR2_X1 U6670 ( .A1(n4266), .A2(n5106), .ZN(n5110) );
  INV_X1 U6671 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5107) );
  OR2_X1 U6672 ( .A1(n6196), .A2(n5107), .ZN(n5109) );
  INV_X1 U6673 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9930) );
  INV_X1 U6674 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6363) );
  OR2_X1 U6675 ( .A1(n5322), .A2(n6363), .ZN(n5118) );
  OR2_X1 U6676 ( .A1(n5112), .A2(n9621), .ZN(n5131) );
  OR2_X1 U6677 ( .A1(n5114), .A2(n5113), .ZN(n5115) );
  NAND2_X1 U6678 ( .A1(n5116), .A2(n5115), .ZN(n6362) );
  NAND2_X1 U6679 ( .A1(n5118), .A2(n5117), .ZN(n5477) );
  NAND2_X1 U6680 ( .A1(n7017), .A2(n5477), .ZN(n5520) );
  INV_X1 U6681 ( .A(n7017), .ZN(n9217) );
  NAND2_X1 U6682 ( .A1(n6193), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5125) );
  OR2_X1 U6683 ( .A1(n5141), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5124) );
  INV_X1 U6684 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5119) );
  OR2_X1 U6685 ( .A1(n4266), .A2(n5119), .ZN(n5123) );
  INV_X1 U6686 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5121) );
  OR2_X1 U6687 ( .A1(n6196), .A2(n5121), .ZN(n5122) );
  OR2_X1 U6688 ( .A1(n5126), .A2(n4867), .ZN(n5127) );
  NAND2_X1 U6689 ( .A1(n5128), .A2(n5127), .ZN(n6350) );
  INV_X1 U6690 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5129) );
  INV_X1 U6691 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5130) );
  NAND2_X1 U6692 ( .A1(n5131), .A2(n5130), .ZN(n5132) );
  NAND2_X1 U6693 ( .A1(n5132), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5133) );
  XNOR2_X1 U6694 ( .A(n5133), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6433) );
  NAND2_X1 U6695 ( .A1(n5256), .A2(n6433), .ZN(n5134) );
  OAI211_X1 U6696 ( .C1(n5287), .C2(n6350), .A(n5135), .B(n5134), .ZN(n9747)
         );
  NAND2_X1 U6697 ( .A1(n6690), .A2(n9747), .ZN(n6084) );
  INV_X2 U6698 ( .A(n9747), .ZN(n7055) );
  NAND2_X1 U6699 ( .A1(n5446), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5145) );
  INV_X1 U6700 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5136) );
  OR2_X1 U6701 ( .A1(n5447), .A2(n5136), .ZN(n5144) );
  INV_X1 U6702 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6992) );
  OR2_X1 U6703 ( .A1(n4266), .A2(n6992), .ZN(n5143) );
  INV_X1 U6704 ( .A(n5138), .ZN(n5158) );
  INV_X1 U6705 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5139) );
  INV_X1 U6706 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9748) );
  NAND2_X1 U6707 ( .A1(n5139), .A2(n9748), .ZN(n5140) );
  NAND2_X1 U6708 ( .A1(n5158), .A2(n5140), .ZN(n6991) );
  OR2_X1 U6709 ( .A1(n5141), .A2(n6991), .ZN(n5142) );
  OR2_X1 U6710 ( .A1(n5146), .A2(n4869), .ZN(n5147) );
  NAND2_X1 U6711 ( .A1(n5148), .A2(n5147), .ZN(n6354) );
  INV_X1 U6712 ( .A(n6354), .ZN(n5149) );
  NAND2_X1 U6713 ( .A1(n5149), .A2(n6191), .ZN(n5154) );
  INV_X1 U6714 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6355) );
  NAND2_X1 U6715 ( .A1(n5150), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5151) );
  XNOR2_X1 U6716 ( .A(n5151), .B(n4973), .ZN(n6501) );
  OAI22_X1 U6717 ( .A1(n5322), .A2(n6355), .B1(n6329), .B2(n6501), .ZN(n5152)
         );
  INV_X1 U6718 ( .A(n5152), .ZN(n5153) );
  NAND2_X1 U6719 ( .A1(n9215), .A2(n7092), .ZN(n6262) );
  NAND2_X1 U6720 ( .A1(n6982), .A2(n6262), .ZN(n7072) );
  NAND2_X1 U6721 ( .A1(n5446), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5164) );
  INV_X1 U6722 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5155) );
  OR2_X1 U6723 ( .A1(n5447), .A2(n5155), .ZN(n5163) );
  INV_X1 U6724 ( .A(n5156), .ZN(n5181) );
  INV_X1 U6725 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5157) );
  NAND2_X1 U6726 ( .A1(n5158), .A2(n5157), .ZN(n5159) );
  NAND2_X1 U6727 ( .A1(n5181), .A2(n5159), .ZN(n7134) );
  OR2_X1 U6728 ( .A1(n5141), .A2(n7134), .ZN(n5162) );
  INV_X1 U6729 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5160) );
  OR2_X1 U6730 ( .A1(n4266), .A2(n5160), .ZN(n5161) );
  OR2_X1 U6731 ( .A1(n5165), .A2(n4870), .ZN(n5166) );
  NAND2_X1 U6732 ( .A1(n5167), .A2(n5166), .ZN(n6364) );
  OR2_X1 U6733 ( .A1(n6364), .A2(n5287), .ZN(n5172) );
  INV_X1 U6734 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6365) );
  NAND2_X1 U6735 ( .A1(n5073), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5169) );
  XNOR2_X1 U6736 ( .A(n5169), .B(n5168), .ZN(n6403) );
  OAI22_X1 U6737 ( .A1(n5322), .A2(n6365), .B1(n6329), .B2(n6403), .ZN(n5170)
         );
  INV_X1 U6738 ( .A(n5170), .ZN(n5171) );
  NAND2_X1 U6739 ( .A1(n5172), .A2(n5171), .ZN(n7131) );
  NAND2_X1 U6740 ( .A1(n7196), .A2(n7131), .ZN(n6087) );
  INV_X1 U6741 ( .A(n7131), .ZN(n7103) );
  NAND2_X1 U6742 ( .A1(n7103), .A2(n9214), .ZN(n6264) );
  NAND2_X1 U6743 ( .A1(n6087), .A2(n6264), .ZN(n7079) );
  NOR2_X1 U6744 ( .A1(n7079), .A2(n5522), .ZN(n5173) );
  NAND2_X1 U6745 ( .A1(n7072), .A2(n5173), .ZN(n7069) );
  NAND2_X1 U6746 ( .A1(n7069), .A2(n6264), .ZN(n7175) );
  OR2_X1 U6747 ( .A1(n5174), .A2(n4868), .ZN(n5175) );
  NAND2_X1 U6748 ( .A1(n5176), .A2(n5175), .ZN(n6356) );
  OR2_X1 U6749 ( .A1(n6356), .A2(n5287), .ZN(n5179) );
  INV_X1 U6750 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6357) );
  OAI21_X1 U6751 ( .B1(n5073), .B2(P1_IR_REG_5__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5191) );
  XNOR2_X1 U6752 ( .A(n5191), .B(n5190), .ZN(n6414) );
  OAI22_X1 U6753 ( .A1(n5322), .A2(n6357), .B1(n6329), .B2(n6414), .ZN(n5177)
         );
  INV_X1 U6754 ( .A(n5177), .ZN(n5178) );
  NAND2_X1 U6755 ( .A1(n5179), .A2(n5178), .ZN(n7210) );
  NAND2_X1 U6756 ( .A1(n5446), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5188) );
  INV_X1 U6757 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6404) );
  OR2_X1 U6758 ( .A1(n5447), .A2(n6404), .ZN(n5187) );
  INV_X1 U6759 ( .A(n5214), .ZN(n5183) );
  INV_X1 U6760 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5180) );
  NAND2_X1 U6761 ( .A1(n5181), .A2(n5180), .ZN(n5182) );
  NAND2_X1 U6762 ( .A1(n5183), .A2(n5182), .ZN(n7192) );
  OR2_X1 U6763 ( .A1(n5141), .A2(n7192), .ZN(n5186) );
  INV_X1 U6764 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5184) );
  OR2_X1 U6765 ( .A1(n4266), .A2(n5184), .ZN(n5185) );
  NAND2_X1 U6766 ( .A1(n7210), .A2(n7211), .ZN(n6236) );
  NAND2_X1 U6767 ( .A1(n6372), .A2(n6191), .ZN(n5197) );
  INV_X1 U6768 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6375) );
  NAND2_X1 U6769 ( .A1(n5191), .A2(n5190), .ZN(n5192) );
  NAND2_X1 U6770 ( .A1(n5192), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5207) );
  NAND2_X1 U6771 ( .A1(n5207), .A2(n10035), .ZN(n5209) );
  NAND2_X1 U6772 ( .A1(n5209), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5194) );
  XNOR2_X1 U6773 ( .A(n5194), .B(n5193), .ZN(n6569) );
  OAI22_X1 U6774 ( .A1(n5322), .A2(n6375), .B1(n6329), .B2(n6569), .ZN(n5195)
         );
  INV_X1 U6775 ( .A(n5195), .ZN(n5196) );
  NAND2_X1 U6776 ( .A1(n6193), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5203) );
  INV_X1 U6777 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5198) );
  OR2_X1 U6778 ( .A1(n4266), .A2(n5198), .ZN(n5202) );
  INV_X1 U6779 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7491) );
  XNOR2_X1 U6780 ( .A(n5224), .B(n7491), .ZN(n7278) );
  OR2_X1 U6781 ( .A1(n5141), .A2(n7278), .ZN(n5201) );
  INV_X1 U6782 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5199) );
  OR2_X1 U6783 ( .A1(n6196), .A2(n5199), .ZN(n5200) );
  NAND2_X1 U6784 ( .A1(n7484), .A2(n7485), .ZN(n6098) );
  OR2_X1 U6785 ( .A1(n5204), .A2(n4865), .ZN(n5205) );
  NAND2_X1 U6786 ( .A1(n5206), .A2(n5205), .ZN(n6358) );
  OR2_X1 U6787 ( .A1(n6358), .A2(n5287), .ZN(n5212) );
  INV_X1 U6788 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6359) );
  OR2_X1 U6789 ( .A1(n5207), .A2(n10035), .ZN(n5208) );
  NAND2_X1 U6790 ( .A1(n5209), .A2(n5208), .ZN(n6454) );
  OAI22_X1 U6791 ( .A1(n5322), .A2(n6359), .B1(n6329), .B2(n6454), .ZN(n5210)
         );
  INV_X1 U6792 ( .A(n5210), .ZN(n5211) );
  NAND2_X1 U6793 ( .A1(n5212), .A2(n5211), .ZN(n7308) );
  NAND2_X1 U6794 ( .A1(n5446), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5218) );
  INV_X1 U6795 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5213) );
  OR2_X1 U6796 ( .A1(n5447), .A2(n5213), .ZN(n5217) );
  OAI21_X1 U6797 ( .B1(n5214), .B2(P1_REG3_REG_7__SCAN_IN), .A(n5224), .ZN(
        n7306) );
  OR2_X1 U6798 ( .A1(n5141), .A2(n7306), .ZN(n5216) );
  INV_X1 U6799 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7183) );
  OR2_X1 U6800 ( .A1(n4266), .A2(n7183), .ZN(n5215) );
  NAND2_X1 U6801 ( .A1(n7308), .A2(n7298), .ZN(n7260) );
  NAND2_X1 U6802 ( .A1(n6098), .A2(n7260), .ZN(n6093) );
  OR2_X1 U6803 ( .A1(n7484), .A2(n7485), .ZN(n7325) );
  NAND2_X1 U6804 ( .A1(n6384), .A2(n6191), .ZN(n5223) );
  OR2_X1 U6805 ( .A1(n5220), .A2(n9621), .ZN(n5221) );
  XNOR2_X1 U6806 ( .A(n5221), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7392) );
  AOI22_X1 U6807 ( .A1(n6190), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5256), .B2(
        n7392), .ZN(n5222) );
  NAND2_X1 U6808 ( .A1(n6193), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5231) );
  INV_X1 U6809 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7332) );
  OR2_X1 U6810 ( .A1(n4266), .A2(n7332), .ZN(n5230) );
  INV_X1 U6811 ( .A(n5224), .ZN(n5225) );
  AOI21_X1 U6812 ( .B1(n5225), .B2(P1_REG3_REG_8__SCAN_IN), .A(
        P1_REG3_REG_9__SCAN_IN), .ZN(n5226) );
  OR2_X1 U6813 ( .A1(n5226), .A2(n5245), .ZN(n7562) );
  OR2_X1 U6814 ( .A1(n5141), .A2(n7562), .ZN(n5229) );
  INV_X1 U6815 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n5227) );
  OR2_X1 U6816 ( .A1(n6196), .A2(n5227), .ZN(n5228) );
  OR2_X1 U6817 ( .A1(n7564), .A2(n7554), .ZN(n6106) );
  NAND2_X1 U6818 ( .A1(n7324), .A2(n6106), .ZN(n5232) );
  NAND2_X1 U6819 ( .A1(n7564), .A2(n7554), .ZN(n6107) );
  INV_X1 U6820 ( .A(n5233), .ZN(n5235) );
  NAND2_X1 U6821 ( .A1(n5235), .A2(n5234), .ZN(n5236) );
  NAND2_X1 U6822 ( .A1(n5237), .A2(n5236), .ZN(n6387) );
  OR2_X1 U6823 ( .A1(n6387), .A2(n5287), .ZN(n5243) );
  NAND2_X1 U6824 ( .A1(n5238), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5240) );
  NAND2_X1 U6825 ( .A1(n5240), .A2(n5239), .ZN(n5254) );
  OR2_X1 U6826 ( .A1(n5240), .A2(n5239), .ZN(n5241) );
  AOI22_X1 U6827 ( .A1(n6190), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5256), .B2(
        n9649), .ZN(n5242) );
  NAND2_X1 U6828 ( .A1(n6193), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5250) );
  INV_X1 U6829 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5244) );
  OR2_X1 U6830 ( .A1(n6196), .A2(n5244), .ZN(n5249) );
  OR2_X1 U6831 ( .A1(n5245), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5246) );
  NAND2_X1 U6832 ( .A1(n5260), .A2(n5246), .ZN(n7598) );
  OR2_X1 U6833 ( .A1(n5141), .A2(n7598), .ZN(n5248) );
  INV_X1 U6834 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7429) );
  OR2_X1 U6835 ( .A1(n4266), .A2(n7429), .ZN(n5247) );
  NAND4_X1 U6836 ( .A1(n5250), .A2(n5249), .A3(n5248), .A4(n5247), .ZN(n9209)
         );
  AND2_X1 U6837 ( .A1(n9792), .A2(n9209), .ZN(n6268) );
  INV_X1 U6838 ( .A(n9209), .ZN(n7644) );
  NAND2_X1 U6839 ( .A1(n7600), .A2(n7644), .ZN(n6110) );
  INV_X1 U6840 ( .A(n6239), .ZN(n5251) );
  OR2_X1 U6841 ( .A1(n7308), .A2(n7298), .ZN(n5523) );
  AND2_X1 U6842 ( .A1(n7325), .A2(n5523), .ZN(n6094) );
  OR2_X1 U6843 ( .A1(n7210), .A2(n7211), .ZN(n6088) );
  NAND3_X1 U6844 ( .A1(n6106), .A2(n6094), .A3(n6088), .ZN(n6240) );
  NAND2_X1 U6845 ( .A1(n7421), .A2(n6110), .ZN(n7642) );
  XNOR2_X1 U6846 ( .A(n5253), .B(n5252), .ZN(n6395) );
  NAND2_X1 U6847 ( .A1(n6395), .A2(n6191), .ZN(n5258) );
  NAND2_X1 U6848 ( .A1(n5254), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5255) );
  XNOR2_X1 U6849 ( .A(n5255), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9677) );
  AOI22_X1 U6850 ( .A1(n6190), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5256), .B2(
        n9677), .ZN(n5257) );
  NAND2_X1 U6851 ( .A1(n5446), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5265) );
  INV_X1 U6852 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7393) );
  OR2_X1 U6853 ( .A1(n5447), .A2(n7393), .ZN(n5264) );
  NAND2_X1 U6854 ( .A1(n5260), .A2(n5259), .ZN(n5261) );
  NAND2_X1 U6855 ( .A1(n5278), .A2(n5261), .ZN(n7678) );
  OR2_X1 U6856 ( .A1(n5141), .A2(n7678), .ZN(n5263) );
  INV_X1 U6857 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7650) );
  OR2_X1 U6858 ( .A1(n4266), .A2(n7650), .ZN(n5262) );
  NAND2_X1 U6859 ( .A1(n7680), .A2(n7669), .ZN(n6111) );
  NAND2_X1 U6860 ( .A1(n6114), .A2(n6111), .ZN(n7643) );
  OR2_X2 U6861 ( .A1(n7642), .A2(n7643), .ZN(n5266) );
  NAND2_X1 U6862 ( .A1(n5268), .A2(n5267), .ZN(n5270) );
  NAND2_X1 U6863 ( .A1(n5270), .A2(n5269), .ZN(n6460) );
  OR2_X1 U6864 ( .A1(n6460), .A2(n5287), .ZN(n5275) );
  INV_X1 U6865 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6461) );
  NAND2_X1 U6866 ( .A1(n5271), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5272) );
  XNOR2_X1 U6867 ( .A(n5272), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9230) );
  INV_X1 U6868 ( .A(n9230), .ZN(n7399) );
  OAI22_X1 U6869 ( .A1(n5322), .A2(n6461), .B1(n6329), .B2(n7399), .ZN(n5273)
         );
  INV_X1 U6870 ( .A(n5273), .ZN(n5274) );
  NAND2_X1 U6871 ( .A1(n5446), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5283) );
  INV_X1 U6872 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5276) );
  OR2_X1 U6873 ( .A1(n5447), .A2(n5276), .ZN(n5282) );
  AND2_X1 U6874 ( .A1(n5278), .A2(n5277), .ZN(n5279) );
  OR2_X1 U6875 ( .A1(n5279), .A2(n5293), .ZN(n7763) );
  OR2_X1 U6876 ( .A1(n5141), .A2(n7763), .ZN(n5281) );
  INV_X1 U6877 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7624) );
  OR2_X1 U6878 ( .A1(n4266), .A2(n7624), .ZN(n5280) );
  OR2_X1 U6879 ( .A1(n7629), .A2(n7755), .ZN(n6115) );
  NAND2_X1 U6880 ( .A1(n7629), .A2(n7755), .ZN(n6273) );
  OR2_X1 U6881 ( .A1(n5284), .A2(n4858), .ZN(n5285) );
  NAND2_X1 U6882 ( .A1(n5286), .A2(n5285), .ZN(n6477) );
  OR2_X1 U6883 ( .A1(n6477), .A2(n5287), .ZN(n5292) );
  INV_X1 U6884 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6478) );
  OR2_X1 U6885 ( .A1(n5288), .A2(n9621), .ZN(n5289) );
  XNOR2_X1 U6886 ( .A(n5289), .B(n9928), .ZN(n9232) );
  OAI22_X1 U6887 ( .A1(n5322), .A2(n6478), .B1(n6329), .B2(n9232), .ZN(n5290)
         );
  INV_X1 U6888 ( .A(n5290), .ZN(n5291) );
  NAND2_X1 U6889 ( .A1(n6193), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5298) );
  INV_X1 U6890 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9231) );
  OR2_X1 U6891 ( .A1(n4266), .A2(n9231), .ZN(n5297) );
  NOR2_X1 U6892 ( .A1(n5293), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5294) );
  OR2_X1 U6893 ( .A1(n5309), .A2(n5294), .ZN(n7870) );
  OR2_X1 U6894 ( .A1(n5141), .A2(n7870), .ZN(n5296) );
  INV_X1 U6895 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10037) );
  OR2_X1 U6896 ( .A1(n6196), .A2(n10037), .ZN(n5295) );
  NAND2_X1 U6897 ( .A1(n7861), .A2(n7863), .ZN(n6272) );
  XNOR2_X1 U6898 ( .A(n5300), .B(SI_14_), .ZN(n5301) );
  XNOR2_X1 U6899 ( .A(n5299), .B(n5301), .ZN(n6709) );
  NAND2_X1 U6900 ( .A1(n6709), .A2(n6191), .ZN(n5308) );
  INV_X1 U6901 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10034) );
  OR2_X1 U6902 ( .A1(n5303), .A2(n5302), .ZN(n5304) );
  INV_X1 U6903 ( .A(n9714), .ZN(n6711) );
  OAI22_X1 U6904 ( .A1(n5322), .A2(n10034), .B1(n6711), .B2(n6329), .ZN(n5306)
         );
  INV_X1 U6905 ( .A(n5306), .ZN(n5307) );
  NAND2_X1 U6906 ( .A1(n5446), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5314) );
  INV_X1 U6907 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7791) );
  OR2_X1 U6908 ( .A1(n5447), .A2(n7791), .ZN(n5313) );
  OR2_X1 U6909 ( .A1(n5309), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5310) );
  NAND2_X1 U6910 ( .A1(n5327), .A2(n5310), .ZN(n9017) );
  OR2_X1 U6911 ( .A1(n5141), .A2(n9017), .ZN(n5312) );
  INV_X1 U6912 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7878) );
  OR2_X1 U6913 ( .A1(n4266), .A2(n7878), .ZN(n5311) );
  NOR2_X1 U6914 ( .A1(n9019), .A2(n8914), .ZN(n6280) );
  INV_X1 U6915 ( .A(n6280), .ZN(n6120) );
  NAND2_X1 U6916 ( .A1(n9019), .A2(n8914), .ZN(n6278) );
  NAND2_X1 U6917 ( .A1(n7785), .A2(n7784), .ZN(n5315) );
  INV_X1 U6918 ( .A(n5318), .ZN(n5319) );
  XNOR2_X1 U6919 ( .A(n5319), .B(SI_16_), .ZN(n5320) );
  XNOR2_X1 U6920 ( .A(n5317), .B(n5320), .ZN(n6964) );
  NAND2_X1 U6921 ( .A1(n6964), .A2(n6191), .ZN(n5325) );
  INV_X1 U6922 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6967) );
  XNOR2_X1 U6923 ( .A(n5321), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9245) );
  INV_X1 U6924 ( .A(n9245), .ZN(n9228) );
  OAI22_X1 U6925 ( .A1(n5322), .A2(n6967), .B1(n6329), .B2(n9228), .ZN(n5323)
         );
  INV_X1 U6926 ( .A(n5323), .ZN(n5324) );
  NAND2_X1 U6927 ( .A1(n5446), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5333) );
  INV_X1 U6928 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9223) );
  OR2_X1 U6929 ( .A1(n5447), .A2(n9223), .ZN(n5332) );
  OAI21_X1 U6930 ( .B1(n5327), .B2(n5326), .A(n9101), .ZN(n5329) );
  NAND2_X1 U6931 ( .A1(n5329), .A2(n5328), .ZN(n9472) );
  OR2_X1 U6932 ( .A1(n5141), .A2(n9472), .ZN(n5331) );
  INV_X1 U6933 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9473) );
  OR2_X1 U6934 ( .A1(n4266), .A2(n9473), .ZN(n5330) );
  NAND2_X1 U6935 ( .A1(n5476), .A2(n9109), .ZN(n6287) );
  OR2_X1 U6936 ( .A1(n9540), .A2(n9154), .ZN(n9424) );
  NAND2_X1 U6937 ( .A1(n9423), .A2(n5334), .ZN(n9426) );
  NAND3_X1 U6938 ( .A1(n9409), .A2(n9407), .A3(n9426), .ZN(n5335) );
  NAND2_X1 U6939 ( .A1(n5336), .A2(n6077), .ZN(n9378) );
  INV_X1 U6940 ( .A(n5337), .ZN(n5338) );
  XNOR2_X1 U6941 ( .A(n5338), .B(SI_21_), .ZN(n5339) );
  NAND2_X1 U6942 ( .A1(n5617), .A2(n6191), .ZN(n5342) );
  NAND2_X1 U6943 ( .A1(n6190), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5341) );
  AND2_X1 U6944 ( .A1(n5344), .A2(n5343), .ZN(n5346) );
  OR2_X1 U6945 ( .A1(n5346), .A2(n5345), .ZN(n9382) );
  AOI22_X1 U6946 ( .A1(n5446), .A2(P1_REG0_REG_21__SCAN_IN), .B1(n6193), .B2(
        P1_REG1_REG_21__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U6947 ( .A1(n5137), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5347) );
  OAI211_X1 U6948 ( .C1(n9382), .C2(n5141), .A(n5348), .B(n5347), .ZN(n9199)
         );
  XNOR2_X1 U6949 ( .A(n9518), .B(n9199), .ZN(n9377) );
  INV_X1 U6950 ( .A(n9199), .ZN(n6075) );
  NAND2_X1 U6951 ( .A1(n9518), .A2(n6075), .ZN(n6144) );
  NAND2_X1 U6952 ( .A1(n9513), .A2(n9079), .ZN(n6073) );
  NAND2_X1 U6953 ( .A1(n5352), .A2(n5351), .ZN(n5367) );
  INV_X1 U6954 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7901) );
  INV_X1 U6955 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n5353) );
  MUX2_X1 U6956 ( .A(n7901), .B(n5353), .S(n6348), .Z(n5355) );
  INV_X1 U6957 ( .A(SI_24_), .ZN(n5354) );
  NAND2_X1 U6958 ( .A1(n5355), .A2(n5354), .ZN(n5368) );
  INV_X1 U6959 ( .A(n5355), .ZN(n5356) );
  NAND2_X1 U6960 ( .A1(n5356), .A2(SI_24_), .ZN(n5357) );
  NAND2_X1 U6961 ( .A1(n7845), .A2(n6191), .ZN(n5359) );
  NAND2_X1 U6962 ( .A1(n6190), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5358) );
  NAND2_X1 U6963 ( .A1(n6193), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5365) );
  INV_X1 U6964 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9962) );
  OR2_X1 U6965 ( .A1(n6196), .A2(n9962), .ZN(n5364) );
  INV_X1 U6966 ( .A(n5376), .ZN(n5377) );
  OAI21_X1 U6967 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n5361), .A(n5377), .ZN(
        n9341) );
  OR2_X1 U6968 ( .A1(n5141), .A2(n9341), .ZN(n5363) );
  INV_X1 U6969 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9342) );
  OR2_X1 U6970 ( .A1(n4266), .A2(n9342), .ZN(n5362) );
  NAND4_X1 U6971 ( .A1(n5365), .A2(n5364), .A3(n5363), .A4(n5362), .ZN(n9196)
         );
  INV_X1 U6972 ( .A(n9196), .ZN(n8979) );
  NAND2_X1 U6973 ( .A1(n9346), .A2(n8979), .ZN(n6216) );
  NAND2_X1 U6974 ( .A1(n5367), .A2(n5366), .ZN(n5369) );
  NAND2_X1 U6975 ( .A1(n5369), .A2(n5368), .ZN(n5387) );
  INV_X1 U6976 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7900) );
  MUX2_X1 U6977 ( .A(n7900), .B(n7904), .S(n6348), .Z(n5371) );
  INV_X1 U6978 ( .A(SI_25_), .ZN(n5370) );
  NAND2_X1 U6979 ( .A1(n5371), .A2(n5370), .ZN(n5388) );
  INV_X1 U6980 ( .A(n5371), .ZN(n5372) );
  NAND2_X1 U6981 ( .A1(n5372), .A2(SI_25_), .ZN(n5373) );
  NAND2_X1 U6982 ( .A1(n7899), .A2(n6191), .ZN(n5375) );
  NAND2_X1 U6983 ( .A1(n6190), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U6984 ( .A1(n5446), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5383) );
  INV_X1 U6985 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9501) );
  OR2_X1 U6986 ( .A1(n5447), .A2(n9501), .ZN(n5382) );
  INV_X1 U6987 ( .A(n5396), .ZN(n5398) );
  INV_X1 U6988 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n10051) );
  NAND2_X1 U6989 ( .A1(n10051), .A2(n5377), .ZN(n5378) );
  NAND2_X1 U6990 ( .A1(n5398), .A2(n5378), .ZN(n9326) );
  OR2_X1 U6991 ( .A1(n5141), .A2(n9326), .ZN(n5381) );
  INV_X1 U6992 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n5379) );
  OR2_X1 U6993 ( .A1(n4266), .A2(n5379), .ZN(n5380) );
  NAND2_X1 U6994 ( .A1(n9500), .A2(n9170), .ZN(n6153) );
  NAND2_X1 U6995 ( .A1(n6221), .A2(n6153), .ZN(n9319) );
  NAND2_X1 U6996 ( .A1(n5387), .A2(n5386), .ZN(n5389) );
  INV_X1 U6997 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7910) );
  INV_X1 U6998 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n5390) );
  MUX2_X1 U6999 ( .A(n7910), .B(n5390), .S(n6348), .Z(n5392) );
  INV_X1 U7000 ( .A(SI_26_), .ZN(n5391) );
  NAND2_X1 U7001 ( .A1(n5392), .A2(n5391), .ZN(n5406) );
  INV_X1 U7002 ( .A(n5392), .ZN(n5393) );
  NAND2_X1 U7003 ( .A1(n5393), .A2(SI_26_), .ZN(n5394) );
  NAND2_X1 U7004 ( .A1(n6193), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5403) );
  INV_X1 U7005 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n5395) );
  OR2_X1 U7006 ( .A1(n6196), .A2(n5395), .ZN(n5402) );
  INV_X1 U7007 ( .A(n5414), .ZN(n5415) );
  INV_X1 U7008 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U7009 ( .A1(n5398), .A2(n5397), .ZN(n5399) );
  NAND2_X1 U7010 ( .A1(n5415), .A2(n5399), .ZN(n9310) );
  OR2_X1 U7011 ( .A1(n5141), .A2(n9310), .ZN(n5401) );
  INV_X1 U7012 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9311) );
  OR2_X1 U7013 ( .A1(n4266), .A2(n9311), .ZN(n5400) );
  NAND4_X1 U7014 ( .A1(n5403), .A2(n5402), .A3(n5401), .A4(n5400), .ZN(n9194)
         );
  INV_X1 U7015 ( .A(n9194), .ZN(n8986) );
  NAND2_X1 U7016 ( .A1(n9315), .A2(n8986), .ZN(n6156) );
  NAND2_X1 U7017 ( .A1(n6154), .A2(n6156), .ZN(n9307) );
  INV_X1 U7018 ( .A(n9307), .ZN(n9303) );
  INV_X1 U7019 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5599) );
  INV_X1 U7020 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5407) );
  MUX2_X1 U7021 ( .A(n5599), .B(n5407), .S(n6348), .Z(n5409) );
  INV_X1 U7022 ( .A(SI_27_), .ZN(n5408) );
  NAND2_X1 U7023 ( .A1(n5409), .A2(n5408), .ZN(n5437) );
  INV_X1 U7024 ( .A(n5409), .ZN(n5410) );
  NAND2_X1 U7025 ( .A1(n5410), .A2(SI_27_), .ZN(n5411) );
  NAND2_X1 U7026 ( .A1(n8897), .A2(n6191), .ZN(n5413) );
  NAND2_X1 U7027 ( .A1(n6190), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U7028 ( .A1(n6193), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5420) );
  INV_X1 U7029 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n6069) );
  OR2_X1 U7030 ( .A1(n6196), .A2(n6069), .ZN(n5419) );
  INV_X1 U7031 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9929) );
  NAND2_X1 U7032 ( .A1(n5415), .A2(n9929), .ZN(n5416) );
  NAND2_X1 U7033 ( .A1(n5430), .A2(n5416), .ZN(n9295) );
  OR2_X1 U7034 ( .A1(n5141), .A2(n9295), .ZN(n5418) );
  INV_X1 U7035 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9296) );
  OR2_X1 U7036 ( .A1(n4266), .A2(n9296), .ZN(n5417) );
  NOR2_X1 U7037 ( .A1(n9010), .A2(n9168), .ZN(n6209) );
  INV_X1 U7038 ( .A(n6209), .ZN(n6163) );
  NAND2_X1 U7039 ( .A1(n9010), .A2(n9168), .ZN(n6158) );
  NAND2_X1 U7040 ( .A1(n6163), .A2(n6158), .ZN(n6251) );
  INV_X1 U7041 ( .A(n6158), .ZN(n5421) );
  NAND2_X1 U7042 ( .A1(n5442), .A2(n5437), .ZN(n5425) );
  INV_X1 U7043 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5573) );
  INV_X1 U7044 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5424) );
  MUX2_X1 U7045 ( .A(n5573), .B(n5424), .S(n6348), .Z(n5436) );
  XNOR2_X1 U7046 ( .A(n5436), .B(SI_28_), .ZN(n5439) );
  NAND2_X1 U7047 ( .A1(n6190), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5426) );
  NAND2_X1 U7048 ( .A1(n5446), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5434) );
  INV_X1 U7049 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9491) );
  OR2_X1 U7050 ( .A1(n5447), .A2(n9491), .ZN(n5433) );
  INV_X1 U7051 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n5428) );
  OR2_X1 U7052 ( .A1(n4266), .A2(n5428), .ZN(n5432) );
  INV_X1 U7053 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5429) );
  XNOR2_X1 U7054 ( .A(n5430), .B(n5429), .ZN(n9287) );
  OR2_X1 U7055 ( .A1(n5141), .A2(n9287), .ZN(n5431) );
  NAND4_X1 U7056 ( .A1(n5434), .A2(n5433), .A3(n5432), .A4(n5431), .ZN(n9192)
         );
  AND2_X1 U7057 ( .A1(n9568), .A2(n9192), .ZN(n6206) );
  INV_X1 U7058 ( .A(n9192), .ZN(n9057) );
  INV_X1 U7059 ( .A(SI_28_), .ZN(n5435) );
  NAND2_X1 U7060 ( .A1(n5436), .A2(n5435), .ZN(n5438) );
  AND2_X1 U7061 ( .A1(n5437), .A2(n5438), .ZN(n5441) );
  INV_X1 U7062 ( .A(n5438), .ZN(n5440) );
  INV_X1 U7063 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7913) );
  INV_X1 U7064 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n5443) );
  MUX2_X1 U7065 ( .A(n7913), .B(n5443), .S(n6348), .Z(n6170) );
  NAND2_X1 U7066 ( .A1(n5946), .A2(n6191), .ZN(n5445) );
  NAND2_X1 U7067 ( .A1(n6190), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U7068 ( .A1(n5446), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5453) );
  INV_X1 U7069 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5552) );
  OR2_X1 U7070 ( .A1(n5447), .A2(n5552), .ZN(n5452) );
  NAND2_X1 U7071 ( .A1(n5448), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n7916) );
  OR2_X1 U7072 ( .A1(n5141), .A2(n7916), .ZN(n5451) );
  INV_X1 U7073 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n5449) );
  OR2_X1 U7074 ( .A1(n4266), .A2(n5449), .ZN(n5450) );
  INV_X1 U7075 ( .A(n6207), .ZN(n5454) );
  NAND2_X1 U7076 ( .A1(n7918), .A2(n9065), .ZN(n6297) );
  INV_X1 U7077 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U7078 ( .A1(n6623), .A2(n6481), .ZN(n5467) );
  NAND2_X1 U7079 ( .A1(n5460), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U7080 ( .A1(n5463), .A2(n5462), .ZN(n5464) );
  XNOR2_X2 U7081 ( .A(n5466), .B(n5465), .ZN(n7551) );
  INV_X1 U7082 ( .A(n7551), .ZN(n6554) );
  AND2_X1 U7083 ( .A1(n6479), .A2(n6554), .ZN(n6205) );
  INV_X1 U7084 ( .A(n6205), .ZN(n6312) );
  INV_X1 U7085 ( .A(n6366), .ZN(n9631) );
  INV_X1 U7086 ( .A(P1_B_REG_SCAN_IN), .ZN(n5468) );
  OR2_X1 U7087 ( .A1(n6489), .A2(n5468), .ZN(n5469) );
  AND2_X1 U7088 ( .A1(n9129), .A2(n5469), .ZN(n9270) );
  INV_X1 U7089 ( .A(n9270), .ZN(n5472) );
  INV_X1 U7090 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9560) );
  NAND2_X1 U7091 ( .A1(n5137), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5471) );
  NAND2_X1 U7092 ( .A1(n6193), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5470) );
  OAI211_X1 U7093 ( .C1(n6196), .C2(n9560), .A(n5471), .B(n5470), .ZN(n9191)
         );
  INV_X1 U7094 ( .A(n9191), .ZN(n6302) );
  INV_X1 U7095 ( .A(n5473), .ZN(n5474) );
  INV_X1 U7096 ( .A(n7564), .ZN(n9787) );
  NAND2_X1 U7097 ( .A1(n6487), .A2(n7051), .ZN(n7008) );
  INV_X1 U7098 ( .A(n7210), .ZN(n9781) );
  NAND2_X1 U7099 ( .A1(n7191), .A2(n9781), .ZN(n7190) );
  OR2_X1 U7100 ( .A1(n7190), .A2(n7308), .ZN(n7264) );
  NAND3_X1 U7101 ( .A1(n9792), .A2(n9787), .A3(n7430), .ZN(n7649) );
  OR2_X1 U7102 ( .A1(n7680), .A2(n7649), .ZN(n7625) );
  OR2_X2 U7103 ( .A1(n7789), .A2(n9019), .ZN(n7886) );
  NOR2_X2 U7104 ( .A1(n9616), .A2(n7886), .ZN(n9476) );
  NAND2_X1 U7105 ( .A1(n9477), .A2(n9476), .ZN(n9475) );
  NAND2_X1 U7106 ( .A1(n9356), .A2(n5480), .ZN(n9343) );
  NOR2_X2 U7107 ( .A1(n9343), .A2(n9500), .ZN(n9325) );
  AND2_X1 U7108 ( .A1(n7918), .A2(n9285), .ZN(n5481) );
  OR3_X2 U7109 ( .A1(n9275), .A2(n5481), .A3(n9443), .ZN(n7920) );
  INV_X1 U7110 ( .A(n7920), .ZN(n5483) );
  NAND2_X1 U7111 ( .A1(n9268), .A2(n7551), .ZN(n6557) );
  NAND2_X1 U7112 ( .A1(n6625), .A2(n6557), .ZN(n9798) );
  NAND2_X1 U7113 ( .A1(n4321), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5485) );
  MUX2_X1 U7114 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5485), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5486) );
  NAND2_X1 U7115 ( .A1(n5486), .A2(n5491), .ZN(n7906) );
  NAND2_X1 U7116 ( .A1(n7906), .A2(P1_B_REG_SCAN_IN), .ZN(n5490) );
  MUX2_X1 U7117 ( .A(n5490), .B(P1_B_REG_SCAN_IN), .S(n7846), .Z(n5493) );
  NAND2_X1 U7118 ( .A1(n5491), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5492) );
  INV_X1 U7119 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n5494) );
  AND2_X1 U7120 ( .A1(n5510), .A2(n7906), .ZN(n6382) );
  NAND2_X1 U7121 ( .A1(n6625), .A2(n6480), .ZN(n6555) );
  INV_X1 U7122 ( .A(n6555), .ZN(n5495) );
  OR2_X1 U7123 ( .A1(n6619), .A2(n5495), .ZN(n5514) );
  NOR2_X1 U7124 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .ZN(
        n9916) );
  NOR4_X1 U7125 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5498) );
  NOR4_X1 U7126 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5497) );
  NOR4_X1 U7127 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n5496) );
  AND4_X1 U7128 ( .A1(n9916), .A2(n5498), .A3(n5497), .A4(n5496), .ZN(n5504)
         );
  NOR4_X1 U7129 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5502) );
  NOR4_X1 U7130 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n5501) );
  NOR4_X1 U7131 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5500) );
  NOR4_X1 U7132 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n5499) );
  AND4_X1 U7133 ( .A1(n5502), .A2(n5501), .A3(n5500), .A4(n5499), .ZN(n5503)
         );
  NAND2_X1 U7134 ( .A1(n5504), .A2(n5503), .ZN(n5505) );
  NAND2_X1 U7135 ( .A1(n6378), .A2(n5505), .ZN(n6519) );
  NAND2_X1 U7136 ( .A1(n5507), .A2(n5506), .ZN(n5508) );
  NAND2_X1 U7137 ( .A1(n5508), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5509) );
  NAND2_X1 U7138 ( .A1(n6549), .A2(n6557), .ZN(n6522) );
  INV_X1 U7139 ( .A(n6522), .ZN(n5512) );
  NOR2_X1 U7140 ( .A1(n6556), .A2(n5512), .ZN(n5513) );
  NAND2_X1 U7141 ( .A1(n6519), .A2(n5513), .ZN(n6618) );
  INV_X1 U7142 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5515) );
  NOR2_X1 U7143 ( .A1(n7846), .A2(n7908), .ZN(n6380) );
  INV_X1 U7144 ( .A(n6520), .ZN(n6621) );
  MUX2_X1 U7145 ( .A(n5516), .B(n5551), .S(n9795), .Z(n5549) );
  INV_X1 U7146 ( .A(n7863), .ZN(n9206) );
  INV_X1 U7147 ( .A(n7211), .ZN(n9213) );
  INV_X1 U7148 ( .A(n7003), .ZN(n5517) );
  INV_X1 U7149 ( .A(n6487), .ZN(n7007) );
  NAND2_X1 U7150 ( .A1(n9219), .A2(n7007), .ZN(n6998) );
  NAND2_X1 U7151 ( .A1(n5517), .A2(n6998), .ZN(n7001) );
  INV_X1 U7152 ( .A(n6559), .ZN(n5518) );
  NAND2_X1 U7153 ( .A1(n7001), .A2(n5519), .ZN(n6922) );
  NAND2_X1 U7154 ( .A1(n6922), .A2(n6921), .ZN(n6920) );
  NAND2_X1 U7155 ( .A1(n6690), .A2(n7055), .ZN(n5521) );
  NAND2_X1 U7156 ( .A1(n7013), .A2(n5521), .ZN(n6988) );
  INV_X1 U7157 ( .A(n5522), .ZN(n7071) );
  INV_X1 U7158 ( .A(n7092), .ZN(n6994) );
  NAND2_X1 U7159 ( .A1(n6986), .A2(n4861), .ZN(n7080) );
  NAND2_X1 U7160 ( .A1(n7080), .A2(n7079), .ZN(n7078) );
  NAND2_X1 U7161 ( .A1(n7078), .A2(n4857), .ZN(n7189) );
  NAND2_X1 U7162 ( .A1(n6088), .A2(n6236), .ZN(n7194) );
  NAND2_X1 U7163 ( .A1(n7189), .A2(n7194), .ZN(n7188) );
  OAI21_X1 U7164 ( .B1(n9213), .B2(n7210), .A(n7188), .ZN(n7174) );
  NAND2_X1 U7165 ( .A1(n5523), .A2(n7260), .ZN(n7176) );
  NAND2_X1 U7166 ( .A1(n7174), .A2(n7176), .ZN(n7173) );
  INV_X1 U7167 ( .A(n7298), .ZN(n9212) );
  NAND2_X1 U7168 ( .A1(n7173), .A2(n4863), .ZN(n7269) );
  NAND2_X1 U7169 ( .A1(n7325), .A2(n6098), .ZN(n7268) );
  INV_X1 U7170 ( .A(n7485), .ZN(n9211) );
  NAND2_X1 U7171 ( .A1(n5524), .A2(n7485), .ZN(n5525) );
  NAND2_X1 U7172 ( .A1(n7267), .A2(n5525), .ZN(n7331) );
  NAND2_X1 U7173 ( .A1(n6106), .A2(n6107), .ZN(n7330) );
  NAND2_X1 U7174 ( .A1(n7331), .A2(n7330), .ZN(n7329) );
  INV_X1 U7175 ( .A(n7554), .ZN(n9210) );
  NAND2_X1 U7176 ( .A1(n7329), .A2(n5526), .ZN(n7428) );
  NAND2_X1 U7177 ( .A1(n7428), .A2(n7427), .ZN(n7426) );
  INV_X1 U7178 ( .A(n7669), .ZN(n9208) );
  INV_X1 U7179 ( .A(n7755), .ZN(n9207) );
  NAND2_X1 U7180 ( .A1(n7621), .A2(n5529), .ZN(n7729) );
  NAND2_X1 U7181 ( .A1(n6276), .A2(n6272), .ZN(n7728) );
  INV_X1 U7182 ( .A(n8914), .ZN(n9205) );
  NAND2_X1 U7183 ( .A1(n9019), .A2(n9205), .ZN(n5530) );
  INV_X1 U7184 ( .A(n9098), .ZN(n9204) );
  INV_X1 U7185 ( .A(n9109), .ZN(n9203) );
  NAND2_X1 U7186 ( .A1(n9540), .A2(n9202), .ZN(n5533) );
  INV_X1 U7187 ( .A(n9540), .ZN(n9445) );
  INV_X1 U7188 ( .A(n9110), .ZN(n9201) );
  NAND2_X1 U7189 ( .A1(n9422), .A2(n5534), .ZN(n5535) );
  INV_X1 U7190 ( .A(n9152), .ZN(n9200) );
  INV_X1 U7191 ( .A(n9529), .ZN(n9419) );
  INV_X1 U7192 ( .A(n9518), .ZN(n9386) );
  NOR2_X1 U7193 ( .A1(n9386), .A2(n6075), .ZN(n5537) );
  OAI22_X2 U7194 ( .A1(n9376), .A2(n5537), .B1(n9518), .B2(n9199), .ZN(n9362)
         );
  INV_X1 U7195 ( .A(n9137), .ZN(n9197) );
  NAND2_X1 U7196 ( .A1(n5480), .A2(n8979), .ZN(n5540) );
  INV_X1 U7197 ( .A(n9170), .ZN(n9195) );
  NAND2_X1 U7198 ( .A1(n9500), .A2(n9195), .ZN(n5541) );
  INV_X1 U7199 ( .A(n9500), .ZN(n9330) );
  NAND2_X1 U7200 ( .A1(n9569), .A2(n8986), .ZN(n5542) );
  NAND2_X1 U7201 ( .A1(n9315), .A2(n9194), .ZN(n5543) );
  INV_X1 U7202 ( .A(n6251), .ZN(n6059) );
  INV_X1 U7203 ( .A(n9168), .ZN(n9193) );
  OAI21_X1 U7204 ( .B1(n9192), .B2(n9289), .A(n9282), .ZN(n5544) );
  XNOR2_X1 U7205 ( .A(n5544), .B(n6167), .ZN(n7925) );
  INV_X1 U7206 ( .A(n7925), .ZN(n5553) );
  INV_X1 U7207 ( .A(n6632), .ZN(n6482) );
  MUX2_X1 U7208 ( .A(n6482), .B(n4681), .S(n6627), .Z(n5546) );
  INV_X1 U7209 ( .A(n6625), .ZN(n5545) );
  NAND2_X1 U7210 ( .A1(n5546), .A2(n5545), .ZN(n7647) );
  NAND2_X1 U7211 ( .A1(n6480), .A2(n4682), .ZN(n7657) );
  NAND2_X1 U7212 ( .A1(n5553), .A2(n5547), .ZN(n5548) );
  NAND2_X1 U7213 ( .A1(n5549), .A2(n5548), .ZN(P1_U3519) );
  MUX2_X1 U7214 ( .A(n5552), .B(n5551), .S(n9811), .Z(n5555) );
  NAND2_X1 U7215 ( .A1(n5553), .A2(n9551), .ZN(n5554) );
  NAND2_X1 U7216 ( .A1(n5555), .A2(n5554), .ZN(P1_U3551) );
  NOR2_X1 U7217 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5562) );
  NAND4_X1 U7218 ( .A1(n5562), .A2(n5848), .A3(n5561), .A4(n5785), .ZN(n5565)
         );
  NAND4_X1 U7219 ( .A1(n5849), .A2(n5854), .A3(n5881), .A4(n5563), .ZN(n5564)
         );
  NAND2_X1 U7220 ( .A1(n6010), .A2(n5569), .ZN(n5587) );
  NAND2_X1 U7221 ( .A1(n5587), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5570) );
  OR2_X1 U7222 ( .A1(n6010), .A2(n8884), .ZN(n5571) );
  MUX2_X1 U7223 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5571), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5572) );
  NAND2_X1 U7224 ( .A1(n5572), .A2(n5587), .ZN(n5992) );
  NAND2_X1 U7226 ( .A1(n8894), .A2(n8113), .ZN(n5575) );
  OR2_X1 U7227 ( .A1(n5656), .A2(n5573), .ZN(n5574) );
  NOR2_X1 U7228 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5698) );
  INV_X1 U7229 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U7230 ( .A1(n5698), .A2(n5576), .ZN(n5721) );
  INV_X1 U7231 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5578) );
  INV_X1 U7232 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8282) );
  INV_X1 U7233 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5579) );
  INV_X1 U7234 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5580) );
  INV_X1 U7235 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5581) );
  INV_X1 U7236 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10054) );
  INV_X1 U7237 ( .A(n5922), .ZN(n5584) );
  INV_X1 U7238 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5583) );
  INV_X1 U7239 ( .A(n5934), .ZN(n5585) );
  INV_X1 U7240 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9978) );
  NAND2_X1 U7241 ( .A1(n5585), .A2(n9978), .ZN(n5603) );
  NAND2_X1 U7242 ( .A1(n5603), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5586) );
  NAND2_X1 U7243 ( .A1(n8522), .A2(n5586), .ZN(n8550) );
  AND2_X2 U7244 ( .A1(n5592), .A2(n5593), .ZN(n5669) );
  INV_X1 U7245 ( .A(n5669), .ZN(n5697) );
  NAND2_X1 U7246 ( .A1(n8550), .A2(n5669), .ZN(n5598) );
  INV_X1 U7247 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8549) );
  NAND2_X1 U7248 ( .A1(n4268), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U7249 ( .A1(n7108), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5594) );
  OAI211_X1 U7250 ( .C1(n8549), .C2(n7111), .A(n5595), .B(n5594), .ZN(n5596)
         );
  INV_X1 U7251 ( .A(n5596), .ZN(n5597) );
  NAND2_X1 U7252 ( .A1(n8897), .A2(n8113), .ZN(n5601) );
  OR2_X1 U7253 ( .A1(n5656), .A2(n5599), .ZN(n5600) );
  INV_X1 U7254 ( .A(n8812), .ZN(n8562) );
  NAND2_X1 U7255 ( .A1(n5934), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5602) );
  NAND2_X1 U7256 ( .A1(n5603), .A2(n5602), .ZN(n8559) );
  NAND2_X1 U7257 ( .A1(n8559), .A2(n5669), .ZN(n5609) );
  INV_X1 U7258 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U7259 ( .A1(n4268), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U7260 ( .A1(n7108), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5604) );
  OAI211_X1 U7261 ( .C1(n5606), .C2(n7111), .A(n5605), .B(n5604), .ZN(n5607)
         );
  INV_X1 U7262 ( .A(n5607), .ZN(n5608) );
  NAND2_X1 U7263 ( .A1(n7497), .A2(n8113), .ZN(n5611) );
  OR2_X1 U7264 ( .A1(n5656), .A2(n7498), .ZN(n5610) );
  INV_X1 U7265 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8645) );
  INV_X1 U7266 ( .A(n5612), .ZN(n5620) );
  INV_X1 U7267 ( .A(n5613), .ZN(n5905) );
  NAND2_X1 U7268 ( .A1(n5905), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5614) );
  NAND2_X1 U7269 ( .A1(n5620), .A2(n5614), .ZN(n8646) );
  NAND2_X1 U7270 ( .A1(n8646), .A2(n5738), .ZN(n5616) );
  AOI22_X1 U7271 ( .A1(n4268), .A2(P2_REG0_REG_20__SCAN_IN), .B1(n7108), .B2(
        P2_REG1_REG_20__SCAN_IN), .ZN(n5615) );
  OAI211_X1 U7272 ( .C1(n5649), .C2(n8645), .A(n5616), .B(n5615), .ZN(n8656)
         );
  AND2_X1 U7273 ( .A1(n7943), .A2(n8656), .ZN(n5979) );
  INV_X1 U7274 ( .A(n8656), .ZN(n8631) );
  NAND2_X1 U7275 ( .A1(n8842), .A2(n8631), .ZN(n8622) );
  NAND2_X1 U7276 ( .A1(n5617), .A2(n8113), .ZN(n5619) );
  INV_X1 U7277 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7580) );
  OR2_X1 U7278 ( .A1(n5656), .A2(n7580), .ZN(n5618) );
  INV_X1 U7279 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8634) );
  NAND2_X1 U7280 ( .A1(n5620), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5621) );
  NAND2_X1 U7281 ( .A1(n5624), .A2(n5621), .ZN(n8633) );
  NAND2_X1 U7282 ( .A1(n8633), .A2(n5738), .ZN(n5623) );
  AOI22_X1 U7283 ( .A1(n4268), .A2(P2_REG0_REG_21__SCAN_IN), .B1(n7108), .B2(
        P2_REG1_REG_21__SCAN_IN), .ZN(n5622) );
  OAI211_X1 U7284 ( .C1(n5649), .C2(n8634), .A(n5623), .B(n5622), .ZN(n8643)
         );
  INV_X1 U7285 ( .A(n8643), .ZN(n8181) );
  NAND2_X1 U7286 ( .A1(n8769), .A2(n8181), .ZN(n7972) );
  INV_X1 U7287 ( .A(n8625), .ZN(n8627) );
  OR2_X1 U7288 ( .A1(n8639), .A2(n8627), .ZN(n8607) );
  NAND2_X1 U7289 ( .A1(n7746), .A2(n8113), .ZN(n8321) );
  OR2_X1 U7290 ( .A1(n5656), .A2(n9968), .ZN(n8320) );
  NAND2_X1 U7291 ( .A1(n5624), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U7292 ( .A1(n5631), .A2(n5625), .ZN(n8617) );
  INV_X1 U7293 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8616) );
  NAND2_X1 U7294 ( .A1(n4268), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U7295 ( .A1(n7108), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5626) );
  OAI211_X1 U7296 ( .C1(n8616), .C2(n5649), .A(n5627), .B(n5626), .ZN(n5628)
         );
  AOI21_X1 U7297 ( .B1(n8617), .B2(n5738), .A(n5628), .ZN(n8632) );
  NOR2_X1 U7298 ( .A1(n5912), .A2(n8632), .ZN(n8076) );
  INV_X1 U7299 ( .A(n8076), .ZN(n5980) );
  NAND2_X1 U7300 ( .A1(n5912), .A2(n8632), .ZN(n8074) );
  INV_X1 U7301 ( .A(n8156), .ZN(n8611) );
  NAND2_X1 U7302 ( .A1(n7750), .A2(n8113), .ZN(n5630) );
  OR2_X1 U7303 ( .A1(n5656), .A2(n7753), .ZN(n5629) );
  NAND2_X1 U7304 ( .A1(n5631), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U7305 ( .A1(n5641), .A2(n5632), .ZN(n8601) );
  NAND2_X1 U7306 ( .A1(n8601), .A2(n5738), .ZN(n5637) );
  INV_X1 U7307 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8600) );
  NAND2_X1 U7308 ( .A1(n7108), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U7309 ( .A1(n4268), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5633) );
  OAI211_X1 U7310 ( .C1(n8600), .C2(n7111), .A(n5634), .B(n5633), .ZN(n5635)
         );
  INV_X1 U7311 ( .A(n5635), .ZN(n5636) );
  NAND2_X1 U7312 ( .A1(n5984), .A2(n8614), .ZN(n5914) );
  INV_X1 U7313 ( .A(n5914), .ZN(n5638) );
  NAND2_X1 U7314 ( .A1(n7845), .A2(n8113), .ZN(n5640) );
  OR2_X1 U7315 ( .A1(n5656), .A2(n7901), .ZN(n5639) );
  NAND2_X1 U7316 ( .A1(n5641), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U7317 ( .A1(n5922), .A2(n5642), .ZN(n8582) );
  NAND2_X1 U7318 ( .A1(n8582), .A2(n5738), .ZN(n5647) );
  INV_X1 U7319 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8589) );
  NAND2_X1 U7320 ( .A1(n4268), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U7321 ( .A1(n7108), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5643) );
  OAI211_X1 U7322 ( .C1(n8589), .C2(n7111), .A(n5644), .B(n5643), .ZN(n5645)
         );
  INV_X1 U7323 ( .A(n5645), .ZN(n5646) );
  NAND2_X1 U7324 ( .A1(n8822), .A2(n8598), .ZN(n5919) );
  INV_X1 U7325 ( .A(n5919), .ZN(n5648) );
  NAND2_X1 U7326 ( .A1(n5668), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U7327 ( .A1(n5669), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5652) );
  NAND2_X1 U7328 ( .A1(n4269), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5651) );
  NAND2_X1 U7329 ( .A1(n5671), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5650) );
  NAND2_X1 U7330 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5654) );
  OR2_X1 U7331 ( .A1(n5656), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5657) );
  INV_X1 U7332 ( .A(n7980), .ZN(n5965) );
  NAND2_X1 U7333 ( .A1(n4269), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5662) );
  NAND2_X1 U7334 ( .A1(n5668), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U7335 ( .A1(n5669), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5659) );
  NAND4_X1 U7336 ( .A1(n5662), .A2(n5661), .A3(n5660), .A4(n5659), .ZN(n5964)
         );
  NAND2_X1 U7337 ( .A1(n6345), .A2(SI_0_), .ZN(n5664) );
  INV_X1 U7338 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5663) );
  XNOR2_X1 U7339 ( .A(n5664), .B(n5663), .ZN(n8902) );
  MUX2_X1 U7340 ( .A(n4807), .B(n8902), .S(n6324), .Z(n6886) );
  INV_X1 U7341 ( .A(n6886), .ZN(n9818) );
  NAND2_X1 U7342 ( .A1(n5964), .A2(n9818), .ZN(n6936) );
  NAND2_X1 U7343 ( .A1(n6932), .A2(n6936), .ZN(n5667) );
  INV_X1 U7344 ( .A(n8383), .ZN(n7242) );
  NAND2_X1 U7345 ( .A1(n7242), .A2(n6941), .ZN(n5666) );
  NAND2_X1 U7346 ( .A1(n5667), .A2(n5666), .ZN(n7240) );
  NAND2_X1 U7347 ( .A1(n5668), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5675) );
  NAND2_X1 U7348 ( .A1(n5669), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U7349 ( .A1(n5670), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U7350 ( .A1(n5671), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5672) );
  OR2_X1 U7351 ( .A1(n5656), .A2(n4886), .ZN(n5682) );
  OR2_X1 U7352 ( .A1(n5676), .A2(n6362), .ZN(n5681) );
  NOR2_X1 U7353 ( .A1(n5677), .A2(n8884), .ZN(n5678) );
  NAND2_X1 U7354 ( .A1(n5897), .A2(n6603), .ZN(n5680) );
  OR2_X1 U7355 ( .A1(n8381), .A2(n6860), .ZN(n7988) );
  NAND2_X1 U7356 ( .A1(n8381), .A2(n6860), .ZN(n7987) );
  NAND2_X1 U7357 ( .A1(n7240), .A2(n8133), .ZN(n5684) );
  NAND2_X1 U7358 ( .A1(n6958), .A2(n6860), .ZN(n5683) );
  NAND2_X1 U7359 ( .A1(n5684), .A2(n5683), .ZN(n6971) );
  NAND2_X1 U7360 ( .A1(n4268), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5688) );
  INV_X1 U7361 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6659) );
  NAND2_X1 U7362 ( .A1(n5669), .A2(n6659), .ZN(n5687) );
  NAND2_X1 U7363 ( .A1(n7108), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5685) );
  INV_X1 U7364 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6346) );
  OR2_X1 U7365 ( .A1(n5656), .A2(n6346), .ZN(n5695) );
  OR2_X1 U7366 ( .A1(n5676), .A2(n6350), .ZN(n5694) );
  NAND2_X1 U7367 ( .A1(n5679), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5689) );
  MUX2_X1 U7368 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5689), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5692) );
  AND2_X1 U7369 ( .A1(n5692), .A2(n5691), .ZN(n6668) );
  NAND2_X1 U7370 ( .A1(n5897), .A2(n6668), .ZN(n5693) );
  NAND2_X1 U7371 ( .A1(n8380), .A2(n7228), .ZN(n8003) );
  NAND2_X1 U7372 ( .A1(n7241), .A2(n7228), .ZN(n5696) );
  NAND2_X1 U7373 ( .A1(n7108), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U7374 ( .A1(n5670), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5702) );
  INV_X1 U7375 ( .A(n5698), .ZN(n5710) );
  NAND2_X1 U7376 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5699) );
  NAND2_X1 U7377 ( .A1(n5710), .A2(n5699), .ZN(n7168) );
  NAND2_X1 U7378 ( .A1(n5738), .A2(n7168), .ZN(n5701) );
  NAND2_X1 U7379 ( .A1(n4268), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5700) );
  INV_X1 U7380 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6347) );
  OR2_X1 U7381 ( .A1(n5656), .A2(n6347), .ZN(n5707) );
  OR2_X1 U7382 ( .A1(n5676), .A2(n6354), .ZN(n5706) );
  NAND2_X1 U7383 ( .A1(n5691), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5704) );
  XNOR2_X1 U7384 ( .A(n5704), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6751) );
  NAND2_X1 U7385 ( .A1(n5897), .A2(n6751), .ZN(n5705) );
  INV_X1 U7386 ( .A(n9827), .ZN(n7169) );
  NOR2_X1 U7387 ( .A1(n8379), .A2(n7169), .ZN(n5708) );
  NAND2_X1 U7388 ( .A1(n8379), .A2(n7169), .ZN(n5709) );
  NAND2_X1 U7389 ( .A1(n4268), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5715) );
  NAND2_X1 U7390 ( .A1(n7108), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5714) );
  INV_X2 U7391 ( .A(n5697), .ZN(n5738) );
  NAND2_X1 U7392 ( .A1(n5710), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U7393 ( .A1(n5721), .A2(n5711), .ZN(n7292) );
  NAND2_X1 U7394 ( .A1(n5738), .A2(n7292), .ZN(n5713) );
  NAND2_X1 U7395 ( .A1(n5670), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5712) );
  NAND4_X1 U7396 ( .A1(n5715), .A2(n5714), .A3(n5713), .A4(n5712), .ZN(n8378)
         );
  OR2_X1 U7397 ( .A1(n5676), .A2(n6364), .ZN(n5719) );
  OR2_X1 U7398 ( .A1(n5656), .A2(n4903), .ZN(n5718) );
  NAND2_X1 U7399 ( .A1(n5727), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5716) );
  NAND2_X1 U7400 ( .A1(n5897), .A2(n6802), .ZN(n5717) );
  INV_X1 U7401 ( .A(n9832), .ZN(n7291) );
  OR2_X1 U7402 ( .A1(n8378), .A2(n7291), .ZN(n7252) );
  NAND2_X1 U7403 ( .A1(n7253), .A2(n7252), .ZN(n5720) );
  NAND2_X1 U7404 ( .A1(n8378), .A2(n7291), .ZN(n7251) );
  NAND2_X1 U7405 ( .A1(n5720), .A2(n7251), .ZN(n7377) );
  NAND2_X1 U7406 ( .A1(n4268), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5726) );
  NAND2_X1 U7407 ( .A1(n7108), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U7408 ( .A1(n5721), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5722) );
  NAND2_X1 U7409 ( .A1(n5736), .A2(n5722), .ZN(n7375) );
  NAND2_X1 U7410 ( .A1(n5738), .A2(n7375), .ZN(n5724) );
  NAND2_X1 U7411 ( .A1(n5670), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5723) );
  NAND4_X1 U7412 ( .A1(n5726), .A2(n5725), .A3(n5724), .A4(n5723), .ZN(n8377)
         );
  INV_X1 U7413 ( .A(n8377), .ZN(n8219) );
  OR2_X1 U7414 ( .A1(n6356), .A2(n5676), .ZN(n5731) );
  OR2_X1 U7415 ( .A1(n5744), .A2(n8884), .ZN(n5728) );
  XNOR2_X1 U7416 ( .A(n5728), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6808) );
  NAND2_X1 U7417 ( .A1(n5897), .A2(n6808), .ZN(n5730) );
  INV_X1 U7418 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6352) );
  OR2_X1 U7419 ( .A1(n5656), .A2(n6352), .ZN(n5729) );
  NAND2_X1 U7420 ( .A1(n8219), .A2(n7360), .ZN(n5732) );
  NAND2_X1 U7421 ( .A1(n7377), .A2(n5732), .ZN(n5734) );
  INV_X1 U7422 ( .A(n7360), .ZN(n9840) );
  NAND2_X1 U7423 ( .A1(n8377), .A2(n9840), .ZN(n5733) );
  NAND2_X1 U7424 ( .A1(n4268), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5742) );
  NAND2_X1 U7425 ( .A1(n7108), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5741) );
  INV_X1 U7426 ( .A(n5735), .ZN(n5753) );
  NAND2_X1 U7427 ( .A1(n5736), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5737) );
  NAND2_X1 U7428 ( .A1(n5753), .A2(n5737), .ZN(n8222) );
  NAND2_X1 U7429 ( .A1(n5738), .A2(n8222), .ZN(n5740) );
  NAND2_X1 U7430 ( .A1(n5670), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5739) );
  NAND4_X1 U7431 ( .A1(n5742), .A2(n5741), .A3(n5740), .A4(n5739), .ZN(n8376)
         );
  OR2_X1 U7432 ( .A1(n6358), .A2(n5676), .ZN(n5747) );
  INV_X1 U7433 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5743) );
  NAND2_X1 U7434 ( .A1(n5744), .A2(n5743), .ZN(n5748) );
  NAND2_X1 U7435 ( .A1(n5748), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5745) );
  XNOR2_X1 U7436 ( .A(n5745), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6813) );
  AOI22_X1 U7437 ( .A1(n5898), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5897), .B2(
        n6813), .ZN(n5746) );
  OR2_X1 U7438 ( .A1(n8376), .A2(n9843), .ZN(n8020) );
  NAND2_X1 U7439 ( .A1(n9843), .A2(n8376), .ZN(n7407) );
  NAND2_X1 U7440 ( .A1(n8020), .A2(n7407), .ZN(n8138) );
  NAND2_X1 U7441 ( .A1(n4878), .A2(n8138), .ZN(n7467) );
  NAND2_X1 U7442 ( .A1(n6372), .A2(n8113), .ZN(n5751) );
  NAND2_X1 U7443 ( .A1(n5761), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5749) );
  XNOR2_X1 U7444 ( .A(n5749), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6902) );
  AOI22_X1 U7445 ( .A1(n5898), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5897), .B2(
        n6902), .ZN(n5750) );
  NAND2_X1 U7446 ( .A1(n5751), .A2(n5750), .ZN(n9850) );
  NAND2_X1 U7447 ( .A1(n4268), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5758) );
  NAND2_X1 U7448 ( .A1(n7108), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5757) );
  INV_X1 U7449 ( .A(n5752), .ZN(n5764) );
  NAND2_X1 U7450 ( .A1(n5753), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5754) );
  NAND2_X1 U7451 ( .A1(n5764), .A2(n5754), .ZN(n7572) );
  NAND2_X1 U7452 ( .A1(n5738), .A2(n7572), .ZN(n5756) );
  NAND2_X1 U7453 ( .A1(n5670), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5755) );
  OR2_X1 U7454 ( .A1(n9850), .A2(n8313), .ZN(n8016) );
  NAND2_X1 U7455 ( .A1(n9850), .A2(n8313), .ZN(n8021) );
  INV_X1 U7456 ( .A(n8376), .ZN(n7569) );
  AND2_X1 U7457 ( .A1(n7569), .A2(n9843), .ZN(n7409) );
  NOR2_X1 U7458 ( .A1(n8141), .A2(n7409), .ZN(n5759) );
  NAND2_X1 U7459 ( .A1(n9850), .A2(n8375), .ZN(n5760) );
  NAND2_X1 U7460 ( .A1(n6384), .A2(n8113), .ZN(n5763) );
  OAI21_X1 U7461 ( .B1(n5761), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5772) );
  INV_X1 U7462 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5771) );
  XNOR2_X1 U7463 ( .A(n5772), .B(n5771), .ZN(n7154) );
  AOI22_X1 U7464 ( .A1(n5898), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5897), .B2(
        n7044), .ZN(n5762) );
  NAND2_X1 U7465 ( .A1(n7108), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U7466 ( .A1(n4268), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5768) );
  NAND2_X1 U7467 ( .A1(n5764), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U7468 ( .A1(n5777), .A2(n5765), .ZN(n8315) );
  NAND2_X1 U7469 ( .A1(n5738), .A2(n8315), .ZN(n5767) );
  NAND2_X1 U7470 ( .A1(n5670), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5766) );
  AND2_X1 U7471 ( .A1(n9856), .A2(n8374), .ZN(n5770) );
  OR2_X1 U7472 ( .A1(n6387), .A2(n5676), .ZN(n5776) );
  NAND2_X1 U7473 ( .A1(n5772), .A2(n5771), .ZN(n5773) );
  NAND2_X1 U7474 ( .A1(n5773), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5774) );
  XNOR2_X1 U7475 ( .A(n5774), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7152) );
  AOI22_X1 U7476 ( .A1(n5898), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5897), .B2(
        n7152), .ZN(n5775) );
  NAND2_X1 U7477 ( .A1(n7108), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5782) );
  NAND2_X1 U7478 ( .A1(n4268), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5781) );
  NAND2_X1 U7479 ( .A1(n5777), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5778) );
  NAND2_X1 U7480 ( .A1(n5789), .A2(n5778), .ZN(n7777) );
  NAND2_X1 U7481 ( .A1(n5738), .A2(n7777), .ZN(n5780) );
  NAND2_X1 U7482 ( .A1(n5670), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5779) );
  NAND2_X1 U7483 ( .A1(n9860), .A2(n8373), .ZN(n7797) );
  NAND2_X1 U7484 ( .A1(n6395), .A2(n8113), .ZN(n5788) );
  NOR2_X1 U7485 ( .A1(n5783), .A2(n8884), .ZN(n5784) );
  MUX2_X1 U7486 ( .A(n8884), .B(n5784), .S(P2_IR_REG_11__SCAN_IN), .Z(n5786)
         );
  AND2_X1 U7487 ( .A1(n5783), .A2(n5785), .ZN(n5809) );
  OR2_X1 U7488 ( .A1(n5786), .A2(n5809), .ZN(n7445) );
  AOI22_X1 U7489 ( .A1(n5898), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5897), .B2(
        n7438), .ZN(n5787) );
  NAND2_X1 U7490 ( .A1(n5788), .A2(n5787), .ZN(n9865) );
  NAND2_X1 U7491 ( .A1(n4268), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U7492 ( .A1(n7108), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5793) );
  NAND2_X1 U7493 ( .A1(n5789), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U7494 ( .A1(n5801), .A2(n5790), .ZN(n7854) );
  NAND2_X1 U7495 ( .A1(n5738), .A2(n7854), .ZN(n5792) );
  NAND2_X1 U7496 ( .A1(n5670), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5791) );
  OR2_X1 U7497 ( .A1(n9865), .A2(n7795), .ZN(n8035) );
  NAND2_X1 U7498 ( .A1(n9865), .A2(n7795), .ZN(n8037) );
  NAND2_X1 U7499 ( .A1(n7706), .A2(n8145), .ZN(n5796) );
  INV_X1 U7500 ( .A(n7795), .ZN(n8372) );
  NAND2_X1 U7501 ( .A1(n9865), .A2(n8372), .ZN(n5795) );
  OR2_X1 U7502 ( .A1(n6460), .A2(n5676), .ZN(n5799) );
  OR2_X1 U7503 ( .A1(n5809), .A2(n8884), .ZN(n5797) );
  XNOR2_X1 U7504 ( .A(n5797), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7687) );
  AOI22_X1 U7505 ( .A1(n5898), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5897), .B2(
        n7687), .ZN(n5798) );
  NAND2_X1 U7506 ( .A1(n7108), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5806) );
  INV_X1 U7507 ( .A(n5800), .ZN(n5813) );
  NAND2_X1 U7508 ( .A1(n5801), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5802) );
  NAND2_X1 U7509 ( .A1(n5813), .A2(n5802), .ZN(n7806) );
  NAND2_X1 U7510 ( .A1(n5738), .A2(n7806), .ZN(n5805) );
  NAND2_X1 U7511 ( .A1(n5670), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U7512 ( .A1(n4268), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5803) );
  INV_X1 U7513 ( .A(n9664), .ZN(n8371) );
  OR2_X1 U7514 ( .A1(n9871), .A2(n8371), .ZN(n5807) );
  OR2_X1 U7515 ( .A1(n6477), .A2(n5676), .ZN(n5811) );
  NAND2_X1 U7516 ( .A1(n5809), .A2(n5808), .ZN(n5851) );
  NAND2_X1 U7517 ( .A1(n5851), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5823) );
  XNOR2_X1 U7518 ( .A(n5823), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7816) );
  AOI22_X1 U7519 ( .A1(n5898), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5897), .B2(
        n7816), .ZN(n5810) );
  INV_X1 U7520 ( .A(n9654), .ZN(n5812) );
  NAND2_X1 U7521 ( .A1(n9660), .A2(n5812), .ZN(n5819) );
  NAND2_X1 U7522 ( .A1(n4268), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5818) );
  NAND2_X1 U7523 ( .A1(n7108), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5817) );
  NAND2_X1 U7524 ( .A1(n5813), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U7525 ( .A1(n5829), .A2(n5814), .ZN(n9655) );
  NAND2_X1 U7526 ( .A1(n5738), .A2(n9655), .ZN(n5816) );
  NAND2_X1 U7527 ( .A1(n5670), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5815) );
  NAND4_X1 U7528 ( .A1(n5818), .A2(n5817), .A3(n5816), .A4(n5815), .ZN(n8724)
         );
  NAND2_X1 U7529 ( .A1(n5819), .A2(n8724), .ZN(n5822) );
  INV_X1 U7530 ( .A(n9660), .ZN(n5820) );
  NAND2_X1 U7531 ( .A1(n5820), .A2(n9654), .ZN(n5821) );
  NAND2_X1 U7532 ( .A1(n5822), .A2(n5821), .ZN(n8721) );
  NAND2_X1 U7533 ( .A1(n6709), .A2(n8113), .ZN(n5828) );
  NAND2_X1 U7534 ( .A1(n5823), .A2(n5848), .ZN(n5824) );
  NAND2_X1 U7535 ( .A1(n5824), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5825) );
  NAND2_X1 U7536 ( .A1(n5825), .A2(n5849), .ZN(n5836) );
  OR2_X1 U7537 ( .A1(n5825), .A2(n5849), .ZN(n5826) );
  AOI22_X1 U7538 ( .A1(n5898), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5897), .B2(
        n8388), .ZN(n5827) );
  NAND2_X1 U7539 ( .A1(n4268), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5834) );
  NAND2_X1 U7540 ( .A1(n7108), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U7541 ( .A1(n5829), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5830) );
  NAND2_X1 U7542 ( .A1(n5841), .A2(n5830), .ZN(n8730) );
  NAND2_X1 U7543 ( .A1(n5738), .A2(n8730), .ZN(n5832) );
  NAND2_X1 U7544 ( .A1(n5670), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5831) );
  OR2_X1 U7545 ( .A1(n8793), .A2(n8705), .ZN(n5835) );
  NAND2_X1 U7546 ( .A1(n8721), .A2(n5835), .ZN(n8716) );
  NAND2_X1 U7547 ( .A1(n8793), .A2(n8705), .ZN(n8717) );
  NAND2_X1 U7548 ( .A1(n6845), .A2(n8113), .ZN(n5839) );
  NAND2_X1 U7549 ( .A1(n5836), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5837) );
  XNOR2_X1 U7550 ( .A(n5837), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8409) );
  AOI22_X1 U7551 ( .A1(n5898), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5897), .B2(
        n8409), .ZN(n5838) );
  NAND2_X1 U7552 ( .A1(n4268), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5846) );
  NAND2_X1 U7553 ( .A1(n7108), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5845) );
  INV_X1 U7554 ( .A(n5840), .ZN(n5860) );
  NAND2_X1 U7555 ( .A1(n5841), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5842) );
  NAND2_X1 U7556 ( .A1(n5860), .A2(n5842), .ZN(n8709) );
  NAND2_X1 U7557 ( .A1(n5738), .A2(n8709), .ZN(n5844) );
  NAND2_X1 U7558 ( .A1(n5670), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5843) );
  NAND4_X1 U7559 ( .A1(n5846), .A2(n5845), .A3(n5844), .A4(n5843), .ZN(n8725)
         );
  AND2_X1 U7560 ( .A1(n8871), .A2(n8725), .ZN(n5847) );
  NAND2_X1 U7561 ( .A1(n6964), .A2(n8113), .ZN(n5858) );
  NAND2_X1 U7562 ( .A1(n4855), .A2(n5561), .ZN(n5850) );
  NOR2_X2 U7563 ( .A1(n5851), .A2(n5850), .ZN(n5855) );
  INV_X1 U7564 ( .A(n5855), .ZN(n5852) );
  NAND2_X1 U7565 ( .A1(n5852), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5853) );
  MUX2_X1 U7566 ( .A(n5853), .B(P2_IR_REG_31__SCAN_IN), .S(n5854), .Z(n5856)
         );
  NAND2_X1 U7567 ( .A1(n5855), .A2(n5854), .ZN(n5877) );
  NAND2_X1 U7568 ( .A1(n5856), .A2(n5877), .ZN(n8443) );
  INV_X1 U7569 ( .A(n8443), .ZN(n8429) );
  AOI22_X1 U7570 ( .A1(n5898), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5897), .B2(
        n8429), .ZN(n5857) );
  NAND2_X1 U7571 ( .A1(n7108), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5865) );
  NAND2_X1 U7572 ( .A1(n5670), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5864) );
  INV_X1 U7573 ( .A(n5859), .ZN(n5869) );
  NAND2_X1 U7574 ( .A1(n5860), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5861) );
  NAND2_X1 U7575 ( .A1(n5869), .A2(n5861), .ZN(n8698) );
  NAND2_X1 U7576 ( .A1(n5738), .A2(n8698), .ZN(n5863) );
  NAND2_X1 U7577 ( .A1(n4268), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U7578 ( .A1(n8699), .A2(n8682), .ZN(n8063) );
  NAND2_X1 U7579 ( .A1(n8060), .A2(n8063), .ZN(n8149) );
  NAND2_X1 U7580 ( .A1(n8699), .A2(n8706), .ZN(n8678) );
  NAND2_X1 U7581 ( .A1(n7202), .A2(n8113), .ZN(n5868) );
  NAND2_X1 U7582 ( .A1(n5877), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5866) );
  XNOR2_X1 U7583 ( .A(n5866), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8470) );
  AOI22_X1 U7584 ( .A1(n5898), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5897), .B2(
        n8470), .ZN(n5867) );
  NAND2_X1 U7585 ( .A1(n7108), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U7586 ( .A1(n5670), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5873) );
  NAND2_X1 U7587 ( .A1(n5869), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5870) );
  NAND2_X1 U7588 ( .A1(n5886), .A2(n5870), .ZN(n8686) );
  NAND2_X1 U7589 ( .A1(n5738), .A2(n8686), .ZN(n5872) );
  NAND2_X1 U7590 ( .A1(n4268), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5871) );
  NAND2_X1 U7591 ( .A1(n8858), .A2(n8668), .ZN(n8059) );
  INV_X1 U7592 ( .A(n8679), .ZN(n5875) );
  INV_X1 U7593 ( .A(n8668), .ZN(n8694) );
  NAND2_X1 U7594 ( .A1(n8858), .A2(n8694), .ZN(n5876) );
  NAND2_X1 U7595 ( .A1(n8681), .A2(n5876), .ZN(n8665) );
  NAND2_X1 U7596 ( .A1(n7296), .A2(n8113), .ZN(n5885) );
  INV_X1 U7597 ( .A(n5877), .ZN(n5879) );
  NAND2_X1 U7598 ( .A1(n5879), .A2(n5878), .ZN(n5880) );
  OR2_X1 U7599 ( .A1(n5882), .A2(n5881), .ZN(n5883) );
  AND2_X1 U7600 ( .A1(n5895), .A2(n5883), .ZN(n8485) );
  AOI22_X1 U7601 ( .A1(n5898), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5897), .B2(
        n8485), .ZN(n5884) );
  NAND2_X1 U7602 ( .A1(n4268), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5891) );
  NAND2_X1 U7603 ( .A1(n7108), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U7604 ( .A1(n5886), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5887) );
  NAND2_X1 U7605 ( .A1(n5903), .A2(n5887), .ZN(n8669) );
  NAND2_X1 U7606 ( .A1(n5669), .A2(n8669), .ZN(n5889) );
  NAND2_X1 U7607 ( .A1(n5670), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5888) );
  OR2_X1 U7608 ( .A1(n8779), .A2(n8655), .ZN(n5892) );
  NAND2_X1 U7609 ( .A1(n8665), .A2(n5892), .ZN(n5894) );
  NAND2_X1 U7610 ( .A1(n8779), .A2(n8655), .ZN(n5893) );
  NAND2_X1 U7611 ( .A1(n5894), .A2(n5893), .ZN(n8654) );
  NAND2_X1 U7612 ( .A1(n7403), .A2(n8113), .ZN(n5900) );
  AOI22_X1 U7613 ( .A1(n5898), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8495), .B2(
        n5897), .ZN(n5899) );
  NAND2_X1 U7614 ( .A1(n4268), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5902) );
  NAND2_X1 U7615 ( .A1(n7108), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5901) );
  AND2_X1 U7616 ( .A1(n5902), .A2(n5901), .ZN(n5908) );
  NAND2_X1 U7617 ( .A1(n5903), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5904) );
  NAND2_X1 U7618 ( .A1(n5905), .A2(n5904), .ZN(n8659) );
  NAND2_X1 U7619 ( .A1(n8659), .A2(n5738), .ZN(n5907) );
  NAND2_X1 U7620 ( .A1(n4269), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U7621 ( .A1(n8848), .A2(n8667), .ZN(n8066) );
  INV_X1 U7622 ( .A(n8653), .ZN(n5909) );
  NAND2_X1 U7623 ( .A1(n8654), .A2(n5909), .ZN(n5911) );
  NAND2_X1 U7624 ( .A1(n8848), .A2(n8642), .ZN(n5910) );
  NAND2_X1 U7625 ( .A1(n8179), .A2(n8181), .ZN(n8610) );
  NAND2_X1 U7626 ( .A1(n7943), .A2(n8631), .ZN(n8626) );
  OR2_X1 U7627 ( .A1(n8627), .A2(n8626), .ZN(n8608) );
  INV_X1 U7628 ( .A(n8632), .ZN(n8597) );
  OR2_X1 U7629 ( .A1(n8597), .A2(n5912), .ZN(n5913) );
  NAND2_X1 U7630 ( .A1(n8593), .A2(n5914), .ZN(n5916) );
  OR2_X1 U7631 ( .A1(n5984), .A2(n8614), .ZN(n5915) );
  NAND2_X1 U7632 ( .A1(n5916), .A2(n5915), .ZN(n8577) );
  INV_X1 U7633 ( .A(n8577), .ZN(n5917) );
  NAND2_X1 U7634 ( .A1(n4876), .A2(n5917), .ZN(n5918) );
  NAND2_X1 U7635 ( .A1(n7899), .A2(n8113), .ZN(n5921) );
  OR2_X1 U7636 ( .A1(n5656), .A2(n7900), .ZN(n5920) );
  NAND2_X1 U7637 ( .A1(n5922), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U7638 ( .A1(n5932), .A2(n5923), .ZN(n8568) );
  NAND2_X1 U7639 ( .A1(n8568), .A2(n5738), .ZN(n5928) );
  INV_X1 U7640 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8572) );
  NAND2_X1 U7641 ( .A1(n7108), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5925) );
  NAND2_X1 U7642 ( .A1(n4268), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5924) );
  OAI211_X1 U7643 ( .C1(n7111), .C2(n8572), .A(n5925), .B(n5924), .ZN(n5926)
         );
  INV_X1 U7644 ( .A(n5926), .ZN(n5927) );
  NAND2_X1 U7645 ( .A1(n8816), .A2(n8580), .ZN(n8084) );
  INV_X1 U7646 ( .A(n8084), .ZN(n5929) );
  OR2_X1 U7647 ( .A1(n8816), .A2(n8580), .ZN(n8085) );
  NAND2_X1 U7648 ( .A1(n7907), .A2(n8113), .ZN(n5931) );
  OR2_X1 U7649 ( .A1(n5656), .A2(n7910), .ZN(n5930) );
  NAND2_X1 U7650 ( .A1(n5932), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5933) );
  NAND2_X1 U7651 ( .A1(n5934), .A2(n5933), .ZN(n8347) );
  NAND2_X1 U7652 ( .A1(n8347), .A2(n5738), .ZN(n5939) );
  INV_X1 U7653 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n7968) );
  NAND2_X1 U7654 ( .A1(n4268), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5936) );
  NAND2_X1 U7655 ( .A1(n7108), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5935) );
  OAI211_X1 U7656 ( .C1(n7968), .C2(n7111), .A(n5936), .B(n5935), .ZN(n5937)
         );
  INV_X1 U7657 ( .A(n5937), .ZN(n5938) );
  NOR2_X1 U7658 ( .A1(n8353), .A2(n8566), .ZN(n5941) );
  NAND2_X1 U7659 ( .A1(n8353), .A2(n8566), .ZN(n5940) );
  OAI21_X1 U7660 ( .B1(n8806), .B2(n5943), .A(n8543), .ZN(n5945) );
  NAND2_X1 U7661 ( .A1(n5945), .A2(n5944), .ZN(n5954) );
  NAND2_X1 U7662 ( .A1(n5946), .A2(n8113), .ZN(n5948) );
  OR2_X1 U7663 ( .A1(n5656), .A2(n7913), .ZN(n5947) );
  INV_X1 U7664 ( .A(n8522), .ZN(n5949) );
  NAND2_X1 U7665 ( .A1(n5949), .A2(n5669), .ZN(n7114) );
  INV_X1 U7666 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n10052) );
  NAND2_X1 U7667 ( .A1(n7108), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5951) );
  NAND2_X1 U7668 ( .A1(n4268), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5950) );
  OAI211_X1 U7669 ( .C1(n7111), .C2(n10052), .A(n5951), .B(n5950), .ZN(n5952)
         );
  INV_X1 U7670 ( .A(n5952), .ZN(n5953) );
  NAND2_X1 U7671 ( .A1(n6040), .A2(n8370), .ZN(n8103) );
  NAND2_X1 U7672 ( .A1(n4297), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U7673 ( .A1(n8495), .A2(n8172), .ZN(n6046) );
  NAND2_X1 U7674 ( .A1(n5956), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5957) );
  MUX2_X1 U7675 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5957), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n5958) );
  INV_X1 U7676 ( .A(n5959), .ZN(n5960) );
  NAND2_X1 U7677 ( .A1(n5960), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5961) );
  NAND2_X1 U7678 ( .A1(n6945), .A2(n8165), .ZN(n5962) );
  NAND2_X1 U7679 ( .A1(n5963), .A2(n8719), .ZN(n6003) );
  NAND2_X1 U7680 ( .A1(n7983), .A2(n7977), .ZN(n6933) );
  NAND2_X1 U7681 ( .A1(n6933), .A2(n5965), .ZN(n7234) );
  NAND2_X1 U7682 ( .A1(n7234), .A2(n7984), .ZN(n7235) );
  NAND2_X1 U7683 ( .A1(n7235), .A2(n7988), .ZN(n6970) );
  INV_X1 U7684 ( .A(n8131), .ZN(n6969) );
  NAND2_X1 U7685 ( .A1(n8379), .A2(n9827), .ZN(n7998) );
  NAND2_X1 U7686 ( .A1(n7167), .A2(n7998), .ZN(n5966) );
  OR2_X1 U7687 ( .A1(n8379), .A2(n9827), .ZN(n8004) );
  NAND2_X1 U7688 ( .A1(n5966), .A2(n8004), .ZN(n7255) );
  OR2_X1 U7689 ( .A1(n8378), .A2(n9832), .ZN(n8005) );
  NAND2_X1 U7690 ( .A1(n8378), .A2(n9832), .ZN(n8009) );
  AND2_X1 U7691 ( .A1(n8377), .A2(n7360), .ZN(n8000) );
  INV_X1 U7692 ( .A(n8000), .ZN(n8008) );
  NAND2_X1 U7693 ( .A1(n8010), .A2(n8008), .ZN(n8137) );
  AND2_X1 U7694 ( .A1(n8016), .A2(n7407), .ZN(n8025) );
  INV_X1 U7695 ( .A(n8021), .ZN(n5967) );
  NAND2_X1 U7696 ( .A1(n9856), .A2(n7773), .ZN(n8022) );
  NAND2_X1 U7697 ( .A1(n7607), .A2(n8142), .ZN(n7606) );
  INV_X1 U7698 ( .A(n8034), .ZN(n5968) );
  NAND2_X1 U7699 ( .A1(n9860), .A2(n8310), .ZN(n8032) );
  XNOR2_X1 U7700 ( .A(n9871), .B(n9664), .ZN(n8044) );
  OR2_X1 U7701 ( .A1(n9871), .A2(n9664), .ZN(n8042) );
  NOR2_X1 U7702 ( .A1(n9654), .A2(n8242), .ZN(n8046) );
  AND2_X1 U7703 ( .A1(n9654), .A2(n8242), .ZN(n8047) );
  XNOR2_X1 U7704 ( .A(n8793), .B(n9662), .ZN(n8722) );
  OR2_X2 U7705 ( .A1(n8732), .A2(n8722), .ZN(n8733) );
  OR2_X1 U7706 ( .A1(n8793), .A2(n9662), .ZN(n8052) );
  INV_X1 U7707 ( .A(n8725), .ZN(n8284) );
  NAND2_X1 U7708 ( .A1(n8871), .A2(n8284), .ZN(n8057) );
  NAND2_X1 U7709 ( .A1(n8702), .A2(n8057), .ZN(n5970) );
  OR2_X1 U7710 ( .A1(n8871), .A2(n8284), .ZN(n8055) );
  NAND2_X1 U7711 ( .A1(n5970), .A2(n8055), .ZN(n8689) );
  NAND2_X1 U7712 ( .A1(n8689), .A2(n8063), .ZN(n5971) );
  NAND2_X1 U7713 ( .A1(n8677), .A2(n8679), .ZN(n8649) );
  INV_X1 U7714 ( .A(n8066), .ZN(n5973) );
  NAND2_X1 U7715 ( .A1(n8069), .A2(n8651), .ZN(n8062) );
  INV_X1 U7716 ( .A(n8062), .ZN(n5972) );
  AND2_X1 U7717 ( .A1(n8650), .A2(n5975), .ZN(n5974) );
  INV_X1 U7718 ( .A(n5975), .ZN(n5977) );
  NAND2_X1 U7719 ( .A1(n8779), .A2(n8683), .ZN(n8067) );
  AND2_X1 U7720 ( .A1(n8664), .A2(n8066), .ZN(n5976) );
  NOR2_X1 U7721 ( .A1(n7973), .A2(n5979), .ZN(n8071) );
  AND2_X1 U7722 ( .A1(n7972), .A2(n8622), .ZN(n8070) );
  NAND2_X1 U7723 ( .A1(n5981), .A2(n5980), .ZN(n8592) );
  INV_X1 U7724 ( .A(n5984), .ZN(n5982) );
  NAND2_X1 U7725 ( .A1(n8822), .A2(n8251), .ZN(n8128) );
  NAND2_X1 U7726 ( .A1(n5984), .A2(n8326), .ZN(n8585) );
  NAND2_X1 U7727 ( .A1(n8128), .A2(n8585), .ZN(n8080) );
  INV_X1 U7728 ( .A(n8080), .ZN(n5985) );
  NOR2_X1 U7729 ( .A1(n8816), .A2(n8303), .ZN(n8087) );
  OR2_X2 U7730 ( .A1(n8570), .A2(n8087), .ZN(n5987) );
  AND2_X1 U7731 ( .A1(n8816), .A2(n8303), .ZN(n8086) );
  INV_X1 U7732 ( .A(n8086), .ZN(n5986) );
  NAND2_X1 U7733 ( .A1(n8353), .A2(n8553), .ZN(n7958) );
  INV_X1 U7734 ( .A(n7958), .ZN(n8536) );
  NAND2_X1 U7735 ( .A1(n8812), .A2(n8350), .ZN(n8539) );
  NAND2_X1 U7736 ( .A1(n8806), .A2(n8554), .ZN(n5988) );
  XNOR2_X1 U7737 ( .A(n8119), .B(n4418), .ZN(n8535) );
  NAND2_X1 U7738 ( .A1(n7404), .A2(n7499), .ZN(n6852) );
  NAND2_X1 U7739 ( .A1(n6783), .A2(n9842), .ZN(n6880) );
  INV_X1 U7740 ( .A(n8172), .ZN(n7976) );
  OR2_X1 U7741 ( .A1(n8495), .A2(n7976), .ZN(n6034) );
  AND2_X1 U7742 ( .A1(n6852), .A2(n6034), .ZN(n5990) );
  OR2_X1 U7743 ( .A1(n5991), .A2(n8474), .ZN(n5993) );
  NAND2_X1 U7744 ( .A1(n5993), .A2(n6324), .ZN(n6766) );
  INV_X1 U7745 ( .A(n6766), .ZN(n6858) );
  INV_X1 U7746 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8527) );
  NAND2_X1 U7747 ( .A1(n4268), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U7748 ( .A1(n7108), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5994) );
  OAI211_X1 U7749 ( .C1(n8527), .C2(n7111), .A(n5995), .B(n5994), .ZN(n5996)
         );
  INV_X1 U7750 ( .A(n5996), .ZN(n5997) );
  AND2_X1 U7751 ( .A1(n7114), .A2(n5997), .ZN(n8102) );
  NAND2_X1 U7752 ( .A1(n6324), .A2(P2_B_REG_SCAN_IN), .ZN(n5998) );
  NAND2_X1 U7753 ( .A1(n8726), .A2(n5998), .ZN(n8520) );
  OAI22_X1 U7754 ( .A1(n8554), .A2(n9665), .B1(n8102), .B2(n8520), .ZN(n5999)
         );
  INV_X1 U7755 ( .A(n5999), .ZN(n6000) );
  NAND2_X1 U7756 ( .A1(n8495), .A2(n7499), .ZN(n7239) );
  INV_X1 U7757 ( .A(n9852), .ZN(n9824) );
  NAND2_X1 U7758 ( .A1(n6031), .A2(n6032), .ZN(n6005) );
  NAND2_X1 U7759 ( .A1(n6005), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6008) );
  INV_X1 U7760 ( .A(n6010), .ZN(n6014) );
  NAND2_X1 U7761 ( .A1(n6011), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6012) );
  INV_X1 U7762 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6020) );
  NOR2_X1 U7763 ( .A1(n6017), .A2(n6018), .ZN(n6019) );
  INV_X1 U7764 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6394) );
  NAND2_X1 U7765 ( .A1(n8881), .A2(n6850), .ZN(n6045) );
  NOR2_X1 U7766 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .ZN(
        n9917) );
  NOR4_X1 U7767 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n6023) );
  NOR4_X1 U7768 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n6022) );
  NOR4_X1 U7769 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6021) );
  NAND4_X1 U7770 ( .A1(n9917), .A2(n6023), .A3(n6022), .A4(n6021), .ZN(n6029)
         );
  NOR4_X1 U7771 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6027) );
  NOR4_X1 U7772 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6026) );
  NOR4_X1 U7773 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n6025) );
  NOR4_X1 U7774 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6024) );
  NAND4_X1 U7775 ( .A1(n6027), .A2(n6026), .A3(n6025), .A4(n6024), .ZN(n6028)
         );
  OAI21_X1 U7776 ( .B1(n6029), .B2(n6028), .A(n6391), .ZN(n6044) );
  NOR2_X1 U7777 ( .A1(n7911), .A2(n7902), .ZN(n6030) );
  NAND2_X1 U7778 ( .A1(n6852), .A2(n8051), .ZN(n6778) );
  AND3_X1 U7779 ( .A1(n6044), .A2(n8880), .A3(n6778), .ZN(n6033) );
  NOR2_X1 U7780 ( .A1(n9852), .A2(n6945), .ZN(n6772) );
  INV_X1 U7781 ( .A(n6850), .ZN(n6036) );
  OR2_X1 U7782 ( .A1(n6034), .A2(n7499), .ZN(n6035) );
  OAI21_X1 U7783 ( .B1(n6772), .B2(n6036), .A(n6874), .ZN(n6038) );
  INV_X1 U7784 ( .A(n8881), .ZN(n6049) );
  INV_X1 U7785 ( .A(n6874), .ZN(n6872) );
  NAND2_X1 U7786 ( .A1(n6049), .A2(n6872), .ZN(n6037) );
  NAND2_X1 U7787 ( .A1(n9890), .A2(n9872), .ZN(n8785) );
  INV_X1 U7788 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6041) );
  OAI21_X1 U7789 ( .B1(n6058), .B2(n8746), .A(n6043), .ZN(P2_U3488) );
  INV_X1 U7790 ( .A(n6044), .ZN(n6048) );
  NOR2_X1 U7791 ( .A1(n6045), .A2(n6048), .ZN(n6775) );
  NAND2_X1 U7792 ( .A1(n6775), .A2(n8880), .ZN(n6771) );
  OR2_X1 U7793 ( .A1(n6046), .A2(n6848), .ZN(n6781) );
  AND2_X1 U7794 ( .A1(n6783), .A2(n6781), .ZN(n6047) );
  NOR2_X1 U7795 ( .A1(n6850), .A2(n6048), .ZN(n6050) );
  NAND2_X1 U7796 ( .A1(n6786), .A2(n8880), .ZN(n6768) );
  AND2_X1 U7797 ( .A1(n9842), .A2(n8110), .ZN(n6051) );
  NAND2_X1 U7798 ( .A1(n6781), .A2(n6051), .ZN(n6767) );
  NAND2_X1 U7799 ( .A1(n7239), .A2(n9872), .ZN(n8714) );
  AND2_X1 U7800 ( .A1(n6767), .A2(n8714), .ZN(n6774) );
  OR2_X1 U7801 ( .A1(n6768), .A2(n6774), .ZN(n6052) );
  NAND2_X1 U7802 ( .A1(n9873), .A2(n9872), .ZN(n8863) );
  INV_X1 U7803 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6054) );
  OR2_X1 U7804 ( .A1(n9873), .A2(n6054), .ZN(n6055) );
  INV_X1 U7805 ( .A(n6056), .ZN(n6057) );
  OAI21_X1 U7806 ( .B1(n6058), .B2(n9875), .A(n6057), .ZN(P2_U3456) );
  XNOR2_X1 U7807 ( .A(n6060), .B(n6059), .ZN(n9294) );
  AOI21_X1 U7808 ( .B1(n6156), .B2(n6251), .A(n6061), .ZN(n6067) );
  OAI21_X1 U7809 ( .B1(n6061), .B2(n6062), .A(n9463), .ZN(n6066) );
  NAND2_X1 U7810 ( .A1(n9192), .A2(n9129), .ZN(n6064) );
  INV_X1 U7811 ( .A(n9169), .ZN(n9138) );
  NAND2_X1 U7812 ( .A1(n9194), .A2(n9138), .ZN(n6063) );
  NAND2_X1 U7813 ( .A1(n6064), .A2(n6063), .ZN(n9007) );
  INV_X1 U7814 ( .A(n9007), .ZN(n6065) );
  OAI21_X1 U7815 ( .B1(n6067), .B2(n6066), .A(n6065), .ZN(n9293) );
  AOI211_X1 U7816 ( .C1(n9010), .C2(n9312), .A(n9443), .B(n4304), .ZN(n9299)
         );
  AOI21_X1 U7817 ( .B1(n9294), .B2(n9801), .A(n6068), .ZN(n6319) );
  OAI21_X1 U7818 ( .B1(n6319), .B2(n9619), .A(n6072), .ZN(P1_U3517) );
  AND2_X1 U7819 ( .A1(n4682), .A2(n6623), .ZN(n6168) );
  NAND2_X1 U7820 ( .A1(n9333), .A2(n6073), .ZN(n6213) );
  OR2_X1 U7821 ( .A1(n9513), .A2(n9079), .ZN(n6074) );
  NAND2_X1 U7822 ( .A1(n6147), .A2(n6074), .ZN(n6210) );
  MUX2_X1 U7823 ( .A(n6213), .B(n6210), .S(n6168), .Z(n6150) );
  NAND2_X1 U7824 ( .A1(n6144), .A2(n6077), .ZN(n6214) );
  AND2_X1 U7825 ( .A1(n6215), .A2(n6078), .ZN(n6211) );
  INV_X1 U7826 ( .A(n6211), .ZN(n6076) );
  MUX2_X1 U7827 ( .A(n6214), .B(n6076), .S(n6310), .Z(n6146) );
  NAND3_X1 U7828 ( .A1(n6077), .A2(n6310), .A3(n9200), .ZN(n6143) );
  NAND2_X1 U7829 ( .A1(n6078), .A2(n6168), .ZN(n6079) );
  OAI21_X1 U7830 ( .B1(n6247), .B2(n9529), .A(n6079), .ZN(n6080) );
  NAND2_X1 U7831 ( .A1(n6080), .A2(n6136), .ZN(n6142) );
  INV_X1 U7832 ( .A(n6265), .ZN(n6081) );
  OAI211_X1 U7833 ( .C1(n6086), .C2(n6081), .A(n6087), .B(n7071), .ZN(n6083)
         );
  AND2_X1 U7834 ( .A1(n6088), .A2(n6264), .ZN(n6082) );
  AOI21_X1 U7835 ( .B1(n6083), .B2(n6082), .A(n4657), .ZN(n6092) );
  INV_X1 U7836 ( .A(n6084), .ZN(n6085) );
  OAI211_X1 U7837 ( .C1(n6086), .C2(n6085), .A(n6264), .B(n6262), .ZN(n6090)
         );
  AND2_X1 U7838 ( .A1(n6236), .A2(n6087), .ZN(n6089) );
  INV_X1 U7839 ( .A(n6088), .ZN(n7177) );
  AOI21_X1 U7840 ( .B1(n6090), .B2(n6089), .A(n7177), .ZN(n6091) );
  MUX2_X1 U7841 ( .A(n6092), .B(n6091), .S(n6168), .Z(n6097) );
  INV_X1 U7842 ( .A(n6093), .ZN(n6095) );
  MUX2_X1 U7843 ( .A(n6095), .B(n6094), .S(n6168), .Z(n6096) );
  OAI21_X1 U7844 ( .B1(n6097), .B2(n7176), .A(n6096), .ZN(n6101) );
  AND2_X1 U7845 ( .A1(n6107), .A2(n6098), .ZN(n6099) );
  MUX2_X1 U7846 ( .A(n7325), .B(n6099), .S(n6168), .Z(n6100) );
  NAND2_X1 U7847 ( .A1(n6101), .A2(n6100), .ZN(n6109) );
  INV_X1 U7848 ( .A(n6110), .ZN(n6102) );
  AOI21_X1 U7849 ( .B1(n6109), .B2(n6106), .A(n6102), .ZN(n6104) );
  NAND2_X1 U7850 ( .A1(n6114), .A2(n6112), .ZN(n6103) );
  OAI211_X1 U7851 ( .C1(n6104), .C2(n6103), .A(n6273), .B(n6111), .ZN(n6105)
         );
  NAND2_X1 U7852 ( .A1(n6105), .A2(n6115), .ZN(n6118) );
  INV_X1 U7853 ( .A(n6106), .ZN(n6108) );
  OAI21_X1 U7854 ( .B1(n6109), .B2(n6108), .A(n6107), .ZN(n6113) );
  NAND2_X1 U7855 ( .A1(n6111), .A2(n6110), .ZN(n6270) );
  AOI21_X1 U7856 ( .B1(n6113), .B2(n6112), .A(n6270), .ZN(n6116) );
  NAND2_X1 U7857 ( .A1(n6115), .A2(n6114), .ZN(n6274) );
  OAI21_X1 U7858 ( .B1(n6116), .B2(n6274), .A(n6273), .ZN(n6117) );
  MUX2_X1 U7859 ( .A(n6118), .B(n6117), .S(n6310), .Z(n6123) );
  NAND2_X1 U7860 ( .A1(n6123), .A2(n6276), .ZN(n6119) );
  NAND3_X1 U7861 ( .A1(n6119), .A2(n6272), .A3(n6278), .ZN(n6121) );
  NAND4_X1 U7862 ( .A1(n6121), .A2(n6284), .A3(n6120), .A4(n6283), .ZN(n6129)
         );
  NAND2_X1 U7863 ( .A1(n6287), .A2(n6279), .ZN(n6130) );
  INV_X1 U7864 ( .A(n6278), .ZN(n6122) );
  NAND2_X1 U7865 ( .A1(n6123), .A2(n6272), .ZN(n6124) );
  NAND3_X1 U7866 ( .A1(n6124), .A2(n7784), .A3(n6276), .ZN(n6128) );
  INV_X1 U7867 ( .A(n6283), .ZN(n6125) );
  NAND2_X1 U7868 ( .A1(n6287), .A2(n6125), .ZN(n6126) );
  NAND2_X1 U7869 ( .A1(n6126), .A2(n6284), .ZN(n6127) );
  NAND3_X1 U7870 ( .A1(n6130), .A2(n6310), .A3(n6284), .ZN(n6131) );
  NAND2_X1 U7871 ( .A1(n9407), .A2(n9424), .ZN(n6285) );
  INV_X1 U7872 ( .A(n6285), .ZN(n6133) );
  NAND2_X1 U7873 ( .A1(n6293), .A2(n6135), .ZN(n6132) );
  AOI21_X1 U7874 ( .B1(n6138), .B2(n6133), .A(n6132), .ZN(n6141) );
  NAND2_X1 U7875 ( .A1(n9540), .A2(n9154), .ZN(n6134) );
  NAND2_X1 U7876 ( .A1(n6135), .A2(n6134), .ZN(n6289) );
  INV_X1 U7877 ( .A(n6289), .ZN(n6139) );
  AND2_X1 U7878 ( .A1(n6136), .A2(n9407), .ZN(n6288) );
  INV_X1 U7879 ( .A(n6288), .ZN(n6137) );
  AOI21_X1 U7880 ( .B1(n6139), .B2(n6138), .A(n6137), .ZN(n6140) );
  MUX2_X1 U7881 ( .A(n6215), .B(n6144), .S(n6310), .Z(n6145) );
  MUX2_X1 U7882 ( .A(n9333), .B(n6147), .S(n6310), .Z(n6148) );
  OAI211_X1 U7883 ( .C1(n6150), .C2(n6149), .A(n9339), .B(n6148), .ZN(n6152)
         );
  MUX2_X1 U7884 ( .A(n6216), .B(n5384), .S(n6168), .Z(n6151) );
  INV_X1 U7885 ( .A(n6153), .ZN(n6155) );
  OAI21_X1 U7886 ( .B1(n9010), .B2(n6310), .A(n6158), .ZN(n6157) );
  INV_X1 U7887 ( .A(n6162), .ZN(n6161) );
  OAI21_X1 U7888 ( .B1(n9193), .B2(n6159), .A(n6223), .ZN(n6160) );
  INV_X1 U7889 ( .A(n6297), .ZN(n6229) );
  INV_X1 U7890 ( .A(SI_29_), .ZN(n6174) );
  INV_X1 U7891 ( .A(n6169), .ZN(n6172) );
  INV_X1 U7892 ( .A(n6170), .ZN(n6171) );
  NAND2_X1 U7893 ( .A1(n6172), .A2(n6171), .ZN(n6173) );
  INV_X1 U7894 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8892) );
  INV_X1 U7895 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n6176) );
  MUX2_X1 U7896 ( .A(n8892), .B(n6176), .S(n6348), .Z(n6178) );
  INV_X1 U7897 ( .A(SI_30_), .ZN(n6177) );
  NAND2_X1 U7898 ( .A1(n6178), .A2(n6177), .ZN(n6183) );
  INV_X1 U7899 ( .A(n6178), .ZN(n6179) );
  NAND2_X1 U7900 ( .A1(n6179), .A2(SI_30_), .ZN(n6180) );
  NAND2_X1 U7901 ( .A1(n6183), .A2(n6180), .ZN(n6184) );
  NAND2_X1 U7902 ( .A1(n8889), .A2(n6191), .ZN(n6182) );
  NAND2_X1 U7903 ( .A1(n6190), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6181) );
  INV_X1 U7904 ( .A(n9562), .ZN(n6301) );
  INV_X1 U7905 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8114) );
  INV_X1 U7906 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6186) );
  MUX2_X1 U7907 ( .A(n8114), .B(n6186), .S(n6348), .Z(n6187) );
  XNOR2_X1 U7908 ( .A(n6187), .B(SI_31_), .ZN(n6188) );
  INV_X1 U7909 ( .A(n9558), .ZN(n6200) );
  NAND3_X1 U7910 ( .A1(n6192), .A2(n6200), .A3(n9191), .ZN(n6204) );
  INV_X1 U7911 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9556) );
  NAND2_X1 U7912 ( .A1(n5137), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U7913 ( .A1(n6193), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6194) );
  OAI211_X1 U7914 ( .C1(n6196), .C2(n9556), .A(n6195), .B(n6194), .ZN(n9271)
         );
  NAND2_X1 U7915 ( .A1(n9271), .A2(n9191), .ZN(n6230) );
  NAND2_X1 U7916 ( .A1(n6314), .A2(n6230), .ZN(n6198) );
  INV_X1 U7917 ( .A(n9271), .ZN(n6199) );
  INV_X1 U7918 ( .A(n6230), .ZN(n6231) );
  NOR2_X1 U7919 ( .A1(n6207), .A2(n6206), .ZN(n6294) );
  INV_X1 U7920 ( .A(n6294), .ZN(n6228) );
  AOI21_X1 U7921 ( .B1(n9333), .B2(n6210), .A(n9320), .ZN(n6212) );
  NAND4_X1 U7922 ( .A1(n6222), .A2(n6211), .A3(n6212), .A4(n6221), .ZN(n6291)
         );
  INV_X1 U7923 ( .A(n6291), .ZN(n6226) );
  INV_X1 U7924 ( .A(n6212), .ZN(n6218) );
  AOI21_X1 U7925 ( .B1(n6215), .B2(n6214), .A(n6213), .ZN(n6217) );
  OAI21_X1 U7926 ( .B1(n6218), .B2(n6217), .A(n6216), .ZN(n6220) );
  AOI21_X1 U7927 ( .B1(n6221), .B2(n6220), .A(n6219), .ZN(n6225) );
  INV_X1 U7928 ( .A(n6222), .ZN(n6224) );
  OAI21_X1 U7929 ( .B1(n6225), .B2(n6224), .A(n6223), .ZN(n6295) );
  AOI21_X1 U7930 ( .B1(n6231), .B2(n9562), .A(n4336), .ZN(n6232) );
  OAI211_X1 U7931 ( .C1(n6232), .C2(n6300), .A(n6549), .B(n6311), .ZN(n6256)
         );
  INV_X1 U7932 ( .A(n6233), .ZN(n7002) );
  NAND2_X1 U7933 ( .A1(n9219), .A2(n6487), .ZN(n6261) );
  NAND2_X1 U7934 ( .A1(n7002), .A2(n6261), .ZN(n6462) );
  NOR2_X1 U7935 ( .A1(n6462), .A2(n6479), .ZN(n6235) );
  INV_X1 U7936 ( .A(n7015), .ZN(n6234) );
  INV_X1 U7937 ( .A(n6921), .ZN(n6919) );
  AND4_X1 U7938 ( .A1(n6235), .A2(n6983), .A3(n6234), .A4(n6919), .ZN(n6237)
         );
  INV_X1 U7939 ( .A(n7079), .ZN(n7070) );
  NAND4_X1 U7940 ( .A1(n6237), .A2(n7070), .A3(n6236), .A4(n7003), .ZN(n6238)
         );
  OR4_X1 U7941 ( .A1(n7427), .A2(n6240), .A3(n6239), .A4(n6238), .ZN(n6241) );
  OR3_X1 U7942 ( .A1(n7622), .A2(n6241), .A3(n7643), .ZN(n6243) );
  INV_X1 U7943 ( .A(n7784), .ZN(n6242) );
  OR4_X1 U7944 ( .A1(n7728), .A2(n6243), .A3(n6242), .A4(n7891), .ZN(n6244) );
  NOR2_X1 U7945 ( .A1(n9468), .A2(n6244), .ZN(n6245) );
  NAND4_X1 U7946 ( .A1(n9409), .A2(n9423), .A3(n6245), .A4(n9452), .ZN(n6246)
         );
  NOR2_X1 U7947 ( .A1(n6247), .A2(n6246), .ZN(n6248) );
  AND2_X1 U7948 ( .A1(n9377), .A2(n6248), .ZN(n6249) );
  NAND4_X1 U7949 ( .A1(n9339), .A2(n9351), .A3(n6249), .A4(n9364), .ZN(n6250)
         );
  OR3_X1 U7950 ( .A1(n9307), .A2(n9319), .A3(n6250), .ZN(n6252) );
  OR3_X1 U7951 ( .A1(n6252), .A2(n9283), .A3(n6251), .ZN(n6253) );
  NOR2_X1 U7952 ( .A1(n4566), .A2(n6253), .ZN(n6255) );
  XNOR2_X1 U7953 ( .A(n6301), .B(n9191), .ZN(n6254) );
  NAND4_X1 U7954 ( .A1(n6314), .A2(n6311), .A3(n6255), .A4(n6254), .ZN(n6258)
         );
  NAND2_X1 U7955 ( .A1(n6258), .A2(n6623), .ZN(n6259) );
  AND3_X1 U7956 ( .A1(n6263), .A2(n6262), .A3(n6261), .ZN(n6267) );
  AOI21_X1 U7957 ( .B1(n6559), .B2(n7051), .A(n7605), .ZN(n6266) );
  NAND4_X1 U7958 ( .A1(n6267), .A2(n6266), .A3(n6265), .A4(n6264), .ZN(n6269)
         );
  AOI211_X1 U7959 ( .C1(n7420), .C2(n6269), .A(n6268), .B(n7419), .ZN(n6271)
         );
  NOR2_X1 U7960 ( .A1(n6271), .A2(n6270), .ZN(n6275) );
  OAI211_X1 U7961 ( .C1(n6275), .C2(n6274), .A(n6273), .B(n6272), .ZN(n6277)
         );
  NAND2_X1 U7962 ( .A1(n6277), .A2(n6276), .ZN(n6281) );
  OAI211_X1 U7963 ( .C1(n6281), .C2(n6280), .A(n6279), .B(n6278), .ZN(n6282)
         );
  NAND3_X1 U7964 ( .A1(n6284), .A2(n6283), .A3(n6282), .ZN(n6286) );
  AOI21_X1 U7965 ( .B1(n6287), .B2(n6286), .A(n6285), .ZN(n6290) );
  OAI21_X1 U7966 ( .B1(n6290), .B2(n6289), .A(n6288), .ZN(n6292) );
  AOI21_X1 U7967 ( .B1(n6293), .B2(n6292), .A(n6291), .ZN(n6296) );
  OAI21_X1 U7968 ( .B1(n6296), .B2(n6295), .A(n6294), .ZN(n6298) );
  AOI22_X1 U7969 ( .A1(n6298), .A2(n6297), .B1(n9562), .B2(n9191), .ZN(n6299)
         );
  AOI211_X1 U7970 ( .C1(n6302), .C2(n6301), .A(n6300), .B(n6299), .ZN(n6304)
         );
  NAND2_X1 U7971 ( .A1(n6305), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6525) );
  NOR2_X1 U7972 ( .A1(n6307), .A2(n6557), .ZN(n6306) );
  AOI211_X1 U7973 ( .C1(n6307), .C2(n6480), .A(n6525), .B(n6306), .ZN(n6308)
         );
  NOR3_X1 U7974 ( .A1(n6525), .A2(n6481), .A3(n6312), .ZN(n6313) );
  NAND2_X1 U7975 ( .A1(n6632), .A2(n9635), .ZN(n6315) );
  OAI21_X1 U7976 ( .B1(n6525), .B2(n6481), .A(P1_B_REG_SCAN_IN), .ZN(n6316) );
  INV_X1 U7977 ( .A(n6316), .ZN(n6317) );
  INV_X1 U7978 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6320) );
  INV_X1 U7979 ( .A(n6521), .ZN(n6484) );
  INV_X1 U7980 ( .A(n6393), .ZN(n6322) );
  NAND2_X1 U7981 ( .A1(n6777), .A2(n8110), .ZN(n6323) );
  NAND2_X1 U7982 ( .A1(n6323), .A2(n6776), .ZN(n6471) );
  NAND2_X1 U7983 ( .A1(n6471), .A2(n6324), .ZN(n6325) );
  NAND2_X1 U7984 ( .A1(n6325), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NAND2_X1 U7985 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n6332) );
  INV_X1 U7986 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6326) );
  MUX2_X1 U7987 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6326), .S(n6401), .Z(n6331)
         );
  NOR3_X1 U7988 ( .A1(n6331), .A2(n6486), .A3(n6327), .ZN(n6402) );
  NAND2_X1 U7989 ( .A1(n6556), .A2(n6525), .ZN(n6337) );
  NAND2_X1 U7990 ( .A1(n6328), .A2(n6549), .ZN(n6330) );
  AND2_X1 U7991 ( .A1(n6330), .A2(n6329), .ZN(n6336) );
  AND2_X1 U7992 ( .A1(n6337), .A2(n6336), .ZN(n6369) );
  NAND2_X1 U7993 ( .A1(n6369), .A2(n6489), .ZN(n9718) );
  AOI211_X1 U7994 ( .C1(n6332), .C2(n6331), .A(n6402), .B(n9718), .ZN(n6344)
         );
  AND2_X1 U7995 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6490) );
  INV_X1 U7996 ( .A(n6490), .ZN(n6335) );
  NOR2_X1 U7997 ( .A1(n6334), .A2(n6335), .ZN(n6407) );
  NOR2_X1 U7998 ( .A1(n6366), .A2(n6489), .ZN(n6333) );
  AOI211_X1 U7999 ( .C1(n6335), .C2(n6334), .A(n6407), .B(n9730), .ZN(n6343)
         );
  NAND2_X1 U8000 ( .A1(n6369), .A2(n6366), .ZN(n9739) );
  NOR2_X1 U8001 ( .A1(n9739), .A2(n6401), .ZN(n6342) );
  INV_X1 U8002 ( .A(n6336), .ZN(n6338) );
  INV_X1 U8003 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6340) );
  OAI22_X1 U8004 ( .A1(n9746), .A2(n6340), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6339), .ZN(n6341) );
  OR4_X1 U8005 ( .A1(n6344), .A2(n6343), .A3(n6342), .A4(n6341), .ZN(P1_U3244)
         );
  AND2_X1 U8006 ( .A1(n6348), .A2(P2_U3151), .ZN(n8899) );
  INV_X2 U8007 ( .A(n8899), .ZN(n8893) );
  INV_X1 U8008 ( .A(n6603), .ZN(n6725) );
  NAND2_X1 U8009 ( .A1(n6345), .A2(P2_U3151), .ZN(n8891) );
  OAI222_X1 U8010 ( .A1(n8893), .A2(n4886), .B1(n6725), .B2(P2_U3151), .C1(
        n8891), .C2(n6362), .ZN(P2_U3293) );
  INV_X1 U8011 ( .A(n6668), .ZN(n6605) );
  OAI222_X1 U8012 ( .A1(n8893), .A2(n6346), .B1(n6605), .B2(P2_U3151), .C1(
        n8891), .C2(n6350), .ZN(P2_U3292) );
  INV_X1 U8013 ( .A(n6751), .ZN(n6749) );
  OAI222_X1 U8014 ( .A1(n8893), .A2(n6347), .B1(n6749), .B2(P2_U3151), .C1(
        n8891), .C2(n6354), .ZN(P2_U3291) );
  NAND2_X1 U8015 ( .A1(n6348), .A2(P1_U3086), .ZN(n9637) );
  CLKBUF_X1 U8016 ( .A(n9637), .Z(n9626) );
  NOR2_X2 U8017 ( .A1(n6348), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9634) );
  AOI22_X1 U8018 ( .A1(n6433), .A2(P1_STATE_REG_SCAN_IN), .B1(n9634), .B2(
        P2_DATAO_REG_3__SCAN_IN), .ZN(n6349) );
  OAI21_X1 U8019 ( .B1(n6350), .B2(n9626), .A(n6349), .ZN(P1_U3352) );
  INV_X1 U8020 ( .A(n8891), .ZN(n7749) );
  INV_X1 U8021 ( .A(n7749), .ZN(n8901) );
  INV_X1 U8022 ( .A(n6802), .ZN(n6754) );
  OAI222_X1 U8023 ( .A1(n8901), .A2(n6364), .B1(n6754), .B2(P2_U3151), .C1(
        n4903), .C2(n8893), .ZN(P2_U3290) );
  INV_X1 U8024 ( .A(n6351), .ZN(n6361) );
  INV_X1 U8025 ( .A(n6651), .ZN(n6592) );
  OAI222_X1 U8026 ( .A1(n8901), .A2(n6361), .B1(n8893), .B2(n4881), .C1(
        P2_U3151), .C2(n6592), .ZN(P2_U3294) );
  INV_X1 U8027 ( .A(n6808), .ZN(n6841) );
  OAI222_X1 U8028 ( .A1(n8901), .A2(n6356), .B1(n6841), .B2(P2_U3151), .C1(
        n6352), .C2(n8893), .ZN(P2_U3289) );
  INV_X1 U8029 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6353) );
  OAI222_X1 U8030 ( .A1(n8901), .A2(n6358), .B1(n4703), .B2(P2_U3151), .C1(
        n6353), .C2(n8893), .ZN(P2_U3288) );
  INV_X1 U8031 ( .A(n9634), .ZN(n8213) );
  OAI222_X1 U8032 ( .A1(n8213), .A2(n6355), .B1(n9626), .B2(n6354), .C1(n6501), 
        .C2(P1_U3086), .ZN(P1_U3351) );
  OAI222_X1 U8033 ( .A1(n8213), .A2(n6357), .B1(n9626), .B2(n6356), .C1(n6414), 
        .C2(P1_U3086), .ZN(P1_U3349) );
  OAI222_X1 U8034 ( .A1(n8213), .A2(n6359), .B1(n9626), .B2(n6358), .C1(n6454), 
        .C2(P1_U3086), .ZN(P1_U3348) );
  OAI222_X1 U8035 ( .A1(P1_U3086), .A2(n6401), .B1(n9626), .B2(n6361), .C1(
        n6360), .C2(n8213), .ZN(P1_U3354) );
  INV_X1 U8036 ( .A(n6409), .ZN(n6512) );
  OAI222_X1 U8037 ( .A1(n8213), .A2(n6363), .B1(n9626), .B2(n6362), .C1(n6512), 
        .C2(P1_U3086), .ZN(P1_U3353) );
  OAI222_X1 U8038 ( .A1(n8213), .A2(n6365), .B1(n9626), .B2(n6364), .C1(n6403), 
        .C2(P1_U3086), .ZN(P1_U3350) );
  INV_X1 U8039 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6371) );
  INV_X1 U8040 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6636) );
  AOI21_X1 U8041 ( .B1(n9635), .B2(n6636), .A(n6366), .ZN(n6491) );
  OAI21_X1 U8042 ( .B1(n9635), .B2(P1_REG1_REG_0__SCAN_IN), .A(n6491), .ZN(
        n6367) );
  XNOR2_X1 U8043 ( .A(n6367), .B(P1_IR_REG_0__SCAN_IN), .ZN(n6368) );
  AOI22_X1 U8044 ( .A1(n6369), .A2(n6368), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n6370) );
  OAI21_X1 U8045 ( .B1(n9746), .B2(n6371), .A(n6370), .ZN(P1_U3243) );
  INV_X1 U8046 ( .A(n9746), .ZN(n9247) );
  NOR2_X1 U8047 ( .A1(n9247), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8048 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6373) );
  INV_X1 U8049 ( .A(n6372), .ZN(n6374) );
  INV_X1 U8050 ( .A(n6902), .ZN(n7041) );
  OAI222_X1 U8051 ( .A1(n8893), .A2(n6373), .B1(n8891), .B2(n6374), .C1(
        P2_U3151), .C2(n7041), .ZN(P2_U3287) );
  OAI222_X1 U8052 ( .A1(n8213), .A2(n6375), .B1(n9626), .B2(n6374), .C1(
        P1_U3086), .C2(n6569), .ZN(P1_U3347) );
  NAND2_X1 U8053 ( .A1(n9271), .A2(P1_U3973), .ZN(n6376) );
  OAI21_X1 U8054 ( .B1(P1_U3973), .B2(n8114), .A(n6376), .ZN(P1_U3585) );
  NAND2_X1 U8055 ( .A1(n6559), .A2(P1_U3973), .ZN(n6377) );
  OAI21_X1 U8056 ( .B1(P1_U3973), .B2(n4881), .A(n6377), .ZN(P1_U3555) );
  NAND2_X1 U8057 ( .A1(n9772), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6379) );
  OAI21_X1 U8058 ( .B1(n9772), .B2(n6380), .A(n6379), .ZN(P1_U3439) );
  NAND2_X1 U8059 ( .A1(n9772), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6381) );
  OAI21_X1 U8060 ( .B1(n9772), .B2(n6382), .A(n6381), .ZN(P1_U3440) );
  AOI22_X1 U8061 ( .A1(n9649), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9634), .ZN(n6383) );
  OAI21_X1 U8062 ( .B1(n6387), .B2(n9626), .A(n6383), .ZN(P1_U3345) );
  INV_X1 U8063 ( .A(n6384), .ZN(n6389) );
  AOI22_X1 U8064 ( .A1(n7392), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9634), .ZN(n6385) );
  OAI21_X1 U8065 ( .B1(n6389), .B2(n9637), .A(n6385), .ZN(P1_U3346) );
  INV_X1 U8066 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6386) );
  OAI222_X1 U8067 ( .A1(n8901), .A2(n6387), .B1(n7340), .B2(P2_U3151), .C1(
        n6386), .C2(n8893), .ZN(P2_U3285) );
  OAI222_X1 U8068 ( .A1(n8901), .A2(n6389), .B1(n7154), .B2(P2_U3151), .C1(
        n6388), .C2(n8893), .ZN(P2_U3286) );
  NAND2_X1 U8069 ( .A1(n9218), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6390) );
  OAI21_X1 U8070 ( .B1(n9078), .B2(n9218), .A(n6390), .ZN(P1_U3574) );
  INV_X1 U8071 ( .A(n6391), .ZN(n6392) );
  NAND2_X1 U8072 ( .A1(n6392), .A2(n8880), .ZN(n6397) );
  AOI22_X1 U8073 ( .A1(n6397), .A2(n6394), .B1(n6393), .B2(n4854), .ZN(
        P2_U3376) );
  AND2_X1 U8074 ( .A1(n6397), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8075 ( .A1(n6397), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8076 ( .A1(n6397), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8077 ( .A1(n6397), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8078 ( .A1(n6397), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8079 ( .A1(n6397), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8080 ( .A1(n6397), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8081 ( .A1(n6397), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8082 ( .A1(n6397), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8083 ( .A1(n6397), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8084 ( .A1(n6397), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8085 ( .A1(n6397), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8086 ( .A1(n6397), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8087 ( .A1(n6397), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8088 ( .A1(n6397), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8089 ( .A1(n6397), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8090 ( .A1(n6397), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8091 ( .A1(n6397), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8092 ( .A1(n6397), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8093 ( .A1(n6397), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8094 ( .A1(n6397), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8095 ( .A1(n6397), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8096 ( .A1(n6397), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8097 ( .A1(n6397), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8098 ( .A1(n6397), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8099 ( .A1(n6397), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  INV_X1 U8100 ( .A(n6395), .ZN(n6399) );
  AOI22_X1 U8101 ( .A1(n9677), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9634), .ZN(n6396) );
  OAI21_X1 U8102 ( .B1(n6399), .B2(n9637), .A(n6396), .ZN(P1_U3344) );
  INV_X1 U8103 ( .A(n6397), .ZN(n6398) );
  INV_X1 U8104 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n9974) );
  NOR2_X1 U8105 ( .A1(n6398), .A2(n9974), .ZN(P2_U3255) );
  INV_X1 U8106 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n10011) );
  NOR2_X1 U8107 ( .A1(n6398), .A2(n10011), .ZN(P2_U3252) );
  INV_X1 U8108 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n10009) );
  NOR2_X1 U8109 ( .A1(n6398), .A2(n10009), .ZN(P2_U3259) );
  INV_X1 U8110 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n9975) );
  NOR2_X1 U8111 ( .A1(n6398), .A2(n9975), .ZN(P2_U3263) );
  INV_X1 U8112 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6400) );
  OAI222_X1 U8113 ( .A1(n8893), .A2(n6400), .B1(n8891), .B2(n6399), .C1(
        P2_U3151), .C2(n7445), .ZN(P2_U3284) );
  INV_X1 U8114 ( .A(n6403), .ZN(n6427) );
  INV_X1 U8115 ( .A(n6501), .ZN(n6410) );
  INV_X1 U8116 ( .A(n6401), .ZN(n6408) );
  XNOR2_X1 U8117 ( .A(n6409), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n6509) );
  NOR2_X1 U8118 ( .A1(n6510), .A2(n6509), .ZN(n6508) );
  AOI21_X1 U8119 ( .B1(n6409), .B2(P1_REG1_REG_2__SCAN_IN), .A(n6508), .ZN(
        n6441) );
  XNOR2_X1 U8120 ( .A(n6433), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n6440) );
  NOR2_X1 U8121 ( .A1(n6441), .A2(n6440), .ZN(n6439) );
  XOR2_X1 U8122 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6501), .Z(n6495) );
  NOR2_X1 U8123 ( .A1(n6496), .A2(n6495), .ZN(n6494) );
  AOI21_X1 U8124 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n6410), .A(n6494), .ZN(
        n6423) );
  XOR2_X1 U8125 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6403), .Z(n6422) );
  NOR2_X1 U8126 ( .A1(n6423), .A2(n6422), .ZN(n6421) );
  MUX2_X1 U8127 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6404), .S(n6414), .Z(n6405)
         );
  NOR2_X1 U8128 ( .A1(n6406), .A2(n6405), .ZN(n6447) );
  AOI211_X1 U8129 ( .C1(n6406), .C2(n6405), .A(n9718), .B(n6447), .ZN(n6420)
         );
  AOI21_X1 U8130 ( .B1(n6408), .B2(P1_REG2_REG_1__SCAN_IN), .A(n6407), .ZN(
        n6507) );
  XNOR2_X1 U8131 ( .A(n6409), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6506) );
  NOR2_X1 U8132 ( .A1(n6507), .A2(n6506), .ZN(n6505) );
  AOI21_X1 U8133 ( .B1(n6409), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6505), .ZN(
        n6438) );
  XNOR2_X1 U8134 ( .A(n6433), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n6437) );
  NOR2_X1 U8135 ( .A1(n6438), .A2(n6437), .ZN(n6436) );
  AOI21_X1 U8136 ( .B1(n6433), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6436), .ZN(
        n6499) );
  XNOR2_X1 U8137 ( .A(n6501), .B(n6992), .ZN(n6498) );
  NOR2_X1 U8138 ( .A1(n6499), .A2(n6498), .ZN(n6497) );
  AOI21_X1 U8139 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n6410), .A(n6497), .ZN(
        n6426) );
  XNOR2_X1 U8140 ( .A(n6427), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n6425) );
  MUX2_X1 U8141 ( .A(n5184), .B(P1_REG2_REG_6__SCAN_IN), .S(n6414), .Z(n6411)
         );
  INV_X1 U8142 ( .A(n6411), .ZN(n6412) );
  AOI211_X1 U8143 ( .C1(n6413), .C2(n6412), .A(n9730), .B(n6450), .ZN(n6419)
         );
  INV_X1 U8144 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6417) );
  INV_X1 U8145 ( .A(n6414), .ZN(n6451) );
  NAND2_X1 U8146 ( .A1(n9726), .A2(n6451), .ZN(n6416) );
  NAND2_X1 U8147 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n6415) );
  OAI211_X1 U8148 ( .C1(n6417), .C2(n9746), .A(n6416), .B(n6415), .ZN(n6418)
         );
  OR3_X1 U8149 ( .A1(n6420), .A2(n6419), .A3(n6418), .ZN(P1_U3249) );
  AOI211_X1 U8150 ( .C1(n6423), .C2(n6422), .A(n9718), .B(n6421), .ZN(n6432)
         );
  AOI211_X1 U8151 ( .C1(n6426), .C2(n6425), .A(n9730), .B(n6424), .ZN(n6431)
         );
  INV_X1 U8152 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6429) );
  NAND2_X1 U8153 ( .A1(n9726), .A2(n6427), .ZN(n6428) );
  NAND2_X1 U8154 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n7128) );
  OAI211_X1 U8155 ( .C1(n6429), .C2(n9746), .A(n6428), .B(n7128), .ZN(n6430)
         );
  OR3_X1 U8156 ( .A1(n6432), .A2(n6431), .A3(n6430), .ZN(P1_U3248) );
  INV_X1 U8157 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7500) );
  NAND2_X1 U8158 ( .A1(n9726), .A2(n6433), .ZN(n6435) );
  NAND2_X1 U8159 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n6434) );
  OAI211_X1 U8160 ( .C1(n7500), .C2(n9746), .A(n6435), .B(n6434), .ZN(n6444)
         );
  AOI211_X1 U8161 ( .C1(n6438), .C2(n6437), .A(n6436), .B(n9730), .ZN(n6443)
         );
  AOI211_X1 U8162 ( .C1(n6441), .C2(n6440), .A(n6439), .B(n9718), .ZN(n6442)
         );
  OR3_X1 U8163 ( .A1(n6444), .A2(n6443), .A3(n6442), .ZN(P1_U3246) );
  NAND2_X1 U8164 ( .A1(n5964), .A2(P2_U3893), .ZN(n6445) );
  OAI21_X1 U8165 ( .B1(P2_U3893), .B2(n5102), .A(n6445), .ZN(P2_U3491) );
  INV_X1 U8166 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6446) );
  OAI222_X1 U8167 ( .A1(n8901), .A2(n6460), .B1(n7684), .B2(P2_U3151), .C1(
        n6446), .C2(n8893), .ZN(P2_U3283) );
  AOI21_X1 U8168 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n6451), .A(n6447), .ZN(
        n6449) );
  XOR2_X1 U8169 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6454), .Z(n6448) );
  NOR2_X1 U8170 ( .A1(n6449), .A2(n6448), .ZN(n6564) );
  AOI211_X1 U8171 ( .C1(n6449), .C2(n6448), .A(n9718), .B(n6564), .ZN(n6459)
         );
  XNOR2_X1 U8172 ( .A(n6454), .B(n7183), .ZN(n6452) );
  NOR2_X1 U8173 ( .A1(n6453), .A2(n6452), .ZN(n6567) );
  AOI211_X1 U8174 ( .C1(n6453), .C2(n6452), .A(n9730), .B(n6567), .ZN(n6458)
         );
  INV_X1 U8175 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7515) );
  INV_X1 U8176 ( .A(n6454), .ZN(n6568) );
  NAND2_X1 U8177 ( .A1(n9726), .A2(n6568), .ZN(n6456) );
  NAND2_X1 U8178 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n6455) );
  OAI211_X1 U8179 ( .C1(n7515), .C2(n9746), .A(n6456), .B(n6455), .ZN(n6457)
         );
  OR3_X1 U8180 ( .A1(n6459), .A2(n6458), .A3(n6457), .ZN(P1_U3250) );
  OAI222_X1 U8181 ( .A1(n8213), .A2(n6461), .B1(n9626), .B2(n6460), .C1(n7399), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  NOR2_X1 U8182 ( .A1(n5518), .A2(n9167), .ZN(n6673) );
  INV_X1 U8183 ( .A(n9801), .ZN(n9525) );
  INV_X1 U8184 ( .A(n6462), .ZN(n6626) );
  AOI21_X1 U8185 ( .B1(n9412), .B2(n9525), .A(n6626), .ZN(n6463) );
  AOI211_X1 U8186 ( .C1(n6625), .C2(n7007), .A(n6673), .B(n6463), .ZN(n6518)
         );
  OR2_X1 U8187 ( .A1(n6518), .A2(n9619), .ZN(n6464) );
  OAI21_X1 U8188 ( .B1(n9804), .B2(n5096), .A(n6464), .ZN(P1_U3453) );
  INV_X1 U8189 ( .A(n6776), .ZN(n7751) );
  NOR2_X1 U8190 ( .A1(n6777), .A2(n7751), .ZN(n6465) );
  OR2_X1 U8191 ( .A1(P2_U3150), .A2(n6465), .ZN(n8506) );
  INV_X1 U8192 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6475) );
  INV_X1 U8193 ( .A(n5991), .ZN(n8169) );
  NOR2_X1 U8194 ( .A1(n5991), .A2(P2_U3151), .ZN(n8895) );
  AND2_X1 U8195 ( .A1(n6471), .A2(n8895), .ZN(n6589) );
  INV_X1 U8196 ( .A(n6589), .ZN(n6611) );
  INV_X1 U8197 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6884) );
  INV_X1 U8198 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6466) );
  MUX2_X1 U8199 ( .A(n6884), .B(n6466), .S(n8474), .Z(n6467) );
  NAND2_X1 U8200 ( .A1(n6467), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6637) );
  INV_X1 U8201 ( .A(n6467), .ZN(n6468) );
  NAND2_X1 U8202 ( .A1(n6468), .A2(n4807), .ZN(n6469) );
  AOI22_X1 U8203 ( .A1(n8481), .A2(n6611), .B1(n6637), .B2(n6469), .ZN(n6470)
         );
  AOI21_X1 U8204 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .A(n6470), .ZN(
        n6474) );
  NOR2_X1 U8205 ( .A1(n8474), .A2(P2_U3151), .ZN(n8898) );
  NAND2_X1 U8206 ( .A1(n6471), .A2(n8898), .ZN(n6472) );
  MUX2_X1 U8207 ( .A(n8382), .B(n6472), .S(n5991), .Z(n8503) );
  NAND2_X1 U8208 ( .A1(n8486), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6473) );
  OAI211_X1 U8209 ( .C1(n8506), .C2(n6475), .A(n6474), .B(n6473), .ZN(P2_U3182) );
  INV_X1 U8210 ( .A(n7816), .ZN(n7823) );
  INV_X1 U8211 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6476) );
  OAI222_X1 U8212 ( .A1(n8901), .A2(n6477), .B1(n7823), .B2(P2_U3151), .C1(
        n6476), .C2(n8893), .ZN(P2_U3282) );
  OAI222_X1 U8213 ( .A1(n8213), .A2(n6478), .B1(n9626), .B2(n6477), .C1(n9232), 
        .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U8214 ( .A(n9219), .ZN(n6483) );
  OAI22_X1 U8215 ( .A1(n6483), .A2(n7121), .B1(n9058), .B2(n6487), .ZN(n6527)
         );
  OAI22_X1 U8216 ( .A1(n6487), .A2(n7121), .B1(n6486), .B2(n6521), .ZN(n6488)
         );
  AOI21_X1 U8217 ( .B1(n9219), .B2(n8988), .A(n6488), .ZN(n6528) );
  XNOR2_X1 U8218 ( .A(n6529), .B(n6528), .ZN(n6676) );
  MUX2_X1 U8219 ( .A(n6490), .B(n6676), .S(n6489), .Z(n6493) );
  OAI21_X1 U8220 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n6491), .A(P1_U3973), .ZN(
        n6492) );
  AOI21_X1 U8221 ( .B1(n6493), .B2(n9631), .A(n6492), .ZN(n6516) );
  AOI211_X1 U8222 ( .C1(n6496), .C2(n6495), .A(n9718), .B(n6494), .ZN(n6504)
         );
  AOI211_X1 U8223 ( .C1(n6499), .C2(n6498), .A(n9730), .B(n6497), .ZN(n6503)
         );
  AND2_X1 U8224 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n6706) );
  AOI21_X1 U8225 ( .B1(n9247), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6706), .ZN(
        n6500) );
  OAI21_X1 U8226 ( .B1(n6501), .B2(n9739), .A(n6500), .ZN(n6502) );
  OR4_X1 U8227 ( .A1(n6516), .A2(n6504), .A3(n6503), .A4(n6502), .ZN(P1_U3247)
         );
  AOI211_X1 U8228 ( .C1(n6507), .C2(n6506), .A(n6505), .B(n9730), .ZN(n6515)
         );
  AOI211_X1 U8229 ( .C1(n6510), .C2(n6509), .A(n6508), .B(n9718), .ZN(n6514)
         );
  AOI22_X1 U8230 ( .A1(n9247), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6511) );
  OAI21_X1 U8231 ( .B1(n6512), .B2(n9739), .A(n6511), .ZN(n6513) );
  OR4_X1 U8232 ( .A1(n6516), .A2(n6515), .A3(n6514), .A4(n6513), .ZN(P1_U3245)
         );
  NAND2_X1 U8233 ( .A1(n9812), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6517) );
  OAI21_X1 U8234 ( .B1(n6518), .B2(n9812), .A(n6517), .ZN(P1_U3522) );
  NAND3_X1 U8235 ( .A1(n6520), .A2(n6619), .A3(n6519), .ZN(n6548) );
  NAND2_X1 U8236 ( .A1(n6548), .A2(n6555), .ZN(n6524) );
  AND2_X1 U8237 ( .A1(n6522), .A2(n6521), .ZN(n6523) );
  NAND2_X1 U8238 ( .A1(n6524), .A2(n6523), .ZN(n6526) );
  INV_X1 U8239 ( .A(n6525), .ZN(n7743) );
  INV_X1 U8240 ( .A(n9157), .ZN(n9144) );
  NOR2_X1 U8241 ( .A1(n9144), .A2(P1_U3086), .ZN(n6672) );
  OAI22_X1 U8242 ( .A1(n6529), .A2(n6528), .B1(n8978), .B2(n6527), .ZN(n6678)
         );
  NAND2_X1 U8243 ( .A1(n5104), .A2(n7593), .ZN(n6530) );
  AND2_X1 U8244 ( .A1(n9761), .A2(n7593), .ZN(n6534) );
  AOI21_X1 U8245 ( .B1(n5104), .B2(n8988), .A(n6534), .ZN(n6535) );
  AND2_X1 U8246 ( .A1(n6536), .A2(n6535), .ZN(n6547) );
  XNOR2_X1 U8247 ( .A(n6537), .B(n6687), .ZN(n6540) );
  OR2_X1 U8248 ( .A1(n7017), .A2(n6689), .ZN(n6539) );
  NAND2_X1 U8249 ( .A1(n5477), .A2(n7593), .ZN(n6538) );
  AND2_X1 U8250 ( .A1(n6539), .A2(n6538), .ZN(n6541) );
  NAND2_X1 U8251 ( .A1(n6540), .A2(n6541), .ZN(n6685) );
  INV_X1 U8252 ( .A(n6540), .ZN(n6543) );
  INV_X1 U8253 ( .A(n6541), .ZN(n6542) );
  NAND2_X1 U8254 ( .A1(n6543), .A2(n6542), .ZN(n6544) );
  INV_X1 U8255 ( .A(n6686), .ZN(n6553) );
  NOR3_X1 U8256 ( .A1(n6545), .A2(n6547), .A3(n6546), .ZN(n6552) );
  INV_X1 U8257 ( .A(n6549), .ZN(n6550) );
  NAND2_X1 U8258 ( .A1(n9798), .A2(n6550), .ZN(n6551) );
  OAI21_X1 U8259 ( .B1(n6553), .B2(n6552), .A(n9165), .ZN(n6563) );
  NAND2_X1 U8260 ( .A1(n6625), .A2(n6554), .ZN(n6624) );
  OR2_X1 U8261 ( .A1(n6558), .A2(n6557), .ZN(n9142) );
  OR2_X1 U8262 ( .A1(n6690), .A2(n9167), .ZN(n6561) );
  NAND2_X1 U8263 ( .A1(n6559), .A2(n9138), .ZN(n6560) );
  NAND2_X1 U8264 ( .A1(n6561), .A2(n6560), .ZN(n6923) );
  AOI22_X1 U8265 ( .A1(n5477), .A2(n4264), .B1(n4270), .B2(n6923), .ZN(n6562)
         );
  OAI211_X1 U8266 ( .C1(n6672), .C2(n9930), .A(n6563), .B(n6562), .ZN(P1_U3237) );
  XOR2_X1 U8267 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6569), .Z(n6565) );
  NOR2_X1 U8268 ( .A1(n6566), .A2(n6565), .ZN(n6730) );
  AOI211_X1 U8269 ( .C1(n6566), .C2(n6565), .A(n9718), .B(n6730), .ZN(n6576)
         );
  INV_X1 U8270 ( .A(n6569), .ZN(n6739) );
  XNOR2_X1 U8271 ( .A(n6739), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n6570) );
  AOI211_X1 U8272 ( .C1(n6571), .C2(n6570), .A(n9730), .B(n6738), .ZN(n6575)
         );
  INV_X1 U8273 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n7519) );
  NAND2_X1 U8274 ( .A1(n9726), .A2(n6739), .ZN(n6573) );
  NAND2_X1 U8275 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n6572) );
  OAI211_X1 U8276 ( .C1(n7519), .C2(n9746), .A(n6573), .B(n6572), .ZN(n6574)
         );
  OR3_X1 U8277 ( .A1(n6576), .A2(n6575), .A3(n6574), .ZN(P1_U3251) );
  MUX2_X1 U8278 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8474), .Z(n6577) );
  XNOR2_X1 U8279 ( .A(n6577), .B(n6651), .ZN(n6638) );
  NAND2_X1 U8280 ( .A1(n6638), .A2(n6637), .ZN(n6579) );
  NAND2_X1 U8281 ( .A1(n6577), .A2(n6592), .ZN(n6578) );
  NAND2_X1 U8282 ( .A1(n6579), .A2(n6578), .ZN(n6713) );
  MUX2_X1 U8283 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8474), .Z(n6580) );
  XNOR2_X1 U8284 ( .A(n6580), .B(n6603), .ZN(n6714) );
  NAND2_X1 U8285 ( .A1(n6713), .A2(n6714), .ZN(n6582) );
  NAND2_X1 U8286 ( .A1(n6580), .A2(n6725), .ZN(n6581) );
  NAND2_X1 U8287 ( .A1(n6582), .A2(n6581), .ZN(n6656) );
  MUX2_X1 U8288 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8474), .Z(n6583) );
  XNOR2_X1 U8289 ( .A(n6583), .B(n6605), .ZN(n6657) );
  OR2_X1 U8290 ( .A1(n6656), .A2(n6657), .ZN(n6654) );
  INV_X1 U8291 ( .A(n6583), .ZN(n6584) );
  NAND2_X1 U8292 ( .A1(n6584), .A2(n6668), .ZN(n6585) );
  AND2_X1 U8293 ( .A1(n6654), .A2(n6585), .ZN(n6588) );
  MUX2_X1 U8294 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8474), .Z(n6745) );
  XNOR2_X1 U8295 ( .A(n6745), .B(n6751), .ZN(n6587) );
  AND2_X1 U8296 ( .A1(n6587), .A2(n6585), .ZN(n6586) );
  NAND2_X1 U8297 ( .A1(n6654), .A2(n6586), .ZN(n6747) );
  OAI211_X1 U8298 ( .C1(n6588), .C2(n6587), .A(n8509), .B(n6747), .ZN(n6616)
         );
  INV_X1 U8299 ( .A(n8516), .ZN(n6916) );
  INV_X1 U8300 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9879) );
  MUX2_X1 U8301 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9879), .S(n6751), .Z(n6596)
         );
  INV_X1 U8302 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9877) );
  MUX2_X1 U8303 ( .A(n9877), .B(P2_REG1_REG_2__SCAN_IN), .S(n6603), .Z(n6717)
         );
  NAND2_X1 U8304 ( .A1(n5677), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6591) );
  INV_X1 U8305 ( .A(n5677), .ZN(n6593) );
  AND2_X1 U8306 ( .A1(n4807), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6590) );
  INV_X1 U8307 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6645) );
  NAND2_X1 U8308 ( .A1(n6717), .A2(n6716), .ZN(n6715) );
  OAI21_X1 U8309 ( .B1(n6603), .B2(n9877), .A(n6715), .ZN(n6594) );
  XNOR2_X1 U8310 ( .A(n6594), .B(n6668), .ZN(n6658) );
  AOI21_X1 U8311 ( .B1(n6596), .B2(n6595), .A(n6748), .ZN(n6597) );
  OAI22_X1 U8312 ( .A1(n6916), .A2(n6597), .B1(n7507), .B2(n8506), .ZN(n6614)
         );
  INV_X1 U8313 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6598) );
  NOR2_X1 U8314 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6598), .ZN(n7065) );
  INV_X1 U8315 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6599) );
  NAND2_X1 U8316 ( .A1(n4807), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6600) );
  NAND2_X1 U8317 ( .A1(n6651), .A2(n6600), .ZN(n6601) );
  NAND2_X1 U8318 ( .A1(n5677), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6602) );
  NAND2_X1 U8319 ( .A1(n6601), .A2(n6602), .ZN(n6641) );
  INV_X1 U8320 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6642) );
  OR2_X1 U8321 ( .A1(n6641), .A2(n6642), .ZN(n6639) );
  NAND2_X1 U8322 ( .A1(n6639), .A2(n6602), .ZN(n6720) );
  NAND2_X1 U8323 ( .A1(n6721), .A2(n6720), .ZN(n6719) );
  OR2_X1 U8324 ( .A1(n6603), .A2(n6599), .ZN(n6604) );
  NAND2_X1 U8325 ( .A1(n6719), .A2(n6604), .ZN(n6606) );
  INV_X1 U8326 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6663) );
  XNOR2_X1 U8327 ( .A(n6751), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n6608) );
  NAND2_X1 U8328 ( .A1(n6607), .A2(n6608), .ZN(n6753) );
  INV_X1 U8329 ( .A(n6608), .ZN(n6610) );
  NAND3_X1 U8330 ( .A1(n6660), .A2(n6610), .A3(n6609), .ZN(n6612) );
  AOI21_X1 U8331 ( .B1(n6753), .B2(n6612), .A(n8519), .ZN(n6613) );
  NOR3_X1 U8332 ( .A1(n6614), .A2(n7065), .A3(n6613), .ZN(n6615) );
  OAI211_X1 U8333 ( .C1(n8503), .C2(n6749), .A(n6616), .B(n6615), .ZN(P2_U3186) );
  NAND2_X1 U8334 ( .A1(n9218), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6617) );
  OAI21_X1 U8335 ( .B1(n9065), .B2(n9218), .A(n6617), .ZN(P1_U3583) );
  INV_X1 U8336 ( .A(n6618), .ZN(n6620) );
  NAND3_X1 U8337 ( .A1(n6621), .A2(n6620), .A3(n6619), .ZN(n6622) );
  NOR2_X1 U8338 ( .A1(n9765), .A2(n9443), .ZN(n9397) );
  OAI21_X1 U8339 ( .B1(n9397), .B2(n9762), .A(n7007), .ZN(n6635) );
  NOR2_X1 U8340 ( .A1(n6626), .A2(n6625), .ZN(n6628) );
  INV_X1 U8341 ( .A(n6628), .ZN(n6631) );
  NAND2_X1 U8342 ( .A1(n6628), .A2(n6627), .ZN(n6630) );
  INV_X1 U8343 ( .A(n9471), .ZN(n9758) );
  AOI21_X1 U8344 ( .B1(n9758), .B2(P1_REG3_REG_0__SCAN_IN), .A(n6673), .ZN(
        n6629) );
  OAI211_X1 U8345 ( .C1(n6632), .C2(n6631), .A(n6630), .B(n6629), .ZN(n6633)
         );
  NAND2_X1 U8346 ( .A1(n6633), .A2(n9474), .ZN(n6634) );
  OAI211_X1 U8347 ( .C1(n6636), .C2(n9474), .A(n6635), .B(n6634), .ZN(P1_U3293) );
  XNOR2_X1 U8348 ( .A(n6638), .B(n6637), .ZN(n6653) );
  INV_X1 U8349 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6644) );
  INV_X1 U8350 ( .A(n6639), .ZN(n6640) );
  AOI21_X1 U8351 ( .B1(n6642), .B2(n6641), .A(n6640), .ZN(n6643) );
  OAI22_X1 U8352 ( .A1(n8506), .A2(n6644), .B1(n8519), .B2(n6643), .ZN(n6650)
         );
  INV_X1 U8353 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6648) );
  NAND2_X1 U8354 ( .A1(n8516), .A2(n6646), .ZN(n6647) );
  OAI21_X1 U8355 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n6648), .A(n6647), .ZN(n6649) );
  AOI211_X1 U8356 ( .C1(n6651), .C2(n8486), .A(n6650), .B(n6649), .ZN(n6652)
         );
  OAI21_X1 U8357 ( .B1(n8481), .B2(n6653), .A(n6652), .ZN(P2_U3183) );
  INV_X1 U8358 ( .A(n6654), .ZN(n6655) );
  AOI21_X1 U8359 ( .B1(n6657), .B2(n6656), .A(n6655), .ZN(n6671) );
  XNOR2_X1 U8360 ( .A(n6658), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n6667) );
  NOR2_X1 U8361 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6659), .ZN(n6960) );
  INV_X1 U8362 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6665) );
  INV_X1 U8363 ( .A(n6660), .ZN(n6661) );
  AOI21_X1 U8364 ( .B1(n6663), .B2(n6662), .A(n6661), .ZN(n6664) );
  OAI22_X1 U8365 ( .A1(n8506), .A2(n6665), .B1(n8519), .B2(n6664), .ZN(n6666)
         );
  AOI211_X1 U8366 ( .C1(n8516), .C2(n6667), .A(n6960), .B(n6666), .ZN(n6670)
         );
  NAND2_X1 U8367 ( .A1(n8486), .A2(n6668), .ZN(n6669) );
  OAI211_X1 U8368 ( .C1(n6671), .C2(n8481), .A(n6670), .B(n6669), .ZN(P2_U3185) );
  INV_X1 U8369 ( .A(n6672), .ZN(n6681) );
  NAND2_X1 U8370 ( .A1(n6681), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6675) );
  AOI22_X1 U8371 ( .A1(n7007), .A2(n4264), .B1(n4270), .B2(n6673), .ZN(n6674)
         );
  OAI211_X1 U8372 ( .C1(n6676), .C2(n9189), .A(n6675), .B(n6674), .ZN(P1_U3232) );
  AOI21_X1 U8373 ( .B1(n6678), .B2(n6677), .A(n6545), .ZN(n6684) );
  OR2_X1 U8374 ( .A1(n7017), .A2(n9167), .ZN(n6680) );
  NAND2_X1 U8375 ( .A1(n9219), .A2(n9138), .ZN(n6679) );
  NAND2_X1 U8376 ( .A1(n6680), .A2(n6679), .ZN(n7006) );
  AOI22_X1 U8377 ( .A1(n9761), .A2(n4264), .B1(n4270), .B2(n7006), .ZN(n6683)
         );
  NAND2_X1 U8378 ( .A1(n6681), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6682) );
  OAI211_X1 U8379 ( .C1(n6684), .C2(n9189), .A(n6683), .B(n6682), .ZN(P1_U3222) );
  XNOR2_X1 U8380 ( .A(n6688), .B(n8978), .ZN(n6695) );
  OR2_X1 U8381 ( .A1(n6690), .A2(n6689), .ZN(n6692) );
  NAND2_X1 U8382 ( .A1(n9747), .A2(n7593), .ZN(n6691) );
  NAND2_X1 U8383 ( .A1(n6692), .A2(n6691), .ZN(n6693) );
  XNOR2_X1 U8384 ( .A(n6695), .B(n6693), .ZN(n9042) );
  INV_X1 U8385 ( .A(n6693), .ZN(n6694) );
  NAND2_X1 U8386 ( .A1(n6695), .A2(n6694), .ZN(n6698) );
  AND2_X1 U8387 ( .A1(n6700), .A2(n6698), .ZN(n6702) );
  NAND2_X1 U8388 ( .A1(n9215), .A2(n7593), .ZN(n6696) );
  OAI21_X1 U8389 ( .B1(n7092), .B2(n9058), .A(n6696), .ZN(n6697) );
  XNOR2_X1 U8390 ( .A(n6697), .B(n8978), .ZN(n7116) );
  AOI22_X1 U8391 ( .A1(n6994), .A2(n7593), .B1(n9215), .B2(n8988), .ZN(n7117)
         );
  XNOR2_X1 U8392 ( .A(n7116), .B(n7117), .ZN(n6701) );
  NAND2_X1 U8393 ( .A1(n6700), .A2(n6699), .ZN(n7120) );
  OAI211_X1 U8394 ( .C1(n6702), .C2(n6701), .A(n9165), .B(n7120), .ZN(n6708)
         );
  OR2_X1 U8395 ( .A1(n7196), .A2(n9167), .ZN(n6704) );
  OR2_X1 U8396 ( .A1(n6690), .A2(n9169), .ZN(n6703) );
  NAND2_X1 U8397 ( .A1(n6704), .A2(n6703), .ZN(n6984) );
  INV_X1 U8398 ( .A(n4264), .ZN(n9147) );
  NOR2_X1 U8399 ( .A1(n9147), .A2(n7092), .ZN(n6705) );
  AOI211_X1 U8400 ( .C1(n4270), .C2(n6984), .A(n6706), .B(n6705), .ZN(n6707)
         );
  OAI211_X1 U8401 ( .C1(n9157), .C2(n6991), .A(n6708), .B(n6707), .ZN(P1_U3230) );
  INV_X1 U8402 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6710) );
  INV_X1 U8403 ( .A(n6709), .ZN(n6712) );
  OAI222_X1 U8404 ( .A1(n8893), .A2(n6710), .B1(n8891), .B2(n6712), .C1(
        P2_U3151), .C2(n8385), .ZN(P2_U3281) );
  OAI222_X1 U8405 ( .A1(n8213), .A2(n10034), .B1(n9626), .B2(n6712), .C1(
        P1_U3086), .C2(n6711), .ZN(P1_U3341) );
  XOR2_X1 U8406 ( .A(n6714), .B(n6713), .Z(n6727) );
  INV_X1 U8407 ( .A(n8506), .ZN(n7838) );
  OAI21_X1 U8408 ( .B1(n6717), .B2(n6716), .A(n6715), .ZN(n6718) );
  AOI22_X1 U8409 ( .A1(n7838), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(n8516), .B2(
        n6718), .ZN(n6724) );
  INV_X1 U8410 ( .A(n8519), .ZN(n6759) );
  OAI21_X1 U8411 ( .B1(n6721), .B2(n6720), .A(n6719), .ZN(n6722) );
  AOI22_X1 U8412 ( .A1(n6759), .A2(n6722), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3151), .ZN(n6723) );
  OAI211_X1 U8413 ( .C1(n6725), .C2(n8503), .A(n6724), .B(n6723), .ZN(n6726)
         );
  AOI21_X1 U8414 ( .B1(n8509), .B2(n6727), .A(n6726), .ZN(n6728) );
  INV_X1 U8415 ( .A(n6728), .ZN(P2_U3184) );
  NOR2_X1 U8416 ( .A1(n7392), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6729) );
  AOI21_X1 U8417 ( .B1(n7392), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6729), .ZN(
        n6732) );
  NAND2_X1 U8418 ( .A1(n6731), .A2(n6732), .ZN(n7391) );
  OAI21_X1 U8419 ( .B1(n6732), .B2(n6731), .A(n7391), .ZN(n6736) );
  INV_X1 U8420 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6734) );
  NAND2_X1 U8421 ( .A1(n9726), .A2(n7392), .ZN(n6733) );
  NAND2_X1 U8422 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7561) );
  OAI211_X1 U8423 ( .C1(n9746), .C2(n6734), .A(n6733), .B(n7561), .ZN(n6735)
         );
  AOI21_X1 U8424 ( .B1(n6736), .B2(n9733), .A(n6735), .ZN(n6744) );
  NOR2_X1 U8425 ( .A1(n7392), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6737) );
  AOI21_X1 U8426 ( .B1(n7392), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6737), .ZN(
        n6741) );
  OAI21_X1 U8427 ( .B1(n6741), .B2(n6740), .A(n7386), .ZN(n6742) );
  INV_X1 U8428 ( .A(n9730), .ZN(n9682) );
  NAND2_X1 U8429 ( .A1(n6742), .A2(n9682), .ZN(n6743) );
  NAND2_X1 U8430 ( .A1(n6744), .A2(n6743), .ZN(P1_U3252) );
  NAND2_X1 U8431 ( .A1(n6745), .A2(n6749), .ZN(n6746) );
  NAND2_X1 U8432 ( .A1(n6747), .A2(n6746), .ZN(n6806) );
  MUX2_X1 U8433 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8474), .Z(n6801) );
  XNOR2_X1 U8434 ( .A(n6801), .B(n6802), .ZN(n6805) );
  XNOR2_X1 U8435 ( .A(n6806), .B(n6805), .ZN(n6765) );
  XOR2_X1 U8436 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6793), .Z(n6763) );
  INV_X1 U8437 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9991) );
  NAND2_X1 U8438 ( .A1(n8486), .A2(n6802), .ZN(n6761) );
  INV_X1 U8439 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6750) );
  OR2_X1 U8440 ( .A1(n6751), .A2(n6750), .ZN(n6752) );
  NAND2_X1 U8441 ( .A1(n6753), .A2(n6752), .ZN(n6755) );
  OAI21_X1 U8442 ( .B1(n6755), .B2(n6754), .A(n6830), .ZN(n6756) );
  INV_X1 U8443 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7257) );
  NAND2_X1 U8444 ( .A1(n6756), .A2(n7257), .ZN(n6757) );
  NAND2_X1 U8445 ( .A1(n6832), .A2(n6757), .ZN(n6758) );
  AND2_X1 U8446 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7290) );
  AOI21_X1 U8447 ( .B1(n6759), .B2(n6758), .A(n7290), .ZN(n6760) );
  OAI211_X1 U8448 ( .C1(n9991), .C2(n8506), .A(n6761), .B(n6760), .ZN(n6762)
         );
  AOI21_X1 U8449 ( .B1(n6763), .B2(n8516), .A(n6762), .ZN(n6764) );
  OAI21_X1 U8450 ( .B1(n6765), .B2(n8481), .A(n6764), .ZN(P2_U3187) );
  NOR2_X1 U8451 ( .A1(n6768), .A2(n6783), .ZN(n6859) );
  OR2_X1 U8452 ( .A1(n6771), .A2(n6767), .ZN(n6770) );
  OR2_X1 U8453 ( .A1(n6768), .A2(n6781), .ZN(n6769) );
  INV_X1 U8454 ( .A(n7977), .ZN(n6935) );
  NAND2_X1 U8455 ( .A1(n5964), .A2(n6886), .ZN(n7982) );
  NAND2_X1 U8456 ( .A1(n6935), .A2(n7982), .ZN(n6879) );
  OR2_X1 U8457 ( .A1(n6771), .A2(n9842), .ZN(n6773) );
  AOI22_X1 U8458 ( .A1(n8336), .A2(n6879), .B1(n9818), .B2(n8352), .ZN(n6790)
         );
  OR2_X1 U8459 ( .A1(n6775), .A2(n6774), .ZN(n6780) );
  AND3_X1 U8460 ( .A1(n6778), .A2(n6777), .A3(n6776), .ZN(n6779) );
  OAI211_X1 U8461 ( .C1(n6786), .C2(n6781), .A(n6780), .B(n6779), .ZN(n6782)
         );
  NAND2_X1 U8462 ( .A1(n6782), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6788) );
  NOR2_X1 U8463 ( .A1(n6784), .A2(n6783), .ZN(n8170) );
  INV_X1 U8464 ( .A(n8170), .ZN(n6785) );
  OR2_X1 U8465 ( .A1(n6786), .A2(n6785), .ZN(n6787) );
  INV_X1 U8466 ( .A(n8365), .ZN(n7372) );
  NAND2_X1 U8467 ( .A1(n7372), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6869) );
  NAND2_X1 U8468 ( .A1(n6869), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6789) );
  OAI211_X1 U8469 ( .C1(n7242), .C2(n8363), .A(n6790), .B(n6789), .ZN(P2_U3172) );
  INV_X1 U8470 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10048) );
  INV_X1 U8471 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6792) );
  OAI22_X1 U8472 ( .A1(n6793), .A2(n6792), .B1(n6802), .B2(n6791), .ZN(n6836)
         );
  MUX2_X1 U8473 ( .A(n10048), .B(P2_REG1_REG_6__SCAN_IN), .S(n6808), .Z(n6837)
         );
  NAND2_X1 U8474 ( .A1(n6836), .A2(n6837), .ZN(n6835) );
  OAI21_X1 U8475 ( .B1(n6808), .B2(n10048), .A(n6835), .ZN(n6887) );
  XNOR2_X1 U8476 ( .A(n6887), .B(n6813), .ZN(n6888) );
  INV_X1 U8477 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6812) );
  XNOR2_X1 U8478 ( .A(n6888), .B(n6812), .ZN(n6825) );
  INV_X1 U8479 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6795) );
  AND2_X1 U8480 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8221) );
  INV_X1 U8481 ( .A(n8221), .ZN(n6794) );
  OAI21_X1 U8482 ( .B1(n8506), .B2(n6795), .A(n6794), .ZN(n6800) );
  INV_X1 U8483 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6807) );
  MUX2_X1 U8484 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6807), .S(n6808), .Z(n6831)
         );
  AOI21_X1 U8485 ( .B1(n4317), .B2(n6813), .A(n6893), .ZN(n6797) );
  INV_X1 U8486 ( .A(n6797), .ZN(n6796) );
  INV_X1 U8487 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7472) );
  NAND2_X1 U8488 ( .A1(n6796), .A2(n7472), .ZN(n6798) );
  AOI21_X1 U8489 ( .B1(n6798), .B2(n6896), .A(n8519), .ZN(n6799) );
  AOI211_X1 U8490 ( .C1(n8486), .C2(n6813), .A(n6800), .B(n6799), .ZN(n6824)
         );
  INV_X1 U8491 ( .A(n6801), .ZN(n6803) );
  NOR2_X1 U8492 ( .A1(n6803), .A2(n6802), .ZN(n6804) );
  AOI21_X1 U8493 ( .B1(n6806), .B2(n6805), .A(n6804), .ZN(n6828) );
  MUX2_X1 U8494 ( .A(n6807), .B(n10048), .S(n8474), .Z(n6809) );
  NAND2_X1 U8495 ( .A1(n6809), .A2(n6808), .ZN(n6819) );
  INV_X1 U8496 ( .A(n6809), .ZN(n6810) );
  NAND2_X1 U8497 ( .A1(n6810), .A2(n6841), .ZN(n6811) );
  AND2_X1 U8498 ( .A1(n6819), .A2(n6811), .ZN(n6827) );
  NAND2_X1 U8499 ( .A1(n6828), .A2(n6827), .ZN(n6826) );
  INV_X1 U8500 ( .A(n6826), .ZN(n6818) );
  INV_X1 U8501 ( .A(n6819), .ZN(n6817) );
  MUX2_X1 U8502 ( .A(n7472), .B(n6812), .S(n8474), .Z(n6814) );
  NAND2_X1 U8503 ( .A1(n6814), .A2(n6813), .ZN(n6908) );
  INV_X1 U8504 ( .A(n6814), .ZN(n6815) );
  NAND2_X1 U8505 ( .A1(n6815), .A2(n4703), .ZN(n6816) );
  AND2_X1 U8506 ( .A1(n6908), .A2(n6816), .ZN(n6820) );
  NOR3_X1 U8507 ( .A1(n6818), .A2(n6817), .A3(n6820), .ZN(n6822) );
  NAND2_X1 U8508 ( .A1(n6826), .A2(n6819), .ZN(n6821) );
  NAND2_X1 U8509 ( .A1(n6821), .A2(n6820), .ZN(n6909) );
  INV_X1 U8510 ( .A(n6909), .ZN(n6907) );
  OAI21_X1 U8511 ( .B1(n6822), .B2(n6907), .A(n8509), .ZN(n6823) );
  OAI211_X1 U8512 ( .C1(n6825), .C2(n6916), .A(n6824), .B(n6823), .ZN(P2_U3189) );
  OAI21_X1 U8513 ( .B1(n6828), .B2(n6827), .A(n6826), .ZN(n6843) );
  INV_X1 U8514 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6829) );
  NOR2_X1 U8515 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6829), .ZN(n7369) );
  NAND3_X1 U8516 ( .A1(n6832), .A2(n6831), .A3(n6830), .ZN(n6833) );
  AOI21_X1 U8517 ( .B1(n4360), .B2(n6833), .A(n8519), .ZN(n6834) );
  AOI211_X1 U8518 ( .C1(n7838), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n7369), .B(
        n6834), .ZN(n6840) );
  OAI21_X1 U8519 ( .B1(n6837), .B2(n6836), .A(n6835), .ZN(n6838) );
  NAND2_X1 U8520 ( .A1(n6838), .A2(n8516), .ZN(n6839) );
  OAI211_X1 U8521 ( .C1(n8503), .C2(n6841), .A(n6840), .B(n6839), .ZN(n6842)
         );
  AOI21_X1 U8522 ( .B1(n6843), .B2(n8509), .A(n6842), .ZN(n6844) );
  INV_X1 U8523 ( .A(n6844), .ZN(P2_U3188) );
  INV_X1 U8524 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6846) );
  INV_X1 U8525 ( .A(n6845), .ZN(n6847) );
  INV_X1 U8526 ( .A(n8409), .ZN(n8416) );
  OAI222_X1 U8527 ( .A1(n8893), .A2(n6846), .B1(n8891), .B2(n6847), .C1(
        P2_U3151), .C2(n8416), .ZN(P2_U3280) );
  OAI222_X1 U8528 ( .A1(n8213), .A2(n9925), .B1(n9626), .B2(n6847), .C1(
        P1_U3086), .C2(n9717), .ZN(P1_U3340) );
  INV_X1 U8529 ( .A(n6848), .ZN(n6849) );
  NAND2_X1 U8530 ( .A1(n6945), .A2(n7499), .ZN(n6851) );
  AOI21_X1 U8531 ( .B1(n8202), .B2(n6886), .A(n6855), .ZN(n6865) );
  XNOR2_X1 U8532 ( .A(n6952), .B(n6958), .ZN(n6954) );
  XOR2_X1 U8533 ( .A(n6955), .B(n6954), .Z(n6864) );
  NAND2_X1 U8534 ( .A1(n6859), .A2(n6858), .ZN(n8341) );
  INV_X1 U8535 ( .A(n6860), .ZN(n7238) );
  AOI22_X1 U8536 ( .A1(n8361), .A2(n8383), .B1(n7238), .B2(n8352), .ZN(n6861)
         );
  OAI21_X1 U8537 ( .B1(n7241), .B2(n8363), .A(n6861), .ZN(n6862) );
  AOI21_X1 U8538 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n6869), .A(n6862), .ZN(
        n6863) );
  OAI21_X1 U8539 ( .B1(n6864), .B2(n8356), .A(n6863), .ZN(P2_U3177) );
  XOR2_X1 U8540 ( .A(n6866), .B(n6865), .Z(n6871) );
  INV_X1 U8541 ( .A(n6941), .ZN(n6948) );
  AOI22_X1 U8542 ( .A1(n8361), .A2(n5964), .B1(n6948), .B2(n8352), .ZN(n6867)
         );
  OAI21_X1 U8543 ( .B1(n6958), .B2(n8363), .A(n6867), .ZN(n6868) );
  AOI21_X1 U8544 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n6869), .A(n6868), .ZN(
        n6870) );
  OAI21_X1 U8545 ( .B1(n8356), .B2(n6871), .A(n6870), .ZN(P2_U3162) );
  OR2_X1 U8546 ( .A1(n6872), .A2(n8881), .ZN(n6873) );
  OAI21_X1 U8547 ( .B1(n6850), .B2(n6874), .A(n6873), .ZN(n6875) );
  INV_X1 U8548 ( .A(n6875), .ZN(n6876) );
  NAND2_X1 U8549 ( .A1(n6877), .A2(n6876), .ZN(n6882) );
  INV_X1 U8550 ( .A(n6882), .ZN(n6878) );
  INV_X1 U8551 ( .A(n8714), .ZN(n8583) );
  NAND2_X1 U8552 ( .A1(n6878), .A2(n8583), .ZN(n8561) );
  NOR2_X1 U8553 ( .A1(n7242), .A2(n9663), .ZN(n9817) );
  INV_X1 U8554 ( .A(n6879), .ZN(n9814) );
  NOR2_X1 U8555 ( .A1(n9814), .A2(n6880), .ZN(n6881) );
  AOI211_X1 U8556 ( .C1(n8731), .C2(P2_REG3_REG_0__SCAN_IN), .A(n9817), .B(
        n6881), .ZN(n6883) );
  MUX2_X1 U8557 ( .A(n6884), .B(n6883), .S(n9668), .Z(n6885) );
  OAI21_X1 U8558 ( .B1(n8561), .B2(n6886), .A(n6885), .ZN(P2_U3233) );
  INV_X1 U8559 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9884) );
  MUX2_X1 U8560 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9884), .S(n6902), .Z(n6890)
         );
  AOI22_X1 U8561 ( .A1(n6888), .A2(P2_REG1_REG_7__SCAN_IN), .B1(n4703), .B2(
        n6887), .ZN(n6889) );
  AOI21_X1 U8562 ( .B1(n6890), .B2(n6889), .A(n7038), .ZN(n6917) );
  INV_X1 U8563 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7518) );
  NOR2_X1 U8564 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6891), .ZN(n7571) );
  INV_X1 U8565 ( .A(n7571), .ZN(n6892) );
  OAI21_X1 U8566 ( .B1(n8506), .B2(n7518), .A(n6892), .ZN(n6900) );
  INV_X1 U8567 ( .A(n6893), .ZN(n6894) );
  INV_X1 U8568 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6901) );
  XNOR2_X1 U8569 ( .A(n6902), .B(n6901), .ZN(n6895) );
  AOI21_X1 U8570 ( .B1(n6896), .B2(n6894), .A(n6895), .ZN(n7040) );
  INV_X1 U8571 ( .A(n7040), .ZN(n6898) );
  NAND3_X1 U8572 ( .A1(n6896), .A2(n6895), .A3(n6894), .ZN(n6897) );
  AOI21_X1 U8573 ( .B1(n6898), .B2(n6897), .A(n8519), .ZN(n6899) );
  AOI211_X1 U8574 ( .C1(n8486), .C2(n6902), .A(n6900), .B(n6899), .ZN(n6915)
         );
  INV_X1 U8575 ( .A(n6908), .ZN(n6906) );
  MUX2_X1 U8576 ( .A(n6901), .B(n9884), .S(n8474), .Z(n6903) );
  NAND2_X1 U8577 ( .A1(n6903), .A2(n6902), .ZN(n7033) );
  INV_X1 U8578 ( .A(n6903), .ZN(n6904) );
  NAND2_X1 U8579 ( .A1(n6904), .A2(n7041), .ZN(n6905) );
  AND2_X1 U8580 ( .A1(n7033), .A2(n6905), .ZN(n6910) );
  NOR3_X1 U8581 ( .A1(n6907), .A2(n6906), .A3(n6910), .ZN(n6913) );
  NAND2_X1 U8582 ( .A1(n6909), .A2(n6908), .ZN(n6911) );
  NAND2_X1 U8583 ( .A1(n6911), .A2(n6910), .ZN(n7036) );
  INV_X1 U8584 ( .A(n7036), .ZN(n6912) );
  OAI21_X1 U8585 ( .B1(n6913), .B2(n6912), .A(n8509), .ZN(n6914) );
  OAI211_X1 U8586 ( .C1(n6917), .C2(n6916), .A(n6915), .B(n6914), .ZN(P2_U3190) );
  XNOR2_X1 U8587 ( .A(n6919), .B(n6918), .ZN(n6925) );
  OAI21_X1 U8588 ( .B1(n6922), .B2(n6921), .A(n6920), .ZN(n9778) );
  INV_X1 U8589 ( .A(n7647), .ZN(n7181) );
  AOI21_X1 U8590 ( .B1(n9778), .B2(n7181), .A(n6923), .ZN(n6924) );
  OAI21_X1 U8591 ( .B1(n9412), .B2(n6925), .A(n6924), .ZN(n9776) );
  INV_X1 U8592 ( .A(n9778), .ZN(n6926) );
  OAI22_X1 U8593 ( .A1(n6926), .A2(n6989), .B1(n9930), .B2(n9471), .ZN(n6927)
         );
  OAI21_X1 U8594 ( .B1(n9776), .B2(n6927), .A(n9474), .ZN(n6931) );
  AOI21_X1 U8595 ( .B1(n7008), .B2(n5477), .A(n9443), .ZN(n6928) );
  INV_X1 U8596 ( .A(n6928), .ZN(n6929) );
  NOR2_X1 U8597 ( .A1(n6929), .A2(n7022), .ZN(n9773) );
  AOI22_X1 U8598 ( .A1(n9450), .A2(n9773), .B1(P1_REG2_REG_2__SCAN_IN), .B2(
        n9749), .ZN(n6930) );
  OAI211_X1 U8599 ( .C1(n9775), .C2(n9444), .A(n6931), .B(n6930), .ZN(P1_U3291) );
  INV_X1 U8600 ( .A(n6933), .ZN(n6934) );
  AOI21_X1 U8601 ( .B1(n6935), .B2(n6932), .A(n6934), .ZN(n6951) );
  INV_X1 U8602 ( .A(n9835), .ZN(n9867) );
  XNOR2_X1 U8603 ( .A(n6932), .B(n6936), .ZN(n6937) );
  AOI222_X1 U8604 ( .A1(n8719), .A2(n6937), .B1(n8381), .B2(n8726), .C1(n5964), 
        .C2(n8723), .ZN(n6947) );
  OAI21_X1 U8605 ( .B1(n6951), .B2(n9867), .A(n6947), .ZN(n6943) );
  OAI22_X1 U8606 ( .A1(n8785), .A2(n6941), .B1(n9890), .B2(n6645), .ZN(n6938)
         );
  AOI21_X1 U8607 ( .B1(n6943), .B2(n9890), .A(n6938), .ZN(n6939) );
  INV_X1 U8608 ( .A(n6939), .ZN(P2_U3460) );
  INV_X1 U8609 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6940) );
  OAI22_X1 U8610 ( .A1(n8863), .A2(n6941), .B1(n6940), .B2(n9873), .ZN(n6942)
         );
  AOI21_X1 U8611 ( .B1(n6943), .B2(n9873), .A(n6942), .ZN(n6944) );
  INV_X1 U8612 ( .A(n6944), .ZN(P2_U3393) );
  INV_X1 U8613 ( .A(n6945), .ZN(n8125) );
  NOR2_X1 U8614 ( .A1(n7239), .A2(n8125), .ZN(n7237) );
  INV_X1 U8615 ( .A(n7237), .ZN(n6946) );
  NAND2_X1 U8616 ( .A1(n7612), .A2(n6946), .ZN(n9667) );
  MUX2_X1 U8617 ( .A(n6642), .B(n6947), .S(n9668), .Z(n6950) );
  AOI22_X1 U8618 ( .A1(n8710), .A2(n6948), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8731), .ZN(n6949) );
  OAI211_X1 U8619 ( .C1(n6951), .C2(n8713), .A(n6950), .B(n6949), .ZN(P2_U3232) );
  INV_X1 U8620 ( .A(n6952), .ZN(n6953) );
  XNOR2_X1 U8621 ( .A(n7059), .B(n7241), .ZN(n6956) );
  OAI211_X1 U8622 ( .C1(n6957), .C2(n6956), .A(n7061), .B(n8336), .ZN(n6963)
         );
  INV_X1 U8623 ( .A(n7228), .ZN(n6961) );
  INV_X1 U8624 ( .A(n8379), .ZN(n7288) );
  OAI22_X1 U8625 ( .A1(n7288), .A2(n8363), .B1(n8341), .B2(n6958), .ZN(n6959)
         );
  AOI211_X1 U8626 ( .C1(n6961), .C2(n8352), .A(n6960), .B(n6959), .ZN(n6962)
         );
  OAI211_X1 U8627 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n7372), .A(n6963), .B(
        n6962), .ZN(P2_U3158) );
  INV_X1 U8628 ( .A(n6964), .ZN(n6966) );
  INV_X1 U8629 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6965) );
  OAI222_X1 U8630 ( .A1(n8901), .A2(n6966), .B1(n8443), .B2(P2_U3151), .C1(
        n6965), .C2(n8893), .ZN(P2_U3279) );
  OAI222_X1 U8631 ( .A1(n8213), .A2(n6967), .B1(n9626), .B2(n6966), .C1(n9228), 
        .C2(P1_U3086), .ZN(P1_U3339) );
  OAI21_X1 U8632 ( .B1(n6970), .B2(n6969), .A(n6968), .ZN(n7232) );
  XNOR2_X1 U8633 ( .A(n6971), .B(n8131), .ZN(n6972) );
  NAND2_X1 U8634 ( .A1(n6972), .A2(n8719), .ZN(n6974) );
  AOI22_X1 U8635 ( .A1(n8726), .A2(n8379), .B1(n8381), .B2(n8723), .ZN(n6973)
         );
  NAND2_X1 U8636 ( .A1(n6974), .A2(n6973), .ZN(n7229) );
  AOI21_X1 U8637 ( .B1(n9835), .B2(n7232), .A(n7229), .ZN(n6981) );
  INV_X1 U8638 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6975) );
  OAI22_X1 U8639 ( .A1(n8863), .A2(n7228), .B1(n6975), .B2(n9873), .ZN(n6976)
         );
  INV_X1 U8640 ( .A(n6976), .ZN(n6977) );
  OAI21_X1 U8641 ( .B1(n6981), .B2(n9875), .A(n6977), .ZN(P2_U3399) );
  INV_X1 U8642 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6978) );
  OAI22_X1 U8643 ( .A1(n8785), .A2(n7228), .B1(n9890), .B2(n6978), .ZN(n6979)
         );
  INV_X1 U8644 ( .A(n6979), .ZN(n6980) );
  OAI21_X1 U8645 ( .B1(n6981), .B2(n8746), .A(n6980), .ZN(P2_U3462) );
  XNOR2_X1 U8646 ( .A(n6983), .B(n6982), .ZN(n6985) );
  AOI21_X1 U8647 ( .B1(n6985), .B2(n9463), .A(n6984), .ZN(n7084) );
  OAI21_X1 U8648 ( .B1(n6988), .B2(n6987), .A(n6986), .ZN(n7094) );
  OR2_X1 U8649 ( .A1(n9405), .A2(n7647), .ZN(n6990) );
  OAI211_X1 U8650 ( .C1(n7020), .C2(n7092), .A(n9521), .B(n7077), .ZN(n7083)
         );
  OAI22_X1 U8651 ( .A1(n9474), .A2(n6992), .B1(n6991), .B2(n9471), .ZN(n6993)
         );
  AOI21_X1 U8652 ( .B1(n9762), .B2(n6994), .A(n6993), .ZN(n6995) );
  OAI21_X1 U8653 ( .B1(n9765), .B2(n7083), .A(n6995), .ZN(n6996) );
  AOI21_X1 U8654 ( .B1(n7094), .B2(n9754), .A(n6996), .ZN(n6997) );
  OAI21_X1 U8655 ( .B1(n9405), .B2(n7084), .A(n6997), .ZN(P1_U3289) );
  INV_X1 U8656 ( .A(n6998), .ZN(n6999) );
  NAND2_X1 U8657 ( .A1(n7003), .A2(n6999), .ZN(n7000) );
  NAND2_X1 U8658 ( .A1(n7001), .A2(n7000), .ZN(n9759) );
  INV_X1 U8659 ( .A(n9759), .ZN(n7010) );
  XNOR2_X1 U8660 ( .A(n7003), .B(n7002), .ZN(n7004) );
  NOR2_X1 U8661 ( .A1(n7004), .A2(n9412), .ZN(n7005) );
  AOI211_X1 U8662 ( .C1(n7181), .C2(n9759), .A(n7006), .B(n7005), .ZN(n9770)
         );
  AOI21_X1 U8663 ( .B1(n7007), .B2(n9761), .A(n9443), .ZN(n7009) );
  NAND2_X1 U8664 ( .A1(n7009), .A2(n7008), .ZN(n9766) );
  OAI211_X1 U8665 ( .C1(n7010), .C2(n7657), .A(n9770), .B(n9766), .ZN(n7053)
         );
  OAI22_X1 U8666 ( .A1(n9537), .A2(n7051), .B1(n9811), .B2(n6326), .ZN(n7011)
         );
  AOI21_X1 U8667 ( .B1(n7053), .B2(n9811), .A(n7011), .ZN(n7012) );
  INV_X1 U8668 ( .A(n7012), .ZN(P1_U3523) );
  OAI21_X1 U8669 ( .B1(n7014), .B2(n7015), .A(n7013), .ZN(n9755) );
  INV_X1 U8670 ( .A(n9755), .ZN(n7023) );
  XNOR2_X1 U8671 ( .A(n7016), .B(n7015), .ZN(n7019) );
  INV_X1 U8672 ( .A(n9215), .ZN(n7018) );
  OAI22_X1 U8673 ( .A1(n7018), .A2(n9167), .B1(n7017), .B2(n9169), .ZN(n9044)
         );
  AOI21_X1 U8674 ( .B1(n7019), .B2(n9463), .A(n9044), .ZN(n9757) );
  INV_X1 U8675 ( .A(n7020), .ZN(n7021) );
  OAI211_X1 U8676 ( .C1(n7055), .C2(n7022), .A(n7021), .B(n9521), .ZN(n9752)
         );
  OAI211_X1 U8677 ( .C1(n7023), .C2(n9525), .A(n9757), .B(n9752), .ZN(n7057)
         );
  INV_X1 U8678 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7024) );
  OAI22_X1 U8679 ( .A1(n9537), .A2(n7055), .B1(n9811), .B2(n7024), .ZN(n7025)
         );
  AOI21_X1 U8680 ( .B1(n7057), .B2(n9811), .A(n7025), .ZN(n7026) );
  INV_X1 U8681 ( .A(n7026), .ZN(P1_U3525) );
  INV_X1 U8682 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7028) );
  INV_X1 U8683 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7027) );
  MUX2_X1 U8684 ( .A(n7028), .B(n7027), .S(n8474), .Z(n7029) );
  NAND2_X1 U8685 ( .A1(n7029), .A2(n7044), .ZN(n7146) );
  INV_X1 U8686 ( .A(n7029), .ZN(n7030) );
  NAND2_X1 U8687 ( .A1(n7030), .A2(n7154), .ZN(n7031) );
  AND2_X1 U8688 ( .A1(n7146), .A2(n7031), .ZN(n7034) );
  INV_X1 U8689 ( .A(n7033), .ZN(n7032) );
  NOR2_X1 U8690 ( .A1(n7034), .A2(n7032), .ZN(n7037) );
  NAND2_X1 U8691 ( .A1(n7036), .A2(n7033), .ZN(n7035) );
  NAND2_X1 U8692 ( .A1(n7035), .A2(n7034), .ZN(n7147) );
  INV_X1 U8693 ( .A(n7147), .ZN(n7145) );
  AOI21_X1 U8694 ( .B1(n7037), .B2(n7036), .A(n7145), .ZN(n7050) );
  NAND2_X1 U8695 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(n7039), .ZN(n7155) );
  OAI21_X1 U8696 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n7039), .A(n7155), .ZN(
        n7048) );
  AOI21_X1 U8697 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n7041), .A(n7040), .ZN(
        n7042) );
  NOR2_X1 U8698 ( .A1(n7042), .A2(n7044), .ZN(n7136) );
  AOI21_X1 U8699 ( .B1(n4298), .B2(n7028), .A(n7135), .ZN(n7046) );
  INV_X1 U8700 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7522) );
  NAND2_X1 U8701 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8311) );
  OAI21_X1 U8702 ( .B1(n8506), .B2(n7522), .A(n8311), .ZN(n7043) );
  AOI21_X1 U8703 ( .B1(n7044), .B2(n8486), .A(n7043), .ZN(n7045) );
  OAI21_X1 U8704 ( .B1(n7046), .B2(n8519), .A(n7045), .ZN(n7047) );
  AOI21_X1 U8705 ( .B1(n8516), .B2(n7048), .A(n7047), .ZN(n7049) );
  OAI21_X1 U8706 ( .B1(n7050), .B2(n8481), .A(n7049), .ZN(P2_U3191) );
  OAI22_X1 U8707 ( .A1(n9604), .A2(n7051), .B1(n9795), .B2(n5086), .ZN(n7052)
         );
  AOI21_X1 U8708 ( .B1(n7053), .B2(n9795), .A(n7052), .ZN(n7054) );
  INV_X1 U8709 ( .A(n7054), .ZN(P1_U3456) );
  OAI22_X1 U8710 ( .A1(n9604), .A2(n7055), .B1(n9795), .B2(n5121), .ZN(n7056)
         );
  AOI21_X1 U8711 ( .B1(n7057), .B2(n9795), .A(n7056), .ZN(n7058) );
  INV_X1 U8712 ( .A(n7058), .ZN(P1_U3462) );
  XNOR2_X1 U8713 ( .A(n8205), .B(n9827), .ZN(n7285) );
  XNOR2_X1 U8714 ( .A(n7285), .B(n8379), .ZN(n7063) );
  INV_X1 U8715 ( .A(n7059), .ZN(n7060) );
  AOI21_X1 U8716 ( .B1(n7063), .B2(n7062), .A(n7286), .ZN(n7068) );
  INV_X1 U8717 ( .A(n8378), .ZN(n7367) );
  OAI22_X1 U8718 ( .A1(n7367), .A2(n8363), .B1(n8341), .B2(n7241), .ZN(n7064)
         );
  AOI211_X1 U8719 ( .C1(n7169), .C2(n8352), .A(n7065), .B(n7064), .ZN(n7067)
         );
  NAND2_X1 U8720 ( .A1(n8365), .A2(n7168), .ZN(n7066) );
  OAI211_X1 U8721 ( .C1(n7068), .C2(n8356), .A(n7067), .B(n7066), .ZN(P2_U3170) );
  NAND2_X1 U8722 ( .A1(n7069), .A2(n9463), .ZN(n7076) );
  AOI21_X1 U8723 ( .B1(n7072), .B2(n7071), .A(n7070), .ZN(n7075) );
  OR2_X1 U8724 ( .A1(n7211), .A2(n9167), .ZN(n7074) );
  NAND2_X1 U8725 ( .A1(n9215), .A2(n9138), .ZN(n7073) );
  AND2_X1 U8726 ( .A1(n7074), .A2(n7073), .ZN(n7129) );
  OAI21_X1 U8727 ( .B1(n7076), .B2(n7075), .A(n7129), .ZN(n7105) );
  AOI211_X1 U8728 ( .C1(n7131), .C2(n7077), .A(n9443), .B(n7191), .ZN(n7099)
         );
  NOR2_X1 U8729 ( .A1(n7105), .A2(n7099), .ZN(n7090) );
  OAI21_X1 U8730 ( .B1(n7080), .B2(n7079), .A(n7078), .ZN(n7098) );
  OAI22_X1 U8731 ( .A1(n9537), .A2(n7103), .B1(n9811), .B2(n5155), .ZN(n7081)
         );
  AOI21_X1 U8732 ( .B1(n7098), .B2(n9551), .A(n7081), .ZN(n7082) );
  OAI21_X1 U8733 ( .B1(n7090), .B2(n9812), .A(n7082), .ZN(P1_U3527) );
  AND2_X1 U8734 ( .A1(n7084), .A2(n7083), .ZN(n7096) );
  OAI22_X1 U8735 ( .A1(n9537), .A2(n7092), .B1(n9811), .B2(n5136), .ZN(n7085)
         );
  AOI21_X1 U8736 ( .B1(n7094), .B2(n9551), .A(n7085), .ZN(n7086) );
  OAI21_X1 U8737 ( .B1(n7096), .B2(n9812), .A(n7086), .ZN(P1_U3526) );
  INV_X1 U8738 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7087) );
  OAI22_X1 U8739 ( .A1(n9604), .A2(n7103), .B1(n9804), .B2(n7087), .ZN(n7088)
         );
  AOI21_X1 U8740 ( .B1(n7098), .B2(n5547), .A(n7088), .ZN(n7089) );
  OAI21_X1 U8741 ( .B1(n7090), .B2(n9619), .A(n7089), .ZN(P1_U3468) );
  INV_X1 U8742 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7091) );
  OAI22_X1 U8743 ( .A1(n9604), .A2(n7092), .B1(n9795), .B2(n7091), .ZN(n7093)
         );
  AOI21_X1 U8744 ( .B1(n7094), .B2(n5547), .A(n7093), .ZN(n7095) );
  OAI21_X1 U8745 ( .B1(n7096), .B2(n9619), .A(n7095), .ZN(P1_U3465) );
  NAND2_X1 U8746 ( .A1(n8382), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7097) );
  OAI21_X1 U8747 ( .B1(n8102), .B2(n8382), .A(n7097), .ZN(P2_U3521) );
  INV_X1 U8748 ( .A(n7098), .ZN(n7107) );
  NAND2_X1 U8749 ( .A1(n7099), .A2(n9450), .ZN(n7102) );
  INV_X1 U8750 ( .A(n7134), .ZN(n7100) );
  AOI22_X1 U8751 ( .A1(n9749), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7100), .B2(
        n9758), .ZN(n7101) );
  OAI211_X1 U8752 ( .C1(n7103), .C2(n9444), .A(n7102), .B(n7101), .ZN(n7104)
         );
  AOI21_X1 U8753 ( .B1(n7105), .B2(n9457), .A(n7104), .ZN(n7106) );
  OAI21_X1 U8754 ( .B1(n7107), .B2(n9460), .A(n7106), .ZN(P1_U3288) );
  INV_X1 U8755 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8524) );
  NAND2_X1 U8756 ( .A1(n4268), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7110) );
  NAND2_X1 U8757 ( .A1(n7108), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n7109) );
  OAI211_X1 U8758 ( .C1(n8524), .C2(n7111), .A(n7110), .B(n7109), .ZN(n7112)
         );
  INV_X1 U8759 ( .A(n7112), .ZN(n7113) );
  NAND2_X1 U8760 ( .A1(n8382), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7115) );
  OAI21_X1 U8761 ( .B1(n8521), .B2(n8382), .A(n7115), .ZN(P2_U3522) );
  CLKBUF_X1 U8762 ( .A(n9157), .Z(n9186) );
  AOI22_X1 U8763 ( .A1(n9214), .A2(n8988), .B1(n7593), .B2(n7131), .ZN(n7126)
         );
  INV_X1 U8764 ( .A(n7117), .ZN(n7118) );
  NAND2_X1 U8765 ( .A1(n7116), .A2(n7118), .ZN(n7119) );
  NAND2_X1 U8766 ( .A1(n7120), .A2(n7119), .ZN(n7124) );
  AOI22_X1 U8767 ( .A1(n9214), .A2(n7593), .B1(n7131), .B2(n4497), .ZN(n7122)
         );
  XOR2_X1 U8768 ( .A(n8978), .B(n7122), .Z(n7123) );
  OAI21_X1 U8769 ( .B1(n7126), .B2(n7125), .A(n7206), .ZN(n7127) );
  NAND2_X1 U8770 ( .A1(n7127), .A2(n9165), .ZN(n7133) );
  OAI21_X1 U8771 ( .B1(n9142), .B2(n7129), .A(n7128), .ZN(n7130) );
  AOI21_X1 U8772 ( .B1(n7131), .B2(n4264), .A(n7130), .ZN(n7132) );
  OAI211_X1 U8773 ( .C1(n9186), .C2(n7134), .A(n7133), .B(n7132), .ZN(P1_U3227) );
  NAND2_X1 U8774 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7340), .ZN(n7137) );
  OAI21_X1 U8775 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7340), .A(n7137), .ZN(
        n7138) );
  AOI21_X1 U8776 ( .B1(n7139), .B2(n7138), .A(n7338), .ZN(n7164) );
  INV_X1 U8777 ( .A(n7146), .ZN(n7144) );
  INV_X1 U8778 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7636) );
  INV_X1 U8779 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7140) );
  MUX2_X1 U8780 ( .A(n7636), .B(n7140), .S(n8474), .Z(n7141) );
  NAND2_X1 U8781 ( .A1(n7141), .A2(n7152), .ZN(n7352) );
  INV_X1 U8782 ( .A(n7141), .ZN(n7142) );
  NAND2_X1 U8783 ( .A1(n7142), .A2(n7340), .ZN(n7143) );
  AND2_X1 U8784 ( .A1(n7352), .A2(n7143), .ZN(n7148) );
  NOR3_X1 U8785 ( .A1(n7145), .A2(n7144), .A3(n7148), .ZN(n7151) );
  NAND2_X1 U8786 ( .A1(n7147), .A2(n7146), .ZN(n7149) );
  NAND2_X1 U8787 ( .A1(n7149), .A2(n7148), .ZN(n7353) );
  INV_X1 U8788 ( .A(n7353), .ZN(n7150) );
  OAI21_X1 U8789 ( .B1(n7151), .B2(n7150), .A(n8509), .ZN(n7163) );
  AOI22_X1 U8790 ( .A1(n7152), .A2(n7140), .B1(P2_REG1_REG_10__SCAN_IN), .B2(
        n7340), .ZN(n7158) );
  NAND2_X1 U8791 ( .A1(n7154), .A2(n7153), .ZN(n7156) );
  OAI21_X1 U8792 ( .B1(n7158), .B2(n7157), .A(n7341), .ZN(n7161) );
  INV_X1 U8793 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9990) );
  NOR2_X1 U8794 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9990), .ZN(n7776) );
  AOI21_X1 U8795 ( .B1(n7838), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7776), .ZN(
        n7159) );
  OAI21_X1 U8796 ( .B1(n7340), .B2(n8503), .A(n7159), .ZN(n7160) );
  AOI21_X1 U8797 ( .B1(n7161), .B2(n8516), .A(n7160), .ZN(n7162) );
  OAI211_X1 U8798 ( .C1(n7164), .C2(n8519), .A(n7163), .B(n7162), .ZN(P2_U3192) );
  NAND2_X1 U8799 ( .A1(n8004), .A2(n7998), .ZN(n8132) );
  XNOR2_X1 U8800 ( .A(n7165), .B(n8132), .ZN(n7166) );
  AOI222_X1 U8801 ( .A1(n8719), .A2(n7166), .B1(n8380), .B2(n8723), .C1(n8378), 
        .C2(n8726), .ZN(n9826) );
  INV_X1 U8802 ( .A(n8132), .ZN(n7995) );
  XNOR2_X1 U8803 ( .A(n7167), .B(n7995), .ZN(n9829) );
  INV_X1 U8804 ( .A(n8713), .ZN(n8736) );
  AOI22_X1 U8805 ( .A1(n8710), .A2(n7169), .B1(n8731), .B2(n7168), .ZN(n7170)
         );
  OAI21_X1 U8806 ( .B1(n6750), .B2(n9668), .A(n7170), .ZN(n7171) );
  AOI21_X1 U8807 ( .B1(n9829), .B2(n8736), .A(n7171), .ZN(n7172) );
  OAI21_X1 U8808 ( .B1(n9826), .B2(n9670), .A(n7172), .ZN(P2_U3229) );
  OAI21_X1 U8809 ( .B1(n7174), .B2(n7176), .A(n7173), .ZN(n7313) );
  OAI22_X1 U8810 ( .A1(n7211), .A2(n9169), .B1(n7485), .B2(n9167), .ZN(n7304)
         );
  INV_X1 U8811 ( .A(n7175), .ZN(n7195) );
  NOR2_X1 U8812 ( .A1(n7195), .A2(n7194), .ZN(n7178) );
  NOR3_X1 U8813 ( .A1(n7178), .A2(n7177), .A3(n7176), .ZN(n7326) );
  INV_X1 U8814 ( .A(n7326), .ZN(n7261) );
  OAI21_X1 U8815 ( .B1(n7178), .B2(n7177), .A(n7176), .ZN(n7179) );
  AOI21_X1 U8816 ( .B1(n7261), .B2(n7179), .A(n9412), .ZN(n7180) );
  AOI211_X1 U8817 ( .C1(n7181), .C2(n7313), .A(n7304), .B(n7180), .ZN(n7315)
         );
  INV_X1 U8818 ( .A(n7655), .ZN(n9760) );
  INV_X1 U8819 ( .A(n7190), .ZN(n7182) );
  INV_X1 U8820 ( .A(n7308), .ZN(n7320) );
  OAI211_X1 U8821 ( .C1(n7182), .C2(n7320), .A(n9521), .B(n7264), .ZN(n7314)
         );
  OAI22_X1 U8822 ( .A1(n9474), .A2(n7183), .B1(n7306), .B2(n9471), .ZN(n7184)
         );
  AOI21_X1 U8823 ( .B1(n9762), .B2(n7308), .A(n7184), .ZN(n7185) );
  OAI21_X1 U8824 ( .B1(n7314), .B2(n9765), .A(n7185), .ZN(n7186) );
  AOI21_X1 U8825 ( .B1(n7313), .B2(n9760), .A(n7186), .ZN(n7187) );
  OAI21_X1 U8826 ( .B1(n7315), .B2(n9749), .A(n7187), .ZN(P1_U3286) );
  OAI21_X1 U8827 ( .B1(n7189), .B2(n7194), .A(n7188), .ZN(n9784) );
  OAI211_X1 U8828 ( .C1(n7191), .C2(n9781), .A(n7190), .B(n9521), .ZN(n9780)
         );
  INV_X1 U8829 ( .A(n7192), .ZN(n7225) );
  AOI22_X1 U8830 ( .A1(n9762), .A2(n7210), .B1(n9758), .B2(n7225), .ZN(n7193)
         );
  OAI21_X1 U8831 ( .B1(n9780), .B2(n9765), .A(n7193), .ZN(n7200) );
  XNOR2_X1 U8832 ( .A(n7195), .B(n7194), .ZN(n7198) );
  OAI22_X1 U8833 ( .A1(n7196), .A2(n9169), .B1(n7298), .B2(n9167), .ZN(n7222)
         );
  INV_X1 U8834 ( .A(n7222), .ZN(n7197) );
  OAI21_X1 U8835 ( .B1(n7198), .B2(n9412), .A(n7197), .ZN(n9782) );
  MUX2_X1 U8836 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9782), .S(n9474), .Z(n7199)
         );
  AOI211_X1 U8837 ( .C1(n9754), .C2(n9784), .A(n7200), .B(n7199), .ZN(n7201)
         );
  INV_X1 U8838 ( .A(n7201), .ZN(P1_U3287) );
  INV_X1 U8839 ( .A(n7202), .ZN(n7204) );
  OAI222_X1 U8840 ( .A1(n8893), .A2(n7203), .B1(n8891), .B2(n7204), .C1(
        P2_U3151), .C2(n8441), .ZN(P2_U3278) );
  OAI222_X1 U8841 ( .A1(n8213), .A2(n7205), .B1(n9637), .B2(n7204), .C1(
        P1_U3086), .C2(n9260), .ZN(P1_U3338) );
  NAND2_X1 U8842 ( .A1(n7210), .A2(n4497), .ZN(n7208) );
  OR2_X1 U8843 ( .A1(n7211), .A2(n9056), .ZN(n7207) );
  NAND2_X1 U8844 ( .A1(n7208), .A2(n7207), .ZN(n7209) );
  XNOR2_X1 U8845 ( .A(n7209), .B(n8978), .ZN(n7214) );
  NAND2_X1 U8846 ( .A1(n7210), .A2(n7593), .ZN(n7213) );
  OR2_X1 U8847 ( .A1(n7211), .A2(n6689), .ZN(n7212) );
  NAND2_X1 U8848 ( .A1(n7213), .A2(n7212), .ZN(n7215) );
  NAND2_X1 U8849 ( .A1(n7214), .A2(n7215), .ZN(n7219) );
  INV_X1 U8850 ( .A(n7303), .ZN(n7221) );
  INV_X1 U8851 ( .A(n7214), .ZN(n7217) );
  INV_X1 U8852 ( .A(n7215), .ZN(n7216) );
  NAND2_X1 U8853 ( .A1(n7217), .A2(n7216), .ZN(n7302) );
  AOI21_X1 U8854 ( .B1(n7219), .B2(n7302), .A(n7218), .ZN(n7220) );
  AOI21_X1 U8855 ( .B1(n7221), .B2(n7302), .A(n7220), .ZN(n7227) );
  AOI22_X1 U8856 ( .A1(n4270), .A2(n7222), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n7223) );
  OAI21_X1 U8857 ( .B1(n9147), .B2(n9781), .A(n7223), .ZN(n7224) );
  AOI21_X1 U8858 ( .B1(n7225), .B2(n9144), .A(n7224), .ZN(n7226) );
  OAI21_X1 U8859 ( .B1(n7227), .B2(n9189), .A(n7226), .ZN(P1_U3239) );
  OAI22_X1 U8860 ( .A1(n8561), .A2(n7228), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9656), .ZN(n7231) );
  MUX2_X1 U8861 ( .A(n7229), .B(P2_REG2_REG_3__SCAN_IN), .S(n9670), .Z(n7230)
         );
  AOI211_X1 U8862 ( .C1(n8736), .C2(n7232), .A(n7231), .B(n7230), .ZN(n7233)
         );
  INV_X1 U8863 ( .A(n7233), .ZN(P2_U3230) );
  OR2_X1 U8864 ( .A1(n7234), .A2(n7984), .ZN(n7236) );
  NAND2_X1 U8865 ( .A1(n7236), .A2(n7235), .ZN(n9823) );
  INV_X1 U8866 ( .A(n9823), .ZN(n7250) );
  NAND2_X1 U8867 ( .A1(n8672), .A2(n7237), .ZN(n8534) );
  NAND2_X1 U8868 ( .A1(n7238), .A2(n9872), .ZN(n9820) );
  INV_X1 U8869 ( .A(n7239), .ZN(n9658) );
  NOR2_X1 U8870 ( .A1(n9820), .A2(n9658), .ZN(n7247) );
  INV_X1 U8871 ( .A(n8719), .ZN(n9815) );
  XNOR2_X1 U8872 ( .A(n7240), .B(n7984), .ZN(n7246) );
  INV_X1 U8873 ( .A(n7612), .ZN(n7244) );
  OAI22_X1 U8874 ( .A1(n7242), .A2(n9665), .B1(n7241), .B2(n9663), .ZN(n7243)
         );
  AOI21_X1 U8875 ( .B1(n9823), .B2(n7244), .A(n7243), .ZN(n7245) );
  OAI21_X1 U8876 ( .B1(n9815), .B2(n7246), .A(n7245), .ZN(n9821) );
  AOI211_X1 U8877 ( .C1(n8731), .C2(P2_REG3_REG_2__SCAN_IN), .A(n7247), .B(
        n9821), .ZN(n7248) );
  MUX2_X1 U8878 ( .A(n6599), .B(n7248), .S(n9668), .Z(n7249) );
  OAI21_X1 U8879 ( .B1(n7250), .B2(n8534), .A(n7249), .ZN(P2_U3231) );
  NAND2_X1 U8880 ( .A1(n7252), .A2(n7251), .ZN(n8134) );
  XNOR2_X1 U8881 ( .A(n7253), .B(n8134), .ZN(n7254) );
  AOI222_X1 U8882 ( .A1(n8719), .A2(n7254), .B1(n8377), .B2(n8726), .C1(n8379), 
        .C2(n8723), .ZN(n9831) );
  XNOR2_X1 U8883 ( .A(n7255), .B(n8134), .ZN(n9834) );
  AOI22_X1 U8884 ( .A1(n8710), .A2(n7291), .B1(n8731), .B2(n7292), .ZN(n7256)
         );
  OAI21_X1 U8885 ( .B1(n7257), .B2(n9668), .A(n7256), .ZN(n7258) );
  AOI21_X1 U8886 ( .B1(n9834), .B2(n8736), .A(n7258), .ZN(n7259) );
  OAI21_X1 U8887 ( .B1(n9831), .B2(n9670), .A(n7259), .ZN(P2_U3228) );
  NAND2_X1 U8888 ( .A1(n7261), .A2(n7260), .ZN(n7262) );
  XNOR2_X1 U8889 ( .A(n7262), .B(n7268), .ZN(n7263) );
  AOI22_X1 U8890 ( .A1(n9138), .A2(n9212), .B1(n9210), .B2(n9129), .ZN(n7492)
         );
  OAI21_X1 U8891 ( .B1(n7263), .B2(n9412), .A(n7492), .ZN(n7282) );
  NAND2_X1 U8892 ( .A1(n7264), .A2(n7484), .ZN(n7265) );
  NAND2_X1 U8893 ( .A1(n7265), .A2(n9521), .ZN(n7266) );
  NOR2_X1 U8894 ( .A1(n7430), .A2(n7266), .ZN(n7277) );
  NOR2_X1 U8895 ( .A1(n7282), .A2(n7277), .ZN(n7275) );
  OAI21_X1 U8896 ( .B1(n7269), .B2(n7268), .A(n7267), .ZN(n7276) );
  INV_X1 U8897 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7270) );
  OAI22_X1 U8898 ( .A1(n5524), .A2(n9537), .B1(n9811), .B2(n7270), .ZN(n7271)
         );
  AOI21_X1 U8899 ( .B1(n7276), .B2(n9551), .A(n7271), .ZN(n7272) );
  OAI21_X1 U8900 ( .B1(n7275), .B2(n9812), .A(n7272), .ZN(P1_U3530) );
  OAI22_X1 U8901 ( .A1(n5524), .A2(n9604), .B1(n9804), .B2(n5199), .ZN(n7273)
         );
  AOI21_X1 U8902 ( .B1(n7276), .B2(n5547), .A(n7273), .ZN(n7274) );
  OAI21_X1 U8903 ( .B1(n7275), .B2(n9619), .A(n7274), .ZN(P1_U3477) );
  INV_X1 U8904 ( .A(n7276), .ZN(n7284) );
  NAND2_X1 U8905 ( .A1(n7277), .A2(n9450), .ZN(n7280) );
  INV_X1 U8906 ( .A(n7278), .ZN(n7494) );
  AOI22_X1 U8907 ( .A1(n9749), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7494), .B2(
        n9758), .ZN(n7279) );
  OAI211_X1 U8908 ( .C1(n5524), .C2(n9444), .A(n7280), .B(n7279), .ZN(n7281)
         );
  AOI21_X1 U8909 ( .B1(n7282), .B2(n9474), .A(n7281), .ZN(n7283) );
  OAI21_X1 U8910 ( .B1(n9460), .B2(n7284), .A(n7283), .ZN(P1_U3285) );
  XNOR2_X1 U8911 ( .A(n8205), .B(n9832), .ZN(n7361) );
  XNOR2_X1 U8912 ( .A(n7361), .B(n8378), .ZN(n7362) );
  INV_X1 U8913 ( .A(n7285), .ZN(n7287) );
  XOR2_X1 U8914 ( .A(n7362), .B(n7363), .Z(n7295) );
  OAI22_X1 U8915 ( .A1(n7288), .A2(n8341), .B1(n8363), .B2(n8219), .ZN(n7289)
         );
  AOI211_X1 U8916 ( .C1(n7291), .C2(n8352), .A(n7290), .B(n7289), .ZN(n7294)
         );
  NAND2_X1 U8917 ( .A1(n8365), .A2(n7292), .ZN(n7293) );
  OAI211_X1 U8918 ( .C1(n7295), .C2(n8356), .A(n7294), .B(n7293), .ZN(P2_U3167) );
  INV_X1 U8919 ( .A(n7296), .ZN(n7311) );
  OAI222_X1 U8920 ( .A1(n8213), .A2(n7297), .B1(n9637), .B2(n7311), .C1(n9738), 
        .C2(P1_U3086), .ZN(P1_U3337) );
  OAI22_X1 U8921 ( .A1(n7320), .A2(n9056), .B1(n7298), .B2(n6689), .ZN(n7479)
         );
  NAND2_X1 U8922 ( .A1(n7308), .A2(n4497), .ZN(n7300) );
  OR2_X1 U8923 ( .A1(n7298), .A2(n9056), .ZN(n7299) );
  NAND2_X1 U8924 ( .A1(n7300), .A2(n7299), .ZN(n7301) );
  XNOR2_X1 U8925 ( .A(n7301), .B(n8978), .ZN(n7478) );
  XOR2_X1 U8926 ( .A(n7479), .B(n7478), .Z(n7482) );
  XOR2_X1 U8927 ( .A(n7482), .B(n7483), .Z(n7310) );
  AOI22_X1 U8928 ( .A1(n4270), .A2(n7304), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n7305) );
  OAI21_X1 U8929 ( .B1(n9186), .B2(n7306), .A(n7305), .ZN(n7307) );
  AOI21_X1 U8930 ( .B1(n7308), .B2(n4264), .A(n7307), .ZN(n7309) );
  OAI21_X1 U8931 ( .B1(n7310), .B2(n9189), .A(n7309), .ZN(P1_U3213) );
  INV_X1 U8932 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7312) );
  INV_X1 U8933 ( .A(n8485), .ZN(n8511) );
  OAI222_X1 U8934 ( .A1(n8893), .A2(n7312), .B1(n8511), .B2(P2_U3151), .C1(
        n8891), .C2(n7311), .ZN(P2_U3277) );
  INV_X1 U8935 ( .A(n7313), .ZN(n7316) );
  OAI211_X1 U8936 ( .C1(n7316), .C2(n7657), .A(n7315), .B(n7314), .ZN(n7322)
         );
  OAI22_X1 U8937 ( .A1(n9537), .A2(n7320), .B1(n9811), .B2(n5213), .ZN(n7317)
         );
  AOI21_X1 U8938 ( .B1(n7322), .B2(n9811), .A(n7317), .ZN(n7318) );
  INV_X1 U8939 ( .A(n7318), .ZN(P1_U3529) );
  INV_X1 U8940 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7319) );
  OAI22_X1 U8941 ( .A1(n9604), .A2(n7320), .B1(n9804), .B2(n7319), .ZN(n7321)
         );
  AOI21_X1 U8942 ( .B1(n7322), .B2(n9795), .A(n7321), .ZN(n7323) );
  INV_X1 U8943 ( .A(n7323), .ZN(P1_U3474) );
  AOI21_X1 U8944 ( .B1(n7326), .B2(n7325), .A(n7324), .ZN(n7327) );
  XNOR2_X1 U8945 ( .A(n7327), .B(n7330), .ZN(n7328) );
  NOR2_X1 U8946 ( .A1(n7485), .A2(n9169), .ZN(n7558) );
  AOI21_X1 U8947 ( .B1(n7328), .B2(n9463), .A(n7558), .ZN(n9786) );
  OAI21_X1 U8948 ( .B1(n7331), .B2(n7330), .A(n7329), .ZN(n9789) );
  NAND2_X1 U8949 ( .A1(n9789), .A2(n9754), .ZN(n7337) );
  OAI22_X1 U8950 ( .A1(n9474), .A2(n7332), .B1(n7562), .B2(n9471), .ZN(n7335)
         );
  XNOR2_X1 U8951 ( .A(n7430), .B(n7564), .ZN(n7333) );
  NOR2_X1 U8952 ( .A1(n7644), .A2(n9167), .ZN(n7559) );
  AOI21_X1 U8953 ( .B1(n7333), .B2(n9521), .A(n7559), .ZN(n9785) );
  NOR2_X1 U8954 ( .A1(n9785), .A2(n9765), .ZN(n7334) );
  AOI211_X1 U8955 ( .C1(n9762), .C2(n7564), .A(n7335), .B(n7334), .ZN(n7336)
         );
  OAI211_X1 U8956 ( .C1(n9749), .C2(n9786), .A(n7337), .B(n7336), .ZN(P1_U3284) );
  INV_X1 U8957 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7709) );
  NOR2_X1 U8958 ( .A1(n7709), .A2(n7339), .ZN(n7439) );
  AOI21_X1 U8959 ( .B1(n7709), .B2(n7339), .A(n7439), .ZN(n7359) );
  NAND2_X1 U8960 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7340), .ZN(n7342) );
  NAND2_X1 U8961 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n7343), .ZN(n7446) );
  OAI21_X1 U8962 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n7343), .A(n7446), .ZN(
        n7357) );
  AND2_X1 U8963 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7853) );
  AOI21_X1 U8964 ( .B1(n7838), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7853), .ZN(
        n7344) );
  OAI21_X1 U8965 ( .B1(n7445), .B2(n8503), .A(n7344), .ZN(n7356) );
  NAND2_X1 U8966 ( .A1(n7353), .A2(n7352), .ZN(n7349) );
  INV_X1 U8967 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7345) );
  MUX2_X1 U8968 ( .A(n7709), .B(n7345), .S(n8474), .Z(n7346) );
  NAND2_X1 U8969 ( .A1(n7346), .A2(n7438), .ZN(n7457) );
  INV_X1 U8970 ( .A(n7346), .ZN(n7347) );
  NAND2_X1 U8971 ( .A1(n7347), .A2(n7445), .ZN(n7348) );
  AND2_X1 U8972 ( .A1(n7457), .A2(n7348), .ZN(n7350) );
  NAND2_X1 U8973 ( .A1(n7349), .A2(n7350), .ZN(n7458) );
  INV_X1 U8974 ( .A(n7350), .ZN(n7351) );
  NAND3_X1 U8975 ( .A1(n7353), .A2(n7352), .A3(n7351), .ZN(n7354) );
  AOI21_X1 U8976 ( .B1(n7458), .B2(n7354), .A(n8481), .ZN(n7355) );
  AOI211_X1 U8977 ( .C1(n7357), .C2(n8516), .A(n7356), .B(n7355), .ZN(n7358)
         );
  OAI21_X1 U8978 ( .B1(n7359), .B2(n8519), .A(n7358), .ZN(P2_U3193) );
  INV_X1 U8979 ( .A(n7375), .ZN(n7373) );
  XNOR2_X1 U8980 ( .A(n7360), .B(n8205), .ZN(n7568) );
  XNOR2_X1 U8981 ( .A(n7568), .B(n8377), .ZN(n7365) );
  AOI211_X1 U8982 ( .C1(n7365), .C2(n7364), .A(n8356), .B(n7567), .ZN(n7366)
         );
  INV_X1 U8983 ( .A(n7366), .ZN(n7371) );
  OAI22_X1 U8984 ( .A1(n7367), .A2(n8341), .B1(n8363), .B2(n7569), .ZN(n7368)
         );
  AOI211_X1 U8985 ( .C1(n9840), .C2(n8352), .A(n7369), .B(n7368), .ZN(n7370)
         );
  OAI211_X1 U8986 ( .C1(n7373), .C2(n7372), .A(n7371), .B(n7370), .ZN(P2_U3179) );
  XOR2_X1 U8987 ( .A(n7374), .B(n8137), .Z(n9837) );
  AOI22_X1 U8988 ( .A1(n8710), .A2(n9840), .B1(n8731), .B2(n7375), .ZN(n7383)
         );
  INV_X1 U8989 ( .A(n8137), .ZN(n7376) );
  XNOR2_X1 U8990 ( .A(n7377), .B(n7376), .ZN(n7378) );
  NAND2_X1 U8991 ( .A1(n7378), .A2(n8719), .ZN(n7380) );
  AOI22_X1 U8992 ( .A1(n8723), .A2(n8378), .B1(n8376), .B2(n8726), .ZN(n7379)
         );
  NAND2_X1 U8993 ( .A1(n7380), .A2(n7379), .ZN(n9839) );
  MUX2_X1 U8994 ( .A(n9839), .B(P2_REG2_REG_6__SCAN_IN), .S(n9670), .Z(n7381)
         );
  INV_X1 U8995 ( .A(n7381), .ZN(n7382) );
  OAI211_X1 U8996 ( .C1(n9837), .C2(n8713), .A(n7383), .B(n7382), .ZN(P2_U3227) );
  NOR2_X1 U8997 ( .A1(n9230), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7384) );
  AOI21_X1 U8998 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9230), .A(n7384), .ZN(
        n7389) );
  NAND2_X1 U8999 ( .A1(n9649), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7385) );
  OAI21_X1 U9000 ( .B1(n9649), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7385), .ZN(
        n9642) );
  OAI21_X1 U9001 ( .B1(n7392), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7386), .ZN(
        n9643) );
  NOR2_X1 U9002 ( .A1(n9642), .A2(n9643), .ZN(n9641) );
  NAND2_X1 U9003 ( .A1(n9677), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7387) );
  OAI21_X1 U9004 ( .B1(n9677), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7387), .ZN(
        n9680) );
  OAI21_X1 U9005 ( .B1(n7389), .B2(n7388), .A(n9229), .ZN(n7401) );
  NAND2_X1 U9006 ( .A1(n9649), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7390) );
  OAI21_X1 U9007 ( .B1(n9649), .B2(P1_REG1_REG_10__SCAN_IN), .A(n7390), .ZN(
        n9645) );
  OAI21_X1 U9008 ( .B1(n7392), .B2(P1_REG1_REG_9__SCAN_IN), .A(n7391), .ZN(
        n9646) );
  NOR2_X1 U9009 ( .A1(n9645), .A2(n9646), .ZN(n9644) );
  MUX2_X1 U9010 ( .A(n7393), .B(P1_REG1_REG_11__SCAN_IN), .S(n9677), .Z(n9685)
         );
  NOR2_X1 U9011 ( .A1(n9684), .A2(n9685), .ZN(n9683) );
  AOI21_X1 U9012 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9677), .A(n9683), .ZN(
        n7395) );
  AOI22_X1 U9013 ( .A1(n9230), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n5276), .B2(
        n7399), .ZN(n7394) );
  NAND2_X1 U9014 ( .A1(n7395), .A2(n7394), .ZN(n9220) );
  OAI21_X1 U9015 ( .B1(n7395), .B2(n7394), .A(n9220), .ZN(n7396) );
  NAND2_X1 U9016 ( .A1(n7396), .A2(n9733), .ZN(n7398) );
  AND2_X1 U9017 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7765) );
  AOI21_X1 U9018 ( .B1(n9247), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n7765), .ZN(
        n7397) );
  OAI211_X1 U9019 ( .C1(n9739), .C2(n7399), .A(n7398), .B(n7397), .ZN(n7400)
         );
  AOI21_X1 U9020 ( .B1(n9682), .B2(n7401), .A(n7400), .ZN(n7402) );
  INV_X1 U9021 ( .A(n7402), .ZN(P1_U3255) );
  INV_X1 U9022 ( .A(n7403), .ZN(n8211) );
  OAI222_X1 U9023 ( .A1(n8893), .A2(n7405), .B1(n8891), .B2(n8211), .C1(n8502), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  NAND2_X1 U9024 ( .A1(n7406), .A2(n7407), .ZN(n7408) );
  XNOR2_X1 U9025 ( .A(n7408), .B(n8141), .ZN(n9847) );
  INV_X1 U9026 ( .A(n7467), .ZN(n7410) );
  OAI21_X1 U9027 ( .B1(n7410), .B2(n7409), .A(n8141), .ZN(n7412) );
  NAND3_X1 U9028 ( .A1(n7412), .A2(n8719), .A3(n7411), .ZN(n7414) );
  AOI22_X1 U9029 ( .A1(n8374), .A2(n8726), .B1(n8723), .B2(n8376), .ZN(n7413)
         );
  NAND2_X1 U9030 ( .A1(n7414), .A2(n7413), .ZN(n9849) );
  INV_X1 U9031 ( .A(n9850), .ZN(n7416) );
  AOI22_X1 U9032 ( .A1(n9670), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n8731), .B2(
        n7572), .ZN(n7415) );
  OAI21_X1 U9033 ( .B1(n7416), .B2(n8561), .A(n7415), .ZN(n7417) );
  AOI21_X1 U9034 ( .B1(n9849), .B2(n8672), .A(n7417), .ZN(n7418) );
  OAI21_X1 U9035 ( .B1(n9847), .B2(n8713), .A(n7418), .ZN(P2_U3225) );
  OAI21_X1 U9036 ( .B1(n7420), .B2(n7419), .A(n7427), .ZN(n7422) );
  AOI21_X1 U9037 ( .B1(n7422), .B2(n7421), .A(n9412), .ZN(n7425) );
  OR2_X1 U9038 ( .A1(n7669), .A2(n9167), .ZN(n7424) );
  OR2_X1 U9039 ( .A1(n7554), .A2(n9169), .ZN(n7423) );
  NAND2_X1 U9040 ( .A1(n7424), .A2(n7423), .ZN(n7596) );
  NOR2_X1 U9041 ( .A1(n7425), .A2(n7596), .ZN(n9791) );
  OAI21_X1 U9042 ( .B1(n7428), .B2(n7427), .A(n7426), .ZN(n9794) );
  NAND2_X1 U9043 ( .A1(n9794), .A2(n9754), .ZN(n7436) );
  OAI22_X1 U9044 ( .A1(n9474), .A2(n7429), .B1(n7598), .B2(n9471), .ZN(n7434)
         );
  INV_X1 U9045 ( .A(n7430), .ZN(n7431) );
  OAI21_X1 U9046 ( .B1(n7431), .B2(n7564), .A(n7600), .ZN(n7432) );
  NAND3_X1 U9047 ( .A1(n7432), .A2(n9521), .A3(n7649), .ZN(n9790) );
  NOR2_X1 U9048 ( .A1(n9790), .A2(n9765), .ZN(n7433) );
  AOI211_X1 U9049 ( .C1(n9762), .C2(n7600), .A(n7434), .B(n7433), .ZN(n7435)
         );
  OAI211_X1 U9050 ( .C1(n9749), .C2(n9791), .A(n7436), .B(n7435), .ZN(P1_U3283) );
  NOR2_X1 U9051 ( .A1(n7438), .A2(n7437), .ZN(n7440) );
  INV_X1 U9052 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7441) );
  AOI22_X1 U9053 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n7687), .B1(n7684), .B2(
        n7441), .ZN(n7442) );
  AOI21_X1 U9054 ( .B1(n7443), .B2(n7442), .A(n7683), .ZN(n7464) );
  INV_X1 U9055 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10012) );
  AOI22_X1 U9056 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n7684), .B1(n7687), .B2(
        n10012), .ZN(n7449) );
  NAND2_X1 U9057 ( .A1(n7445), .A2(n7444), .ZN(n7447) );
  OAI21_X1 U9058 ( .B1(n7449), .B2(n7448), .A(n7686), .ZN(n7462) );
  INV_X1 U9059 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10057) );
  NOR2_X1 U9060 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10057), .ZN(n7805) );
  AOI21_X1 U9061 ( .B1(n7838), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7805), .ZN(
        n7450) );
  OAI21_X1 U9062 ( .B1(n7684), .B2(n8503), .A(n7450), .ZN(n7461) );
  NAND2_X1 U9063 ( .A1(n7458), .A2(n7457), .ZN(n7454) );
  MUX2_X1 U9064 ( .A(n7441), .B(n10012), .S(n8474), .Z(n7451) );
  NAND2_X1 U9065 ( .A1(n7451), .A2(n7687), .ZN(n7696) );
  INV_X1 U9066 ( .A(n7451), .ZN(n7452) );
  NAND2_X1 U9067 ( .A1(n7452), .A2(n7684), .ZN(n7453) );
  AND2_X1 U9068 ( .A1(n7696), .A2(n7453), .ZN(n7455) );
  NAND2_X1 U9069 ( .A1(n7454), .A2(n7455), .ZN(n7697) );
  INV_X1 U9070 ( .A(n7455), .ZN(n7456) );
  NAND3_X1 U9071 ( .A1(n7458), .A2(n7457), .A3(n7456), .ZN(n7459) );
  AOI21_X1 U9072 ( .B1(n7697), .B2(n7459), .A(n8481), .ZN(n7460) );
  AOI211_X1 U9073 ( .C1(n7462), .C2(n8516), .A(n7461), .B(n7460), .ZN(n7463)
         );
  OAI21_X1 U9074 ( .B1(n7464), .B2(n8519), .A(n7463), .ZN(P2_U3194) );
  OAI21_X1 U9075 ( .B1(n7466), .B2(n7465), .A(n7406), .ZN(n9844) );
  OAI21_X1 U9076 ( .B1(n4878), .B2(n8138), .A(n7467), .ZN(n7469) );
  OAI22_X1 U9077 ( .A1(n8219), .A2(n9665), .B1(n8313), .B2(n9663), .ZN(n7468)
         );
  AOI21_X1 U9078 ( .B1(n7469), .B2(n8719), .A(n7468), .ZN(n7470) );
  OAI21_X1 U9079 ( .B1(n9844), .B2(n7612), .A(n7470), .ZN(n9846) );
  NAND2_X1 U9080 ( .A1(n9846), .A2(n8672), .ZN(n7475) );
  INV_X1 U9081 ( .A(n9843), .ZN(n8218) );
  INV_X1 U9082 ( .A(n8222), .ZN(n7471) );
  OAI22_X1 U9083 ( .A1(n9668), .A2(n7472), .B1(n7471), .B2(n9656), .ZN(n7473)
         );
  AOI21_X1 U9084 ( .B1(n8710), .B2(n8218), .A(n7473), .ZN(n7474) );
  OAI211_X1 U9085 ( .C1(n9844), .C2(n8534), .A(n7475), .B(n7474), .ZN(P2_U3226) );
  NAND2_X1 U9086 ( .A1(n7484), .A2(n7593), .ZN(n7477) );
  OR2_X1 U9087 ( .A1(n7485), .A2(n6689), .ZN(n7476) );
  NAND2_X1 U9088 ( .A1(n7477), .A2(n7476), .ZN(n7583) );
  INV_X1 U9089 ( .A(n7583), .ZN(n7582) );
  INV_X1 U9090 ( .A(n7478), .ZN(n7481) );
  INV_X1 U9091 ( .A(n7479), .ZN(n7480) );
  NAND2_X1 U9092 ( .A1(n7484), .A2(n4497), .ZN(n7487) );
  INV_X2 U9093 ( .A(n7593), .ZN(n9056) );
  OR2_X1 U9094 ( .A1(n7485), .A2(n9056), .ZN(n7486) );
  NAND2_X1 U9095 ( .A1(n7487), .A2(n7486), .ZN(n7488) );
  XNOR2_X1 U9096 ( .A(n7488), .B(n8978), .ZN(n7584) );
  INV_X1 U9097 ( .A(n7584), .ZN(n7581) );
  XNOR2_X1 U9098 ( .A(n7591), .B(n7581), .ZN(n7489) );
  NAND2_X1 U9099 ( .A1(n7489), .A2(n7582), .ZN(n7552) );
  OAI21_X1 U9100 ( .B1(n7582), .B2(n7489), .A(n7552), .ZN(n7490) );
  NAND2_X1 U9101 ( .A1(n7490), .A2(n9165), .ZN(n7496) );
  OAI22_X1 U9102 ( .A1(n9142), .A2(n7492), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7491), .ZN(n7493) );
  AOI21_X1 U9103 ( .B1(n7494), .B2(n9144), .A(n7493), .ZN(n7495) );
  OAI211_X1 U9104 ( .C1(n5524), .C2(n9147), .A(n7496), .B(n7495), .ZN(P1_U3221) );
  INV_X1 U9105 ( .A(n7497), .ZN(n7550) );
  OAI222_X1 U9106 ( .A1(n8901), .A2(n7550), .B1(P2_U3151), .B2(n7499), .C1(
        n7498), .C2(n8893), .ZN(P2_U3275) );
  INV_X1 U9107 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8455) );
  INV_X1 U9108 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9947) );
  NOR2_X1 U9109 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7543) );
  NOR2_X1 U9110 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7540) );
  INV_X1 U9111 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7538) );
  INV_X1 U9112 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9965) );
  NOR2_X1 U9113 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7536) );
  NOR2_X1 U9114 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7533) );
  NOR2_X1 U9115 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7529) );
  NOR2_X1 U9116 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7526) );
  NOR2_X1 U9117 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7524) );
  NOR2_X1 U9118 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7521) );
  NOR2_X1 U9119 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(P2_ADDR_REG_7__SCAN_IN), 
        .ZN(n7517) );
  NOR2_X1 U9120 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7514) );
  NOR2_X1 U9121 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7511) );
  NOR2_X1 U9122 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7509) );
  NAND2_X1 U9123 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7506) );
  XNOR2_X1 U9124 ( .A(n7500), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(n10084) );
  NAND2_X1 U9125 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7504) );
  AOI21_X1 U9126 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9891) );
  NAND2_X1 U9127 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7501) );
  NOR2_X1 U9128 ( .A1(n6340), .A2(n7501), .ZN(n9892) );
  NOR2_X1 U9129 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n9892), .ZN(n7502) );
  NOR2_X1 U9130 ( .A1(n9891), .A2(n7502), .ZN(n10082) );
  XOR2_X1 U9131 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10081) );
  NAND2_X1 U9132 ( .A1(n10082), .A2(n10081), .ZN(n7503) );
  NAND2_X1 U9133 ( .A1(n7504), .A2(n7503), .ZN(n10083) );
  NAND2_X1 U9134 ( .A1(n10084), .A2(n10083), .ZN(n7505) );
  NAND2_X1 U9135 ( .A1(n7506), .A2(n7505), .ZN(n10086) );
  XOR2_X1 U9136 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n7507), .Z(n10085) );
  NOR2_X1 U9137 ( .A1(n10086), .A2(n10085), .ZN(n7508) );
  NOR2_X1 U9138 ( .A1(n7509), .A2(n7508), .ZN(n10074) );
  XOR2_X1 U9139 ( .A(n9991), .B(P1_ADDR_REG_5__SCAN_IN), .Z(n10073) );
  NOR2_X1 U9140 ( .A1(n10074), .A2(n10073), .ZN(n7510) );
  NOR2_X1 U9141 ( .A1(n7511), .A2(n7510), .ZN(n10072) );
  INV_X1 U9142 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7512) );
  XOR2_X1 U9143 ( .A(n7512), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10071) );
  NOR2_X1 U9144 ( .A1(n10072), .A2(n10071), .ZN(n7513) );
  NOR2_X1 U9145 ( .A1(n7514), .A2(n7513), .ZN(n10080) );
  XOR2_X1 U9146 ( .A(n7515), .B(P2_ADDR_REG_7__SCAN_IN), .Z(n10079) );
  NOR2_X1 U9147 ( .A1(n10080), .A2(n10079), .ZN(n7516) );
  NOR2_X1 U9148 ( .A1(n7517), .A2(n7516), .ZN(n10078) );
  AOI22_X1 U9149 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n7519), .B1(
        P1_ADDR_REG_8__SCAN_IN), .B2(n7518), .ZN(n10077) );
  NOR2_X1 U9150 ( .A1(n10078), .A2(n10077), .ZN(n7520) );
  NOR2_X1 U9151 ( .A1(n7521), .A2(n7520), .ZN(n10076) );
  AOI22_X1 U9152 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n6734), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n7522), .ZN(n10075) );
  NOR2_X1 U9153 ( .A1(n10076), .A2(n10075), .ZN(n7523) );
  NOR2_X1 U9154 ( .A1(n7524), .A2(n7523), .ZN(n9912) );
  INV_X1 U9155 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9652) );
  INV_X1 U9156 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n9997) );
  AOI22_X1 U9157 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n9652), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n9997), .ZN(n9911) );
  NOR2_X1 U9158 ( .A1(n9912), .A2(n9911), .ZN(n7525) );
  NOR2_X1 U9159 ( .A1(n7526), .A2(n7525), .ZN(n9910) );
  INV_X1 U9160 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9693) );
  INV_X1 U9161 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7527) );
  AOI22_X1 U9162 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n9693), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n7527), .ZN(n9909) );
  NOR2_X1 U9163 ( .A1(n9910), .A2(n9909), .ZN(n7528) );
  NOR2_X1 U9164 ( .A1(n7529), .A2(n7528), .ZN(n9908) );
  INV_X1 U9165 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7531) );
  INV_X1 U9166 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7530) );
  AOI22_X1 U9167 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n7531), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n7530), .ZN(n9907) );
  NOR2_X1 U9168 ( .A1(n9908), .A2(n9907), .ZN(n7532) );
  NOR2_X1 U9169 ( .A1(n7533), .A2(n7532), .ZN(n9906) );
  INV_X1 U9170 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9705) );
  INV_X1 U9171 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7534) );
  AOI22_X1 U9172 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n9705), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n7534), .ZN(n9905) );
  NOR2_X1 U9173 ( .A1(n9906), .A2(n9905), .ZN(n7535) );
  NOR2_X1 U9174 ( .A1(n7536), .A2(n7535), .ZN(n9904) );
  AOI22_X1 U9175 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n9965), .B1(
        P1_ADDR_REG_14__SCAN_IN), .B2(n7538), .ZN(n9903) );
  NOR2_X1 U9176 ( .A1(n9904), .A2(n9903), .ZN(n7537) );
  AOI21_X1 U9177 ( .B1(n7538), .B2(n9965), .A(n7537), .ZN(n9902) );
  INV_X1 U9178 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9729) );
  INV_X1 U9179 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8402) );
  AOI22_X1 U9180 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n9729), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n8402), .ZN(n9901) );
  NOR2_X1 U9181 ( .A1(n9902), .A2(n9901), .ZN(n7539) );
  NOR2_X1 U9182 ( .A1(n7540), .A2(n7539), .ZN(n9900) );
  INV_X1 U9183 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7541) );
  INV_X1 U9184 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8433) );
  AOI22_X1 U9185 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n7541), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n8433), .ZN(n9899) );
  NOR2_X1 U9186 ( .A1(n9900), .A2(n9899), .ZN(n7542) );
  NOR2_X1 U9187 ( .A1(n7543), .A2(n7542), .ZN(n9898) );
  AOI22_X1 U9188 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n9947), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n8455), .ZN(n9897) );
  NOR2_X1 U9189 ( .A1(n9898), .A2(n9897), .ZN(n7544) );
  AOI21_X1 U9190 ( .B1(n8455), .B2(n9947), .A(n7544), .ZN(n7545) );
  AND2_X1 U9191 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7545), .ZN(n9894) );
  NOR2_X1 U9192 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n9894), .ZN(n7546) );
  NOR2_X1 U9193 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7545), .ZN(n9895) );
  NOR2_X1 U9194 ( .A1(n7546), .A2(n9895), .ZN(n7548) );
  XNOR2_X1 U9195 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7547) );
  XNOR2_X1 U9196 ( .A(n7548), .B(n7547), .ZN(ADD_1068_U4) );
  OAI222_X1 U9197 ( .A1(P1_U3086), .A2(n7551), .B1(n9637), .B2(n7550), .C1(
        n7549), .C2(n8213), .ZN(P1_U3335) );
  OAI21_X1 U9198 ( .B1(n7591), .B2(n7584), .A(n7552), .ZN(n7557) );
  OAI22_X1 U9199 ( .A1(n9787), .A2(n9058), .B1(n7554), .B2(n9056), .ZN(n7553)
         );
  XOR2_X1 U9200 ( .A(n8978), .B(n7553), .Z(n7585) );
  NOR2_X1 U9201 ( .A1(n7554), .A2(n6689), .ZN(n7555) );
  AOI21_X1 U9202 ( .B1(n7564), .B2(n7593), .A(n7555), .ZN(n7586) );
  XNOR2_X1 U9203 ( .A(n7585), .B(n7586), .ZN(n7556) );
  XNOR2_X1 U9204 ( .A(n7557), .B(n7556), .ZN(n7566) );
  OAI21_X1 U9205 ( .B1(n7559), .B2(n7558), .A(n4270), .ZN(n7560) );
  OAI211_X1 U9206 ( .C1(n9186), .C2(n7562), .A(n7561), .B(n7560), .ZN(n7563)
         );
  AOI21_X1 U9207 ( .B1(n7564), .B2(n4264), .A(n7563), .ZN(n7565) );
  OAI21_X1 U9208 ( .B1(n7566), .B2(n9189), .A(n7565), .ZN(P1_U3231) );
  XNOR2_X1 U9209 ( .A(n9843), .B(n8205), .ZN(n7570) );
  XNOR2_X1 U9210 ( .A(n7570), .B(n7569), .ZN(n8216) );
  XNOR2_X1 U9211 ( .A(n9850), .B(n8205), .ZN(n7769) );
  XNOR2_X1 U9212 ( .A(n7769), .B(n8375), .ZN(n7771) );
  XNOR2_X1 U9213 ( .A(n7772), .B(n7771), .ZN(n7578) );
  AOI21_X1 U9214 ( .B1(n8361), .B2(n8376), .A(n7571), .ZN(n7576) );
  NAND2_X1 U9215 ( .A1(n8352), .A2(n9850), .ZN(n7575) );
  NAND2_X1 U9216 ( .A1(n8365), .A2(n7572), .ZN(n7574) );
  OR2_X1 U9217 ( .A1(n8363), .A2(n7773), .ZN(n7573) );
  NAND4_X1 U9218 ( .A1(n7576), .A2(n7575), .A3(n7574), .A4(n7573), .ZN(n7577)
         );
  AOI21_X1 U9219 ( .B1(n7578), .B2(n8336), .A(n7577), .ZN(n7579) );
  INV_X1 U9220 ( .A(n7579), .ZN(P2_U3161) );
  INV_X1 U9221 ( .A(n5617), .ZN(n7604) );
  OAI222_X1 U9222 ( .A1(n8901), .A2(n7604), .B1(P2_U3151), .B2(n8125), .C1(
        n7580), .C2(n8893), .ZN(P2_U3274) );
  AOI22_X1 U9223 ( .A1(n7585), .A2(n7586), .B1(n7582), .B2(n7581), .ZN(n7590)
         );
  NAND2_X1 U9224 ( .A1(n7584), .A2(n7583), .ZN(n7587) );
  AOI21_X1 U9225 ( .B1(n7586), .B2(n7587), .A(n7585), .ZN(n7589) );
  NOR2_X1 U9226 ( .A1(n7587), .A2(n7586), .ZN(n7588) );
  OAI22_X1 U9227 ( .A1(n9792), .A2(n9058), .B1(n7644), .B2(n9056), .ZN(n7592)
         );
  OAI22_X1 U9228 ( .A1(n9792), .A2(n9056), .B1(n7644), .B2(n6689), .ZN(n7594)
         );
  AOI21_X1 U9229 ( .B1(n7595), .B2(n7594), .A(n7668), .ZN(n7602) );
  AOI22_X1 U9230 ( .A1(n4270), .A2(n7596), .B1(P1_REG3_REG_10__SCAN_IN), .B2(
        P1_U3086), .ZN(n7597) );
  OAI21_X1 U9231 ( .B1(n9186), .B2(n7598), .A(n7597), .ZN(n7599) );
  AOI21_X1 U9232 ( .B1(n7600), .B2(n4264), .A(n7599), .ZN(n7601) );
  OAI21_X1 U9233 ( .B1(n7602), .B2(n9189), .A(n7601), .ZN(P1_U3217) );
  INV_X1 U9234 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7603) );
  OAI222_X1 U9235 ( .A1(P1_U3086), .A2(n7605), .B1(n9626), .B2(n7604), .C1(
        n7603), .C2(n8213), .ZN(P1_U3334) );
  OAI21_X1 U9236 ( .B1(n7607), .B2(n8142), .A(n7606), .ZN(n9853) );
  AOI22_X1 U9237 ( .A1(n8726), .A2(n8373), .B1(n8375), .B2(n8723), .ZN(n7611)
         );
  XNOR2_X1 U9238 ( .A(n7608), .B(n8142), .ZN(n7609) );
  NAND2_X1 U9239 ( .A1(n7609), .A2(n8719), .ZN(n7610) );
  OAI211_X1 U9240 ( .C1(n9853), .C2(n7612), .A(n7611), .B(n7610), .ZN(n9854)
         );
  NAND2_X1 U9241 ( .A1(n9854), .A2(n8672), .ZN(n7616) );
  INV_X1 U9242 ( .A(n8315), .ZN(n7613) );
  OAI22_X1 U9243 ( .A1(n9668), .A2(n7028), .B1(n7613), .B2(n9656), .ZN(n7614)
         );
  AOI21_X1 U9244 ( .B1(n8710), .B2(n9856), .A(n7614), .ZN(n7615) );
  OAI211_X1 U9245 ( .C1(n9853), .C2(n8534), .A(n7616), .B(n7615), .ZN(P2_U3224) );
  XNOR2_X1 U9246 ( .A(n7617), .B(n7622), .ZN(n7620) );
  OR2_X1 U9247 ( .A1(n7863), .A2(n9167), .ZN(n7619) );
  OR2_X1 U9248 ( .A1(n7669), .A2(n9169), .ZN(n7618) );
  NAND2_X1 U9249 ( .A1(n7619), .A2(n7618), .ZN(n7766) );
  AOI21_X1 U9250 ( .B1(n7620), .B2(n9463), .A(n7766), .ZN(n9797) );
  OAI21_X1 U9251 ( .B1(n7623), .B2(n7622), .A(n7621), .ZN(n9802) );
  NAND2_X1 U9252 ( .A1(n9802), .A2(n9754), .ZN(n7631) );
  OAI22_X1 U9253 ( .A1(n9474), .A2(n7624), .B1(n7763), .B2(n9471), .ZN(n7628)
         );
  INV_X1 U9254 ( .A(n7625), .ZN(n7648) );
  INV_X1 U9255 ( .A(n7626), .ZN(n7730) );
  OAI211_X1 U9256 ( .C1(n9799), .C2(n7648), .A(n9521), .B(n7730), .ZN(n9796)
         );
  NOR2_X1 U9257 ( .A1(n9796), .A2(n9765), .ZN(n7627) );
  AOI211_X1 U9258 ( .C1(n9762), .C2(n7629), .A(n7628), .B(n7627), .ZN(n7630)
         );
  OAI211_X1 U9259 ( .C1(n9749), .C2(n9797), .A(n7631), .B(n7630), .ZN(P1_U3281) );
  XNOR2_X1 U9260 ( .A(n7632), .B(n8143), .ZN(n9857) );
  XNOR2_X1 U9261 ( .A(n7633), .B(n8143), .ZN(n7634) );
  OAI222_X1 U9262 ( .A1(n9663), .A2(n7795), .B1(n9665), .B2(n7773), .C1(n9815), 
        .C2(n7634), .ZN(n9858) );
  NAND2_X1 U9263 ( .A1(n9858), .A2(n8672), .ZN(n7639) );
  INV_X1 U9264 ( .A(n7777), .ZN(n7635) );
  OAI22_X1 U9265 ( .A1(n9668), .A2(n7636), .B1(n7635), .B2(n9656), .ZN(n7637)
         );
  AOI21_X1 U9266 ( .B1(n9860), .B2(n8710), .A(n7637), .ZN(n7638) );
  OAI211_X1 U9267 ( .C1(n9857), .C2(n8713), .A(n7639), .B(n7638), .ZN(P2_U3223) );
  OAI21_X1 U9268 ( .B1(n7641), .B2(n7643), .A(n7640), .ZN(n7660) );
  INV_X1 U9269 ( .A(n7660), .ZN(n7656) );
  XOR2_X1 U9270 ( .A(n7642), .B(n7643), .Z(n7645) );
  OAI22_X1 U9271 ( .A1(n7644), .A2(n9169), .B1(n7755), .B2(n9167), .ZN(n7676)
         );
  AOI21_X1 U9272 ( .B1(n7645), .B2(n9463), .A(n7676), .ZN(n7646) );
  OAI21_X1 U9273 ( .B1(n7656), .B2(n7647), .A(n7646), .ZN(n7658) );
  NAND2_X1 U9274 ( .A1(n7658), .A2(n9474), .ZN(n7654) );
  AOI211_X1 U9275 ( .C1(n7680), .C2(n7649), .A(n9443), .B(n7648), .ZN(n7659)
         );
  INV_X1 U9276 ( .A(n7680), .ZN(n7670) );
  NOR2_X1 U9277 ( .A1(n7670), .A2(n9444), .ZN(n7652) );
  OAI22_X1 U9278 ( .A1(n9474), .A2(n7650), .B1(n7678), .B2(n9471), .ZN(n7651)
         );
  AOI211_X1 U9279 ( .C1(n7659), .C2(n9450), .A(n7652), .B(n7651), .ZN(n7653)
         );
  OAI211_X1 U9280 ( .C1(n7656), .C2(n7655), .A(n7654), .B(n7653), .ZN(P1_U3282) );
  INV_X1 U9281 ( .A(n7657), .ZN(n9779) );
  AOI211_X1 U9282 ( .C1(n9779), .C2(n7660), .A(n7659), .B(n7658), .ZN(n7665)
         );
  INV_X1 U9283 ( .A(n9537), .ZN(n9552) );
  AOI22_X1 U9284 ( .A1(n7680), .A2(n9552), .B1(n9812), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7661) );
  OAI21_X1 U9285 ( .B1(n7665), .B2(n9812), .A(n7661), .ZN(P1_U3533) );
  INV_X1 U9286 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7662) );
  OAI22_X1 U9287 ( .A1(n7670), .A2(n9604), .B1(n9804), .B2(n7662), .ZN(n7663)
         );
  INV_X1 U9288 ( .A(n7663), .ZN(n7664) );
  OAI21_X1 U9289 ( .B1(n7665), .B2(n9619), .A(n7664), .ZN(P1_U3486) );
  AND2_X1 U9290 ( .A1(n7666), .A2(n4296), .ZN(n7667) );
  OAI22_X1 U9291 ( .A1(n7670), .A2(n9058), .B1(n7669), .B2(n9056), .ZN(n7671)
         );
  XOR2_X1 U9292 ( .A(n8978), .B(n7671), .Z(n7673) );
  AOI22_X1 U9293 ( .A1(n7680), .A2(n7593), .B1(n8988), .B2(n9208), .ZN(n7672)
         );
  NOR2_X1 U9294 ( .A1(n7673), .A2(n7672), .ZN(n7759) );
  NAND2_X1 U9295 ( .A1(n7673), .A2(n7672), .ZN(n7758) );
  INV_X1 U9296 ( .A(n7758), .ZN(n7674) );
  NOR2_X1 U9297 ( .A1(n7759), .A2(n7674), .ZN(n7675) );
  XNOR2_X1 U9298 ( .A(n4345), .B(n7675), .ZN(n7682) );
  AOI22_X1 U9299 ( .A1(n4270), .A2(n7676), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n7677) );
  OAI21_X1 U9300 ( .B1(n9157), .B2(n7678), .A(n7677), .ZN(n7679) );
  AOI21_X1 U9301 ( .B1(n7680), .B2(n4264), .A(n7679), .ZN(n7681) );
  OAI21_X1 U9302 ( .B1(n7682), .B2(n9189), .A(n7681), .ZN(P1_U3236) );
  INV_X1 U9303 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n9964) );
  NOR2_X1 U9304 ( .A1(n9964), .A2(n7685), .ZN(n7817) );
  AOI21_X1 U9305 ( .B1(n9964), .B2(n7685), .A(n7817), .ZN(n7704) );
  NAND2_X1 U9306 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n7688), .ZN(n7824) );
  OAI21_X1 U9307 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n7688), .A(n7824), .ZN(
        n7702) );
  NAND2_X1 U9308 ( .A1(n7697), .A2(n7696), .ZN(n7693) );
  INV_X1 U9309 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7689) );
  MUX2_X1 U9310 ( .A(n9964), .B(n7689), .S(n8474), .Z(n7690) );
  NAND2_X1 U9311 ( .A1(n7690), .A2(n7816), .ZN(n7834) );
  INV_X1 U9312 ( .A(n7690), .ZN(n7691) );
  NAND2_X1 U9313 ( .A1(n7691), .A2(n7823), .ZN(n7692) );
  AND2_X1 U9314 ( .A1(n7834), .A2(n7692), .ZN(n7694) );
  NAND2_X1 U9315 ( .A1(n7693), .A2(n7694), .ZN(n7835) );
  INV_X1 U9316 ( .A(n7694), .ZN(n7695) );
  NAND3_X1 U9317 ( .A1(n7697), .A2(n7696), .A3(n7695), .ZN(n7698) );
  AOI21_X1 U9318 ( .B1(n7835), .B2(n7698), .A(n8481), .ZN(n7701) );
  AND2_X1 U9319 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7951) );
  AOI21_X1 U9320 ( .B1(n7838), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n7951), .ZN(
        n7699) );
  OAI21_X1 U9321 ( .B1(n8503), .B2(n7823), .A(n7699), .ZN(n7700) );
  AOI211_X1 U9322 ( .C1(n7702), .C2(n8516), .A(n7701), .B(n7700), .ZN(n7703)
         );
  OAI21_X1 U9323 ( .B1(n7704), .B2(n8519), .A(n7703), .ZN(P2_U3195) );
  XNOR2_X1 U9324 ( .A(n7705), .B(n8145), .ZN(n9862) );
  XNOR2_X1 U9325 ( .A(n7706), .B(n8145), .ZN(n7707) );
  OAI222_X1 U9326 ( .A1(n9663), .A2(n9664), .B1(n9665), .B2(n8310), .C1(n7707), 
        .C2(n9815), .ZN(n9864) );
  NAND2_X1 U9327 ( .A1(n9864), .A2(n8672), .ZN(n7712) );
  INV_X1 U9328 ( .A(n7854), .ZN(n7708) );
  OAI22_X1 U9329 ( .A1(n9668), .A2(n7709), .B1(n7708), .B2(n9656), .ZN(n7710)
         );
  AOI21_X1 U9330 ( .B1(n9865), .B2(n8710), .A(n7710), .ZN(n7711) );
  OAI211_X1 U9331 ( .C1(n8713), .C2(n9862), .A(n7712), .B(n7711), .ZN(P2_U3222) );
  OAI21_X1 U9332 ( .B1(n4347), .B2(n4622), .A(n7713), .ZN(n9868) );
  INV_X1 U9333 ( .A(n7806), .ZN(n7714) );
  OAI22_X1 U9334 ( .A1(n9668), .A2(n7441), .B1(n7714), .B2(n9656), .ZN(n7715)
         );
  AOI21_X1 U9335 ( .B1(n9871), .B2(n8710), .A(n7715), .ZN(n7721) );
  XNOR2_X1 U9336 ( .A(n7716), .B(n4622), .ZN(n7717) );
  NAND2_X1 U9337 ( .A1(n7717), .A2(n8719), .ZN(n7719) );
  AOI22_X1 U9338 ( .A1(n8372), .A2(n8723), .B1(n8726), .B2(n8724), .ZN(n7718)
         );
  NAND2_X1 U9339 ( .A1(n7719), .A2(n7718), .ZN(n9870) );
  NAND2_X1 U9340 ( .A1(n9870), .A2(n8672), .ZN(n7720) );
  OAI211_X1 U9341 ( .C1(n9868), .C2(n8713), .A(n7721), .B(n7720), .ZN(P2_U3221) );
  INV_X1 U9342 ( .A(n7728), .ZN(n7722) );
  XNOR2_X1 U9343 ( .A(n7723), .B(n7722), .ZN(n7726) );
  OR2_X1 U9344 ( .A1(n8914), .A2(n9167), .ZN(n7725) );
  OR2_X1 U9345 ( .A1(n7755), .A2(n9169), .ZN(n7724) );
  NAND2_X1 U9346 ( .A1(n7725), .A2(n7724), .ZN(n7873) );
  AOI21_X1 U9347 ( .B1(n7726), .B2(n9463), .A(n7873), .ZN(n7736) );
  OAI21_X1 U9348 ( .B1(n7729), .B2(n7728), .A(n7727), .ZN(n7739) );
  NAND2_X1 U9349 ( .A1(n7739), .A2(n9754), .ZN(n7734) );
  OAI22_X1 U9350 ( .A1(n9474), .A2(n9231), .B1(n7870), .B2(n9471), .ZN(n7732)
         );
  OAI211_X1 U9351 ( .C1(n5478), .C2(n7626), .A(n9521), .B(n7789), .ZN(n7735)
         );
  NOR2_X1 U9352 ( .A1(n7735), .A2(n9765), .ZN(n7731) );
  AOI211_X1 U9353 ( .C1(n9762), .C2(n7861), .A(n7732), .B(n7731), .ZN(n7733)
         );
  OAI211_X1 U9354 ( .C1(n9749), .C2(n7736), .A(n7734), .B(n7733), .ZN(P1_U3280) );
  AND2_X1 U9355 ( .A1(n7736), .A2(n7735), .ZN(n7742) );
  NAND2_X1 U9356 ( .A1(n7739), .A2(n9551), .ZN(n7738) );
  AOI22_X1 U9357 ( .A1(n7861), .A2(n9552), .B1(P1_REG1_REG_13__SCAN_IN), .B2(
        n9812), .ZN(n7737) );
  OAI211_X1 U9358 ( .C1(n7742), .C2(n9812), .A(n7738), .B(n7737), .ZN(P1_U3535) );
  NAND2_X1 U9359 ( .A1(n7739), .A2(n5547), .ZN(n7741) );
  AOI22_X1 U9360 ( .A1(n7861), .A2(n6071), .B1(P1_REG0_REG_13__SCAN_IN), .B2(
        n9619), .ZN(n7740) );
  OAI211_X1 U9361 ( .C1(n7742), .C2(n9619), .A(n7741), .B(n7740), .ZN(P1_U3492) );
  INV_X1 U9362 ( .A(n7750), .ZN(n7745) );
  AOI21_X1 U9363 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9634), .A(n7743), .ZN(
        n7744) );
  OAI21_X1 U9364 ( .B1(n7745), .B2(n9626), .A(n7744), .ZN(P1_U3332) );
  INV_X1 U9365 ( .A(n7746), .ZN(n7747) );
  OAI222_X1 U9366 ( .A1(n8893), .A2(n9968), .B1(n8891), .B2(n7747), .C1(n7976), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  OAI222_X1 U9367 ( .A1(n8213), .A2(n7748), .B1(n9626), .B2(n7747), .C1(
        P1_U3086), .C2(n4682), .ZN(P1_U3333) );
  NAND2_X1 U9368 ( .A1(n7750), .A2(n7749), .ZN(n7752) );
  NAND2_X1 U9369 ( .A1(n7751), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8174) );
  OAI211_X1 U9370 ( .C1(n7753), .C2(n8893), .A(n7752), .B(n8174), .ZN(P2_U3272) );
  OAI22_X1 U9371 ( .A1(n9799), .A2(n9058), .B1(n7755), .B2(n9056), .ZN(n7754)
         );
  XNOR2_X1 U9372 ( .A(n7754), .B(n8978), .ZN(n7757) );
  OAI22_X1 U9373 ( .A1(n9799), .A2(n9056), .B1(n7755), .B2(n6689), .ZN(n7756)
         );
  NOR2_X1 U9374 ( .A1(n7757), .A2(n7756), .ZN(n7864) );
  AOI21_X1 U9375 ( .B1(n7757), .B2(n7756), .A(n7864), .ZN(n7761) );
  NAND2_X1 U9376 ( .A1(n7760), .A2(n7761), .ZN(n7866) );
  OAI21_X1 U9377 ( .B1(n7761), .B2(n7760), .A(n7866), .ZN(n7762) );
  NAND2_X1 U9378 ( .A1(n7762), .A2(n9165), .ZN(n7768) );
  NOR2_X1 U9379 ( .A1(n9186), .A2(n7763), .ZN(n7764) );
  AOI211_X1 U9380 ( .C1(n4270), .C2(n7766), .A(n7765), .B(n7764), .ZN(n7767)
         );
  OAI211_X1 U9381 ( .C1(n9799), .C2(n9147), .A(n7768), .B(n7767), .ZN(P1_U3224) );
  XOR2_X1 U9382 ( .A(n8205), .B(n9860), .Z(n7849) );
  XNOR2_X1 U9383 ( .A(n9856), .B(n8205), .ZN(n7774) );
  XNOR2_X1 U9384 ( .A(n7774), .B(n8374), .ZN(n8308) );
  XNOR2_X1 U9385 ( .A(n7848), .B(n8373), .ZN(n7850) );
  XOR2_X1 U9386 ( .A(n7849), .B(n7850), .Z(n7782) );
  AOI21_X1 U9387 ( .B1(n8361), .B2(n8374), .A(n7776), .ZN(n7779) );
  NAND2_X1 U9388 ( .A1(n8365), .A2(n7777), .ZN(n7778) );
  OAI211_X1 U9389 ( .C1(n7795), .C2(n8363), .A(n7779), .B(n7778), .ZN(n7780)
         );
  AOI21_X1 U9390 ( .B1(n9860), .B2(n8352), .A(n7780), .ZN(n7781) );
  OAI21_X1 U9391 ( .B1(n7782), .B2(n8356), .A(n7781), .ZN(P2_U3157) );
  XNOR2_X1 U9392 ( .A(n7783), .B(n7784), .ZN(n7876) );
  XNOR2_X1 U9393 ( .A(n7785), .B(n7784), .ZN(n7788) );
  OR2_X1 U9394 ( .A1(n9098), .A2(n9167), .ZN(n7787) );
  OR2_X1 U9395 ( .A1(n7863), .A2(n9169), .ZN(n7786) );
  NAND2_X1 U9396 ( .A1(n7787), .A2(n7786), .ZN(n9015) );
  AOI21_X1 U9397 ( .B1(n7788), .B2(n9463), .A(n9015), .ZN(n7884) );
  INV_X1 U9398 ( .A(n7789), .ZN(n7790) );
  OAI211_X1 U9399 ( .C1(n8915), .C2(n7790), .A(n9521), .B(n7886), .ZN(n7879)
         );
  NAND2_X1 U9400 ( .A1(n7884), .A2(n7879), .ZN(n7812) );
  OAI22_X1 U9401 ( .A1(n8915), .A2(n9537), .B1(n9811), .B2(n7791), .ZN(n7792)
         );
  AOI21_X1 U9402 ( .B1(n7812), .B2(n9811), .A(n7792), .ZN(n7793) );
  OAI21_X1 U9403 ( .B1(n7876), .B2(n9548), .A(n7793), .ZN(P1_U3536) );
  XNOR2_X1 U9404 ( .A(n7798), .B(n8205), .ZN(n7852) );
  NAND2_X1 U9405 ( .A1(n7848), .A2(n4877), .ZN(n7803) );
  NOR2_X1 U9406 ( .A1(n7795), .A2(n8205), .ZN(n7796) );
  AOI211_X1 U9407 ( .C1(n5968), .C2(n8205), .A(n7796), .B(n8145), .ZN(n7801)
         );
  NOR2_X1 U9408 ( .A1(n7797), .A2(n8205), .ZN(n7799) );
  AOI211_X1 U9409 ( .C1(n8372), .C2(n8205), .A(n7799), .B(n7798), .ZN(n7800)
         );
  XOR2_X1 U9410 ( .A(n8205), .B(n9871), .Z(n7926) );
  XNOR2_X1 U9411 ( .A(n7926), .B(n9664), .ZN(n7804) );
  XNOR2_X1 U9412 ( .A(n7927), .B(n7804), .ZN(n7811) );
  AOI21_X1 U9413 ( .B1(n8361), .B2(n8372), .A(n7805), .ZN(n7808) );
  NAND2_X1 U9414 ( .A1(n8365), .A2(n7806), .ZN(n7807) );
  OAI211_X1 U9415 ( .C1(n8242), .C2(n8363), .A(n7808), .B(n7807), .ZN(n7809)
         );
  AOI21_X1 U9416 ( .B1(n9871), .B2(n8352), .A(n7809), .ZN(n7810) );
  OAI21_X1 U9417 ( .B1(n7811), .B2(n8356), .A(n7810), .ZN(P2_U3164) );
  AOI22_X1 U9418 ( .A1(n9019), .A2(n6071), .B1(P1_REG0_REG_14__SCAN_IN), .B2(
        n9619), .ZN(n7814) );
  NAND2_X1 U9419 ( .A1(n7812), .A2(n9795), .ZN(n7813) );
  OAI211_X1 U9420 ( .C1(n7876), .C2(n9613), .A(n7814), .B(n7813), .ZN(P1_U3495) );
  NOR2_X1 U9421 ( .A1(n7816), .A2(n7815), .ZN(n7818) );
  INV_X1 U9422 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7819) );
  AOI22_X1 U9423 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8388), .B1(n8385), .B2(
        n7819), .ZN(n7820) );
  AOI21_X1 U9424 ( .B1(n7821), .B2(n7820), .A(n8384), .ZN(n7844) );
  INV_X1 U9425 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8794) );
  AOI22_X1 U9426 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8385), .B1(n8388), .B2(
        n8794), .ZN(n7827) );
  NAND2_X1 U9427 ( .A1(n7823), .A2(n7822), .ZN(n7825) );
  NAND2_X1 U9428 ( .A1(n7825), .A2(n7824), .ZN(n7826) );
  NAND2_X1 U9429 ( .A1(n7827), .A2(n7826), .ZN(n8387) );
  OAI21_X1 U9430 ( .B1(n7827), .B2(n7826), .A(n8387), .ZN(n7842) );
  NAND2_X1 U9431 ( .A1(n7835), .A2(n7834), .ZN(n7831) );
  MUX2_X1 U9432 ( .A(n7819), .B(n8794), .S(n8474), .Z(n7828) );
  NAND2_X1 U9433 ( .A1(n7828), .A2(n8388), .ZN(n8396) );
  INV_X1 U9434 ( .A(n7828), .ZN(n7829) );
  NAND2_X1 U9435 ( .A1(n7829), .A2(n8385), .ZN(n7830) );
  AND2_X1 U9436 ( .A1(n8396), .A2(n7830), .ZN(n7832) );
  NAND2_X1 U9437 ( .A1(n7831), .A2(n7832), .ZN(n8397) );
  INV_X1 U9438 ( .A(n7832), .ZN(n7833) );
  NAND3_X1 U9439 ( .A1(n7835), .A2(n7834), .A3(n7833), .ZN(n7836) );
  AOI21_X1 U9440 ( .B1(n8397), .B2(n7836), .A(n8481), .ZN(n7841) );
  INV_X1 U9441 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7837) );
  NOR2_X1 U9442 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7837), .ZN(n8240) );
  AOI21_X1 U9443 ( .B1(n7838), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n8240), .ZN(
        n7839) );
  OAI21_X1 U9444 ( .B1(n8503), .B2(n8385), .A(n7839), .ZN(n7840) );
  AOI211_X1 U9445 ( .C1(n7842), .C2(n8516), .A(n7841), .B(n7840), .ZN(n7843)
         );
  OAI21_X1 U9446 ( .B1(n7844), .B2(n8519), .A(n7843), .ZN(P2_U3196) );
  INV_X1 U9447 ( .A(n7845), .ZN(n7903) );
  AOI22_X1 U9448 ( .A1(n7846), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n9634), .ZN(n7847) );
  OAI21_X1 U9449 ( .B1(n7903), .B2(n9637), .A(n7847), .ZN(P1_U3331) );
  OAI22_X1 U9450 ( .A1(n7850), .A2(n7849), .B1(n8373), .B2(n7848), .ZN(n7851)
         );
  XOR2_X1 U9451 ( .A(n7852), .B(n7851), .Z(n7859) );
  AOI21_X1 U9452 ( .B1(n8361), .B2(n8373), .A(n7853), .ZN(n7856) );
  NAND2_X1 U9453 ( .A1(n8365), .A2(n7854), .ZN(n7855) );
  OAI211_X1 U9454 ( .C1(n9664), .C2(n8363), .A(n7856), .B(n7855), .ZN(n7857)
         );
  AOI21_X1 U9455 ( .B1(n9865), .B2(n8352), .A(n7857), .ZN(n7858) );
  OAI21_X1 U9456 ( .B1(n7859), .B2(n8356), .A(n7858), .ZN(P2_U3176) );
  NOR2_X1 U9457 ( .A1(n7863), .A2(n9056), .ZN(n7860) );
  AOI21_X1 U9458 ( .B1(n7861), .B2(n4497), .A(n7860), .ZN(n7862) );
  XNOR2_X1 U9459 ( .A(n7862), .B(n8978), .ZN(n8906) );
  OAI22_X1 U9460 ( .A1(n5478), .A2(n9056), .B1(n7863), .B2(n6689), .ZN(n8904)
         );
  XNOR2_X1 U9461 ( .A(n8906), .B(n8904), .ZN(n7868) );
  INV_X1 U9462 ( .A(n7864), .ZN(n7865) );
  NAND2_X1 U9463 ( .A1(n7866), .A2(n7865), .ZN(n7867) );
  NAND2_X1 U9464 ( .A1(n7867), .A2(n7868), .ZN(n8908) );
  OAI21_X1 U9465 ( .B1(n7868), .B2(n7867), .A(n8908), .ZN(n7869) );
  NAND2_X1 U9466 ( .A1(n7869), .A2(n9165), .ZN(n7875) );
  NAND2_X1 U9467 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9703) );
  INV_X1 U9468 ( .A(n9703), .ZN(n7872) );
  NOR2_X1 U9469 ( .A1(n9186), .A2(n7870), .ZN(n7871) );
  AOI211_X1 U9470 ( .C1(n4270), .C2(n7873), .A(n7872), .B(n7871), .ZN(n7874)
         );
  OAI211_X1 U9471 ( .C1(n5478), .C2(n9147), .A(n7875), .B(n7874), .ZN(P1_U3234) );
  INV_X1 U9472 ( .A(n7876), .ZN(n7877) );
  NAND2_X1 U9473 ( .A1(n7877), .A2(n9754), .ZN(n7883) );
  OAI22_X1 U9474 ( .A1(n9474), .A2(n7878), .B1(n9017), .B2(n9471), .ZN(n7881)
         );
  NOR2_X1 U9475 ( .A1(n7879), .A2(n9765), .ZN(n7880) );
  AOI211_X1 U9476 ( .C1(n9762), .C2(n9019), .A(n7881), .B(n7880), .ZN(n7882)
         );
  OAI211_X1 U9477 ( .C1(n9749), .C2(n7884), .A(n7883), .B(n7882), .ZN(P1_U3279) );
  XOR2_X1 U9478 ( .A(n7885), .B(n7891), .Z(n9615) );
  INV_X1 U9479 ( .A(n9615), .ZN(n7898) );
  AOI211_X1 U9480 ( .C1(n9616), .C2(n7886), .A(n9443), .B(n9476), .ZN(n9550)
         );
  NOR2_X1 U9481 ( .A1(n8919), .A2(n9444), .ZN(n7889) );
  OAI22_X1 U9482 ( .A1(n9474), .A2(n7887), .B1(n9185), .B2(n9471), .ZN(n7888)
         );
  AOI211_X1 U9483 ( .C1(n9550), .C2(n9450), .A(n7889), .B(n7888), .ZN(n7897)
         );
  XNOR2_X1 U9484 ( .A(n7891), .B(n7890), .ZN(n7895) );
  OR2_X1 U9485 ( .A1(n8914), .A2(n9169), .ZN(n7893) );
  OR2_X1 U9486 ( .A1(n9109), .A2(n9167), .ZN(n7892) );
  NAND2_X1 U9487 ( .A1(n7893), .A2(n7892), .ZN(n9183) );
  INV_X1 U9488 ( .A(n9183), .ZN(n7894) );
  OAI21_X1 U9489 ( .B1(n7895), .B2(n9412), .A(n7894), .ZN(n9549) );
  NAND2_X1 U9490 ( .A1(n9549), .A2(n9474), .ZN(n7896) );
  OAI211_X1 U9491 ( .C1(n7898), .C2(n9460), .A(n7897), .B(n7896), .ZN(P1_U3278) );
  INV_X1 U9492 ( .A(n7899), .ZN(n7905) );
  OAI222_X1 U9493 ( .A1(n7906), .A2(P1_U3086), .B1(n9626), .B2(n7905), .C1(
        n7904), .C2(n8213), .ZN(P1_U3330) );
  INV_X1 U9494 ( .A(n7907), .ZN(n7912) );
  AOI22_X1 U9495 ( .A1(n7908), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n9634), .ZN(n7909) );
  OAI21_X1 U9496 ( .B1(n7912), .B2(n9637), .A(n7909), .ZN(P1_U3329) );
  OAI222_X1 U9497 ( .A1(n8891), .A2(n7912), .B1(P2_U3151), .B2(n7911), .C1(
        n7910), .C2(n8893), .ZN(P2_U3269) );
  INV_X1 U9498 ( .A(n5946), .ZN(n9630) );
  OAI222_X1 U9499 ( .A1(n8901), .A2(n9630), .B1(n7914), .B2(P2_U3151), .C1(
        n7913), .C2(n8893), .ZN(P2_U3266) );
  NAND2_X1 U9500 ( .A1(n9405), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n7915) );
  OAI21_X1 U9501 ( .B1(n9471), .B2(n7916), .A(n7915), .ZN(n7917) );
  AOI21_X1 U9502 ( .B1(n7918), .B2(n9762), .A(n7917), .ZN(n7919) );
  OAI21_X1 U9503 ( .B1(n7920), .B2(n9765), .A(n7919), .ZN(n7921) );
  INV_X1 U9504 ( .A(n7921), .ZN(n7924) );
  NAND2_X1 U9505 ( .A1(n7922), .A2(n9457), .ZN(n7923) );
  OAI211_X1 U9506 ( .C1(n7925), .C2(n9460), .A(n7924), .B(n7923), .ZN(P1_U3356) );
  XNOR2_X1 U9507 ( .A(n8793), .B(n8205), .ZN(n7930) );
  INV_X1 U9508 ( .A(n7930), .ZN(n7931) );
  XNOR2_X1 U9509 ( .A(n9654), .B(n8205), .ZN(n7928) );
  NAND2_X1 U9510 ( .A1(n7928), .A2(n8242), .ZN(n7929) );
  OAI21_X1 U9511 ( .B1(n7928), .B2(n8242), .A(n7929), .ZN(n7950) );
  INV_X1 U9512 ( .A(n7929), .ZN(n8236) );
  XNOR2_X1 U9513 ( .A(n7930), .B(n8705), .ZN(n8235) );
  OAI21_X1 U9514 ( .B1(n7931), .B2(n8705), .A(n8234), .ZN(n8358) );
  XNOR2_X1 U9515 ( .A(n8871), .B(n8205), .ZN(n7933) );
  XNOR2_X1 U9516 ( .A(n7933), .B(n8284), .ZN(n8357) );
  XNOR2_X1 U9517 ( .A(n8699), .B(n8202), .ZN(n7932) );
  NOR2_X1 U9518 ( .A1(n7932), .A2(n8706), .ZN(n8289) );
  AOI21_X1 U9519 ( .B1(n7932), .B2(n8706), .A(n8289), .ZN(n8279) );
  INV_X1 U9520 ( .A(n7933), .ZN(n7934) );
  NAND2_X1 U9521 ( .A1(n7934), .A2(n8725), .ZN(n8280) );
  XNOR2_X1 U9522 ( .A(n8858), .B(n8205), .ZN(n7936) );
  NAND2_X1 U9523 ( .A1(n7936), .A2(n8668), .ZN(n8331) );
  INV_X1 U9524 ( .A(n7936), .ZN(n7937) );
  NAND2_X1 U9525 ( .A1(n7937), .A2(n8694), .ZN(n7938) );
  AND2_X1 U9526 ( .A1(n8331), .A2(n7938), .ZN(n8288) );
  NAND2_X1 U9527 ( .A1(n8290), .A2(n8331), .ZN(n7939) );
  XNOR2_X1 U9528 ( .A(n8779), .B(n8205), .ZN(n7940) );
  XNOR2_X1 U9529 ( .A(n7940), .B(n8655), .ZN(n8332) );
  NAND2_X1 U9530 ( .A1(n7939), .A2(n8332), .ZN(n8335) );
  NAND2_X1 U9531 ( .A1(n7940), .A2(n8683), .ZN(n7941) );
  XNOR2_X1 U9532 ( .A(n8848), .B(n8202), .ZN(n7942) );
  NAND2_X1 U9533 ( .A1(n7942), .A2(n8642), .ZN(n8255) );
  XNOR2_X1 U9534 ( .A(n7943), .B(n8205), .ZN(n8176) );
  XNOR2_X1 U9535 ( .A(n8176), .B(n8656), .ZN(n8177) );
  XOR2_X1 U9536 ( .A(n8178), .B(n8177), .Z(n7948) );
  AOI22_X1 U9537 ( .A1(n8339), .A2(n8643), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n7945) );
  NAND2_X1 U9538 ( .A1(n8365), .A2(n8646), .ZN(n7944) );
  OAI211_X1 U9539 ( .C1(n8667), .C2(n8341), .A(n7945), .B(n7944), .ZN(n7946)
         );
  AOI21_X1 U9540 ( .B1(n8842), .B2(n8352), .A(n7946), .ZN(n7947) );
  OAI21_X1 U9541 ( .B1(n7948), .B2(n8356), .A(n7947), .ZN(P2_U3173) );
  AOI21_X1 U9542 ( .B1(n7950), .B2(n7949), .A(n8237), .ZN(n7956) );
  AOI21_X1 U9543 ( .B1(n8361), .B2(n8371), .A(n7951), .ZN(n7953) );
  NAND2_X1 U9544 ( .A1(n8365), .A2(n9655), .ZN(n7952) );
  OAI211_X1 U9545 ( .C1(n9662), .C2(n8363), .A(n7953), .B(n7952), .ZN(n7954)
         );
  AOI21_X1 U9546 ( .B1(n9654), .B2(n8352), .A(n7954), .ZN(n7955) );
  OAI21_X1 U9547 ( .B1(n7956), .B2(n8356), .A(n7955), .ZN(P2_U3174) );
  NAND2_X1 U9548 ( .A1(n8537), .A2(n7958), .ZN(n8159) );
  XNOR2_X1 U9549 ( .A(n7957), .B(n8159), .ZN(n7971) );
  INV_X1 U9550 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n7961) );
  XNOR2_X1 U9551 ( .A(n7959), .B(n8159), .ZN(n7960) );
  AOI222_X1 U9552 ( .A1(n8719), .A2(n7960), .B1(n8580), .B2(n8723), .C1(n8546), 
        .C2(n8726), .ZN(n7967) );
  MUX2_X1 U9553 ( .A(n7961), .B(n7967), .S(n9873), .Z(n7963) );
  NAND2_X1 U9554 ( .A1(n8353), .A2(n8870), .ZN(n7962) );
  OAI211_X1 U9555 ( .C1(n7971), .C2(n8878), .A(n7963), .B(n7962), .ZN(P2_U3453) );
  INV_X1 U9556 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n7964) );
  MUX2_X1 U9557 ( .A(n7964), .B(n7967), .S(n9890), .Z(n7966) );
  NAND2_X1 U9558 ( .A1(n8353), .A2(n8789), .ZN(n7965) );
  OAI211_X1 U9559 ( .C1(n8796), .C2(n7971), .A(n7966), .B(n7965), .ZN(P2_U3485) );
  MUX2_X1 U9560 ( .A(n7968), .B(n7967), .S(n9668), .Z(n7970) );
  AOI22_X1 U9561 ( .A1(n8353), .A2(n8710), .B1(n8731), .B2(n8347), .ZN(n7969)
         );
  OAI211_X1 U9562 ( .C1(n7971), .C2(n8713), .A(n7970), .B(n7969), .ZN(P2_U3207) );
  INV_X1 U9563 ( .A(n7972), .ZN(n7974) );
  MUX2_X1 U9564 ( .A(n7974), .B(n7973), .S(n8110), .Z(n7975) );
  NOR2_X1 U9565 ( .A1(n8156), .A2(n7975), .ZN(n8079) );
  INV_X1 U9566 ( .A(n8622), .ZN(n8073) );
  AND2_X1 U9567 ( .A1(n7982), .A2(n7976), .ZN(n7978) );
  MUX2_X1 U9568 ( .A(n7978), .B(n7977), .S(n8125), .Z(n7986) );
  AOI21_X1 U9569 ( .B1(n7986), .B2(n7979), .A(n8051), .ZN(n7981) );
  MUX2_X1 U9570 ( .A(n7981), .B(n8051), .S(n7980), .Z(n7994) );
  NAND2_X1 U9571 ( .A1(n7983), .A2(n7982), .ZN(n7985) );
  OAI21_X1 U9572 ( .B1(n7986), .B2(n7985), .A(n7984), .ZN(n7993) );
  NAND2_X1 U9573 ( .A1(n8003), .A2(n7987), .ZN(n7990) );
  NAND2_X1 U9574 ( .A1(n7997), .A2(n7988), .ZN(n7989) );
  MUX2_X1 U9575 ( .A(n7990), .B(n7989), .S(n8110), .Z(n7991) );
  INV_X1 U9576 ( .A(n7991), .ZN(n7992) );
  OAI21_X1 U9577 ( .B1(n7994), .B2(n7993), .A(n7992), .ZN(n7996) );
  NAND2_X1 U9578 ( .A1(n7996), .A2(n7995), .ZN(n8007) );
  INV_X1 U9579 ( .A(n7997), .ZN(n7999) );
  OAI211_X1 U9580 ( .C1(n8007), .C2(n7999), .A(n8009), .B(n7998), .ZN(n8002)
         );
  AND2_X1 U9581 ( .A1(n8010), .A2(n8005), .ZN(n8001) );
  AOI21_X1 U9582 ( .B1(n8002), .B2(n8001), .A(n8000), .ZN(n8015) );
  INV_X1 U9583 ( .A(n8003), .ZN(n8006) );
  OAI211_X1 U9584 ( .C1(n8007), .C2(n8006), .A(n8005), .B(n8004), .ZN(n8013)
         );
  AND2_X1 U9585 ( .A1(n8009), .A2(n8008), .ZN(n8012) );
  INV_X1 U9586 ( .A(n8010), .ZN(n8011) );
  AOI21_X1 U9587 ( .B1(n8013), .B2(n8012), .A(n8011), .ZN(n8014) );
  MUX2_X1 U9588 ( .A(n8015), .B(n8014), .S(n8110), .Z(n8019) );
  NAND2_X1 U9589 ( .A1(n8017), .A2(n8022), .ZN(n8026) );
  NOR2_X1 U9590 ( .A1(n8026), .A2(n8138), .ZN(n8018) );
  NAND2_X1 U9591 ( .A1(n8019), .A2(n8018), .ZN(n8031) );
  AND2_X1 U9592 ( .A1(n8021), .A2(n8020), .ZN(n8023) );
  OAI211_X1 U9593 ( .C1(n8026), .C2(n8023), .A(n8022), .B(n8032), .ZN(n8028)
         );
  OAI211_X1 U9594 ( .C1(n8026), .C2(n8025), .A(n8034), .B(n8024), .ZN(n8027)
         );
  MUX2_X1 U9595 ( .A(n8028), .B(n8027), .S(n8110), .Z(n8029) );
  INV_X1 U9596 ( .A(n8029), .ZN(n8030) );
  NAND2_X1 U9597 ( .A1(n8031), .A2(n8030), .ZN(n8036) );
  NAND3_X1 U9598 ( .A1(n8036), .A2(n8032), .A3(n8037), .ZN(n8033) );
  NAND2_X1 U9599 ( .A1(n8033), .A2(n8035), .ZN(n8040) );
  NAND3_X1 U9600 ( .A1(n8036), .A2(n8035), .A3(n8034), .ZN(n8038) );
  NAND2_X1 U9601 ( .A1(n8038), .A2(n8037), .ZN(n8039) );
  MUX2_X1 U9602 ( .A(n8040), .B(n8039), .S(n8051), .Z(n8045) );
  NAND2_X1 U9603 ( .A1(n9871), .A2(n9664), .ZN(n8041) );
  MUX2_X1 U9604 ( .A(n8042), .B(n8041), .S(n8110), .Z(n8043) );
  XNOR2_X1 U9605 ( .A(n9654), .B(n8724), .ZN(n9659) );
  OAI211_X1 U9606 ( .C1(n8045), .C2(n8044), .A(n8043), .B(n9659), .ZN(n8050)
         );
  MUX2_X1 U9607 ( .A(n8047), .B(n8046), .S(n8110), .Z(n8048) );
  NOR2_X1 U9608 ( .A1(n8722), .A2(n8048), .ZN(n8049) );
  XNOR2_X1 U9609 ( .A(n8871), .B(n8725), .ZN(n8703) );
  NAND2_X1 U9610 ( .A1(n8793), .A2(n9662), .ZN(n8053) );
  MUX2_X1 U9611 ( .A(n8053), .B(n8052), .S(n8051), .Z(n8054) );
  AND2_X1 U9612 ( .A1(n8060), .A2(n8055), .ZN(n8056) );
  MUX2_X1 U9613 ( .A(n8057), .B(n8056), .S(n8110), .Z(n8058) );
  INV_X1 U9614 ( .A(n8065), .ZN(n8061) );
  NAND2_X1 U9615 ( .A1(n8067), .A2(n8059), .ZN(n8151) );
  INV_X1 U9616 ( .A(n8063), .ZN(n8064) );
  NOR2_X1 U9617 ( .A1(n8065), .A2(n8064), .ZN(n8068) );
  NAND2_X1 U9618 ( .A1(n8651), .A2(n8650), .ZN(n8130) );
  MUX2_X1 U9619 ( .A(n8071), .B(n8070), .S(n8110), .Z(n8072) );
  NAND2_X1 U9620 ( .A1(n8585), .A2(n8074), .ZN(n8075) );
  MUX2_X1 U9621 ( .A(n8076), .B(n8075), .S(n8110), .Z(n8077) );
  NAND2_X1 U9622 ( .A1(n8129), .A2(n5983), .ZN(n8082) );
  NAND2_X1 U9623 ( .A1(n8085), .A2(n8084), .ZN(n8571) );
  MUX2_X1 U9624 ( .A(n8087), .B(n8086), .S(n8110), .Z(n8088) );
  INV_X1 U9625 ( .A(n8537), .ZN(n8089) );
  MUX2_X1 U9626 ( .A(n8536), .B(n8089), .S(n8110), .Z(n8090) );
  NAND2_X1 U9627 ( .A1(n8540), .A2(n8539), .ZN(n8557) );
  INV_X1 U9628 ( .A(n8540), .ZN(n8092) );
  INV_X1 U9629 ( .A(n8539), .ZN(n8091) );
  MUX2_X1 U9630 ( .A(n8092), .B(n8091), .S(n8110), .Z(n8093) );
  MUX2_X1 U9631 ( .A(n8554), .B(n8095), .S(n8110), .Z(n8097) );
  MUX2_X1 U9632 ( .A(n8806), .B(n5943), .S(n8110), .Z(n8096) );
  OR2_X1 U9633 ( .A1(n5656), .A2(n8892), .ZN(n8100) );
  AND2_X1 U9634 ( .A1(n8105), .A2(n8118), .ZN(n8163) );
  NAND2_X1 U9635 ( .A1(n8120), .A2(n8102), .ZN(n8108) );
  INV_X1 U9636 ( .A(n8117), .ZN(n8162) );
  INV_X1 U9637 ( .A(n8105), .ZN(n8122) );
  NAND2_X1 U9638 ( .A1(n8109), .A2(n8108), .ZN(n8111) );
  NAND2_X1 U9639 ( .A1(n8882), .A2(n8113), .ZN(n8116) );
  OR2_X1 U9640 ( .A1(n5656), .A2(n8114), .ZN(n8115) );
  NOR2_X1 U9641 ( .A1(n8797), .A2(n8521), .ZN(n8127) );
  INV_X1 U9642 ( .A(n8120), .ZN(n8744) );
  NAND3_X1 U9643 ( .A1(n8121), .A2(n8521), .A3(n8744), .ZN(n8124) );
  INV_X1 U9644 ( .A(n8797), .ZN(n8741) );
  AOI22_X1 U9645 ( .A1(n8124), .A2(n8741), .B1(n8123), .B2(n8105), .ZN(n8126)
         );
  INV_X1 U9646 ( .A(n8127), .ZN(n8164) );
  INV_X1 U9647 ( .A(n8130), .ZN(n8153) );
  INV_X1 U9648 ( .A(n8703), .ZN(n8148) );
  INV_X1 U9649 ( .A(n8722), .ZN(n8734) );
  NOR2_X1 U9650 ( .A1(n8132), .A2(n8131), .ZN(n8136) );
  NOR2_X1 U9651 ( .A1(n8133), .A2(n6932), .ZN(n8135) );
  NAND4_X1 U9652 ( .A1(n8136), .A2(n8135), .A3(n9814), .A4(n8134), .ZN(n8139)
         );
  NOR3_X1 U9653 ( .A1(n8139), .A2(n8138), .A3(n8137), .ZN(n8140) );
  NAND4_X1 U9654 ( .A1(n8143), .A2(n8142), .A3(n8141), .A4(n8140), .ZN(n8144)
         );
  NOR2_X1 U9655 ( .A1(n8145), .A2(n8144), .ZN(n8146) );
  NAND4_X1 U9656 ( .A1(n8734), .A2(n8146), .A3(n4622), .A4(n9659), .ZN(n8147)
         );
  OR3_X1 U9657 ( .A1(n8149), .A2(n8148), .A3(n8147), .ZN(n8150) );
  NOR2_X1 U9658 ( .A1(n8151), .A2(n8150), .ZN(n8152) );
  NAND4_X1 U9659 ( .A1(n8639), .A2(n8153), .A3(n8653), .A4(n8152), .ZN(n8154)
         );
  OR2_X1 U9660 ( .A1(n8154), .A2(n8625), .ZN(n8155) );
  NOR2_X1 U9661 ( .A1(n8156), .A2(n8155), .ZN(n8157) );
  NAND4_X1 U9662 ( .A1(n8571), .A2(n8588), .A3(n8596), .A4(n8157), .ZN(n8158)
         );
  OR3_X1 U9663 ( .A1(n8557), .A2(n8159), .A3(n8158), .ZN(n8160) );
  NOR2_X1 U9664 ( .A1(n8544), .A2(n8160), .ZN(n8161) );
  NAND4_X1 U9665 ( .A1(n8164), .A2(n8163), .A3(n8162), .A4(n8161), .ZN(n8166)
         );
  NAND3_X1 U9666 ( .A1(n8170), .A2(n8169), .A3(n8474), .ZN(n8171) );
  OAI211_X1 U9667 ( .C1(n8172), .C2(n8174), .A(n8171), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8173) );
  OAI21_X1 U9668 ( .B1(n8175), .B2(n8174), .A(n8173), .ZN(P2_U3296) );
  XNOR2_X1 U9669 ( .A(n8179), .B(n8205), .ZN(n8180) );
  XNOR2_X1 U9670 ( .A(n8180), .B(n8181), .ZN(n8263) );
  INV_X1 U9671 ( .A(n8180), .ZN(n8182) );
  XNOR2_X1 U9672 ( .A(n5912), .B(n8205), .ZN(n8183) );
  XNOR2_X1 U9673 ( .A(n8183), .B(n8597), .ZN(n8323) );
  INV_X1 U9674 ( .A(n8183), .ZN(n8184) );
  NAND2_X1 U9675 ( .A1(n8184), .A2(n8597), .ZN(n8185) );
  XNOR2_X1 U9676 ( .A(n5984), .B(n8205), .ZN(n8187) );
  INV_X1 U9677 ( .A(n8186), .ZN(n8188) );
  XNOR2_X1 U9678 ( .A(n8822), .B(n8205), .ZN(n8191) );
  NAND2_X1 U9679 ( .A1(n8191), .A2(n8251), .ZN(n8190) );
  NAND2_X1 U9680 ( .A1(n8297), .A2(n8189), .ZN(n8271) );
  INV_X1 U9681 ( .A(n8190), .ZN(n8192) );
  XNOR2_X1 U9682 ( .A(n8191), .B(n8598), .ZN(n8300) );
  OR2_X1 U9683 ( .A1(n8192), .A2(n8300), .ZN(n8270) );
  XNOR2_X1 U9684 ( .A(n8816), .B(n8205), .ZN(n8194) );
  XNOR2_X1 U9685 ( .A(n8194), .B(n8580), .ZN(n8273) );
  AND2_X1 U9686 ( .A1(n8270), .A2(n8273), .ZN(n8193) );
  NAND2_X1 U9687 ( .A1(n8271), .A2(n8193), .ZN(n8196) );
  NAND2_X1 U9688 ( .A1(n8194), .A2(n8303), .ZN(n8195) );
  XNOR2_X1 U9689 ( .A(n8353), .B(n8202), .ZN(n8198) );
  INV_X1 U9690 ( .A(n8198), .ZN(n8199) );
  NAND2_X1 U9691 ( .A1(n8197), .A2(n8199), .ZN(n8200) );
  XNOR2_X1 U9692 ( .A(n8812), .B(n8202), .ZN(n8203) );
  NAND2_X1 U9693 ( .A1(n8203), .A2(n8546), .ZN(n8204) );
  OAI21_X1 U9694 ( .B1(n8203), .B2(n8546), .A(n8204), .ZN(n8227) );
  NOR2_X1 U9695 ( .A1(n8370), .A2(n8363), .ZN(n8209) );
  AOI22_X1 U9696 ( .A1(n8550), .A2(n8365), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8207) );
  OAI21_X1 U9697 ( .B1(n8350), .B2(n8341), .A(n8207), .ZN(n8208) );
  AOI211_X1 U9698 ( .C1(n8806), .C2(n8352), .A(n8209), .B(n8208), .ZN(n8210)
         );
  OAI222_X1 U9699 ( .A1(n8213), .A2(n8212), .B1(n9637), .B2(n8211), .C1(
        P1_U3086), .C2(n9268), .ZN(P1_U3336) );
  OAI21_X1 U9700 ( .B1(n8214), .B2(n8216), .A(n8215), .ZN(n8217) );
  NAND2_X1 U9701 ( .A1(n8217), .A2(n8336), .ZN(n8225) );
  AOI22_X1 U9702 ( .A1(n8339), .A2(n8375), .B1(n8218), .B2(n8352), .ZN(n8224)
         );
  NOR2_X1 U9703 ( .A1(n8341), .A2(n8219), .ZN(n8220) );
  AOI211_X1 U9704 ( .C1(n8222), .C2(n8365), .A(n8221), .B(n8220), .ZN(n8223)
         );
  NAND3_X1 U9705 ( .A1(n8225), .A2(n8224), .A3(n8223), .ZN(P2_U3153) );
  AOI21_X1 U9706 ( .B1(n8226), .B2(n8227), .A(n8356), .ZN(n8229) );
  NAND2_X1 U9707 ( .A1(n8229), .A2(n8228), .ZN(n8233) );
  AOI22_X1 U9708 ( .A1(n8559), .A2(n8365), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8230) );
  OAI21_X1 U9709 ( .B1(n8553), .B2(n8341), .A(n8230), .ZN(n8231) );
  AOI21_X1 U9710 ( .B1(n5943), .B2(n8339), .A(n8231), .ZN(n8232) );
  OAI211_X1 U9711 ( .C1(n8562), .C2(n8368), .A(n8233), .B(n8232), .ZN(P2_U3154) );
  INV_X1 U9712 ( .A(n8793), .ZN(n8715) );
  INV_X1 U9713 ( .A(n8234), .ZN(n8239) );
  NOR3_X1 U9714 ( .A1(n8237), .A2(n8236), .A3(n8235), .ZN(n8238) );
  OAI21_X1 U9715 ( .B1(n8239), .B2(n8238), .A(n8336), .ZN(n8245) );
  AOI21_X1 U9716 ( .B1(n8339), .B2(n8725), .A(n8240), .ZN(n8241) );
  OAI21_X1 U9717 ( .B1(n8242), .B2(n8341), .A(n8241), .ZN(n8243) );
  AOI21_X1 U9718 ( .B1(n8730), .B2(n8365), .A(n8243), .ZN(n8244) );
  OAI211_X1 U9719 ( .C1(n8715), .C2(n8368), .A(n8245), .B(n8244), .ZN(P2_U3155) );
  XNOR2_X1 U9720 ( .A(n8246), .B(n8614), .ZN(n8254) );
  INV_X1 U9721 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8247) );
  OAI22_X1 U9722 ( .A1(n8632), .A2(n8341), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8247), .ZN(n8248) );
  INV_X1 U9723 ( .A(n8248), .ZN(n8250) );
  NAND2_X1 U9724 ( .A1(n8365), .A2(n8601), .ZN(n8249) );
  OAI211_X1 U9725 ( .C1(n8251), .C2(n8363), .A(n8250), .B(n8249), .ZN(n8252)
         );
  AOI21_X1 U9726 ( .B1(n5984), .B2(n8352), .A(n8252), .ZN(n8253) );
  OAI21_X1 U9727 ( .B1(n8254), .B2(n8356), .A(n8253), .ZN(P2_U3156) );
  NAND2_X1 U9728 ( .A1(n4358), .A2(n8255), .ZN(n8256) );
  XNOR2_X1 U9729 ( .A(n8257), .B(n8256), .ZN(n8262) );
  NAND2_X1 U9730 ( .A1(n8361), .A2(n8655), .ZN(n8258) );
  NAND2_X1 U9731 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8504) );
  OAI211_X1 U9732 ( .C1(n8631), .C2(n8363), .A(n8258), .B(n8504), .ZN(n8259)
         );
  AOI21_X1 U9733 ( .B1(n8659), .B2(n8365), .A(n8259), .ZN(n8261) );
  NAND2_X1 U9734 ( .A1(n8848), .A2(n8352), .ZN(n8260) );
  OAI211_X1 U9735 ( .C1(n8262), .C2(n8356), .A(n8261), .B(n8260), .ZN(P2_U3159) );
  XOR2_X1 U9736 ( .A(n8264), .B(n8263), .Z(n8269) );
  AOI22_X1 U9737 ( .A1(n8597), .A2(n8339), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8266) );
  NAND2_X1 U9738 ( .A1(n8365), .A2(n8633), .ZN(n8265) );
  OAI211_X1 U9739 ( .C1(n8631), .C2(n8341), .A(n8266), .B(n8265), .ZN(n8267)
         );
  AOI21_X1 U9740 ( .B1(n8769), .B2(n8352), .A(n8267), .ZN(n8268) );
  OAI21_X1 U9741 ( .B1(n8269), .B2(n8356), .A(n8268), .ZN(P2_U3163) );
  AND2_X1 U9742 ( .A1(n4272), .A2(n8270), .ZN(n8272) );
  XOR2_X1 U9743 ( .A(n8273), .B(n8272), .Z(n8278) );
  AOI22_X1 U9744 ( .A1(n8598), .A2(n8361), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8275) );
  NAND2_X1 U9745 ( .A1(n8568), .A2(n8365), .ZN(n8274) );
  OAI211_X1 U9746 ( .C1(n8553), .C2(n8363), .A(n8275), .B(n8274), .ZN(n8276)
         );
  AOI21_X1 U9747 ( .B1(n8816), .B2(n8352), .A(n8276), .ZN(n8277) );
  OAI21_X1 U9748 ( .B1(n8278), .B2(n8356), .A(n8277), .ZN(P2_U3165) );
  INV_X1 U9749 ( .A(n8699), .ZN(n8864) );
  AOI21_X1 U9750 ( .B1(n8359), .B2(n8280), .A(n8279), .ZN(n8281) );
  OAI21_X1 U9751 ( .B1(n4342), .B2(n8281), .A(n8336), .ZN(n8287) );
  NOR2_X1 U9752 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8282), .ZN(n8430) );
  AOI21_X1 U9753 ( .B1(n8339), .B2(n8694), .A(n8430), .ZN(n8283) );
  OAI21_X1 U9754 ( .B1(n8284), .B2(n8341), .A(n8283), .ZN(n8285) );
  AOI21_X1 U9755 ( .B1(n8698), .B2(n8365), .A(n8285), .ZN(n8286) );
  OAI211_X1 U9756 ( .C1(n8864), .C2(n8368), .A(n8287), .B(n8286), .ZN(P2_U3166) );
  INV_X1 U9757 ( .A(n8858), .ZN(n8296) );
  NOR3_X1 U9758 ( .A1(n4342), .A2(n8289), .A3(n8288), .ZN(n8291) );
  INV_X1 U9759 ( .A(n8290), .ZN(n8334) );
  OAI21_X1 U9760 ( .B1(n8291), .B2(n8334), .A(n8336), .ZN(n8295) );
  NAND2_X1 U9761 ( .A1(n8339), .A2(n8655), .ZN(n8292) );
  NAND2_X1 U9762 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8453) );
  OAI211_X1 U9763 ( .C1(n8682), .C2(n8341), .A(n8292), .B(n8453), .ZN(n8293)
         );
  AOI21_X1 U9764 ( .B1(n8686), .B2(n8365), .A(n8293), .ZN(n8294) );
  OAI211_X1 U9765 ( .C1(n8296), .C2(n8368), .A(n8295), .B(n8294), .ZN(P2_U3168) );
  NAND2_X1 U9766 ( .A1(n8297), .A2(n8298), .ZN(n8299) );
  XOR2_X1 U9767 ( .A(n8300), .B(n8299), .Z(n8306) );
  AOI22_X1 U9768 ( .A1(n8614), .A2(n8361), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8302) );
  NAND2_X1 U9769 ( .A1(n8582), .A2(n8365), .ZN(n8301) );
  OAI211_X1 U9770 ( .C1(n8303), .C2(n8363), .A(n8302), .B(n8301), .ZN(n8304)
         );
  AOI21_X1 U9771 ( .B1(n8822), .B2(n8352), .A(n8304), .ZN(n8305) );
  OAI21_X1 U9772 ( .B1(n8306), .B2(n8356), .A(n8305), .ZN(P2_U3169) );
  OAI211_X1 U9773 ( .C1(n8309), .C2(n8308), .A(n8307), .B(n8336), .ZN(n8319)
         );
  OR2_X1 U9774 ( .A1(n8363), .A2(n8310), .ZN(n8312) );
  OAI211_X1 U9775 ( .C1(n8341), .C2(n8313), .A(n8312), .B(n8311), .ZN(n8314)
         );
  INV_X1 U9776 ( .A(n8314), .ZN(n8318) );
  NAND2_X1 U9777 ( .A1(n9856), .A2(n8352), .ZN(n8317) );
  NAND2_X1 U9778 ( .A1(n8365), .A2(n8315), .ZN(n8316) );
  NAND4_X1 U9779 ( .A1(n8319), .A2(n8318), .A3(n8317), .A4(n8316), .ZN(
        P2_U3171) );
  AND2_X1 U9780 ( .A1(n8321), .A2(n8320), .ZN(n8330) );
  OAI211_X1 U9781 ( .C1(n8324), .C2(n8323), .A(n8322), .B(n8336), .ZN(n8329)
         );
  AOI22_X1 U9782 ( .A1(n8361), .A2(n8643), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8325) );
  OAI21_X1 U9783 ( .B1(n8326), .B2(n8363), .A(n8325), .ZN(n8327) );
  AOI21_X1 U9784 ( .B1(n8617), .B2(n8365), .A(n8327), .ZN(n8328) );
  OAI211_X1 U9785 ( .C1(n8330), .C2(n8368), .A(n8329), .B(n8328), .ZN(P2_U3175) );
  INV_X1 U9786 ( .A(n8779), .ZN(n8345) );
  INV_X1 U9787 ( .A(n8331), .ZN(n8333) );
  NOR3_X1 U9788 ( .A1(n8334), .A2(n8333), .A3(n8332), .ZN(n8338) );
  INV_X1 U9789 ( .A(n8335), .ZN(n8337) );
  OAI21_X1 U9790 ( .B1(n8338), .B2(n8337), .A(n8336), .ZN(n8344) );
  NAND2_X1 U9791 ( .A1(n8339), .A2(n8642), .ZN(n8340) );
  NAND2_X1 U9792 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8479) );
  OAI211_X1 U9793 ( .C1(n8668), .C2(n8341), .A(n8340), .B(n8479), .ZN(n8342)
         );
  AOI21_X1 U9794 ( .B1(n8669), .B2(n8365), .A(n8342), .ZN(n8343) );
  OAI211_X1 U9795 ( .C1(n8345), .C2(n8368), .A(n8344), .B(n8343), .ZN(P2_U3178) );
  XNOR2_X1 U9796 ( .A(n8346), .B(n8566), .ZN(n8355) );
  AOI22_X1 U9797 ( .A1(n8580), .A2(n8361), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8349) );
  NAND2_X1 U9798 ( .A1(n8347), .A2(n8365), .ZN(n8348) );
  OAI211_X1 U9799 ( .C1(n8350), .C2(n8363), .A(n8349), .B(n8348), .ZN(n8351)
         );
  AOI21_X1 U9800 ( .B1(n8353), .B2(n8352), .A(n8351), .ZN(n8354) );
  OAI21_X1 U9801 ( .B1(n8355), .B2(n8356), .A(n8354), .ZN(P2_U3180) );
  INV_X1 U9802 ( .A(n8871), .ZN(n8369) );
  AOI21_X1 U9803 ( .B1(n8358), .B2(n8357), .A(n8356), .ZN(n8360) );
  NAND2_X1 U9804 ( .A1(n8360), .A2(n8359), .ZN(n8367) );
  AND2_X1 U9805 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8399) );
  AOI21_X1 U9806 ( .B1(n8361), .B2(n8705), .A(n8399), .ZN(n8362) );
  OAI21_X1 U9807 ( .B1(n8682), .B2(n8363), .A(n8362), .ZN(n8364) );
  AOI21_X1 U9808 ( .B1(n8709), .B2(n8365), .A(n8364), .ZN(n8366) );
  OAI211_X1 U9809 ( .C1(n8369), .C2(n8368), .A(n8367), .B(n8366), .ZN(P2_U3181) );
  INV_X1 U9810 ( .A(n8370), .ZN(n8545) );
  MUX2_X1 U9811 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8545), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9812 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n5943), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9813 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8546), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9814 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8566), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9815 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8580), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9816 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8598), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9817 ( .A(n8614), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8382), .Z(
        P2_U3514) );
  MUX2_X1 U9818 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8597), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9819 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8643), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9820 ( .A(n8656), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8382), .Z(
        P2_U3511) );
  MUX2_X1 U9821 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8642), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9822 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8655), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9823 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8694), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9824 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8706), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9825 ( .A(n8725), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8382), .Z(
        P2_U3506) );
  MUX2_X1 U9826 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8705), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U9827 ( .A(n8724), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8382), .Z(
        P2_U3504) );
  MUX2_X1 U9828 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8371), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U9829 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8372), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U9830 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8373), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U9831 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8374), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U9832 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8375), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U9833 ( .A(n8376), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8382), .Z(
        P2_U3498) );
  MUX2_X1 U9834 ( .A(n8377), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8382), .Z(
        P2_U3497) );
  MUX2_X1 U9835 ( .A(n8378), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8382), .Z(
        P2_U3496) );
  MUX2_X1 U9836 ( .A(n8379), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8382), .Z(
        P2_U3495) );
  MUX2_X1 U9837 ( .A(n8380), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8382), .Z(
        P2_U3494) );
  MUX2_X1 U9838 ( .A(n8381), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8382), .Z(
        P2_U3493) );
  MUX2_X1 U9839 ( .A(n8383), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8382), .Z(
        P2_U3492) );
  INV_X1 U9840 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8708) );
  NOR2_X1 U9841 ( .A1(n8708), .A2(n8386), .ZN(n8410) );
  AOI21_X1 U9842 ( .B1(n8708), .B2(n8386), .A(n8410), .ZN(n8407) );
  OAI21_X1 U9843 ( .B1(n8388), .B2(n8794), .A(n8387), .ZN(n8415) );
  XNOR2_X1 U9844 ( .A(n8409), .B(n8415), .ZN(n8389) );
  NAND2_X1 U9845 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8389), .ZN(n8417) );
  OAI21_X1 U9846 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n8389), .A(n8417), .ZN(
        n8405) );
  NAND2_X1 U9847 ( .A1(n8397), .A2(n8396), .ZN(n8393) );
  INV_X1 U9848 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8788) );
  MUX2_X1 U9849 ( .A(n8708), .B(n8788), .S(n8474), .Z(n8390) );
  NAND2_X1 U9850 ( .A1(n8390), .A2(n8409), .ZN(n8426) );
  INV_X1 U9851 ( .A(n8390), .ZN(n8391) );
  NAND2_X1 U9852 ( .A1(n8391), .A2(n8416), .ZN(n8392) );
  AND2_X1 U9853 ( .A1(n8426), .A2(n8392), .ZN(n8394) );
  NAND2_X1 U9854 ( .A1(n8393), .A2(n8394), .ZN(n8427) );
  INV_X1 U9855 ( .A(n8394), .ZN(n8395) );
  NAND3_X1 U9856 ( .A1(n8397), .A2(n8396), .A3(n8395), .ZN(n8398) );
  AOI21_X1 U9857 ( .B1(n8427), .B2(n8398), .A(n8481), .ZN(n8404) );
  NAND2_X1 U9858 ( .A1(n8486), .A2(n8409), .ZN(n8401) );
  INV_X1 U9859 ( .A(n8399), .ZN(n8400) );
  OAI211_X1 U9860 ( .C1(n8402), .C2(n8506), .A(n8401), .B(n8400), .ZN(n8403)
         );
  AOI211_X1 U9861 ( .C1(n8405), .C2(n8516), .A(n8404), .B(n8403), .ZN(n8406)
         );
  OAI21_X1 U9862 ( .B1(n8407), .B2(n8519), .A(n8406), .ZN(P2_U3197) );
  XNOR2_X1 U9863 ( .A(n8443), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n8414) );
  NOR2_X1 U9864 ( .A1(n8409), .A2(n8408), .ZN(n8411) );
  INV_X1 U9865 ( .A(n8440), .ZN(n8412) );
  AOI21_X1 U9866 ( .B1(n8414), .B2(n8413), .A(n8412), .ZN(n8438) );
  NAND2_X1 U9867 ( .A1(n8416), .A2(n8415), .ZN(n8418) );
  INV_X1 U9868 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9960) );
  XNOR2_X1 U9869 ( .A(n8443), .B(n9960), .ZN(n8444) );
  XNOR2_X1 U9870 ( .A(n8445), .B(n8444), .ZN(n8436) );
  NAND2_X1 U9871 ( .A1(n8427), .A2(n8426), .ZN(n8423) );
  INV_X1 U9872 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8419) );
  MUX2_X1 U9873 ( .A(n8419), .B(n9960), .S(n8474), .Z(n8420) );
  NAND2_X1 U9874 ( .A1(n8420), .A2(n8429), .ZN(n8449) );
  INV_X1 U9875 ( .A(n8420), .ZN(n8421) );
  NAND2_X1 U9876 ( .A1(n8421), .A2(n8443), .ZN(n8422) );
  AND2_X1 U9877 ( .A1(n8449), .A2(n8422), .ZN(n8424) );
  NAND2_X1 U9878 ( .A1(n8423), .A2(n8424), .ZN(n8451) );
  INV_X1 U9879 ( .A(n8424), .ZN(n8425) );
  NAND3_X1 U9880 ( .A1(n8427), .A2(n8426), .A3(n8425), .ZN(n8428) );
  AOI21_X1 U9881 ( .B1(n8451), .B2(n8428), .A(n8481), .ZN(n8435) );
  NAND2_X1 U9882 ( .A1(n8486), .A2(n8429), .ZN(n8432) );
  INV_X1 U9883 ( .A(n8430), .ZN(n8431) );
  OAI211_X1 U9884 ( .C1(n8433), .C2(n8506), .A(n8432), .B(n8431), .ZN(n8434)
         );
  AOI211_X1 U9885 ( .C1(n8436), .C2(n8516), .A(n8435), .B(n8434), .ZN(n8437)
         );
  OAI21_X1 U9886 ( .B1(n8438), .B2(n8519), .A(n8437), .ZN(P2_U3198) );
  INV_X1 U9887 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9951) );
  NAND2_X1 U9888 ( .A1(n8443), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8439) );
  NOR2_X1 U9889 ( .A1(n9951), .A2(n8442), .ZN(n8463) );
  AOI21_X1 U9890 ( .B1(n9951), .B2(n8442), .A(n8463), .ZN(n8460) );
  NAND2_X1 U9891 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n8446), .ZN(n8467) );
  OAI21_X1 U9892 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8446), .A(n8467), .ZN(
        n8458) );
  NAND2_X1 U9893 ( .A1(n8451), .A2(n8449), .ZN(n8447) );
  MUX2_X1 U9894 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8474), .Z(n8469) );
  XNOR2_X1 U9895 ( .A(n8469), .B(n8470), .ZN(n8448) );
  NAND2_X1 U9896 ( .A1(n8447), .A2(n8448), .ZN(n8473) );
  INV_X1 U9897 ( .A(n8448), .ZN(n8450) );
  NAND3_X1 U9898 ( .A1(n8451), .A2(n8450), .A3(n8449), .ZN(n8452) );
  AOI21_X1 U9899 ( .B1(n8473), .B2(n8452), .A(n8481), .ZN(n8457) );
  NAND2_X1 U9900 ( .A1(n8486), .A2(n8470), .ZN(n8454) );
  OAI211_X1 U9901 ( .C1(n8455), .C2(n8506), .A(n8454), .B(n8453), .ZN(n8456)
         );
  AOI211_X1 U9902 ( .C1(n8458), .C2(n8516), .A(n8457), .B(n8456), .ZN(n8459)
         );
  OAI21_X1 U9903 ( .B1(n8460), .B2(n8519), .A(n8459), .ZN(P2_U3199) );
  NAND2_X1 U9904 ( .A1(n8511), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8493) );
  OAI21_X1 U9905 ( .B1(n8511), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8493), .ZN(
        n8464) );
  NAND2_X1 U9906 ( .A1(n8441), .A2(n8466), .ZN(n8468) );
  NAND2_X1 U9907 ( .A1(n8468), .A2(n8467), .ZN(n8513) );
  XNOR2_X1 U9908 ( .A(n8485), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8512) );
  XNOR2_X1 U9909 ( .A(n8513), .B(n8512), .ZN(n8490) );
  INV_X1 U9910 ( .A(n8469), .ZN(n8471) );
  NAND2_X1 U9911 ( .A1(n8471), .A2(n8470), .ZN(n8472) );
  AND2_X1 U9912 ( .A1(n8473), .A2(n8472), .ZN(n8475) );
  MUX2_X1 U9913 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8474), .Z(n8476) );
  NAND2_X1 U9914 ( .A1(n8475), .A2(n8476), .ZN(n8482) );
  NAND2_X1 U9915 ( .A1(n8482), .A2(n8485), .ZN(n8497) );
  INV_X1 U9916 ( .A(n8475), .ZN(n8478) );
  INV_X1 U9917 ( .A(n8476), .ZN(n8477) );
  NAND2_X1 U9918 ( .A1(n8478), .A2(n8477), .ZN(n8496) );
  NAND2_X1 U9919 ( .A1(n8496), .A2(P2_U3893), .ZN(n8488) );
  INV_X1 U9920 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8480) );
  OAI21_X1 U9921 ( .B1(n8506), .B2(n8480), .A(n8479), .ZN(n8484) );
  AOI211_X1 U9922 ( .C1(n8482), .C2(n8496), .A(n8485), .B(n8481), .ZN(n8483)
         );
  AOI211_X1 U9923 ( .C1(n8486), .C2(n8485), .A(n8484), .B(n8483), .ZN(n8487)
         );
  OAI21_X1 U9924 ( .B1(n8497), .B2(n8488), .A(n8487), .ZN(n8489) );
  AOI21_X1 U9925 ( .B1(n8490), .B2(n8516), .A(n8489), .ZN(n8491) );
  OAI21_X1 U9926 ( .B1(n8492), .B2(n8519), .A(n8491), .ZN(P2_U3200) );
  INV_X1 U9927 ( .A(n8493), .ZN(n8494) );
  XNOR2_X1 U9928 ( .A(n8495), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8499) );
  NAND2_X1 U9929 ( .A1(n8497), .A2(n8496), .ZN(n8501) );
  XNOR2_X1 U9930 ( .A(n8502), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8514) );
  INV_X1 U9931 ( .A(n8514), .ZN(n8498) );
  MUX2_X1 U9932 ( .A(n8499), .B(n8498), .S(n8474), .Z(n8500) );
  XNOR2_X1 U9933 ( .A(n8501), .B(n8500), .ZN(n8510) );
  NOR2_X1 U9934 ( .A1(n8503), .A2(n8502), .ZN(n8508) );
  OAI21_X1 U9935 ( .B1(n8506), .B2(n8505), .A(n8504), .ZN(n8507) );
  AOI211_X1 U9936 ( .C1(n8510), .C2(n8509), .A(n8508), .B(n8507), .ZN(n8518)
         );
  AOI22_X1 U9937 ( .A1(n8513), .A2(n8512), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8511), .ZN(n8515) );
  XNOR2_X1 U9938 ( .A(n8515), .B(n8514), .ZN(n8517) );
  NAND2_X1 U9939 ( .A1(n8797), .A2(n8710), .ZN(n8523) );
  NOR2_X1 U9940 ( .A1(n8521), .A2(n8520), .ZN(n8798) );
  NOR2_X1 U9941 ( .A1(n8522), .A2(n9656), .ZN(n8531) );
  AOI21_X1 U9942 ( .B1(n8798), .B2(n8672), .A(n8531), .ZN(n8525) );
  OAI211_X1 U9943 ( .C1(n9668), .C2(n8524), .A(n8523), .B(n8525), .ZN(P2_U3202) );
  NAND2_X1 U9944 ( .A1(n8120), .A2(n8710), .ZN(n8526) );
  OAI211_X1 U9945 ( .C1(n9668), .C2(n8527), .A(n8526), .B(n8525), .ZN(P2_U3203) );
  NAND2_X1 U9946 ( .A1(n8528), .A2(n8672), .ZN(n8533) );
  NOR2_X1 U9947 ( .A1(n8529), .A2(n8561), .ZN(n8530) );
  AOI211_X1 U9948 ( .C1(n9670), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8531), .B(
        n8530), .ZN(n8532) );
  OAI211_X1 U9949 ( .C1(n8535), .C2(n8534), .A(n8533), .B(n8532), .ZN(P2_U3204) );
  OR2_X1 U9950 ( .A1(n7957), .A2(n8536), .ZN(n8538) );
  NAND2_X1 U9951 ( .A1(n8538), .A2(n8537), .ZN(n8558) );
  NAND2_X1 U9952 ( .A1(n8558), .A2(n8539), .ZN(n8541) );
  NAND2_X1 U9953 ( .A1(n8541), .A2(n8540), .ZN(n8542) );
  XOR2_X1 U9954 ( .A(n8544), .B(n8542), .Z(n8809) );
  NAND2_X1 U9955 ( .A1(n8545), .A2(n8726), .ZN(n8548) );
  NAND2_X1 U9956 ( .A1(n8546), .A2(n8723), .ZN(n8547) );
  AOI22_X1 U9957 ( .A1(n8806), .A2(n8710), .B1(n8731), .B2(n8550), .ZN(n8551)
         );
  XNOR2_X1 U9958 ( .A(n8552), .B(n4443), .ZN(n8556) );
  OAI22_X1 U9959 ( .A1(n8554), .A2(n9663), .B1(n8553), .B2(n9665), .ZN(n8555)
         );
  AOI21_X1 U9960 ( .B1(n8556), .B2(n8719), .A(n8555), .ZN(n8753) );
  XNOR2_X1 U9961 ( .A(n8558), .B(n8557), .ZN(n8751) );
  AOI22_X1 U9962 ( .A1(n8559), .A2(n8731), .B1(n9670), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8560) );
  OAI21_X1 U9963 ( .B1(n8562), .B2(n8561), .A(n8560), .ZN(n8563) );
  AOI21_X1 U9964 ( .B1(n8751), .B2(n8736), .A(n8563), .ZN(n8564) );
  OAI21_X1 U9965 ( .B1(n8753), .B2(n9670), .A(n8564), .ZN(P2_U3206) );
  XNOR2_X1 U9966 ( .A(n8565), .B(n8571), .ZN(n8567) );
  AOI222_X1 U9967 ( .A1(n8719), .A2(n8567), .B1(n8598), .B2(n8723), .C1(n8566), 
        .C2(n8726), .ZN(n8814) );
  AOI22_X1 U9968 ( .A1(n8816), .A2(n8583), .B1(n8731), .B2(n8568), .ZN(n8569)
         );
  AOI21_X1 U9969 ( .B1(n8814), .B2(n8569), .A(n9670), .ZN(n8574) );
  XNOR2_X1 U9970 ( .A(n8570), .B(n8571), .ZN(n8819) );
  OAI22_X1 U9971 ( .A1(n8819), .A2(n8713), .B1(n8572), .B2(n8672), .ZN(n8573)
         );
  OR2_X1 U9972 ( .A1(n8574), .A2(n8573), .ZN(P2_U3208) );
  NOR2_X1 U9973 ( .A1(n8575), .A2(n8576), .ZN(n8578) );
  OR2_X1 U9974 ( .A1(n8578), .A2(n8577), .ZN(n8579) );
  XOR2_X1 U9975 ( .A(n8588), .B(n8579), .Z(n8581) );
  AOI222_X1 U9976 ( .A1(n8719), .A2(n8581), .B1(n8580), .B2(n8726), .C1(n8614), 
        .C2(n8723), .ZN(n8820) );
  AOI22_X1 U9977 ( .A1(n8822), .A2(n8583), .B1(n8731), .B2(n8582), .ZN(n8584)
         );
  AOI21_X1 U9978 ( .B1(n8820), .B2(n8584), .A(n9670), .ZN(n8591) );
  NAND2_X1 U9979 ( .A1(n8586), .A2(n8585), .ZN(n8587) );
  XOR2_X1 U9980 ( .A(n8588), .B(n8587), .Z(n8825) );
  OAI22_X1 U9981 ( .A1(n8825), .A2(n8713), .B1(n8589), .B2(n8672), .ZN(n8590)
         );
  OR2_X1 U9982 ( .A1(n8591), .A2(n8590), .ZN(P2_U3209) );
  XNOR2_X1 U9983 ( .A(n8592), .B(n8596), .ZN(n8830) );
  NOR2_X1 U9984 ( .A1(n8575), .A2(n8604), .ZN(n8594) );
  OR2_X1 U9985 ( .A1(n8594), .A2(n8593), .ZN(n8595) );
  XOR2_X1 U9986 ( .A(n8596), .B(n8595), .Z(n8599) );
  AOI222_X1 U9987 ( .A1(n8719), .A2(n8599), .B1(n8598), .B2(n8726), .C1(n8597), 
        .C2(n8723), .ZN(n8826) );
  MUX2_X1 U9988 ( .A(n8600), .B(n8826), .S(n9668), .Z(n8603) );
  AOI22_X1 U9989 ( .A1(n5984), .A2(n8710), .B1(n8731), .B2(n8601), .ZN(n8602)
         );
  OAI211_X1 U9990 ( .C1(n8830), .C2(n8713), .A(n8603), .B(n8602), .ZN(P2_U3210) );
  XOR2_X1 U9991 ( .A(n4354), .B(n8156), .Z(n8835) );
  OR2_X1 U9992 ( .A1(n8575), .A2(n8604), .ZN(n8605) );
  AND2_X1 U9993 ( .A1(n8606), .A2(n8605), .ZN(n8613) );
  OR2_X1 U9994 ( .A1(n8575), .A2(n8607), .ZN(n8609) );
  AND2_X1 U9995 ( .A1(n8609), .A2(n8608), .ZN(n8629) );
  NAND3_X1 U9996 ( .A1(n8629), .A2(n8611), .A3(n8610), .ZN(n8612) );
  NAND2_X1 U9997 ( .A1(n8613), .A2(n8612), .ZN(n8615) );
  AOI222_X1 U9998 ( .A1(n8719), .A2(n8615), .B1(n8614), .B2(n8726), .C1(n8643), 
        .C2(n8723), .ZN(n8831) );
  MUX2_X1 U9999 ( .A(n8616), .B(n8831), .S(n9668), .Z(n8619) );
  AOI22_X1 U10000 ( .A1(n5912), .A2(n8710), .B1(n8731), .B2(n8617), .ZN(n8618)
         );
  OAI211_X1 U10001 ( .C1(n8835), .C2(n8713), .A(n8619), .B(n8618), .ZN(
        P2_U3211) );
  NAND2_X1 U10002 ( .A1(n8620), .A2(n8621), .ZN(n8623) );
  NAND2_X1 U10003 ( .A1(n8623), .A2(n8622), .ZN(n8624) );
  XNOR2_X1 U10004 ( .A(n8625), .B(n8624), .ZN(n8839) );
  NAND3_X1 U10005 ( .A1(n8640), .A2(n8627), .A3(n8626), .ZN(n8628) );
  AND2_X1 U10006 ( .A1(n8629), .A2(n8628), .ZN(n8630) );
  OAI222_X1 U10007 ( .A1(n9663), .A2(n8632), .B1(n9665), .B2(n8631), .C1(n9815), .C2(n8630), .ZN(n8768) );
  NAND2_X1 U10008 ( .A1(n8768), .A2(n8672), .ZN(n8638) );
  INV_X1 U10009 ( .A(n8633), .ZN(n8635) );
  OAI22_X1 U10010 ( .A1(n8635), .A2(n9656), .B1(n9668), .B2(n8634), .ZN(n8636)
         );
  AOI21_X1 U10011 ( .B1(n8769), .B2(n8710), .A(n8636), .ZN(n8637) );
  OAI211_X1 U10012 ( .C1(n8839), .C2(n8713), .A(n8638), .B(n8637), .ZN(
        P2_U3212) );
  XOR2_X1 U10013 ( .A(n8620), .B(n8639), .Z(n8845) );
  INV_X1 U10014 ( .A(n8639), .ZN(n8641) );
  OAI21_X1 U10015 ( .B1(n4477), .B2(n8641), .A(n8640), .ZN(n8644) );
  AOI222_X1 U10016 ( .A1(n8719), .A2(n8644), .B1(n8643), .B2(n8726), .C1(n8642), .C2(n8723), .ZN(n8840) );
  MUX2_X1 U10017 ( .A(n8645), .B(n8840), .S(n9668), .Z(n8648) );
  AOI22_X1 U10018 ( .A1(n8842), .A2(n8710), .B1(n8731), .B2(n8646), .ZN(n8647)
         );
  OAI211_X1 U10019 ( .C1(n8845), .C2(n8713), .A(n8648), .B(n8647), .ZN(
        P2_U3213) );
  NAND2_X1 U10020 ( .A1(n8676), .A2(n8650), .ZN(n8663) );
  NAND2_X1 U10021 ( .A1(n8663), .A2(n8664), .ZN(n8662) );
  NAND2_X1 U10022 ( .A1(n8662), .A2(n8651), .ZN(n8652) );
  XNOR2_X1 U10023 ( .A(n8652), .B(n8653), .ZN(n8851) );
  INV_X1 U10024 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8658) );
  XNOR2_X1 U10025 ( .A(n8654), .B(n8653), .ZN(n8657) );
  AOI222_X1 U10026 ( .A1(n8719), .A2(n8657), .B1(n8656), .B2(n8726), .C1(n8655), .C2(n8723), .ZN(n8846) );
  MUX2_X1 U10027 ( .A(n8658), .B(n8846), .S(n9668), .Z(n8661) );
  AOI22_X1 U10028 ( .A1(n8848), .A2(n8710), .B1(n8731), .B2(n8659), .ZN(n8660)
         );
  OAI211_X1 U10029 ( .C1(n8851), .C2(n8713), .A(n8661), .B(n8660), .ZN(
        P2_U3214) );
  OAI21_X1 U10030 ( .B1(n8663), .B2(n8664), .A(n8662), .ZN(n8855) );
  XOR2_X1 U10031 ( .A(n8665), .B(n8664), .Z(n8666) );
  OAI222_X1 U10032 ( .A1(n9665), .A2(n8668), .B1(n9663), .B2(n8667), .C1(n8666), .C2(n9815), .ZN(n8778) );
  NAND2_X1 U10033 ( .A1(n8778), .A2(n8672), .ZN(n8675) );
  INV_X1 U10034 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8671) );
  INV_X1 U10035 ( .A(n8669), .ZN(n8670) );
  OAI22_X1 U10036 ( .A1(n8672), .A2(n8671), .B1(n8670), .B2(n9656), .ZN(n8673)
         );
  AOI21_X1 U10037 ( .B1(n8779), .B2(n8710), .A(n8673), .ZN(n8674) );
  OAI211_X1 U10038 ( .C1(n8855), .C2(n8713), .A(n8675), .B(n8674), .ZN(
        P2_U3215) );
  OAI21_X1 U10039 ( .B1(n8677), .B2(n8679), .A(n8676), .ZN(n8861) );
  NAND3_X1 U10040 ( .A1(n8693), .A2(n8679), .A3(n8678), .ZN(n8680) );
  AND3_X1 U10041 ( .A1(n8681), .A2(n8719), .A3(n8680), .ZN(n8685) );
  OAI22_X1 U10042 ( .A1(n8683), .A2(n9663), .B1(n8682), .B2(n9665), .ZN(n8684)
         );
  NOR2_X1 U10043 ( .A1(n8685), .A2(n8684), .ZN(n8856) );
  MUX2_X1 U10044 ( .A(n9951), .B(n8856), .S(n9668), .Z(n8688) );
  AOI22_X1 U10045 ( .A1(n8858), .A2(n8710), .B1(n8731), .B2(n8686), .ZN(n8687)
         );
  OAI211_X1 U10046 ( .C1(n8861), .C2(n8713), .A(n8688), .B(n8687), .ZN(
        P2_U3216) );
  XNOR2_X1 U10047 ( .A(n8689), .B(n8690), .ZN(n8865) );
  NAND2_X1 U10048 ( .A1(n8691), .A2(n8690), .ZN(n8692) );
  NAND3_X1 U10049 ( .A1(n8693), .A2(n8719), .A3(n8692), .ZN(n8696) );
  AOI22_X1 U10050 ( .A1(n8694), .A2(n8726), .B1(n8723), .B2(n8725), .ZN(n8695)
         );
  NAND2_X1 U10051 ( .A1(n8696), .A2(n8695), .ZN(n8862) );
  MUX2_X1 U10052 ( .A(n8862), .B(P2_REG2_REG_16__SCAN_IN), .S(n9670), .Z(n8697) );
  INV_X1 U10053 ( .A(n8697), .ZN(n8701) );
  AOI22_X1 U10054 ( .A1(n8699), .A2(n8710), .B1(n8731), .B2(n8698), .ZN(n8700)
         );
  OAI211_X1 U10055 ( .C1(n8865), .C2(n8713), .A(n8701), .B(n8700), .ZN(
        P2_U3217) );
  XNOR2_X1 U10056 ( .A(n8702), .B(n8703), .ZN(n8874) );
  XNOR2_X1 U10057 ( .A(n8704), .B(n8703), .ZN(n8707) );
  AOI222_X1 U10058 ( .A1(n8719), .A2(n8707), .B1(n8706), .B2(n8726), .C1(n8705), .C2(n8723), .ZN(n8868) );
  MUX2_X1 U10059 ( .A(n8708), .B(n8868), .S(n9668), .Z(n8712) );
  AOI22_X1 U10060 ( .A1(n8871), .A2(n8710), .B1(n8731), .B2(n8709), .ZN(n8711)
         );
  OAI211_X1 U10061 ( .C1(n8874), .C2(n8713), .A(n8712), .B(n8711), .ZN(
        P2_U3218) );
  NOR2_X1 U10062 ( .A1(n8715), .A2(n8714), .ZN(n8729) );
  INV_X1 U10063 ( .A(n8716), .ZN(n8718) );
  NAND2_X1 U10064 ( .A1(n8718), .A2(n8717), .ZN(n8720) );
  OAI211_X1 U10065 ( .C1(n8722), .C2(n8721), .A(n8720), .B(n8719), .ZN(n8728)
         );
  AOI22_X1 U10066 ( .A1(n8726), .A2(n8725), .B1(n8724), .B2(n8723), .ZN(n8727)
         );
  NAND2_X1 U10067 ( .A1(n8728), .A2(n8727), .ZN(n8792) );
  AOI211_X1 U10068 ( .C1(n8731), .C2(n8730), .A(n8729), .B(n8792), .ZN(n8739)
         );
  INV_X1 U10069 ( .A(n8732), .ZN(n8735) );
  OAI21_X1 U10070 ( .B1(n8735), .B2(n8734), .A(n8733), .ZN(n8879) );
  INV_X1 U10071 ( .A(n8879), .ZN(n8737) );
  AOI22_X1 U10072 ( .A1(n8737), .A2(n8736), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n9670), .ZN(n8738) );
  OAI21_X1 U10073 ( .B1(n8739), .B2(n9670), .A(n8738), .ZN(P2_U3219) );
  NAND2_X1 U10074 ( .A1(n8798), .A2(n9890), .ZN(n8742) );
  NAND2_X1 U10075 ( .A1(n8746), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8740) );
  OAI211_X1 U10076 ( .C1(n8741), .C2(n8785), .A(n8742), .B(n8740), .ZN(
        P2_U3490) );
  NAND2_X1 U10077 ( .A1(n8746), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8743) );
  OAI211_X1 U10078 ( .C1(n8744), .C2(n8785), .A(n8743), .B(n8742), .ZN(
        P2_U3489) );
  INV_X1 U10079 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8745) );
  NAND2_X1 U10080 ( .A1(n8806), .A2(n8789), .ZN(n8749) );
  OAI211_X1 U10081 ( .C1(n8809), .C2(n8796), .A(n8750), .B(n8749), .ZN(
        P2_U3487) );
  NAND2_X1 U10082 ( .A1(n8751), .A2(n9835), .ZN(n8752) );
  NAND2_X1 U10083 ( .A1(n8753), .A2(n8752), .ZN(n8810) );
  MUX2_X1 U10084 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8810), .S(n9890), .Z(n8754) );
  AOI21_X1 U10085 ( .B1(n8789), .B2(n8812), .A(n8754), .ZN(n8755) );
  INV_X1 U10086 ( .A(n8755), .ZN(P2_U3486) );
  INV_X1 U10087 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8756) );
  MUX2_X1 U10088 ( .A(n8756), .B(n8814), .S(n9890), .Z(n8758) );
  NAND2_X1 U10089 ( .A1(n8816), .A2(n8789), .ZN(n8757) );
  OAI211_X1 U10090 ( .C1(n8796), .C2(n8819), .A(n8758), .B(n8757), .ZN(
        P2_U3484) );
  INV_X1 U10091 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8759) );
  MUX2_X1 U10092 ( .A(n8759), .B(n8820), .S(n9890), .Z(n8761) );
  NAND2_X1 U10093 ( .A1(n8822), .A2(n8789), .ZN(n8760) );
  OAI211_X1 U10094 ( .C1(n8796), .C2(n8825), .A(n8761), .B(n8760), .ZN(
        P2_U3483) );
  INV_X1 U10095 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8762) );
  MUX2_X1 U10096 ( .A(n8762), .B(n8826), .S(n9890), .Z(n8764) );
  NAND2_X1 U10097 ( .A1(n5984), .A2(n8789), .ZN(n8763) );
  OAI211_X1 U10098 ( .C1(n8830), .C2(n8796), .A(n8764), .B(n8763), .ZN(
        P2_U3482) );
  INV_X1 U10099 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8765) );
  MUX2_X1 U10100 ( .A(n8765), .B(n8831), .S(n9890), .Z(n8767) );
  NAND2_X1 U10101 ( .A1(n5912), .A2(n8789), .ZN(n8766) );
  OAI211_X1 U10102 ( .C1(n8835), .C2(n8796), .A(n8767), .B(n8766), .ZN(
        P2_U3481) );
  INV_X1 U10103 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8770) );
  AOI21_X1 U10104 ( .B1(n9872), .B2(n8769), .A(n8768), .ZN(n8836) );
  MUX2_X1 U10105 ( .A(n8770), .B(n8836), .S(n9890), .Z(n8771) );
  OAI21_X1 U10106 ( .B1(n8796), .B2(n8839), .A(n8771), .ZN(P2_U3480) );
  INV_X1 U10107 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8772) );
  MUX2_X1 U10108 ( .A(n8772), .B(n8840), .S(n9890), .Z(n8774) );
  NAND2_X1 U10109 ( .A1(n8842), .A2(n8789), .ZN(n8773) );
  OAI211_X1 U10110 ( .C1(n8796), .C2(n8845), .A(n8774), .B(n8773), .ZN(
        P2_U3479) );
  INV_X1 U10111 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8775) );
  MUX2_X1 U10112 ( .A(n8775), .B(n8846), .S(n9890), .Z(n8777) );
  NAND2_X1 U10113 ( .A1(n8848), .A2(n8789), .ZN(n8776) );
  OAI211_X1 U10114 ( .C1(n8851), .C2(n8796), .A(n8777), .B(n8776), .ZN(
        P2_U3478) );
  INV_X1 U10115 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8780) );
  AOI21_X1 U10116 ( .B1(n9872), .B2(n8779), .A(n8778), .ZN(n8852) );
  MUX2_X1 U10117 ( .A(n8780), .B(n8852), .S(n9890), .Z(n8781) );
  OAI21_X1 U10118 ( .B1(n8796), .B2(n8855), .A(n8781), .ZN(P2_U3477) );
  INV_X1 U10119 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8782) );
  MUX2_X1 U10120 ( .A(n8782), .B(n8856), .S(n9890), .Z(n8784) );
  NAND2_X1 U10121 ( .A1(n8858), .A2(n8789), .ZN(n8783) );
  OAI211_X1 U10122 ( .C1(n8796), .C2(n8861), .A(n8784), .B(n8783), .ZN(
        P2_U3476) );
  MUX2_X1 U10123 ( .A(n8862), .B(P2_REG1_REG_16__SCAN_IN), .S(n8746), .Z(n8787) );
  OAI22_X1 U10124 ( .A1(n8865), .A2(n8796), .B1(n8864), .B2(n8785), .ZN(n8786)
         );
  OR2_X1 U10125 ( .A1(n8787), .A2(n8786), .ZN(P2_U3475) );
  MUX2_X1 U10126 ( .A(n8788), .B(n8868), .S(n9890), .Z(n8791) );
  NAND2_X1 U10127 ( .A1(n8871), .A2(n8789), .ZN(n8790) );
  OAI211_X1 U10128 ( .C1(n8796), .C2(n8874), .A(n8791), .B(n8790), .ZN(
        P2_U3474) );
  AOI21_X1 U10129 ( .B1(n9872), .B2(n8793), .A(n8792), .ZN(n8875) );
  MUX2_X1 U10130 ( .A(n8794), .B(n8875), .S(n9890), .Z(n8795) );
  OAI21_X1 U10131 ( .B1(n8796), .B2(n8879), .A(n8795), .ZN(P2_U3473) );
  INV_X1 U10132 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8800) );
  NAND2_X1 U10133 ( .A1(n8797), .A2(n8870), .ZN(n8799) );
  NAND2_X1 U10134 ( .A1(n8798), .A2(n9873), .ZN(n8801) );
  OAI211_X1 U10135 ( .C1(n8800), .C2(n9873), .A(n8799), .B(n8801), .ZN(
        P2_U3458) );
  INV_X1 U10136 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8803) );
  NAND2_X1 U10137 ( .A1(n8120), .A2(n8870), .ZN(n8802) );
  OAI211_X1 U10138 ( .C1(n8803), .C2(n9873), .A(n8802), .B(n8801), .ZN(
        P2_U3457) );
  INV_X1 U10139 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8805) );
  MUX2_X1 U10140 ( .A(n8805), .B(n8804), .S(n9873), .Z(n8808) );
  NAND2_X1 U10141 ( .A1(n8806), .A2(n8870), .ZN(n8807) );
  OAI211_X1 U10142 ( .C1(n8809), .C2(n8878), .A(n8808), .B(n8807), .ZN(
        P2_U3455) );
  MUX2_X1 U10143 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8810), .S(n9873), .Z(n8811) );
  AOI21_X1 U10144 ( .B1(n8870), .B2(n8812), .A(n8811), .ZN(n8813) );
  INV_X1 U10145 ( .A(n8813), .ZN(P2_U3454) );
  INV_X1 U10146 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8815) );
  MUX2_X1 U10147 ( .A(n8815), .B(n8814), .S(n9873), .Z(n8818) );
  NAND2_X1 U10148 ( .A1(n8816), .A2(n8870), .ZN(n8817) );
  OAI211_X1 U10149 ( .C1(n8819), .C2(n8878), .A(n8818), .B(n8817), .ZN(
        P2_U3452) );
  INV_X1 U10150 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8821) );
  MUX2_X1 U10151 ( .A(n8821), .B(n8820), .S(n9873), .Z(n8824) );
  NAND2_X1 U10152 ( .A1(n8822), .A2(n8870), .ZN(n8823) );
  OAI211_X1 U10153 ( .C1(n8825), .C2(n8878), .A(n8824), .B(n8823), .ZN(
        P2_U3451) );
  INV_X1 U10154 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8827) );
  MUX2_X1 U10155 ( .A(n8827), .B(n8826), .S(n9873), .Z(n8829) );
  NAND2_X1 U10156 ( .A1(n5984), .A2(n8870), .ZN(n8828) );
  OAI211_X1 U10157 ( .C1(n8830), .C2(n8878), .A(n8829), .B(n8828), .ZN(
        P2_U3450) );
  INV_X1 U10158 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8832) );
  MUX2_X1 U10159 ( .A(n8832), .B(n8831), .S(n9873), .Z(n8834) );
  NAND2_X1 U10160 ( .A1(n5912), .A2(n8870), .ZN(n8833) );
  OAI211_X1 U10161 ( .C1(n8835), .C2(n8878), .A(n8834), .B(n8833), .ZN(
        P2_U3449) );
  INV_X1 U10162 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8837) );
  MUX2_X1 U10163 ( .A(n8837), .B(n8836), .S(n9873), .Z(n8838) );
  OAI21_X1 U10164 ( .B1(n8839), .B2(n8878), .A(n8838), .ZN(P2_U3448) );
  INV_X1 U10165 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8841) );
  MUX2_X1 U10166 ( .A(n8841), .B(n8840), .S(n9873), .Z(n8844) );
  NAND2_X1 U10167 ( .A1(n8842), .A2(n8870), .ZN(n8843) );
  OAI211_X1 U10168 ( .C1(n8845), .C2(n8878), .A(n8844), .B(n8843), .ZN(
        P2_U3447) );
  INV_X1 U10169 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8847) );
  MUX2_X1 U10170 ( .A(n8847), .B(n8846), .S(n9873), .Z(n8850) );
  NAND2_X1 U10171 ( .A1(n8848), .A2(n8870), .ZN(n8849) );
  OAI211_X1 U10172 ( .C1(n8851), .C2(n8878), .A(n8850), .B(n8849), .ZN(
        P2_U3446) );
  INV_X1 U10173 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8853) );
  MUX2_X1 U10174 ( .A(n8853), .B(n8852), .S(n9873), .Z(n8854) );
  OAI21_X1 U10175 ( .B1(n8855), .B2(n8878), .A(n8854), .ZN(P2_U3444) );
  INV_X1 U10176 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8857) );
  MUX2_X1 U10177 ( .A(n8857), .B(n8856), .S(n9873), .Z(n8860) );
  NAND2_X1 U10178 ( .A1(n8858), .A2(n8870), .ZN(n8859) );
  OAI211_X1 U10179 ( .C1(n8861), .C2(n8878), .A(n8860), .B(n8859), .ZN(
        P2_U3441) );
  MUX2_X1 U10180 ( .A(n8862), .B(P2_REG0_REG_16__SCAN_IN), .S(n9875), .Z(n8867) );
  OAI22_X1 U10181 ( .A1(n8865), .A2(n8878), .B1(n8864), .B2(n8863), .ZN(n8866)
         );
  OR2_X1 U10182 ( .A1(n8867), .A2(n8866), .ZN(P2_U3438) );
  INV_X1 U10183 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8869) );
  MUX2_X1 U10184 ( .A(n8869), .B(n8868), .S(n9873), .Z(n8873) );
  NAND2_X1 U10185 ( .A1(n8871), .A2(n8870), .ZN(n8872) );
  OAI211_X1 U10186 ( .C1(n8874), .C2(n8878), .A(n8873), .B(n8872), .ZN(
        P2_U3435) );
  INV_X1 U10187 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8876) );
  MUX2_X1 U10188 ( .A(n8876), .B(n8875), .S(n9873), .Z(n8877) );
  OAI21_X1 U10189 ( .B1(n8879), .B2(n8878), .A(n8877), .ZN(P2_U3432) );
  MUX2_X1 U10190 ( .A(P2_D_REG_1__SCAN_IN), .B(n8881), .S(n8880), .Z(P2_U3377)
         );
  INV_X1 U10191 ( .A(n8882), .ZN(n9624) );
  INV_X1 U10192 ( .A(n8883), .ZN(n8886) );
  NOR4_X1 U10193 ( .A1(n8886), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n8884), .ZN(n8887) );
  AOI21_X1 U10194 ( .B1(n8899), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8887), .ZN(
        n8888) );
  OAI21_X1 U10195 ( .B1(n9624), .B2(n8891), .A(n8888), .ZN(P2_U3264) );
  INV_X1 U10196 ( .A(n8889), .ZN(n9627) );
  OAI222_X1 U10197 ( .A1(n8893), .A2(n8892), .B1(n8891), .B2(n9627), .C1(
        P2_U3151), .C2(n8890), .ZN(P2_U3265) );
  INV_X1 U10198 ( .A(n8894), .ZN(n9633) );
  AOI21_X1 U10199 ( .B1(n8899), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8895), .ZN(
        n8896) );
  OAI21_X1 U10200 ( .B1(n9633), .B2(n8901), .A(n8896), .ZN(P2_U3267) );
  INV_X1 U10201 ( .A(n8897), .ZN(n9638) );
  AOI21_X1 U10202 ( .B1(n8899), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n8898), .ZN(
        n8900) );
  OAI21_X1 U10203 ( .B1(n9638), .B2(n8901), .A(n8900), .ZN(P2_U3268) );
  INV_X1 U10204 ( .A(n8902), .ZN(n8903) );
  MUX2_X1 U10205 ( .A(n8903), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10206 ( .A(n8904), .ZN(n8905) );
  NAND2_X1 U10207 ( .A1(n8906), .A2(n8905), .ZN(n8907) );
  NAND2_X1 U10208 ( .A1(n8908), .A2(n8907), .ZN(n8910) );
  OAI22_X1 U10209 ( .A1(n8915), .A2(n9058), .B1(n8914), .B2(n9056), .ZN(n8909)
         );
  XOR2_X1 U10210 ( .A(n6532), .B(n8909), .Z(n8911) );
  INV_X1 U10211 ( .A(n8910), .ZN(n8913) );
  INV_X1 U10212 ( .A(n8911), .ZN(n8912) );
  OAI22_X1 U10213 ( .A1(n8915), .A2(n9056), .B1(n8914), .B2(n6689), .ZN(n9014)
         );
  OAI22_X1 U10214 ( .A1(n8919), .A2(n9058), .B1(n9098), .B2(n9056), .ZN(n8916)
         );
  XOR2_X1 U10215 ( .A(n6532), .B(n8916), .Z(n8917) );
  INV_X1 U10216 ( .A(n8917), .ZN(n8918) );
  OAI22_X1 U10217 ( .A1(n8919), .A2(n9056), .B1(n9098), .B2(n6689), .ZN(n9180)
         );
  NAND2_X1 U10218 ( .A1(n9178), .A2(n8920), .ZN(n9094) );
  OAI22_X1 U10219 ( .A1(n9477), .A2(n9056), .B1(n9109), .B2(n6689), .ZN(n8924)
         );
  NAND2_X1 U10220 ( .A1(n5476), .A2(n4497), .ZN(n8922) );
  OR2_X1 U10221 ( .A1(n9109), .A2(n9056), .ZN(n8921) );
  NAND2_X1 U10222 ( .A1(n8922), .A2(n8921), .ZN(n8923) );
  XNOR2_X1 U10223 ( .A(n8923), .B(n8978), .ZN(n8925) );
  XOR2_X1 U10224 ( .A(n8924), .B(n8925), .Z(n9096) );
  NAND2_X1 U10225 ( .A1(n9540), .A2(n4497), .ZN(n8928) );
  OR2_X1 U10226 ( .A1(n9154), .A2(n9056), .ZN(n8927) );
  NAND2_X1 U10227 ( .A1(n8928), .A2(n8927), .ZN(n8929) );
  XNOR2_X1 U10228 ( .A(n8929), .B(n6687), .ZN(n8932) );
  NOR2_X1 U10229 ( .A1(n9154), .A2(n6689), .ZN(n8930) );
  AOI21_X1 U10230 ( .B1(n9540), .B2(n7593), .A(n8930), .ZN(n8931) );
  OR2_X1 U10231 ( .A1(n8932), .A2(n8931), .ZN(n9107) );
  NAND2_X1 U10232 ( .A1(n8932), .A2(n8931), .ZN(n9106) );
  OAI22_X1 U10233 ( .A1(n9605), .A2(n9058), .B1(n9110), .B2(n9056), .ZN(n8933)
         );
  XNOR2_X1 U10234 ( .A(n8933), .B(n6532), .ZN(n9150) );
  OAI22_X1 U10235 ( .A1(n9605), .A2(n9056), .B1(n9110), .B2(n6689), .ZN(n9149)
         );
  NAND2_X1 U10236 ( .A1(n9150), .A2(n9149), .ZN(n8934) );
  NAND2_X1 U10237 ( .A1(n9529), .A2(n4497), .ZN(n8936) );
  OR2_X1 U10238 ( .A1(n9152), .A2(n9056), .ZN(n8935) );
  NAND2_X1 U10239 ( .A1(n8936), .A2(n8935), .ZN(n8937) );
  XNOR2_X1 U10240 ( .A(n8937), .B(n6687), .ZN(n8940) );
  NOR2_X1 U10241 ( .A1(n9152), .A2(n6689), .ZN(n8938) );
  AOI21_X1 U10242 ( .B1(n9529), .B2(n7593), .A(n8938), .ZN(n8939) );
  NAND2_X1 U10243 ( .A1(n8940), .A2(n8939), .ZN(n9050) );
  OAI22_X1 U10244 ( .A1(n9401), .A2(n9056), .B1(n9078), .B2(n6485), .ZN(n8963)
         );
  NAND2_X1 U10245 ( .A1(n9520), .A2(n4497), .ZN(n8942) );
  OR2_X1 U10246 ( .A1(n9078), .A2(n9056), .ZN(n8941) );
  NAND2_X1 U10247 ( .A1(n8942), .A2(n8941), .ZN(n8943) );
  XNOR2_X1 U10248 ( .A(n8943), .B(n6532), .ZN(n8962) );
  XOR2_X1 U10249 ( .A(n8963), .B(n8962), .Z(n9126) );
  NAND2_X1 U10250 ( .A1(n9513), .A2(n7593), .ZN(n8945) );
  OR2_X1 U10251 ( .A1(n9079), .A2(n6485), .ZN(n8944) );
  NAND2_X1 U10252 ( .A1(n8945), .A2(n8944), .ZN(n8969) );
  NAND2_X1 U10253 ( .A1(n9513), .A2(n4497), .ZN(n8947) );
  OR2_X1 U10254 ( .A1(n9079), .A2(n9056), .ZN(n8946) );
  NAND2_X1 U10255 ( .A1(n8947), .A2(n8946), .ZN(n8948) );
  XNOR2_X1 U10256 ( .A(n8948), .B(n8978), .ZN(n9026) );
  NAND2_X1 U10257 ( .A1(n5475), .A2(n4497), .ZN(n8950) );
  OR2_X1 U10258 ( .A1(n9137), .A2(n9056), .ZN(n8949) );
  NAND2_X1 U10259 ( .A1(n8950), .A2(n8949), .ZN(n8951) );
  XNOR2_X1 U10260 ( .A(n8951), .B(n6687), .ZN(n9030) );
  NOR2_X1 U10261 ( .A1(n9137), .A2(n6689), .ZN(n8952) );
  AOI21_X1 U10262 ( .B1(n5475), .B2(n7593), .A(n8952), .ZN(n9029) );
  NOR2_X1 U10263 ( .A1(n9030), .A2(n9029), .ZN(n9028) );
  AOI21_X1 U10264 ( .B1(n8969), .B2(n9026), .A(n9028), .ZN(n8960) );
  NAND2_X1 U10265 ( .A1(n9518), .A2(n4497), .ZN(n8954) );
  NAND2_X1 U10266 ( .A1(n9199), .A2(n7593), .ZN(n8953) );
  NAND2_X1 U10267 ( .A1(n8954), .A2(n8953), .ZN(n8955) );
  XNOR2_X1 U10268 ( .A(n8955), .B(n6532), .ZN(n8958) );
  INV_X1 U10269 ( .A(n8958), .ZN(n8956) );
  AOI22_X1 U10270 ( .A1(n9518), .A2(n7593), .B1(n8988), .B2(n9199), .ZN(n8957)
         );
  NAND2_X1 U10271 ( .A1(n8956), .A2(n8957), .ZN(n8966) );
  INV_X1 U10272 ( .A(n8966), .ZN(n8959) );
  XNOR2_X1 U10273 ( .A(n8958), .B(n8957), .ZN(n9077) );
  AND2_X1 U10274 ( .A1(n8960), .A2(n9022), .ZN(n8961) );
  AND2_X1 U10275 ( .A1(n9126), .A2(n8961), .ZN(n8968) );
  INV_X1 U10276 ( .A(n8961), .ZN(n8967) );
  INV_X1 U10277 ( .A(n8962), .ZN(n8965) );
  INV_X1 U10278 ( .A(n8963), .ZN(n8964) );
  NAND2_X1 U10279 ( .A1(n8965), .A2(n8964), .ZN(n9075) );
  AND2_X1 U10280 ( .A1(n9075), .A2(n8966), .ZN(n9024) );
  AOI21_X1 U10281 ( .B1(n9125), .B2(n8968), .A(n4860), .ZN(n8976) );
  INV_X1 U10282 ( .A(n9026), .ZN(n8970) );
  AOI21_X1 U10283 ( .B1(n8970), .B2(n9135), .A(n9029), .ZN(n8973) );
  INV_X1 U10284 ( .A(n9030), .ZN(n8972) );
  NAND3_X1 U10285 ( .A1(n9029), .A2(n9135), .A3(n8970), .ZN(n8971) );
  OAI21_X1 U10286 ( .B1(n8973), .B2(n8972), .A(n8971), .ZN(n8974) );
  INV_X1 U10287 ( .A(n8974), .ZN(n8975) );
  NAND2_X1 U10288 ( .A1(n8976), .A2(n8975), .ZN(n9116) );
  AOI22_X1 U10289 ( .A1(n9346), .A2(n4497), .B1(n7593), .B2(n9196), .ZN(n8977)
         );
  XOR2_X1 U10290 ( .A(n8978), .B(n8977), .Z(n8981) );
  OAI22_X1 U10291 ( .A1(n5480), .A2(n9056), .B1(n8979), .B2(n6485), .ZN(n8980)
         );
  NOR2_X1 U10292 ( .A1(n8981), .A2(n8980), .ZN(n8982) );
  AOI21_X1 U10293 ( .B1(n8981), .B2(n8980), .A(n8982), .ZN(n9117) );
  NAND2_X1 U10294 ( .A1(n9116), .A2(n9117), .ZN(n9115) );
  INV_X1 U10295 ( .A(n8982), .ZN(n8983) );
  NAND2_X1 U10296 ( .A1(n9115), .A2(n8983), .ZN(n9085) );
  OAI22_X1 U10297 ( .A1(n9330), .A2(n9058), .B1(n9170), .B2(n9056), .ZN(n8984)
         );
  XNOR2_X1 U10298 ( .A(n8984), .B(n6532), .ZN(n8991) );
  NOR2_X1 U10299 ( .A1(n9170), .A2(n6485), .ZN(n8985) );
  AOI21_X1 U10300 ( .B1(n9500), .B2(n7593), .A(n8985), .ZN(n8992) );
  XNOR2_X1 U10301 ( .A(n8991), .B(n8992), .ZN(n9086) );
  NAND2_X1 U10302 ( .A1(n9085), .A2(n9086), .ZN(n9084) );
  OAI22_X1 U10303 ( .A1(n9569), .A2(n9058), .B1(n8986), .B2(n9056), .ZN(n8987)
         );
  XNOR2_X1 U10304 ( .A(n8987), .B(n6532), .ZN(n8996) );
  OR2_X1 U10305 ( .A1(n9569), .A2(n9056), .ZN(n8990) );
  NAND2_X1 U10306 ( .A1(n9194), .A2(n8988), .ZN(n8989) );
  NAND2_X1 U10307 ( .A1(n8990), .A2(n8989), .ZN(n8995) );
  XNOR2_X1 U10308 ( .A(n8996), .B(n8995), .ZN(n9161) );
  INV_X1 U10309 ( .A(n8991), .ZN(n8993) );
  AND2_X1 U10310 ( .A1(n8993), .A2(n8992), .ZN(n9162) );
  NOR2_X1 U10311 ( .A1(n9161), .A2(n9162), .ZN(n8994) );
  NAND2_X1 U10312 ( .A1(n9084), .A2(n8994), .ZN(n9164) );
  NAND2_X1 U10313 ( .A1(n8996), .A2(n8995), .ZN(n9002) );
  AOI22_X1 U10314 ( .A1(n9010), .A2(n4497), .B1(n7593), .B2(n9193), .ZN(n8998)
         );
  XOR2_X1 U10315 ( .A(n6532), .B(n8998), .Z(n9000) );
  OAI22_X1 U10316 ( .A1(n4394), .A2(n9056), .B1(n9168), .B2(n6485), .ZN(n8999)
         );
  NOR2_X1 U10317 ( .A1(n9000), .A2(n8999), .ZN(n9068) );
  AOI21_X1 U10318 ( .B1(n9000), .B2(n8999), .A(n9068), .ZN(n9001) );
  AOI21_X1 U10319 ( .B1(n9164), .B2(n9002), .A(n9001), .ZN(n9006) );
  INV_X1 U10320 ( .A(n9001), .ZN(n9004) );
  INV_X1 U10321 ( .A(n9002), .ZN(n9003) );
  NOR2_X1 U10322 ( .A1(n9004), .A2(n9003), .ZN(n9005) );
  AND2_X2 U10323 ( .A1(n9164), .A2(n9005), .ZN(n9064) );
  OAI21_X1 U10324 ( .B1(n9006), .B2(n9064), .A(n9165), .ZN(n9012) );
  AOI22_X1 U10325 ( .A1(n4270), .A2(n9007), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n9008) );
  OAI21_X1 U10326 ( .B1(n9157), .B2(n9295), .A(n9008), .ZN(n9009) );
  AOI21_X1 U10327 ( .B1(n9010), .B2(n4264), .A(n9009), .ZN(n9011) );
  NAND2_X1 U10328 ( .A1(n9012), .A2(n9011), .ZN(P1_U3214) );
  AOI21_X1 U10329 ( .B1(n9014), .B2(n9013), .A(n4293), .ZN(n9021) );
  NAND2_X1 U10330 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9715) );
  NAND2_X1 U10331 ( .A1(n4270), .A2(n9015), .ZN(n9016) );
  OAI211_X1 U10332 ( .C1(n9186), .C2(n9017), .A(n9715), .B(n9016), .ZN(n9018)
         );
  AOI21_X1 U10333 ( .B1(n9019), .B2(n4264), .A(n9018), .ZN(n9020) );
  OAI21_X1 U10334 ( .B1(n9021), .B2(n9189), .A(n9020), .ZN(P1_U3215) );
  NAND2_X1 U10335 ( .A1(n9125), .A2(n9126), .ZN(n9074) );
  AOI21_X2 U10336 ( .B1(n9074), .B2(n9024), .A(n9023), .ZN(n9025) );
  XNOR2_X1 U10337 ( .A(n9025), .B(n9026), .ZN(n9134) );
  NAND2_X1 U10338 ( .A1(n9134), .A2(n9135), .ZN(n9133) );
  INV_X1 U10339 ( .A(n9025), .ZN(n9027) );
  AOI21_X1 U10340 ( .B1(n9030), .B2(n9029), .A(n9028), .ZN(n9031) );
  INV_X1 U10341 ( .A(n9357), .ZN(n9037) );
  OR2_X1 U10342 ( .A1(n9079), .A2(n9169), .ZN(n9035) );
  NAND2_X1 U10343 ( .A1(n9196), .A2(n9129), .ZN(n9034) );
  NAND2_X1 U10344 ( .A1(n9035), .A2(n9034), .ZN(n9353) );
  AOI22_X1 U10345 ( .A1(n9353), .A2(n4270), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9036) );
  OAI21_X1 U10346 ( .B1(n9157), .B2(n9037), .A(n9036), .ZN(n9038) );
  AOI21_X1 U10347 ( .B1(n5475), .B2(n4264), .A(n9038), .ZN(n9039) );
  OAI21_X1 U10348 ( .B1(n9040), .B2(n9189), .A(n9039), .ZN(P1_U3216) );
  OAI21_X1 U10349 ( .B1(n9042), .B2(n9041), .A(n6700), .ZN(n9043) );
  NAND2_X1 U10350 ( .A1(n9043), .A2(n9165), .ZN(n9047) );
  AOI22_X1 U10351 ( .A1(n9747), .A2(n4264), .B1(n4270), .B2(n9044), .ZN(n9046)
         );
  MUX2_X1 U10352 ( .A(P1_STATE_REG_SCAN_IN), .B(n9157), .S(n9748), .Z(n9045)
         );
  NAND3_X1 U10353 ( .A1(n9047), .A2(n9046), .A3(n9045), .ZN(P1_U3218) );
  NAND2_X1 U10354 ( .A1(n4852), .A2(n9050), .ZN(n9048) );
  AOI22_X1 U10355 ( .A1(n4311), .A2(n9050), .B1(n9049), .B2(n9048), .ZN(n9054)
         );
  OAI22_X1 U10356 ( .A1(n9078), .A2(n9167), .B1(n9110), .B2(n9169), .ZN(n9410)
         );
  AOI22_X1 U10357 ( .A1(n9410), .A2(n4270), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3086), .ZN(n9051) );
  OAI21_X1 U10358 ( .B1(n9186), .B2(n9415), .A(n9051), .ZN(n9052) );
  AOI21_X1 U10359 ( .B1(n9529), .B2(n4264), .A(n9052), .ZN(n9053) );
  OAI21_X1 U10360 ( .B1(n9054), .B2(n9189), .A(n9053), .ZN(P1_U3219) );
  INV_X1 U10361 ( .A(n9064), .ZN(n9063) );
  OAI22_X1 U10362 ( .A1(n9568), .A2(n9056), .B1(n9057), .B2(n6485), .ZN(n9055)
         );
  XNOR2_X1 U10363 ( .A(n9055), .B(n6687), .ZN(n9060) );
  OAI22_X1 U10364 ( .A1(n9568), .A2(n9058), .B1(n9057), .B2(n9056), .ZN(n9059)
         );
  XNOR2_X1 U10365 ( .A(n9060), .B(n9059), .ZN(n9069) );
  INV_X1 U10366 ( .A(n9069), .ZN(n9062) );
  INV_X1 U10367 ( .A(n9068), .ZN(n9061) );
  NAND3_X1 U10368 ( .A1(n9064), .A2(n9165), .A3(n9069), .ZN(n9072) );
  OAI22_X1 U10369 ( .A1(n9168), .A2(n9169), .B1(n9065), .B2(n9167), .ZN(n9280)
         );
  AOI22_X1 U10370 ( .A1(n4270), .A2(n9280), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n9066) );
  OAI21_X1 U10371 ( .B1(n9157), .B2(n9287), .A(n9066), .ZN(n9067) );
  AOI21_X1 U10372 ( .B1(n9289), .B2(n4264), .A(n9067), .ZN(n9071) );
  NAND3_X1 U10373 ( .A1(n9069), .A2(n9165), .A3(n9068), .ZN(n9070) );
  NAND4_X1 U10374 ( .A1(n9073), .A2(n9072), .A3(n9071), .A4(n9070), .ZN(
        P1_U3220) );
  NAND2_X1 U10375 ( .A1(n9074), .A2(n9075), .ZN(n9076) );
  XOR2_X1 U10376 ( .A(n9077), .B(n9076), .Z(n9083) );
  OAI22_X1 U10377 ( .A1(n9079), .A2(n9167), .B1(n9078), .B2(n9169), .ZN(n9379)
         );
  AOI22_X1 U10378 ( .A1(n9379), .A2(n4270), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9080) );
  OAI21_X1 U10379 ( .B1(n9186), .B2(n9382), .A(n9080), .ZN(n9081) );
  AOI21_X1 U10380 ( .B1(n9518), .B2(n4264), .A(n9081), .ZN(n9082) );
  OAI21_X1 U10381 ( .B1(n9083), .B2(n9189), .A(n9082), .ZN(P1_U3223) );
  OAI21_X1 U10382 ( .B1(n9086), .B2(n9085), .A(n9084), .ZN(n9092) );
  NAND2_X1 U10383 ( .A1(n9500), .A2(n4264), .ZN(n9090) );
  NAND2_X1 U10384 ( .A1(n9196), .A2(n9138), .ZN(n9088) );
  NAND2_X1 U10385 ( .A1(n9194), .A2(n9129), .ZN(n9087) );
  NAND2_X1 U10386 ( .A1(n9088), .A2(n9087), .ZN(n9323) );
  AOI22_X1 U10387 ( .A1(n4270), .A2(n9323), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9089) );
  OAI211_X1 U10388 ( .C1(n9186), .C2(n9326), .A(n9090), .B(n9089), .ZN(n9091)
         );
  AOI21_X1 U10389 ( .B1(n9092), .B2(n9165), .A(n9091), .ZN(n9093) );
  INV_X1 U10390 ( .A(n9093), .ZN(P1_U3225) );
  OAI21_X1 U10391 ( .B1(n9096), .B2(n9094), .A(n9095), .ZN(n9097) );
  NAND2_X1 U10392 ( .A1(n9097), .A2(n9165), .ZN(n9104) );
  OR2_X1 U10393 ( .A1(n9154), .A2(n9167), .ZN(n9100) );
  OR2_X1 U10394 ( .A1(n9098), .A2(n9169), .ZN(n9099) );
  NAND2_X1 U10395 ( .A1(n9100), .A2(n9099), .ZN(n9465) );
  NOR2_X1 U10396 ( .A1(n9101), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9226) );
  NOR2_X1 U10397 ( .A1(n9186), .A2(n9472), .ZN(n9102) );
  AOI211_X1 U10398 ( .C1(n4270), .C2(n9465), .A(n9226), .B(n9102), .ZN(n9103)
         );
  OAI211_X1 U10399 ( .C1(n9477), .C2(n9147), .A(n9104), .B(n9103), .ZN(
        P1_U3226) );
  NAND2_X1 U10400 ( .A1(n9107), .A2(n9106), .ZN(n9108) );
  XNOR2_X1 U10401 ( .A(n9105), .B(n9108), .ZN(n9114) );
  OAI22_X1 U10402 ( .A1(n9110), .A2(n9167), .B1(n9109), .B2(n9169), .ZN(n9454)
         );
  NOR2_X1 U10403 ( .A1(n9967), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9246) );
  AOI21_X1 U10404 ( .B1(n4270), .B2(n9454), .A(n9246), .ZN(n9111) );
  OAI21_X1 U10405 ( .B1(n9157), .B2(n9446), .A(n9111), .ZN(n9112) );
  AOI21_X1 U10406 ( .B1(n9540), .B2(n4264), .A(n9112), .ZN(n9113) );
  OAI21_X1 U10407 ( .B1(n9114), .B2(n9189), .A(n9113), .ZN(P1_U3228) );
  OAI21_X1 U10408 ( .B1(n9117), .B2(n9116), .A(n9115), .ZN(n9123) );
  NAND2_X1 U10409 ( .A1(n9346), .A2(n4264), .ZN(n9121) );
  OR2_X1 U10410 ( .A1(n9137), .A2(n9169), .ZN(n9119) );
  OR2_X1 U10411 ( .A1(n9170), .A2(n9167), .ZN(n9118) );
  NAND2_X1 U10412 ( .A1(n9119), .A2(n9118), .ZN(n9336) );
  AOI22_X1 U10413 ( .A1(n9336), .A2(n4270), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n9120) );
  OAI211_X1 U10414 ( .C1(n9157), .C2(n9341), .A(n9121), .B(n9120), .ZN(n9122)
         );
  AOI21_X1 U10415 ( .B1(n9123), .B2(n9165), .A(n9122), .ZN(n9124) );
  INV_X1 U10416 ( .A(n9124), .ZN(P1_U3229) );
  OAI21_X1 U10417 ( .B1(n9126), .B2(n9125), .A(n9074), .ZN(n9127) );
  NAND2_X1 U10418 ( .A1(n9127), .A2(n9165), .ZN(n9132) );
  NOR2_X1 U10419 ( .A1(n9152), .A2(n9169), .ZN(n9128) );
  AOI21_X1 U10420 ( .B1(n9199), .B2(n9129), .A(n9128), .ZN(n9390) );
  OAI22_X1 U10421 ( .A1(n9390), .A2(n9142), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9996), .ZN(n9130) );
  AOI21_X1 U10422 ( .B1(n9398), .B2(n9144), .A(n9130), .ZN(n9131) );
  OAI211_X1 U10423 ( .C1(n9401), .C2(n9147), .A(n9132), .B(n9131), .ZN(
        P1_U3233) );
  OAI21_X1 U10424 ( .B1(n9135), .B2(n9134), .A(n9133), .ZN(n9136) );
  NAND2_X1 U10425 ( .A1(n9136), .A2(n9165), .ZN(n9146) );
  OR2_X1 U10426 ( .A1(n9137), .A2(n9167), .ZN(n9140) );
  NAND2_X1 U10427 ( .A1(n9199), .A2(n9138), .ZN(n9139) );
  AND2_X1 U10428 ( .A1(n9140), .A2(n9139), .ZN(n9366) );
  INV_X1 U10429 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9141) );
  OAI22_X1 U10430 ( .A1(n9366), .A2(n9142), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9141), .ZN(n9143) );
  AOI21_X1 U10431 ( .B1(n9371), .B2(n9144), .A(n9143), .ZN(n9145) );
  OAI211_X1 U10432 ( .C1(n5479), .C2(n9147), .A(n9146), .B(n9145), .ZN(
        P1_U3235) );
  XNOR2_X1 U10433 ( .A(n9150), .B(n9149), .ZN(n9151) );
  XNOR2_X1 U10434 ( .A(n9148), .B(n9151), .ZN(n9160) );
  INV_X1 U10435 ( .A(n9435), .ZN(n9156) );
  OR2_X1 U10436 ( .A1(n9152), .A2(n9167), .ZN(n9153) );
  OAI21_X1 U10437 ( .B1(n9154), .B2(n9169), .A(n9153), .ZN(n9428) );
  AOI22_X1 U10438 ( .A1(n4270), .A2(n9428), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n9155) );
  OAI21_X1 U10439 ( .B1(n9157), .B2(n9156), .A(n9155), .ZN(n9158) );
  AOI21_X1 U10440 ( .B1(n9434), .B2(n4264), .A(n9158), .ZN(n9159) );
  OAI21_X1 U10441 ( .B1(n9160), .B2(n9189), .A(n9159), .ZN(P1_U3238) );
  INV_X1 U10442 ( .A(n9084), .ZN(n9163) );
  NAND3_X1 U10443 ( .A1(n9166), .A2(n9165), .A3(n9164), .ZN(n9177) );
  OR2_X1 U10444 ( .A1(n9168), .A2(n9167), .ZN(n9172) );
  OR2_X1 U10445 ( .A1(n9170), .A2(n9169), .ZN(n9171) );
  NAND2_X1 U10446 ( .A1(n9172), .A2(n9171), .ZN(n9305) );
  AOI22_X1 U10447 ( .A1(n4270), .A2(n9305), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9173) );
  OAI21_X1 U10448 ( .B1(n9186), .B2(n9310), .A(n9173), .ZN(n9174) );
  AOI21_X1 U10449 ( .B1(n9315), .B2(n4264), .A(n9174), .ZN(n9176) );
  NAND2_X1 U10450 ( .A1(n9177), .A2(n9176), .ZN(P1_U3240) );
  INV_X1 U10451 ( .A(n9178), .ZN(n9179) );
  AOI21_X1 U10452 ( .B1(n9181), .B2(n9180), .A(n9179), .ZN(n9190) );
  NAND2_X1 U10453 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9727) );
  NAND2_X1 U10454 ( .A1(n4270), .A2(n9183), .ZN(n9184) );
  OAI211_X1 U10455 ( .C1(n9186), .C2(n9185), .A(n9727), .B(n9184), .ZN(n9187)
         );
  AOI21_X1 U10456 ( .B1(n9616), .B2(n4264), .A(n9187), .ZN(n9188) );
  OAI21_X1 U10457 ( .B1(n9190), .B2(n9189), .A(n9188), .ZN(P1_U3241) );
  MUX2_X1 U10458 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9191), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10459 ( .A(n9192), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9218), .Z(
        P1_U3582) );
  MUX2_X1 U10460 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9193), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10461 ( .A(n9194), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9218), .Z(
        P1_U3580) );
  MUX2_X1 U10462 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9195), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10463 ( .A(n9196), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9218), .Z(
        P1_U3578) );
  MUX2_X1 U10464 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9197), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10465 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9198), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10466 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9199), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10467 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9200), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10468 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9201), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10469 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9202), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10470 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9203), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10471 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9204), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10472 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9205), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10473 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9206), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10474 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9207), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10475 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9208), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10476 ( .A(n9209), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9218), .Z(
        P1_U3564) );
  MUX2_X1 U10477 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9210), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10478 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9211), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10479 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9212), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10480 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9213), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10481 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9214), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10482 ( .A(n9215), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9218), .Z(
        P1_U3558) );
  MUX2_X1 U10483 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9216), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10484 ( .A(n9217), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9218), .Z(
        P1_U3556) );
  MUX2_X1 U10485 ( .A(n9219), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9218), .Z(
        P1_U3554) );
  INV_X1 U10486 ( .A(n9232), .ZN(n9702) );
  OAI21_X1 U10487 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n9230), .A(n9220), .ZN(
        n9695) );
  XNOR2_X1 U10488 ( .A(n9702), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9696) );
  NOR2_X1 U10489 ( .A1(n9695), .A2(n9696), .ZN(n9694) );
  XNOR2_X1 U10490 ( .A(n9714), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9710) );
  NOR2_X1 U10491 ( .A1(n9711), .A2(n9710), .ZN(n9709) );
  NOR2_X1 U10492 ( .A1(n9221), .A2(n9717), .ZN(n9222) );
  XNOR2_X1 U10493 ( .A(n9717), .B(n9221), .ZN(n9720) );
  NOR2_X1 U10494 ( .A1(n10024), .A2(n9720), .ZN(n9719) );
  NOR2_X1 U10495 ( .A1(n9222), .A2(n9719), .ZN(n9225) );
  AOI22_X1 U10496 ( .A1(n9245), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9223), .B2(
        n9228), .ZN(n9224) );
  NAND2_X1 U10497 ( .A1(n9224), .A2(n9225), .ZN(n9244) );
  OAI21_X1 U10498 ( .B1(n9225), .B2(n9224), .A(n9244), .ZN(n9241) );
  AOI21_X1 U10499 ( .B1(n9247), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n9226), .ZN(
        n9227) );
  OAI21_X1 U10500 ( .B1(n9228), .B2(n9739), .A(n9227), .ZN(n9240) );
  OAI21_X1 U10501 ( .B1(n9230), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9229), .ZN(
        n9699) );
  XNOR2_X1 U10502 ( .A(n9232), .B(n9231), .ZN(n9698) );
  NOR2_X1 U10503 ( .A1(n9699), .A2(n9698), .ZN(n9697) );
  NAND2_X1 U10504 ( .A1(n9714), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9233) );
  OAI21_X1 U10505 ( .B1(n9714), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9233), .ZN(
        n9707) );
  NOR2_X1 U10506 ( .A1(n9234), .A2(n9717), .ZN(n9235) );
  NOR2_X1 U10507 ( .A1(n7887), .A2(n9722), .ZN(n9721) );
  NOR2_X1 U10508 ( .A1(n9235), .A2(n9721), .ZN(n9238) );
  NAND2_X1 U10509 ( .A1(n9245), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9236) );
  OAI21_X1 U10510 ( .B1(n9245), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9236), .ZN(
        n9237) );
  NOR2_X1 U10511 ( .A1(n9238), .A2(n9237), .ZN(n9243) );
  AOI211_X1 U10512 ( .C1(n9238), .C2(n9237), .A(n9243), .B(n9730), .ZN(n9239)
         );
  AOI211_X1 U10513 ( .C1(n9733), .C2(n9241), .A(n9240), .B(n9239), .ZN(n9242)
         );
  INV_X1 U10514 ( .A(n9242), .ZN(P1_U3259) );
  XNOR2_X1 U10515 ( .A(n9260), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n9253) );
  XOR2_X1 U10516 ( .A(n9253), .B(n9254), .Z(n9252) );
  XNOR2_X1 U10517 ( .A(n9260), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9261) );
  XNOR2_X1 U10518 ( .A(n9262), .B(n9261), .ZN(n9250) );
  AOI21_X1 U10519 ( .B1(n9247), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n9246), .ZN(
        n9248) );
  OAI21_X1 U10520 ( .B1(n9260), .B2(n9739), .A(n9248), .ZN(n9249) );
  AOI21_X1 U10521 ( .B1(n9250), .B2(n9733), .A(n9249), .ZN(n9251) );
  OAI21_X1 U10522 ( .B1(n9252), .B2(n9730), .A(n9251), .ZN(P1_U3260) );
  INV_X1 U10523 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9447) );
  NAND2_X1 U10524 ( .A1(n9260), .A2(n9447), .ZN(n9255) );
  INV_X1 U10525 ( .A(n9738), .ZN(n9256) );
  NAND2_X1 U10526 ( .A1(n9256), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9258) );
  NAND2_X1 U10527 ( .A1(n9738), .A2(n10055), .ZN(n9257) );
  NAND2_X1 U10528 ( .A1(n9258), .A2(n9257), .ZN(n9731) );
  NAND2_X1 U10529 ( .A1(n9741), .A2(n9258), .ZN(n9259) );
  NOR2_X1 U10530 ( .A1(n9738), .A2(n9534), .ZN(n9263) );
  AOI21_X1 U10531 ( .B1(n9534), .B2(n9738), .A(n9263), .ZN(n9735) );
  NAND2_X1 U10532 ( .A1(n9736), .A2(n9735), .ZN(n9734) );
  INV_X1 U10533 ( .A(n9263), .ZN(n9264) );
  NAND2_X1 U10534 ( .A1(n9734), .A2(n9264), .ZN(n9265) );
  XNOR2_X1 U10535 ( .A(n9265), .B(n9530), .ZN(n9267) );
  OAI21_X1 U10536 ( .B1(n9267), .B2(n9718), .A(n9739), .ZN(n9266) );
  NAND2_X1 U10537 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9269) );
  NAND2_X1 U10538 ( .A1(n9275), .A2(n9562), .ZN(n9274) );
  NAND2_X1 U10539 ( .A1(n9271), .A2(n9270), .ZN(n9485) );
  NOR2_X1 U10540 ( .A1(n9749), .A2(n9485), .ZN(n9277) );
  NOR2_X1 U10541 ( .A1(n9558), .A2(n9444), .ZN(n9272) );
  AOI211_X1 U10542 ( .C1(n9405), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9277), .B(
        n9272), .ZN(n9273) );
  OAI21_X1 U10543 ( .B1(n9482), .B2(n9765), .A(n9273), .ZN(P1_U3263) );
  OAI211_X1 U10544 ( .C1(n9275), .C2(n9562), .A(n9521), .B(n9274), .ZN(n9486)
         );
  NOR2_X1 U10545 ( .A1(n9562), .A2(n9444), .ZN(n9276) );
  AOI211_X1 U10546 ( .C1(n9405), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9277), .B(
        n9276), .ZN(n9278) );
  OAI21_X1 U10547 ( .B1(n9486), .B2(n9765), .A(n9278), .ZN(P1_U3264) );
  XNOR2_X1 U10548 ( .A(n9279), .B(n9283), .ZN(n9281) );
  AOI21_X1 U10549 ( .B1(n9281), .B2(n9463), .A(n9280), .ZN(n9490) );
  OAI21_X1 U10550 ( .B1(n9284), .B2(n9283), .A(n9282), .ZN(n9563) );
  OAI211_X1 U10551 ( .C1(n9568), .C2(n4304), .A(n9521), .B(n9285), .ZN(n9489)
         );
  NAND2_X1 U10552 ( .A1(n9405), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9286) );
  OAI21_X1 U10553 ( .B1(n9471), .B2(n9287), .A(n9286), .ZN(n9288) );
  AOI21_X1 U10554 ( .B1(n9289), .B2(n9762), .A(n9288), .ZN(n9290) );
  OAI21_X1 U10555 ( .B1(n9489), .B2(n9765), .A(n9290), .ZN(n9291) );
  AOI21_X1 U10556 ( .B1(n9563), .B2(n9754), .A(n9291), .ZN(n9292) );
  OAI21_X1 U10557 ( .B1(n9405), .B2(n9490), .A(n9292), .ZN(P1_U3265) );
  INV_X1 U10558 ( .A(n9293), .ZN(n9302) );
  NAND2_X1 U10559 ( .A1(n9294), .A2(n9754), .ZN(n9301) );
  NOR2_X1 U10560 ( .A1(n4394), .A2(n9444), .ZN(n9298) );
  OAI22_X1 U10561 ( .A1(n9457), .A2(n9296), .B1(n9295), .B2(n9471), .ZN(n9297)
         );
  AOI211_X1 U10562 ( .C1(n9299), .C2(n9450), .A(n9298), .B(n9297), .ZN(n9300)
         );
  OAI211_X1 U10563 ( .C1(n9749), .C2(n9302), .A(n9301), .B(n9300), .ZN(
        P1_U3266) );
  XNOR2_X1 U10564 ( .A(n9304), .B(n9303), .ZN(n9306) );
  AOI21_X1 U10565 ( .B1(n9306), .B2(n9463), .A(n9305), .ZN(n9495) );
  XNOR2_X1 U10566 ( .A(n9308), .B(n9307), .ZN(n9570) );
  INV_X1 U10567 ( .A(n9570), .ZN(n9309) );
  NAND2_X1 U10568 ( .A1(n9309), .A2(n9754), .ZN(n9317) );
  OAI22_X1 U10569 ( .A1(n9457), .A2(n9311), .B1(n9310), .B2(n9471), .ZN(n9314)
         );
  OAI211_X1 U10570 ( .C1(n9569), .C2(n9325), .A(n9521), .B(n9312), .ZN(n9494)
         );
  NOR2_X1 U10571 ( .A1(n9494), .A2(n9765), .ZN(n9313) );
  AOI211_X1 U10572 ( .C1(n9762), .C2(n9315), .A(n9314), .B(n9313), .ZN(n9316)
         );
  OAI211_X1 U10573 ( .C1(n9749), .C2(n9495), .A(n9317), .B(n9316), .ZN(
        P1_U3267) );
  XOR2_X1 U10574 ( .A(n9319), .B(n9318), .Z(n9577) );
  OAI21_X1 U10575 ( .B1(n9334), .B2(n9320), .A(n9319), .ZN(n9322) );
  AOI21_X1 U10576 ( .B1(n9322), .B2(n9321), .A(n9412), .ZN(n9324) );
  AOI211_X1 U10577 ( .C1(n9500), .C2(n9343), .A(n9443), .B(n9325), .ZN(n9498)
         );
  NAND2_X1 U10578 ( .A1(n9498), .A2(n9450), .ZN(n9329) );
  NOR2_X1 U10579 ( .A1(n9471), .A2(n9326), .ZN(n9327) );
  AOI21_X1 U10580 ( .B1(n9405), .B2(P1_REG2_REG_25__SCAN_IN), .A(n9327), .ZN(
        n9328) );
  OAI211_X1 U10581 ( .C1(n9330), .C2(n9444), .A(n9329), .B(n9328), .ZN(n9331)
         );
  AOI21_X1 U10582 ( .B1(n9457), .B2(n9499), .A(n9331), .ZN(n9332) );
  OAI21_X1 U10583 ( .B1(n9577), .B2(n9460), .A(n9332), .ZN(P1_U3268) );
  AOI21_X1 U10584 ( .B1(n9333), .B2(n9349), .A(n9339), .ZN(n9335) );
  NOR3_X1 U10585 ( .A1(n9335), .A2(n9334), .A3(n9412), .ZN(n9337) );
  NOR2_X1 U10586 ( .A1(n9337), .A2(n9336), .ZN(n9504) );
  XOR2_X1 U10587 ( .A(n9339), .B(n9338), .Z(n9578) );
  INV_X1 U10588 ( .A(n9578), .ZN(n9340) );
  NAND2_X1 U10589 ( .A1(n9340), .A2(n9754), .ZN(n9348) );
  OAI22_X1 U10590 ( .A1(n9474), .A2(n9342), .B1(n9341), .B2(n9471), .ZN(n9345)
         );
  OAI211_X1 U10591 ( .C1(n9356), .C2(n5480), .A(n9521), .B(n9343), .ZN(n9503)
         );
  NOR2_X1 U10592 ( .A1(n9503), .A2(n9765), .ZN(n9344) );
  AOI211_X1 U10593 ( .C1(n9762), .C2(n9346), .A(n9345), .B(n9344), .ZN(n9347)
         );
  OAI211_X1 U10594 ( .C1(n9749), .C2(n9504), .A(n9348), .B(n9347), .ZN(
        P1_U3269) );
  XNOR2_X1 U10595 ( .A(n4330), .B(n9351), .ZN(n9585) );
  OAI21_X1 U10596 ( .B1(n9351), .B2(n9350), .A(n9349), .ZN(n9352) );
  NAND2_X1 U10597 ( .A1(n9352), .A2(n9463), .ZN(n9355) );
  INV_X1 U10598 ( .A(n9353), .ZN(n9354) );
  NAND2_X1 U10599 ( .A1(n9355), .A2(n9354), .ZN(n9508) );
  AOI211_X1 U10600 ( .C1(n5475), .C2(n9369), .A(n9443), .B(n9356), .ZN(n9507)
         );
  NAND2_X1 U10601 ( .A1(n9507), .A2(n9450), .ZN(n9359) );
  AOI22_X1 U10602 ( .A1(n9357), .A2(n9758), .B1(n9405), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n9358) );
  OAI211_X1 U10603 ( .C1(n4395), .C2(n9444), .A(n9359), .B(n9358), .ZN(n9360)
         );
  AOI21_X1 U10604 ( .B1(n9457), .B2(n9508), .A(n9360), .ZN(n9361) );
  OAI21_X1 U10605 ( .B1(n9585), .B2(n9460), .A(n9361), .ZN(P1_U3270) );
  XNOR2_X1 U10606 ( .A(n9362), .B(n9364), .ZN(n9589) );
  XNOR2_X1 U10607 ( .A(n9363), .B(n9364), .ZN(n9365) );
  NAND2_X1 U10608 ( .A1(n9365), .A2(n9463), .ZN(n9367) );
  NAND2_X1 U10609 ( .A1(n9367), .A2(n9366), .ZN(n9512) );
  INV_X1 U10610 ( .A(n9369), .ZN(n9370) );
  AOI211_X1 U10611 ( .C1(n9513), .C2(n4399), .A(n9443), .B(n9370), .ZN(n9511)
         );
  NAND2_X1 U10612 ( .A1(n9511), .A2(n9450), .ZN(n9373) );
  AOI22_X1 U10613 ( .A1(n9371), .A2(n9758), .B1(n9405), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9372) );
  OAI211_X1 U10614 ( .C1(n5479), .C2(n9444), .A(n9373), .B(n9372), .ZN(n9374)
         );
  AOI21_X1 U10615 ( .B1(n9474), .B2(n9512), .A(n9374), .ZN(n9375) );
  OAI21_X1 U10616 ( .B1(n9589), .B2(n9460), .A(n9375), .ZN(P1_U3271) );
  XOR2_X1 U10617 ( .A(n9377), .B(n9376), .Z(n9593) );
  XOR2_X1 U10618 ( .A(n9378), .B(n9377), .Z(n9381) );
  INV_X1 U10619 ( .A(n9379), .ZN(n9380) );
  OAI21_X1 U10620 ( .B1(n9381), .B2(n9412), .A(n9380), .ZN(n9516) );
  AOI211_X1 U10621 ( .C1(n9518), .C2(n9396), .A(n9443), .B(n9368), .ZN(n9517)
         );
  NAND2_X1 U10622 ( .A1(n9517), .A2(n9450), .ZN(n9385) );
  INV_X1 U10623 ( .A(n9382), .ZN(n9383) );
  AOI22_X1 U10624 ( .A1(n9749), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9383), .B2(
        n9758), .ZN(n9384) );
  OAI211_X1 U10625 ( .C1(n9386), .C2(n9444), .A(n9385), .B(n9384), .ZN(n9387)
         );
  AOI21_X1 U10626 ( .B1(n9457), .B2(n9516), .A(n9387), .ZN(n9388) );
  OAI21_X1 U10627 ( .B1(n9593), .B2(n9460), .A(n9388), .ZN(P1_U3272) );
  XNOR2_X1 U10628 ( .A(n9389), .B(n9394), .ZN(n9392) );
  INV_X1 U10629 ( .A(n9390), .ZN(n9391) );
  AOI21_X1 U10630 ( .B1(n9392), .B2(n9463), .A(n9391), .ZN(n9524) );
  AOI21_X1 U10631 ( .B1(n9394), .B2(n9393), .A(n4314), .ZN(n9526) );
  INV_X1 U10632 ( .A(n9526), .ZN(n9403) );
  OR2_X1 U10633 ( .A1(n9401), .A2(n9414), .ZN(n9395) );
  AND2_X1 U10634 ( .A1(n9396), .A2(n9395), .ZN(n9522) );
  NAND2_X1 U10635 ( .A1(n9522), .A2(n9397), .ZN(n9400) );
  AOI22_X1 U10636 ( .A1(n9749), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9398), .B2(
        n9758), .ZN(n9399) );
  OAI211_X1 U10637 ( .C1(n9401), .C2(n9444), .A(n9400), .B(n9399), .ZN(n9402)
         );
  AOI21_X1 U10638 ( .B1(n9403), .B2(n9754), .A(n9402), .ZN(n9404) );
  OAI21_X1 U10639 ( .B1(n9405), .B2(n9524), .A(n9404), .ZN(P1_U3273) );
  XOR2_X1 U10640 ( .A(n9406), .B(n9409), .Z(n9598) );
  NAND2_X1 U10641 ( .A1(n9426), .A2(n9407), .ZN(n9408) );
  XNOR2_X1 U10642 ( .A(n9409), .B(n9408), .ZN(n9413) );
  INV_X1 U10643 ( .A(n9410), .ZN(n9411) );
  OAI21_X1 U10644 ( .B1(n9413), .B2(n9412), .A(n9411), .ZN(n9528) );
  AOI211_X1 U10645 ( .C1(n9529), .C2(n9432), .A(n9443), .B(n9414), .ZN(n9527)
         );
  NAND2_X1 U10646 ( .A1(n9527), .A2(n9450), .ZN(n9418) );
  INV_X1 U10647 ( .A(n9415), .ZN(n9416) );
  AOI22_X1 U10648 ( .A1(n9749), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9416), .B2(
        n9758), .ZN(n9417) );
  OAI211_X1 U10649 ( .C1(n9419), .C2(n9444), .A(n9418), .B(n9417), .ZN(n9420)
         );
  AOI21_X1 U10650 ( .B1(n9457), .B2(n9528), .A(n9420), .ZN(n9421) );
  OAI21_X1 U10651 ( .B1(n9598), .B2(n9460), .A(n9421), .ZN(P1_U3274) );
  XNOR2_X1 U10652 ( .A(n9422), .B(n9423), .ZN(n9599) );
  INV_X1 U10653 ( .A(n9599), .ZN(n9440) );
  INV_X1 U10654 ( .A(n9423), .ZN(n9425) );
  NAND3_X1 U10655 ( .A1(n9425), .A2(n9424), .A3(n9451), .ZN(n9427) );
  NAND3_X1 U10656 ( .A1(n9427), .A2(n9426), .A3(n9463), .ZN(n9430) );
  INV_X1 U10657 ( .A(n9428), .ZN(n9429) );
  NAND2_X1 U10658 ( .A1(n9430), .A2(n9429), .ZN(n9532) );
  INV_X1 U10659 ( .A(n9431), .ZN(n9442) );
  INV_X1 U10660 ( .A(n9432), .ZN(n9433) );
  AOI211_X1 U10661 ( .C1(n9434), .C2(n9442), .A(n9443), .B(n9433), .ZN(n9533)
         );
  NAND2_X1 U10662 ( .A1(n9533), .A2(n9450), .ZN(n9437) );
  AOI22_X1 U10663 ( .A1(n9749), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9435), .B2(
        n9758), .ZN(n9436) );
  OAI211_X1 U10664 ( .C1(n9605), .C2(n9444), .A(n9437), .B(n9436), .ZN(n9438)
         );
  AOI21_X1 U10665 ( .B1(n9457), .B2(n9532), .A(n9438), .ZN(n9439) );
  OAI21_X1 U10666 ( .B1(n9440), .B2(n9460), .A(n9439), .ZN(P1_U3275) );
  XNOR2_X1 U10667 ( .A(n9441), .B(n9452), .ZN(n9609) );
  AOI211_X1 U10668 ( .C1(n9540), .C2(n9475), .A(n9443), .B(n9431), .ZN(n9538)
         );
  NOR2_X1 U10669 ( .A1(n9445), .A2(n9444), .ZN(n9449) );
  OAI22_X1 U10670 ( .A1(n9457), .A2(n9447), .B1(n9446), .B2(n9471), .ZN(n9448)
         );
  AOI211_X1 U10671 ( .C1(n9538), .C2(n9450), .A(n9449), .B(n9448), .ZN(n9459)
         );
  OAI211_X1 U10672 ( .C1(n9453), .C2(n9452), .A(n9451), .B(n9463), .ZN(n9456)
         );
  INV_X1 U10673 ( .A(n9454), .ZN(n9455) );
  NAND2_X1 U10674 ( .A1(n9456), .A2(n9455), .ZN(n9539) );
  NAND2_X1 U10675 ( .A1(n9539), .A2(n9457), .ZN(n9458) );
  OAI211_X1 U10676 ( .C1(n9609), .C2(n9460), .A(n9459), .B(n9458), .ZN(
        P1_U3276) );
  NAND2_X1 U10677 ( .A1(n9461), .A2(n9468), .ZN(n9462) );
  NAND3_X1 U10678 ( .A1(n9464), .A2(n9463), .A3(n9462), .ZN(n9467) );
  INV_X1 U10679 ( .A(n9465), .ZN(n9466) );
  AND2_X1 U10680 ( .A1(n9467), .A2(n9466), .ZN(n9545) );
  XNOR2_X1 U10681 ( .A(n9469), .B(n9468), .ZN(n9614) );
  INV_X1 U10682 ( .A(n9614), .ZN(n9470) );
  NAND2_X1 U10683 ( .A1(n9470), .A2(n9754), .ZN(n9481) );
  OAI22_X1 U10684 ( .A1(n9474), .A2(n9473), .B1(n9472), .B2(n9471), .ZN(n9479)
         );
  OAI211_X1 U10685 ( .C1(n9477), .C2(n9476), .A(n9521), .B(n9475), .ZN(n9544)
         );
  NOR2_X1 U10686 ( .A1(n9544), .A2(n9765), .ZN(n9478) );
  AOI211_X1 U10687 ( .C1(n9762), .C2(n5476), .A(n9479), .B(n9478), .ZN(n9480)
         );
  OAI211_X1 U10688 ( .C1(n9749), .C2(n9545), .A(n9481), .B(n9480), .ZN(
        P1_U3277) );
  INV_X1 U10689 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9483) );
  MUX2_X1 U10690 ( .A(n9483), .B(n9555), .S(n9811), .Z(n9484) );
  OAI21_X1 U10691 ( .B1(n9558), .B2(n9537), .A(n9484), .ZN(P1_U3553) );
  INV_X1 U10692 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9487) );
  AND2_X1 U10693 ( .A1(n9486), .A2(n9485), .ZN(n9559) );
  MUX2_X1 U10694 ( .A(n9487), .B(n9559), .S(n9811), .Z(n9488) );
  OAI21_X1 U10695 ( .B1(n9562), .B2(n9537), .A(n9488), .ZN(P1_U3552) );
  NAND2_X1 U10696 ( .A1(n9563), .A2(n9551), .ZN(n9493) );
  AND2_X1 U10697 ( .A1(n9490), .A2(n9489), .ZN(n9564) );
  MUX2_X1 U10698 ( .A(n9491), .B(n9564), .S(n9811), .Z(n9492) );
  OAI211_X1 U10699 ( .C1(n9568), .C2(n9537), .A(n9493), .B(n9492), .ZN(
        P1_U3550) );
  OAI22_X1 U10700 ( .A1(n9570), .A2(n9548), .B1(n9569), .B2(n9537), .ZN(n9497)
         );
  NAND2_X1 U10701 ( .A1(n9495), .A2(n9494), .ZN(n9571) );
  MUX2_X1 U10702 ( .A(n9571), .B(P1_REG1_REG_26__SCAN_IN), .S(n9812), .Z(n9496) );
  OR2_X1 U10703 ( .A1(n9497), .A2(n9496), .ZN(P1_U3548) );
  AOI211_X1 U10704 ( .C1(n9541), .C2(n9500), .A(n9499), .B(n9498), .ZN(n9574)
         );
  MUX2_X1 U10705 ( .A(n9501), .B(n9574), .S(n9811), .Z(n9502) );
  OAI21_X1 U10706 ( .B1(n9577), .B2(n9548), .A(n9502), .ZN(P1_U3547) );
  OAI22_X1 U10707 ( .A1(n9578), .A2(n9548), .B1(n5480), .B2(n9537), .ZN(n9506)
         );
  NAND2_X1 U10708 ( .A1(n9504), .A2(n9503), .ZN(n9579) );
  MUX2_X1 U10709 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9579), .S(n9811), .Z(n9505) );
  OR2_X1 U10710 ( .A1(n9506), .A2(n9505), .ZN(P1_U3546) );
  INV_X1 U10711 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9509) );
  AOI211_X1 U10712 ( .C1(n9541), .C2(n5475), .A(n9508), .B(n9507), .ZN(n9582)
         );
  MUX2_X1 U10713 ( .A(n9509), .B(n9582), .S(n9811), .Z(n9510) );
  OAI21_X1 U10714 ( .B1(n9585), .B2(n9548), .A(n9510), .ZN(P1_U3545) );
  INV_X1 U10715 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9514) );
  AOI211_X1 U10716 ( .C1(n9541), .C2(n9513), .A(n9512), .B(n9511), .ZN(n9586)
         );
  MUX2_X1 U10717 ( .A(n9514), .B(n9586), .S(n9811), .Z(n9515) );
  OAI21_X1 U10718 ( .B1(n9589), .B2(n9548), .A(n9515), .ZN(P1_U3544) );
  INV_X1 U10719 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10021) );
  AOI211_X1 U10720 ( .C1(n9541), .C2(n9518), .A(n9517), .B(n9516), .ZN(n9590)
         );
  MUX2_X1 U10721 ( .A(n10021), .B(n9590), .S(n9811), .Z(n9519) );
  OAI21_X1 U10722 ( .B1(n9593), .B2(n9548), .A(n9519), .ZN(P1_U3543) );
  AOI22_X1 U10723 ( .A1(n9522), .A2(n9521), .B1(n9541), .B2(n9520), .ZN(n9523)
         );
  OAI211_X1 U10724 ( .C1(n9526), .C2(n9525), .A(n9524), .B(n9523), .ZN(n9594)
         );
  MUX2_X1 U10725 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9594), .S(n9811), .Z(
        P1_U3542) );
  AOI211_X1 U10726 ( .C1(n9541), .C2(n9529), .A(n9528), .B(n9527), .ZN(n9595)
         );
  MUX2_X1 U10727 ( .A(n9530), .B(n9595), .S(n9811), .Z(n9531) );
  OAI21_X1 U10728 ( .B1(n9598), .B2(n9548), .A(n9531), .ZN(P1_U3541) );
  NAND2_X1 U10729 ( .A1(n9599), .A2(n9551), .ZN(n9536) );
  NOR2_X1 U10730 ( .A1(n9533), .A2(n9532), .ZN(n9600) );
  MUX2_X1 U10731 ( .A(n9534), .B(n9600), .S(n9811), .Z(n9535) );
  OAI211_X1 U10732 ( .C1(n9605), .C2(n9537), .A(n9536), .B(n9535), .ZN(
        P1_U3540) );
  AOI211_X1 U10733 ( .C1(n9541), .C2(n9540), .A(n9539), .B(n9538), .ZN(n9606)
         );
  MUX2_X1 U10734 ( .A(n9542), .B(n9606), .S(n9811), .Z(n9543) );
  OAI21_X1 U10735 ( .B1(n9609), .B2(n9548), .A(n9543), .ZN(P1_U3539) );
  AOI22_X1 U10736 ( .A1(n5476), .A2(n9552), .B1(P1_REG1_REG_16__SCAN_IN), .B2(
        n9812), .ZN(n9547) );
  NAND2_X1 U10737 ( .A1(n9545), .A2(n9544), .ZN(n9610) );
  NAND2_X1 U10738 ( .A1(n9610), .A2(n9811), .ZN(n9546) );
  OAI211_X1 U10739 ( .C1(n9614), .C2(n9548), .A(n9547), .B(n9546), .ZN(
        P1_U3538) );
  NOR2_X1 U10740 ( .A1(n9550), .A2(n9549), .ZN(n9620) );
  NAND2_X1 U10741 ( .A1(n9615), .A2(n9551), .ZN(n9554) );
  AOI22_X1 U10742 ( .A1(n9616), .A2(n9552), .B1(P1_REG1_REG_15__SCAN_IN), .B2(
        n9812), .ZN(n9553) );
  OAI211_X1 U10743 ( .C1(n9620), .C2(n9812), .A(n9554), .B(n9553), .ZN(
        P1_U3537) );
  OAI21_X1 U10744 ( .B1(n9558), .B2(n9604), .A(n9557), .ZN(P1_U3521) );
  MUX2_X1 U10745 ( .A(n9560), .B(n9559), .S(n9795), .Z(n9561) );
  OAI21_X1 U10746 ( .B1(n9562), .B2(n9604), .A(n9561), .ZN(P1_U3520) );
  NAND2_X1 U10747 ( .A1(n9563), .A2(n5547), .ZN(n9567) );
  INV_X1 U10748 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9565) );
  MUX2_X1 U10749 ( .A(n9565), .B(n9564), .S(n9795), .Z(n9566) );
  OAI211_X1 U10750 ( .C1(n9568), .C2(n9604), .A(n9567), .B(n9566), .ZN(
        P1_U3518) );
  OAI22_X1 U10751 ( .A1(n9570), .A2(n9613), .B1(n9569), .B2(n9604), .ZN(n9573)
         );
  MUX2_X1 U10752 ( .A(n9571), .B(P1_REG0_REG_26__SCAN_IN), .S(n9619), .Z(n9572) );
  OR2_X1 U10753 ( .A1(n9573), .A2(n9572), .ZN(P1_U3516) );
  INV_X1 U10754 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9575) );
  MUX2_X1 U10755 ( .A(n9575), .B(n9574), .S(n9795), .Z(n9576) );
  OAI21_X1 U10756 ( .B1(n9577), .B2(n9613), .A(n9576), .ZN(P1_U3515) );
  OAI22_X1 U10757 ( .A1(n9578), .A2(n9613), .B1(n5480), .B2(n9604), .ZN(n9581)
         );
  MUX2_X1 U10758 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9579), .S(n9804), .Z(n9580) );
  OR2_X1 U10759 ( .A1(n9581), .A2(n9580), .ZN(P1_U3514) );
  MUX2_X1 U10760 ( .A(n9583), .B(n9582), .S(n9795), .Z(n9584) );
  OAI21_X1 U10761 ( .B1(n9585), .B2(n9613), .A(n9584), .ZN(P1_U3513) );
  MUX2_X1 U10762 ( .A(n9587), .B(n9586), .S(n9795), .Z(n9588) );
  OAI21_X1 U10763 ( .B1(n9589), .B2(n9613), .A(n9588), .ZN(P1_U3512) );
  INV_X1 U10764 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9591) );
  MUX2_X1 U10765 ( .A(n9591), .B(n9590), .S(n9804), .Z(n9592) );
  OAI21_X1 U10766 ( .B1(n9593), .B2(n9613), .A(n9592), .ZN(P1_U3511) );
  MUX2_X1 U10767 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9594), .S(n9804), .Z(
        P1_U3510) );
  MUX2_X1 U10768 ( .A(n9596), .B(n9595), .S(n9804), .Z(n9597) );
  OAI21_X1 U10769 ( .B1(n9598), .B2(n9613), .A(n9597), .ZN(P1_U3509) );
  NAND2_X1 U10770 ( .A1(n9599), .A2(n5547), .ZN(n9603) );
  INV_X1 U10771 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9601) );
  MUX2_X1 U10772 ( .A(n9601), .B(n9600), .S(n9804), .Z(n9602) );
  OAI211_X1 U10773 ( .C1(n9605), .C2(n9604), .A(n9603), .B(n9602), .ZN(
        P1_U3507) );
  MUX2_X1 U10774 ( .A(n9607), .B(n9606), .S(n9804), .Z(n9608) );
  OAI21_X1 U10775 ( .B1(n9609), .B2(n9613), .A(n9608), .ZN(P1_U3504) );
  AOI22_X1 U10776 ( .A1(n5476), .A2(n6071), .B1(P1_REG0_REG_16__SCAN_IN), .B2(
        n9619), .ZN(n9612) );
  NAND2_X1 U10777 ( .A1(n9610), .A2(n9795), .ZN(n9611) );
  OAI211_X1 U10778 ( .C1(n9614), .C2(n9613), .A(n9612), .B(n9611), .ZN(
        P1_U3501) );
  NAND2_X1 U10779 ( .A1(n9615), .A2(n5547), .ZN(n9618) );
  AOI22_X1 U10780 ( .A1(n9616), .A2(n6071), .B1(P1_REG0_REG_15__SCAN_IN), .B2(
        n9619), .ZN(n9617) );
  OAI211_X1 U10781 ( .C1(n9620), .C2(n9619), .A(n9618), .B(n9617), .ZN(
        P1_U3498) );
  NOR4_X1 U10782 ( .A1(n4994), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9621), .A4(
        P1_U3086), .ZN(n9622) );
  AOI21_X1 U10783 ( .B1(n9634), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9622), .ZN(
        n9623) );
  OAI21_X1 U10784 ( .B1(n9624), .B2(n9637), .A(n9623), .ZN(P1_U3324) );
  AOI22_X1 U10785 ( .A1(n4799), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9634), .ZN(n9625) );
  OAI21_X1 U10786 ( .B1(n9627), .B2(n9626), .A(n9625), .ZN(P1_U3325) );
  AOI22_X1 U10787 ( .A1(n9628), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n9634), .ZN(n9629) );
  OAI21_X1 U10788 ( .B1(n9630), .B2(n9637), .A(n9629), .ZN(P1_U3326) );
  AOI22_X1 U10789 ( .A1(n9631), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n9634), .ZN(n9632) );
  OAI21_X1 U10790 ( .B1(n9633), .B2(n9637), .A(n9632), .ZN(P1_U3327) );
  AOI22_X1 U10791 ( .A1(n9635), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n9634), .ZN(n9636) );
  OAI21_X1 U10792 ( .B1(n9638), .B2(n9637), .A(n9636), .ZN(P1_U3328) );
  INV_X1 U10793 ( .A(n9639), .ZN(n9640) );
  MUX2_X1 U10794 ( .A(n9640), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI211_X1 U10795 ( .C1(n9643), .C2(n9642), .A(n9641), .B(n9730), .ZN(n9648)
         );
  AOI211_X1 U10796 ( .C1(n9646), .C2(n9645), .A(n9644), .B(n9718), .ZN(n9647)
         );
  AOI211_X1 U10797 ( .C1(n9726), .C2(n9649), .A(n9648), .B(n9647), .ZN(n9651)
         );
  NAND2_X1 U10798 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n9650) );
  OAI211_X1 U10799 ( .C1(n9746), .C2(n9652), .A(n9651), .B(n9650), .ZN(
        P1_U3253) );
  XOR2_X1 U10800 ( .A(n9659), .B(n9653), .Z(n9674) );
  NAND2_X1 U10801 ( .A1(n9654), .A2(n9872), .ZN(n9671) );
  INV_X1 U10802 ( .A(n9655), .ZN(n9657) );
  OAI22_X1 U10803 ( .A1(n9671), .A2(n9658), .B1(n9657), .B2(n9656), .ZN(n9666)
         );
  XNOR2_X1 U10804 ( .A(n9660), .B(n9659), .ZN(n9661) );
  OAI222_X1 U10805 ( .A1(n9665), .A2(n9664), .B1(n9663), .B2(n9662), .C1(n9661), .C2(n9815), .ZN(n9672) );
  AOI211_X1 U10806 ( .C1(n9674), .C2(n9667), .A(n9666), .B(n9672), .ZN(n9669)
         );
  AOI22_X1 U10807 ( .A1(n9670), .A2(n9964), .B1(n9669), .B2(n9668), .ZN(
        P2_U3220) );
  INV_X1 U10808 ( .A(n9671), .ZN(n9673) );
  AOI211_X1 U10809 ( .C1(n9674), .C2(n9835), .A(n9673), .B(n9672), .ZN(n9675)
         );
  AOI22_X1 U10810 ( .A1(n9890), .A2(n9675), .B1(n7689), .B2(n8746), .ZN(
        P2_U3472) );
  INV_X1 U10811 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9676) );
  AOI22_X1 U10812 ( .A1(n9875), .A2(n9676), .B1(n9675), .B2(n9873), .ZN(
        P2_U3429) );
  XNOR2_X1 U10813 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X1 U10814 ( .A(n9677), .ZN(n9689) );
  AOI21_X1 U10815 ( .B1(n9680), .B2(n9679), .A(n9678), .ZN(n9681) );
  NAND2_X1 U10816 ( .A1(n9682), .A2(n9681), .ZN(n9688) );
  AOI21_X1 U10817 ( .B1(n9685), .B2(n9684), .A(n9683), .ZN(n9686) );
  NAND2_X1 U10818 ( .A1(n9733), .A2(n9686), .ZN(n9687) );
  OAI211_X1 U10819 ( .C1(n9739), .C2(n9689), .A(n9688), .B(n9687), .ZN(n9690)
         );
  INV_X1 U10820 ( .A(n9690), .ZN(n9692) );
  NAND2_X1 U10821 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9691) );
  OAI211_X1 U10822 ( .C1(n9746), .C2(n9693), .A(n9692), .B(n9691), .ZN(
        P1_U3254) );
  AOI211_X1 U10823 ( .C1(n9696), .C2(n9695), .A(n9718), .B(n9694), .ZN(n9701)
         );
  AOI211_X1 U10824 ( .C1(n9699), .C2(n9698), .A(n9730), .B(n9697), .ZN(n9700)
         );
  AOI211_X1 U10825 ( .C1(n9726), .C2(n9702), .A(n9701), .B(n9700), .ZN(n9704)
         );
  OAI211_X1 U10826 ( .C1(n9746), .C2(n9705), .A(n9704), .B(n9703), .ZN(
        P1_U3256) );
  AOI211_X1 U10827 ( .C1(n9708), .C2(n9707), .A(n9706), .B(n9730), .ZN(n9713)
         );
  AOI211_X1 U10828 ( .C1(n9711), .C2(n9710), .A(n9718), .B(n9709), .ZN(n9712)
         );
  AOI211_X1 U10829 ( .C1(n9726), .C2(n9714), .A(n9713), .B(n9712), .ZN(n9716)
         );
  OAI211_X1 U10830 ( .C1(n9746), .C2(n9965), .A(n9716), .B(n9715), .ZN(
        P1_U3257) );
  INV_X1 U10831 ( .A(n9717), .ZN(n9725) );
  AOI211_X1 U10832 ( .C1(n9720), .C2(n10024), .A(n9719), .B(n9718), .ZN(n9724)
         );
  AOI211_X1 U10833 ( .C1(n9722), .C2(n7887), .A(n9721), .B(n9730), .ZN(n9723)
         );
  AOI211_X1 U10834 ( .C1(n9726), .C2(n9725), .A(n9724), .B(n9723), .ZN(n9728)
         );
  OAI211_X1 U10835 ( .C1(n9746), .C2(n9729), .A(n9728), .B(n9727), .ZN(
        P1_U3258) );
  INV_X1 U10836 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9745) );
  AOI21_X1 U10837 ( .B1(n9732), .B2(n9731), .A(n9730), .ZN(n9742) );
  OAI211_X1 U10838 ( .C1(n9736), .C2(n9735), .A(n9734), .B(n9733), .ZN(n9737)
         );
  OAI21_X1 U10839 ( .B1(n9739), .B2(n9738), .A(n9737), .ZN(n9740) );
  AOI21_X1 U10840 ( .B1(n9742), .B2(n9741), .A(n9740), .ZN(n9744) );
  NAND2_X1 U10841 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9743) );
  OAI211_X1 U10842 ( .C1(n9746), .C2(n9745), .A(n9744), .B(n9743), .ZN(
        P1_U3261) );
  NAND2_X1 U10843 ( .A1(n9762), .A2(n9747), .ZN(n9751) );
  AOI22_X1 U10844 ( .A1(n9749), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9758), .B2(
        n9748), .ZN(n9750) );
  OAI211_X1 U10845 ( .C1(n9752), .C2(n9765), .A(n9751), .B(n9750), .ZN(n9753)
         );
  AOI21_X1 U10846 ( .B1(n9755), .B2(n9754), .A(n9753), .ZN(n9756) );
  OAI21_X1 U10847 ( .B1(n9749), .B2(n9757), .A(n9756), .ZN(P1_U3290) );
  AOI22_X1 U10848 ( .A1(n9758), .A2(P1_REG3_REG_1__SCAN_IN), .B1(
        P1_REG2_REG_1__SCAN_IN), .B2(n9749), .ZN(n9769) );
  NAND2_X1 U10849 ( .A1(n9760), .A2(n9759), .ZN(n9764) );
  NAND2_X1 U10850 ( .A1(n9762), .A2(n9761), .ZN(n9763) );
  OAI211_X1 U10851 ( .C1(n9766), .C2(n9765), .A(n9764), .B(n9763), .ZN(n9767)
         );
  INV_X1 U10852 ( .A(n9767), .ZN(n9768) );
  OAI211_X1 U10853 ( .C1(n9749), .C2(n9770), .A(n9769), .B(n9768), .ZN(
        P1_U3292) );
  AND2_X1 U10854 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9772), .ZN(P1_U3294) );
  AND2_X1 U10855 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9772), .ZN(P1_U3295) );
  INV_X1 U10856 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n9977) );
  NOR2_X1 U10857 ( .A1(n9771), .A2(n9977), .ZN(P1_U3296) );
  AND2_X1 U10858 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9772), .ZN(P1_U3297) );
  AND2_X1 U10859 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9772), .ZN(P1_U3298) );
  INV_X1 U10860 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10022) );
  NOR2_X1 U10861 ( .A1(n9771), .A2(n10022), .ZN(P1_U3299) );
  AND2_X1 U10862 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9772), .ZN(P1_U3300) );
  AND2_X1 U10863 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9772), .ZN(P1_U3301) );
  INV_X1 U10864 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n9981) );
  NOR2_X1 U10865 ( .A1(n9771), .A2(n9981), .ZN(P1_U3302) );
  AND2_X1 U10866 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9772), .ZN(P1_U3303) );
  INV_X1 U10867 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10049) );
  NOR2_X1 U10868 ( .A1(n9771), .A2(n10049), .ZN(P1_U3304) );
  INV_X1 U10869 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9984) );
  NOR2_X1 U10870 ( .A1(n9771), .A2(n9984), .ZN(P1_U3305) );
  AND2_X1 U10871 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9772), .ZN(P1_U3306) );
  AND2_X1 U10872 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9772), .ZN(P1_U3307) );
  AND2_X1 U10873 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9772), .ZN(P1_U3308) );
  AND2_X1 U10874 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9772), .ZN(P1_U3309) );
  AND2_X1 U10875 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9772), .ZN(P1_U3310) );
  AND2_X1 U10876 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9772), .ZN(P1_U3311) );
  AND2_X1 U10877 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9772), .ZN(P1_U3312) );
  AND2_X1 U10878 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9772), .ZN(P1_U3313) );
  AND2_X1 U10879 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9772), .ZN(P1_U3314) );
  AND2_X1 U10880 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9772), .ZN(P1_U3315) );
  AND2_X1 U10881 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9772), .ZN(P1_U3316) );
  INV_X1 U10882 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n9952) );
  NOR2_X1 U10883 ( .A1(n9771), .A2(n9952), .ZN(P1_U3317) );
  AND2_X1 U10884 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9772), .ZN(P1_U3318) );
  AND2_X1 U10885 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9772), .ZN(P1_U3319) );
  AND2_X1 U10886 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9772), .ZN(P1_U3320) );
  AND2_X1 U10887 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9772), .ZN(P1_U3321) );
  AND2_X1 U10888 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9772), .ZN(P1_U3322) );
  AND2_X1 U10889 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9772), .ZN(P1_U3323) );
  INV_X1 U10890 ( .A(n9773), .ZN(n9774) );
  OAI21_X1 U10891 ( .B1(n9775), .B2(n9798), .A(n9774), .ZN(n9777) );
  AOI211_X1 U10892 ( .C1(n9779), .C2(n9778), .A(n9777), .B(n9776), .ZN(n9806)
         );
  AOI22_X1 U10893 ( .A1(n9804), .A2(n9806), .B1(n5107), .B2(n9619), .ZN(
        P1_U3459) );
  OAI21_X1 U10894 ( .B1(n9781), .B2(n9798), .A(n9780), .ZN(n9783) );
  AOI211_X1 U10895 ( .C1(n9801), .C2(n9784), .A(n9783), .B(n9782), .ZN(n9807)
         );
  INV_X1 U10896 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9993) );
  AOI22_X1 U10897 ( .A1(n9795), .A2(n9807), .B1(n9993), .B2(n9619), .ZN(
        P1_U3471) );
  OAI211_X1 U10898 ( .C1(n9787), .C2(n9798), .A(n9786), .B(n9785), .ZN(n9788)
         );
  AOI21_X1 U10899 ( .B1(n9801), .B2(n9789), .A(n9788), .ZN(n9809) );
  AOI22_X1 U10900 ( .A1(n9795), .A2(n9809), .B1(n5227), .B2(n9619), .ZN(
        P1_U3480) );
  OAI211_X1 U10901 ( .C1(n9792), .C2(n9798), .A(n9791), .B(n9790), .ZN(n9793)
         );
  AOI21_X1 U10902 ( .B1(n9794), .B2(n9801), .A(n9793), .ZN(n9810) );
  AOI22_X1 U10903 ( .A1(n9795), .A2(n9810), .B1(n5244), .B2(n9619), .ZN(
        P1_U3483) );
  OAI211_X1 U10904 ( .C1(n9799), .C2(n9798), .A(n9797), .B(n9796), .ZN(n9800)
         );
  AOI21_X1 U10905 ( .B1(n9802), .B2(n9801), .A(n9800), .ZN(n9813) );
  INV_X1 U10906 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9803) );
  AOI22_X1 U10907 ( .A1(n9804), .A2(n9813), .B1(n9803), .B2(n9619), .ZN(
        P1_U3489) );
  INV_X1 U10908 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9805) );
  AOI22_X1 U10909 ( .A1(n9811), .A2(n9806), .B1(n9805), .B2(n9812), .ZN(
        P1_U3524) );
  AOI22_X1 U10910 ( .A1(n9811), .A2(n9807), .B1(n6404), .B2(n9812), .ZN(
        P1_U3528) );
  INV_X1 U10911 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9808) );
  AOI22_X1 U10912 ( .A1(n9811), .A2(n9809), .B1(n9808), .B2(n9812), .ZN(
        P1_U3531) );
  INV_X1 U10913 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9949) );
  AOI22_X1 U10914 ( .A1(n9811), .A2(n9810), .B1(n9949), .B2(n9812), .ZN(
        P1_U3532) );
  AOI22_X1 U10915 ( .A1(n9811), .A2(n9813), .B1(n5276), .B2(n9812), .ZN(
        P1_U3534) );
  INV_X1 U10916 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9819) );
  AOI21_X1 U10917 ( .B1(n9815), .B2(n9867), .A(n9814), .ZN(n9816) );
  AOI211_X1 U10918 ( .C1(n9872), .C2(n9818), .A(n9817), .B(n9816), .ZN(n9876)
         );
  AOI22_X1 U10919 ( .A1(n9875), .A2(n9819), .B1(n9876), .B2(n9873), .ZN(
        P2_U3390) );
  INV_X1 U10920 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9825) );
  INV_X1 U10921 ( .A(n9820), .ZN(n9822) );
  AOI211_X1 U10922 ( .C1(n9824), .C2(n9823), .A(n9822), .B(n9821), .ZN(n9878)
         );
  AOI22_X1 U10923 ( .A1(n9875), .A2(n9825), .B1(n9878), .B2(n9873), .ZN(
        P2_U3396) );
  INV_X1 U10924 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9830) );
  OAI21_X1 U10925 ( .B1(n9827), .B2(n9842), .A(n9826), .ZN(n9828) );
  AOI21_X1 U10926 ( .B1(n9829), .B2(n9835), .A(n9828), .ZN(n9880) );
  AOI22_X1 U10927 ( .A1(n9875), .A2(n9830), .B1(n9880), .B2(n9873), .ZN(
        P2_U3402) );
  INV_X1 U10928 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9836) );
  OAI21_X1 U10929 ( .B1(n9832), .B2(n9842), .A(n9831), .ZN(n9833) );
  AOI21_X1 U10930 ( .B1(n9835), .B2(n9834), .A(n9833), .ZN(n9881) );
  AOI22_X1 U10931 ( .A1(n9875), .A2(n9836), .B1(n9881), .B2(n9873), .ZN(
        P2_U3405) );
  INV_X1 U10932 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9841) );
  NOR2_X1 U10933 ( .A1(n9837), .A2(n9867), .ZN(n9838) );
  AOI211_X1 U10934 ( .C1(n9872), .C2(n9840), .A(n9839), .B(n9838), .ZN(n9882)
         );
  AOI22_X1 U10935 ( .A1(n9875), .A2(n9841), .B1(n9882), .B2(n9873), .ZN(
        P2_U3408) );
  INV_X1 U10936 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9983) );
  OAI22_X1 U10937 ( .A1(n9844), .A2(n9852), .B1(n9843), .B2(n9842), .ZN(n9845)
         );
  NOR2_X1 U10938 ( .A1(n9846), .A2(n9845), .ZN(n9883) );
  AOI22_X1 U10939 ( .A1(n9875), .A2(n9983), .B1(n9883), .B2(n9873), .ZN(
        P2_U3411) );
  INV_X1 U10940 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9851) );
  NOR2_X1 U10941 ( .A1(n9847), .A2(n9867), .ZN(n9848) );
  AOI211_X1 U10942 ( .C1(n9872), .C2(n9850), .A(n9849), .B(n9848), .ZN(n9885)
         );
  AOI22_X1 U10943 ( .A1(n9875), .A2(n9851), .B1(n9885), .B2(n9873), .ZN(
        P2_U3414) );
  INV_X1 U10944 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10039) );
  NOR2_X1 U10945 ( .A1(n9853), .A2(n9852), .ZN(n9855) );
  AOI211_X1 U10946 ( .C1(n9872), .C2(n9856), .A(n9855), .B(n9854), .ZN(n9886)
         );
  AOI22_X1 U10947 ( .A1(n9875), .A2(n10039), .B1(n9886), .B2(n9873), .ZN(
        P2_U3417) );
  INV_X1 U10948 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9861) );
  NOR2_X1 U10949 ( .A1(n9857), .A2(n9867), .ZN(n9859) );
  AOI211_X1 U10950 ( .C1(n9872), .C2(n9860), .A(n9859), .B(n9858), .ZN(n9887)
         );
  AOI22_X1 U10951 ( .A1(n9875), .A2(n9861), .B1(n9887), .B2(n9873), .ZN(
        P2_U3420) );
  INV_X1 U10952 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9866) );
  NOR2_X1 U10953 ( .A1(n9862), .A2(n9867), .ZN(n9863) );
  AOI211_X1 U10954 ( .C1(n9872), .C2(n9865), .A(n9864), .B(n9863), .ZN(n9888)
         );
  AOI22_X1 U10955 ( .A1(n9875), .A2(n9866), .B1(n9888), .B2(n9873), .ZN(
        P2_U3423) );
  INV_X1 U10956 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9874) );
  NOR2_X1 U10957 ( .A1(n9868), .A2(n9867), .ZN(n9869) );
  AOI211_X1 U10958 ( .C1(n9872), .C2(n9871), .A(n9870), .B(n9869), .ZN(n9889)
         );
  AOI22_X1 U10959 ( .A1(n9875), .A2(n9874), .B1(n9889), .B2(n9873), .ZN(
        P2_U3426) );
  AOI22_X1 U10960 ( .A1(n9890), .A2(n9876), .B1(n6466), .B2(n8746), .ZN(
        P2_U3459) );
  AOI22_X1 U10961 ( .A1(n9890), .A2(n9878), .B1(n9877), .B2(n8746), .ZN(
        P2_U3461) );
  AOI22_X1 U10962 ( .A1(n9890), .A2(n9880), .B1(n9879), .B2(n8746), .ZN(
        P2_U3463) );
  AOI22_X1 U10963 ( .A1(n9890), .A2(n9881), .B1(n6792), .B2(n8746), .ZN(
        P2_U3464) );
  AOI22_X1 U10964 ( .A1(n9890), .A2(n9882), .B1(n10048), .B2(n8746), .ZN(
        P2_U3465) );
  AOI22_X1 U10965 ( .A1(n9890), .A2(n9883), .B1(n6812), .B2(n8746), .ZN(
        P2_U3466) );
  AOI22_X1 U10966 ( .A1(n9890), .A2(n9885), .B1(n9884), .B2(n8746), .ZN(
        P2_U3467) );
  AOI22_X1 U10967 ( .A1(n9890), .A2(n9886), .B1(n7027), .B2(n8746), .ZN(
        P2_U3468) );
  AOI22_X1 U10968 ( .A1(n9890), .A2(n9887), .B1(n7140), .B2(n8746), .ZN(
        P2_U3469) );
  AOI22_X1 U10969 ( .A1(n9890), .A2(n9888), .B1(n7345), .B2(n8746), .ZN(
        P2_U3470) );
  AOI22_X1 U10970 ( .A1(n9890), .A2(n9889), .B1(n10012), .B2(n8746), .ZN(
        P2_U3471) );
  NOR2_X1 U10971 ( .A1(n9892), .A2(n9891), .ZN(n9893) );
  XOR2_X1 U10972 ( .A(n9893), .B(P2_ADDR_REG_1__SCAN_IN), .Z(ADD_1068_U5) );
  XOR2_X1 U10973 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U10974 ( .A1(n9895), .A2(n9894), .ZN(n9896) );
  XOR2_X1 U10975 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n9896), .Z(ADD_1068_U55) );
  XNOR2_X1 U10976 ( .A(n9898), .B(n9897), .ZN(ADD_1068_U56) );
  XNOR2_X1 U10977 ( .A(n9900), .B(n9899), .ZN(ADD_1068_U57) );
  XNOR2_X1 U10978 ( .A(n9902), .B(n9901), .ZN(ADD_1068_U58) );
  XNOR2_X1 U10979 ( .A(n9904), .B(n9903), .ZN(ADD_1068_U59) );
  XNOR2_X1 U10980 ( .A(n9906), .B(n9905), .ZN(ADD_1068_U60) );
  XNOR2_X1 U10981 ( .A(n9908), .B(n9907), .ZN(ADD_1068_U61) );
  XNOR2_X1 U10982 ( .A(n9910), .B(n9909), .ZN(ADD_1068_U62) );
  XNOR2_X1 U10983 ( .A(n9912), .B(n9911), .ZN(ADD_1068_U63) );
  NAND4_X1 U10984 ( .A1(P1_REG0_REG_17__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .A3(P2_REG1_REG_6__SCAN_IN), .A4(n10052), .ZN(n9915) );
  NAND3_X1 U10985 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(P1_REG2_REG_18__SCAN_IN), 
        .A3(n10057), .ZN(n9914) );
  NAND4_X1 U10986 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(SI_17_), .A3(
        P2_REG0_REG_9__SCAN_IN), .A4(n10037), .ZN(n9913) );
  NOR4_X1 U10987 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n9915), .A3(n9914), .A4(
        n9913), .ZN(n9944) );
  NOR4_X1 U10988 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), 
        .A3(P2_REG1_REG_1__SCAN_IN), .A4(n4881), .ZN(n9943) );
  AND2_X1 U10989 ( .A1(n9917), .A2(n9916), .ZN(n9942) );
  NAND4_X1 U10990 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P2_REG2_REG_4__SCAN_IN), 
        .A3(n9951), .A4(n9947), .ZN(n9919) );
  NAND4_X1 U10991 ( .A1(P1_REG0_REG_24__SCAN_IN), .A2(P2_REG1_REG_16__SCAN_IN), 
        .A3(n8247), .A4(n8114), .ZN(n9918) );
  NOR2_X1 U10992 ( .A1(n9919), .A2(n9918), .ZN(n9936) );
  NAND4_X1 U10993 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), .A3(P2_REG2_REG_13__SCAN_IN), .A4(P1_ADDR_REG_14__SCAN_IN), .ZN(n9920) );
  NOR2_X1 U10994 ( .A1(n9991), .A2(n9920), .ZN(n9935) );
  NAND4_X1 U10995 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .A3(
        P2_DATAO_REG_14__SCAN_IN), .A4(P2_REG3_REG_22__SCAN_IN), .ZN(n9921) );
  NOR2_X1 U10996 ( .A1(n10012), .A2(n9921), .ZN(n9922) );
  AND2_X1 U10997 ( .A1(n9922), .A2(n9949), .ZN(n9923) );
  NAND4_X1 U10998 ( .A1(n9925), .A2(n9924), .A3(SI_3_), .A4(n9923), .ZN(n9927)
         );
  NAND4_X1 U10999 ( .A1(n4806), .A2(n9978), .A3(P2_IR_REG_16__SCAN_IN), .A4(
        P2_REG1_REG_10__SCAN_IN), .ZN(n9926) );
  NOR2_X1 U11000 ( .A1(n9927), .A2(n9926), .ZN(n9934) );
  INV_X1 U11001 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10025) );
  NAND4_X1 U11002 ( .A1(n9929), .A2(n10025), .A3(n9928), .A4(
        P2_REG3_REG_10__SCAN_IN), .ZN(n9932) );
  NAND4_X1 U11003 ( .A1(n10021), .A2(n10024), .A3(n9930), .A4(
        P1_REG0_REG_3__SCAN_IN), .ZN(n9931) );
  NOR2_X1 U11004 ( .A1(n9932), .A2(n9931), .ZN(n9933) );
  NAND4_X1 U11005 ( .A1(n9936), .A2(n9935), .A3(n9934), .A4(n9933), .ZN(n9940)
         );
  AND4_X1 U11006 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_REG0_REG_20__SCAN_IN), 
        .A3(P2_REG0_REG_7__SCAN_IN), .A4(n9977), .ZN(n9938) );
  INV_X1 U11007 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9994) );
  AND4_X1 U11008 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .A3(n9994), .A4(n9993), .ZN(n9937) );
  NAND4_X1 U11009 ( .A1(n9938), .A2(n9937), .A3(P2_D_REG_6__SCAN_IN), .A4(
        n10022), .ZN(n9939) );
  NOR2_X1 U11010 ( .A1(n9940), .A2(n9939), .ZN(n9941) );
  AND4_X1 U11011 ( .A1(n9944), .A2(n9943), .A3(n9942), .A4(n9941), .ZN(n9945)
         );
  XOR2_X1 U11012 ( .A(P2_RD_REG_SCAN_IN), .B(n9945), .Z(n10069) );
  AOI22_X1 U11013 ( .A1(n6750), .A2(keyinput57), .B1(keyinput19), .B2(n9947), 
        .ZN(n9946) );
  OAI221_X1 U11014 ( .B1(n6750), .B2(keyinput57), .C1(n9947), .C2(keyinput19), 
        .A(n9946), .ZN(n9958) );
  AOI22_X1 U11015 ( .A1(n7140), .A2(keyinput46), .B1(n9949), .B2(keyinput42), 
        .ZN(n9948) );
  OAI221_X1 U11016 ( .B1(n7140), .B2(keyinput46), .C1(n9949), .C2(keyinput42), 
        .A(n9948), .ZN(n9957) );
  AOI22_X1 U11017 ( .A1(n9952), .A2(keyinput16), .B1(keyinput17), .B2(n9951), 
        .ZN(n9950) );
  OAI221_X1 U11018 ( .B1(n9952), .B2(keyinput16), .C1(n9951), .C2(keyinput17), 
        .A(n9950), .ZN(n9956) );
  XOR2_X1 U11019 ( .A(n5121), .B(keyinput44), .Z(n9954) );
  XNOR2_X1 U11020 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput48), .ZN(n9953) );
  NAND2_X1 U11021 ( .A1(n9954), .A2(n9953), .ZN(n9955) );
  NOR4_X1 U11022 ( .A1(n9958), .A2(n9957), .A3(n9956), .A4(n9955), .ZN(n10007)
         );
  AOI22_X1 U11023 ( .A1(n8114), .A2(keyinput33), .B1(n9960), .B2(keyinput55), 
        .ZN(n9959) );
  OAI221_X1 U11024 ( .B1(n8114), .B2(keyinput33), .C1(n9960), .C2(keyinput55), 
        .A(n9959), .ZN(n9972) );
  AOI22_X1 U11025 ( .A1(n9962), .A2(keyinput56), .B1(keyinput43), .B2(n8247), 
        .ZN(n9961) );
  OAI221_X1 U11026 ( .B1(n9962), .B2(keyinput56), .C1(n8247), .C2(keyinput43), 
        .A(n9961), .ZN(n9971) );
  AOI22_X1 U11027 ( .A1(n9965), .A2(keyinput36), .B1(n9964), .B2(keyinput59), 
        .ZN(n9963) );
  OAI221_X1 U11028 ( .B1(n9965), .B2(keyinput36), .C1(n9964), .C2(keyinput59), 
        .A(n9963), .ZN(n9970) );
  AOI22_X1 U11029 ( .A1(n9968), .A2(keyinput62), .B1(keyinput45), .B2(n9967), 
        .ZN(n9966) );
  OAI221_X1 U11030 ( .B1(n9968), .B2(keyinput62), .C1(n9967), .C2(keyinput45), 
        .A(n9966), .ZN(n9969) );
  NOR4_X1 U11031 ( .A1(n9972), .A2(n9971), .A3(n9970), .A4(n9969), .ZN(n10006)
         );
  AOI22_X1 U11032 ( .A1(n9975), .A2(keyinput24), .B1(keyinput10), .B2(n9974), 
        .ZN(n9973) );
  OAI221_X1 U11033 ( .B1(n9975), .B2(keyinput24), .C1(n9974), .C2(keyinput10), 
        .A(n9973), .ZN(n9988) );
  AOI22_X1 U11034 ( .A1(n9978), .A2(keyinput54), .B1(n9977), .B2(keyinput23), 
        .ZN(n9976) );
  OAI221_X1 U11035 ( .B1(n9978), .B2(keyinput54), .C1(n9977), .C2(keyinput23), 
        .A(n9976), .ZN(n9987) );
  INV_X1 U11036 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9980) );
  AOI22_X1 U11037 ( .A1(n9981), .A2(keyinput9), .B1(keyinput63), .B2(n9980), 
        .ZN(n9979) );
  OAI221_X1 U11038 ( .B1(n9981), .B2(keyinput9), .C1(n9980), .C2(keyinput63), 
        .A(n9979), .ZN(n9986) );
  AOI22_X1 U11039 ( .A1(n9984), .A2(keyinput7), .B1(keyinput2), .B2(n9983), 
        .ZN(n9982) );
  OAI221_X1 U11040 ( .B1(n9984), .B2(keyinput7), .C1(n9983), .C2(keyinput2), 
        .A(n9982), .ZN(n9985) );
  NOR4_X1 U11041 ( .A1(n9988), .A2(n9987), .A3(n9986), .A4(n9985), .ZN(n10005)
         );
  AOI22_X1 U11042 ( .A1(n9991), .A2(keyinput47), .B1(n9990), .B2(keyinput35), 
        .ZN(n9989) );
  OAI221_X1 U11043 ( .B1(n9991), .B2(keyinput47), .C1(n9990), .C2(keyinput35), 
        .A(n9989), .ZN(n10003) );
  AOI22_X1 U11044 ( .A1(n9994), .A2(keyinput28), .B1(n9993), .B2(keyinput58), 
        .ZN(n9992) );
  OAI221_X1 U11045 ( .B1(n9994), .B2(keyinput28), .C1(n9993), .C2(keyinput58), 
        .A(n9992), .ZN(n10002) );
  AOI22_X1 U11046 ( .A1(n9997), .A2(keyinput32), .B1(n9996), .B2(keyinput1), 
        .ZN(n9995) );
  OAI221_X1 U11047 ( .B1(n9997), .B2(keyinput32), .C1(n9996), .C2(keyinput1), 
        .A(n9995), .ZN(n10001) );
  XNOR2_X1 U11048 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput12), .ZN(n9999)
         );
  XNOR2_X1 U11049 ( .A(SI_2_), .B(keyinput5), .ZN(n9998) );
  NAND2_X1 U11050 ( .A1(n9999), .A2(n9998), .ZN(n10000) );
  NOR4_X1 U11051 ( .A1(n10003), .A2(n10002), .A3(n10001), .A4(n10000), .ZN(
        n10004) );
  NAND4_X1 U11052 ( .A1(n10007), .A2(n10006), .A3(n10005), .A4(n10004), .ZN(
        n10067) );
  AOI22_X1 U11053 ( .A1(n6645), .A2(keyinput26), .B1(n10009), .B2(keyinput14), 
        .ZN(n10008) );
  OAI221_X1 U11054 ( .B1(n6645), .B2(keyinput26), .C1(n10009), .C2(keyinput14), 
        .A(n10008), .ZN(n10019) );
  AOI22_X1 U11055 ( .A1(n5581), .A2(keyinput39), .B1(n10011), .B2(keyinput31), 
        .ZN(n10010) );
  OAI221_X1 U11056 ( .B1(n5581), .B2(keyinput39), .C1(n10011), .C2(keyinput31), 
        .A(n10010), .ZN(n10018) );
  XOR2_X1 U11057 ( .A(n10012), .B(keyinput34), .Z(n10016) );
  XNOR2_X1 U11058 ( .A(P1_REG0_REG_17__SCAN_IN), .B(keyinput6), .ZN(n10015) );
  XNOR2_X1 U11059 ( .A(P1_REG3_REG_2__SCAN_IN), .B(keyinput3), .ZN(n10014) );
  XNOR2_X1 U11060 ( .A(SI_3_), .B(keyinput37), .ZN(n10013) );
  NAND4_X1 U11061 ( .A1(n10016), .A2(n10015), .A3(n10014), .A4(n10013), .ZN(
        n10017) );
  NOR3_X1 U11062 ( .A1(n10019), .A2(n10018), .A3(n10017), .ZN(n10065) );
  AOI22_X1 U11063 ( .A1(n10022), .A2(keyinput29), .B1(keyinput20), .B2(n10021), 
        .ZN(n10020) );
  OAI221_X1 U11064 ( .B1(n10022), .B2(keyinput29), .C1(n10021), .C2(keyinput20), .A(n10020), .ZN(n10032) );
  AOI22_X1 U11065 ( .A1(n10025), .A2(keyinput4), .B1(keyinput38), .B2(n10024), 
        .ZN(n10023) );
  OAI221_X1 U11066 ( .B1(n10025), .B2(keyinput4), .C1(n10024), .C2(keyinput38), 
        .A(n10023), .ZN(n10031) );
  XOR2_X1 U11067 ( .A(n4881), .B(keyinput25), .Z(n10029) );
  XNOR2_X1 U11068 ( .A(P1_REG3_REG_27__SCAN_IN), .B(keyinput0), .ZN(n10028) );
  XNOR2_X1 U11069 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput40), .ZN(n10027) );
  NAND4_X1 U11070 ( .A1(n10029), .A2(n10028), .A3(n10027), .A4(n10026), .ZN(
        n10030) );
  NOR3_X1 U11071 ( .A1(n10032), .A2(n10031), .A3(n10030), .ZN(n10064) );
  AOI22_X1 U11072 ( .A1(n10035), .A2(keyinput13), .B1(keyinput52), .B2(n10034), 
        .ZN(n10033) );
  OAI221_X1 U11073 ( .B1(n10035), .B2(keyinput13), .C1(n10034), .C2(keyinput52), .A(n10033), .ZN(n10046) );
  AOI22_X1 U11074 ( .A1(n10038), .A2(keyinput11), .B1(keyinput22), .B2(n10037), 
        .ZN(n10036) );
  OAI221_X1 U11075 ( .B1(n10038), .B2(keyinput11), .C1(n10037), .C2(keyinput22), .A(n10036), .ZN(n10045) );
  XOR2_X1 U11076 ( .A(n10039), .B(keyinput21), .Z(n10043) );
  XNOR2_X1 U11077 ( .A(P1_REG3_REG_4__SCAN_IN), .B(keyinput15), .ZN(n10042) );
  XNOR2_X1 U11078 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput49), .ZN(n10041)
         );
  XNOR2_X1 U11079 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput8), .ZN(n10040) );
  NAND4_X1 U11080 ( .A1(n10043), .A2(n10042), .A3(n10041), .A4(n10040), .ZN(
        n10044) );
  NOR3_X1 U11081 ( .A1(n10046), .A2(n10045), .A3(n10044), .ZN(n10063) );
  AOI22_X1 U11082 ( .A1(n10049), .A2(keyinput18), .B1(keyinput53), .B2(n10048), 
        .ZN(n10047) );
  OAI221_X1 U11083 ( .B1(n10049), .B2(keyinput18), .C1(n10048), .C2(keyinput53), .A(n10047), .ZN(n10061) );
  AOI22_X1 U11084 ( .A1(n10052), .A2(keyinput61), .B1(n10051), .B2(keyinput50), 
        .ZN(n10050) );
  OAI221_X1 U11085 ( .B1(n10052), .B2(keyinput61), .C1(n10051), .C2(keyinput50), .A(n10050), .ZN(n10060) );
  AOI22_X1 U11086 ( .A1(n10055), .A2(keyinput30), .B1(keyinput41), .B2(n10054), 
        .ZN(n10053) );
  OAI221_X1 U11087 ( .B1(n10055), .B2(keyinput30), .C1(n10054), .C2(keyinput41), .A(n10053), .ZN(n10059) );
  AOI22_X1 U11088 ( .A1(n5276), .A2(keyinput60), .B1(keyinput51), .B2(n10057), 
        .ZN(n10056) );
  OAI221_X1 U11089 ( .B1(n5276), .B2(keyinput60), .C1(n10057), .C2(keyinput51), 
        .A(n10056), .ZN(n10058) );
  NOR4_X1 U11090 ( .A1(n10061), .A2(n10060), .A3(n10059), .A4(n10058), .ZN(
        n10062) );
  NAND4_X1 U11091 ( .A1(n10065), .A2(n10064), .A3(n10063), .A4(n10062), .ZN(
        n10066) );
  NOR2_X1 U11092 ( .A1(n10067), .A2(n10066), .ZN(n10068) );
  XOR2_X1 U11093 ( .A(n10069), .B(n10068), .Z(n10070) );
  XNOR2_X1 U11094 ( .A(P1_RD_REG_SCAN_IN), .B(n10070), .ZN(U126) );
  XNOR2_X1 U11095 ( .A(n10072), .B(n10071), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11096 ( .A(n10074), .B(n10073), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11097 ( .A(n10076), .B(n10075), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11098 ( .A(n10078), .B(n10077), .ZN(ADD_1068_U48) );
  XNOR2_X1 U11099 ( .A(n10080), .B(n10079), .ZN(ADD_1068_U49) );
  XOR2_X1 U11100 ( .A(n10082), .B(n10081), .Z(ADD_1068_U54) );
  XOR2_X1 U11101 ( .A(n10084), .B(n10083), .Z(ADD_1068_U53) );
  XNOR2_X1 U11102 ( .A(n10086), .B(n10085), .ZN(ADD_1068_U52) );
  INV_X1 U4781 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8884) );
  NAND2_X1 U4812 ( .A1(n5665), .A2(n6345), .ZN(n5676) );
  NAND4_X1 U4814 ( .A1(n5556), .A2(n4714), .A3(n4807), .A4(n4806), .ZN(n5690)
         );
  NAND2_X1 U4824 ( .A1(n4994), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4993) );
  INV_X1 U5807 ( .A(n5035), .ZN(n6193) );
  NAND2_X1 U6177 ( .A1(n7606), .A2(n8024), .ZN(n7632) );
  NAND2_X1 U6208 ( .A1(n4997), .A2(n4996), .ZN(n6196) );
  CLKBUF_X1 U7225 ( .A(n9457), .Z(n9474) );
endmodule

