

module b15_C_AntiSAT_k_256_6 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
         keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
         keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
         keyinput139, keyinput140, keyinput141, keyinput142, keyinput143,
         keyinput144, keyinput145, keyinput146, keyinput147, keyinput148,
         keyinput149, keyinput150, keyinput151, keyinput152, keyinput153,
         keyinput154, keyinput155, keyinput156, keyinput157, keyinput158,
         keyinput159, keyinput160, keyinput161, keyinput162, keyinput163,
         keyinput164, keyinput165, keyinput166, keyinput167, keyinput168,
         keyinput169, keyinput170, keyinput171, keyinput172, keyinput173,
         keyinput174, keyinput175, keyinput176, keyinput177, keyinput178,
         keyinput179, keyinput180, keyinput181, keyinput182, keyinput183,
         keyinput184, keyinput185, keyinput186, keyinput187, keyinput188,
         keyinput189, keyinput190, keyinput191, keyinput192, keyinput193,
         keyinput194, keyinput195, keyinput196, keyinput197, keyinput198,
         keyinput199, keyinput200, keyinput201, keyinput202, keyinput203,
         keyinput204, keyinput205, keyinput206, keyinput207, keyinput208,
         keyinput209, keyinput210, keyinput211, keyinput212, keyinput213,
         keyinput214, keyinput215, keyinput216, keyinput217, keyinput218,
         keyinput219, keyinput220, keyinput221, keyinput222, keyinput223,
         keyinput224, keyinput225, keyinput226, keyinput227, keyinput228,
         keyinput229, keyinput230, keyinput231, keyinput232, keyinput233,
         keyinput234, keyinput235, keyinput236, keyinput237, keyinput238,
         keyinput239, keyinput240, keyinput241, keyinput242, keyinput243,
         keyinput244, keyinput245, keyinput246, keyinput247, keyinput248,
         keyinput249, keyinput250, keyinput251, keyinput252, keyinput253,
         keyinput254, keyinput255;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189;

  OAI22_X1 U3631 ( .A1(n5707), .A2(n7149), .B1(n6498), .B2(n5238), .ZN(n5708)
         );
  OR2_X1 U3632 ( .A1(n4299), .A2(n5413), .ZN(n5623) );
  OAI221_X1 U3633 ( .B1(n4904), .B2(keyinput25), .C1(n7149), .C2(keyinput31), 
        .A(n7148), .ZN(n7161) );
  OAI221_X1 U3634 ( .B1(n6943), .B2(keyinput182), .C1(n7098), .C2(keyinput140), 
        .A(n6942), .ZN(n6955) );
  NAND2_X1 U3635 ( .A1(n4119), .A2(n4118), .ZN(n5560) );
  NAND2_X1 U3636 ( .A1(n4052), .A2(n4051), .ZN(n5406) );
  NAND2_X1 U3637 ( .A1(n4808), .A2(n3245), .ZN(n5146) );
  INV_X1 U3638 ( .A(n4406), .ZN(n5395) );
  OR2_X1 U3639 ( .A1(n3598), .A2(n3597), .ZN(n3330) );
  CLKBUF_X2 U3640 ( .A(n3546), .Z(n3222) );
  CLKBUF_X2 U3641 ( .A(n3528), .Z(n4251) );
  CLKBUF_X2 U3642 ( .A(n3428), .Z(n4281) );
  CLKBUF_X2 U3643 ( .A(n3641), .Z(n3216) );
  AND2_X1 U3644 ( .A1(n5495), .A2(n4589), .ZN(n3511) );
  AND2_X1 U3645 ( .A1(n3339), .A2(n4581), .ZN(n3545) );
  AND2_X1 U3646 ( .A1(n5495), .A2(n4581), .ZN(n3428) );
  CLKBUF_X2 U3647 ( .A(n3527), .Z(n3183) );
  AND2_X2 U3648 ( .A1(n4593), .A2(n3339), .ZN(n3546) );
  INV_X2 U3649 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4621) );
  AOI22_X1 U3650 ( .A1(n6994), .A2(keyinput133), .B1(keyinput159), .B2(n7149), 
        .ZN(n6993) );
  AOI22_X1 U3651 ( .A1(n7089), .A2(keyinput238), .B1(n6969), .B2(keyinput212), 
        .ZN(n6968) );
  AOI22_X1 U3652 ( .A1(n6943), .A2(keyinput182), .B1(n7098), .B2(keyinput140), 
        .ZN(n6942) );
  AND2_X1 U3653 ( .A1(n4588), .A2(n4581), .ZN(n3231) );
  AOI22_X1 U3654 ( .A1(n4904), .A2(keyinput25), .B1(keyinput31), .B2(n7149), 
        .ZN(n7148) );
  OAI221_X1 U3655 ( .B1(n6994), .B2(keyinput133), .C1(n7149), .C2(keyinput159), 
        .A(n6993), .ZN(n7004) );
  OAI221_X1 U3656 ( .B1(n7089), .B2(keyinput238), .C1(n6969), .C2(keyinput212), 
        .A(n6968), .ZN(n6978) );
  INV_X2 U3657 ( .A(n4322), .ZN(n4391) );
  AND4_X1 U3660 ( .A1(n3359), .A2(n3358), .A3(n3357), .A4(n3356), .ZN(n3375)
         );
  OR2_X1 U3661 ( .A1(n3967), .A2(n3968), .ZN(n3969) );
  OAI21_X1 U3662 ( .B1(n3904), .B2(n3269), .A(n3711), .ZN(n3712) );
  INV_X1 U3663 ( .A(n3728), .ZN(n5663) );
  INV_X4 U3664 ( .A(n5663), .ZN(n3184) );
  NOR2_X1 U3665 ( .A1(n5300), .A2(n5301), .ZN(n5299) );
  INV_X1 U3666 ( .A(n4469), .ZN(n4742) );
  INV_X1 U3667 ( .A(n6278), .ZN(n6254) );
  AND2_X1 U3668 ( .A1(n6296), .A2(n4417), .ZN(n6302) );
  AND2_X1 U3669 ( .A1(n5553), .A2(n3297), .ZN(n5413) );
  NAND2_X2 U3670 ( .A1(n3444), .A2(n3202), .ZN(n4318) );
  INV_X1 U3672 ( .A(n6302), .ZN(n6319) );
  AOI211_X1 U3673 ( .C1(n5490), .C2(n5489), .A(n5488), .B(n5624), .ZN(n5491)
         );
  INV_X1 U3674 ( .A(n3511), .ZN(n3186) );
  AND4_X1 U3675 ( .A1(n3421), .A2(n3420), .A3(n3419), .A4(n3418), .ZN(n3181)
         );
  NAND2_X2 U3676 ( .A1(n5184), .A2(n5183), .ZN(n5182) );
  NAND2_X2 U3677 ( .A1(n3970), .A2(n3969), .ZN(n5184) );
  NOR2_X2 U3678 ( .A1(n5334), .A2(n5335), .ZN(n5333) );
  NAND2_X2 U3679 ( .A1(n3261), .A2(n3593), .ZN(n3657) );
  AND2_X4 U3680 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4588) );
  CLKBUF_X3 U3681 ( .A(n3527), .Z(n3182) );
  AND2_X1 U3682 ( .A1(n4589), .A2(n4588), .ZN(n3527) );
  NAND2_X1 U3683 ( .A1(n5431), .A2(n3187), .ZN(n5654) );
  NAND2_X1 U3684 ( .A1(n5591), .A2(n5594), .ZN(n5592) );
  NOR2_X2 U3685 ( .A1(n5146), .A2(n5147), .ZN(n5169) );
  AOI21_X1 U3686 ( .B1(n3802), .B2(n3801), .A(n3800), .ZN(n4648) );
  BUF_X1 U3687 ( .A(n3910), .Z(n3230) );
  AND4_X1 U3688 ( .A1(n3432), .A2(n3431), .A3(n3430), .A4(n3429), .ZN(n3445)
         );
  BUF_X2 U3690 ( .A(n4279), .Z(n3220) );
  BUF_X2 U3691 ( .A(n3545), .Z(n4274) );
  INV_X1 U3692 ( .A(n3186), .ZN(n3185) );
  CLKBUF_X2 U3693 ( .A(n3526), .Z(n4595) );
  INV_X2 U3694 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3332) );
  NOR2_X2 U3695 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4644) );
  INV_X1 U3696 ( .A(n5433), .ZN(n5665) );
  NOR2_X1 U3697 ( .A1(n3246), .A2(n5485), .ZN(n5486) );
  NAND2_X1 U3698 ( .A1(n5654), .A2(n5432), .ZN(n5433) );
  NOR2_X1 U3699 ( .A1(n4441), .A2(n3739), .ZN(n3741) );
  AND2_X1 U3700 ( .A1(n5640), .A2(n3237), .ZN(n4441) );
  AND2_X1 U3701 ( .A1(n3243), .A2(n5537), .ZN(n6016) );
  AND2_X1 U3702 ( .A1(n3193), .A2(n3194), .ZN(n5431) );
  XNOR2_X1 U3703 ( .A(n5418), .B(n5417), .ZN(n5595) );
  AND2_X1 U3704 ( .A1(n5544), .A2(n5543), .ZN(n6027) );
  NAND2_X1 U3705 ( .A1(n5764), .A2(n5766), .ZN(n5765) );
  CLKBUF_X1 U3706 ( .A(n5683), .Z(n5684) );
  NAND2_X1 U3707 ( .A1(n3302), .A2(n4150), .ZN(n5561) );
  NAND2_X1 U3708 ( .A1(n5683), .A2(n3250), .ZN(n5655) );
  AOI21_X1 U3709 ( .B1(n3266), .B2(n3268), .A(n3248), .ZN(n3263) );
  NAND2_X1 U3710 ( .A1(n3702), .A2(n3701), .ZN(n5109) );
  OR2_X1 U3711 ( .A1(n4464), .A2(n4411), .ZN(n5534) );
  OAI21_X1 U3712 ( .B1(n3242), .B2(n3268), .A(n5307), .ZN(n3267) );
  OAI21_X1 U3713 ( .B1(n5465), .B2(n5466), .A(n5464), .ZN(n5532) );
  NAND2_X1 U3714 ( .A1(n3950), .A2(n5008), .ZN(n3967) );
  AND2_X1 U3715 ( .A1(n5385), .A2(n3730), .ZN(n3200) );
  AND2_X1 U3716 ( .A1(n5110), .A2(n5082), .ZN(n3192) );
  OAI21_X1 U3717 ( .B1(n3904), .B2(n3987), .A(n3903), .ZN(n5108) );
  NAND2_X1 U3718 ( .A1(n3715), .A2(n3717), .ZN(n3728) );
  NAND2_X1 U3719 ( .A1(n3289), .A2(n4578), .ZN(n4665) );
  NAND2_X1 U3720 ( .A1(n4816), .A2(n3593), .ZN(n4757) );
  CLKBUF_X1 U3721 ( .A(n4650), .Z(n5863) );
  AND2_X1 U3722 ( .A1(n3572), .A2(n3571), .ZN(n3598) );
  XNOR2_X1 U3723 ( .A(n3618), .B(n3617), .ZN(n4650) );
  NAND2_X1 U3724 ( .A1(n3610), .A2(n3609), .ZN(n5862) );
  NOR2_X1 U3725 ( .A1(n4743), .A2(n3474), .ZN(n6605) );
  NOR2_X1 U3726 ( .A1(n4743), .A2(n5594), .ZN(n6620) );
  NOR2_X1 U3727 ( .A1(n4743), .A2(n4722), .ZN(n6593) );
  NOR2_X1 U3728 ( .A1(n4743), .A2(n4716), .ZN(n6562) );
  AND2_X2 U3729 ( .A1(n6438), .A2(n3816), .ZN(n6442) );
  NAND2_X2 U3730 ( .A1(n4556), .A2(n4515), .ZN(n6438) );
  NAND2_X1 U3731 ( .A1(n4556), .A2(n6655), .ZN(n6794) );
  NAND2_X1 U3732 ( .A1(n5169), .A2(n5170), .ZN(n5300) );
  NAND2_X1 U3733 ( .A1(n3525), .A2(n3524), .ZN(n3615) );
  CLKBUF_X1 U3734 ( .A(n4652), .Z(n5317) );
  AND2_X1 U3735 ( .A1(n3544), .A2(n3543), .ZN(n3510) );
  NOR2_X1 U3736 ( .A1(n4680), .A2(n3282), .ZN(n3281) );
  NAND2_X1 U3737 ( .A1(n3325), .A2(n3457), .ZN(n4475) );
  NAND3_X1 U3738 ( .A1(n3806), .A2(n3451), .A3(n3328), .ZN(n3452) );
  OR2_X1 U3739 ( .A1(n4446), .A2(n4722), .ZN(n3465) );
  AND2_X1 U3740 ( .A1(n4378), .A2(n4323), .ZN(n4325) );
  INV_X1 U3741 ( .A(n4562), .ZN(n4387) );
  NAND2_X1 U3742 ( .A1(n3377), .A2(n3376), .ZN(n3323) );
  AND2_X1 U3743 ( .A1(n4572), .A2(n4509), .ZN(n4553) );
  NAND2_X1 U3744 ( .A1(n4391), .A2(n4349), .ZN(n4378) );
  AND2_X1 U3745 ( .A1(n3387), .A2(n4576), .ZN(n3458) );
  AND2_X1 U3746 ( .A1(n3290), .A2(n3474), .ZN(n4572) );
  OR2_X2 U3747 ( .A1(n4319), .A2(n4716), .ZN(n4322) );
  OR2_X2 U3748 ( .A1(n3397), .A2(n3396), .ZN(n4319) );
  INV_X1 U3749 ( .A(n3409), .ZN(n3376) );
  OR2_X1 U3750 ( .A1(n3557), .A2(n3556), .ZN(n3621) );
  AND4_X2 U3751 ( .A1(n3446), .A2(n3445), .A3(n3444), .A4(n3443), .ZN(n4716)
         );
  NAND2_X2 U3752 ( .A1(n3406), .A2(n3326), .ZN(n4469) );
  NAND2_X2 U3753 ( .A1(n3386), .A2(n3241), .ZN(n4576) );
  AND4_X1 U3754 ( .A1(n3371), .A2(n3370), .A3(n3369), .A4(n3368), .ZN(n3372)
         );
  AND4_X1 U3755 ( .A1(n3337), .A2(n3336), .A3(n3335), .A4(n3334), .ZN(n3345)
         );
  AND4_X1 U3756 ( .A1(n3405), .A2(n3404), .A3(n3403), .A4(n3402), .ZN(n3326)
         );
  AND4_X1 U3757 ( .A1(n3401), .A2(n3400), .A3(n3399), .A4(n3398), .ZN(n3406)
         );
  AND4_X1 U3758 ( .A1(n3381), .A2(n3380), .A3(n3379), .A4(n3378), .ZN(n3386)
         );
  AND4_X1 U3759 ( .A1(n3349), .A2(n3348), .A3(n3347), .A4(n3346), .ZN(n3355)
         );
  AND4_X1 U3760 ( .A1(n3426), .A2(n3425), .A3(n3424), .A4(n3423), .ZN(n3446)
         );
  AND4_X1 U3761 ( .A1(n3343), .A2(n3342), .A3(n3341), .A4(n3340), .ZN(n3344)
         );
  AND4_X1 U3762 ( .A1(n3442), .A2(n3441), .A3(n3440), .A4(n3439), .ZN(n3443)
         );
  AND4_X1 U3763 ( .A1(n3363), .A2(n3362), .A3(n3361), .A4(n3360), .ZN(n3374)
         );
  AND4_X1 U3764 ( .A1(n3367), .A2(n3366), .A3(n3365), .A4(n3364), .ZN(n3373)
         );
  AND4_X1 U3765 ( .A1(n3353), .A2(n3352), .A3(n3351), .A4(n3350), .ZN(n3354)
         );
  BUF_X4 U3766 ( .A(n3434), .Z(n3215) );
  BUF_X2 U3767 ( .A(n3492), .Z(n3225) );
  AND2_X2 U3768 ( .A1(n3338), .A2(n4588), .ZN(n3526) );
  AND2_X2 U3769 ( .A1(n3339), .A2(n4589), .ZN(n3433) );
  AND2_X2 U3770 ( .A1(n3338), .A2(n3223), .ZN(n3234) );
  AND2_X2 U3771 ( .A1(n4644), .A2(n4589), .ZN(n3434) );
  AND2_X2 U3772 ( .A1(n5495), .A2(n4593), .ZN(n3492) );
  CLKBUF_X2 U3773 ( .A(n4644), .Z(n3224) );
  AND2_X2 U3774 ( .A1(n3332), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4593)
         );
  AND2_X2 U3775 ( .A1(n4588), .A2(n4581), .ZN(n3232) );
  CLKBUF_X2 U3776 ( .A(n4644), .Z(n3223) );
  AND2_X2 U3777 ( .A1(n4621), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3338)
         );
  AND2_X1 U3778 ( .A1(n5499), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5495)
         );
  AND2_X2 U3779 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4581) );
  NOR2_X2 U3780 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6564) );
  AND2_X1 U3781 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4592) );
  NOR2_X1 U3782 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3333) );
  INV_X2 U3783 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6780) );
  AOI21_X1 U3784 ( .B1(n6036), .B2(n6035), .A(n6034), .ZN(n6037) );
  NAND2_X2 U3785 ( .A1(n3330), .A2(n3599), .ZN(n4656) );
  OAI22_X2 U3786 ( .A1(n4622), .A2(STATE2_REG_0__SCAN_IN), .B1(n3601), .B2(
        n3579), .ZN(n3507) );
  NOR2_X2 U3787 ( .A1(n5560), .A2(n3300), .ZN(n5514) );
  OR2_X2 U3788 ( .A1(n5182), .A2(n3305), .ZN(n5374) );
  XNOR2_X1 U3789 ( .A(n3967), .B(n3968), .ZN(n5177) );
  INV_X1 U3790 ( .A(n3269), .ZN(n3786) );
  AND2_X2 U3791 ( .A1(n4801), .A2(n5009), .ZN(n5008) );
  AND2_X1 U3792 ( .A1(n5430), .A2(n3188), .ZN(n3187) );
  INV_X1 U3793 ( .A(n5672), .ZN(n3188) );
  NAND2_X1 U3794 ( .A1(n5109), .A2(n3192), .ZN(n3189) );
  AND2_X1 U3795 ( .A1(n3189), .A2(n3190), .ZN(n3724) );
  OR2_X1 U3796 ( .A1(n3191), .A2(n3713), .ZN(n3190) );
  INV_X1 U3797 ( .A(n5082), .ZN(n3191) );
  NAND2_X1 U3798 ( .A1(n5764), .A2(n3196), .ZN(n3193) );
  OR2_X1 U3799 ( .A1(n3195), .A2(n5427), .ZN(n3194) );
  INV_X1 U3800 ( .A(n5429), .ZN(n3195) );
  AND2_X1 U3801 ( .A1(n5766), .A2(n5429), .ZN(n3196) );
  NAND2_X1 U3802 ( .A1(n5383), .A2(n3200), .ZN(n3197) );
  AND2_X1 U3803 ( .A1(n3197), .A2(n3198), .ZN(n3732) );
  OR2_X1 U3804 ( .A1(n3199), .A2(n3729), .ZN(n3198) );
  INV_X1 U3805 ( .A(n3730), .ZN(n3199) );
  NAND2_X1 U3806 ( .A1(n3657), .A2(n3594), .ZN(n3201) );
  AND3_X2 U3807 ( .A1(n3443), .A2(n3446), .A3(n3445), .ZN(n3202) );
  OAI21_X1 U3808 ( .B1(n3483), .B2(n3331), .A(n3453), .ZN(n3203) );
  OAI21_X1 U3809 ( .B1(n3483), .B2(n3331), .A(n3453), .ZN(n3204) );
  AND2_X1 U3810 ( .A1(n3452), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3205) );
  INV_X1 U3812 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3207) );
  NAND2_X1 U3813 ( .A1(n3657), .A2(n3594), .ZN(n3920) );
  AND4_X1 U3814 ( .A1(n3438), .A2(n3437), .A3(n3436), .A4(n3435), .ZN(n3444)
         );
  OAI21_X1 U3815 ( .B1(n3483), .B2(n3331), .A(n3453), .ZN(n3544) );
  NAND2_X2 U3816 ( .A1(n3452), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3483) );
  AND2_X1 U3817 ( .A1(n3224), .A2(n4581), .ZN(n3208) );
  AND2_X2 U3818 ( .A1(n3224), .A2(n4581), .ZN(n3528) );
  NAND2_X1 U3819 ( .A1(n3482), .A2(n3240), .ZN(n3491) );
  NAND2_X1 U3820 ( .A1(n4301), .A2(n3475), .ZN(n4636) );
  AND2_X1 U3821 ( .A1(n4593), .A2(n4588), .ZN(n3209) );
  AND2_X1 U3822 ( .A1(n4593), .A2(n4588), .ZN(n3210) );
  AND2_X1 U3823 ( .A1(n4593), .A2(n4588), .ZN(n4279) );
  AND2_X1 U3824 ( .A1(n4593), .A2(n3223), .ZN(n3211) );
  AND2_X1 U3825 ( .A1(n4593), .A2(n3223), .ZN(n3422) );
  AND4_X2 U3826 ( .A1(n3413), .A2(n3412), .A3(n3411), .A4(n3410), .ZN(n4301)
         );
  AND2_X1 U3827 ( .A1(n3503), .A2(n3409), .ZN(n3795) );
  INV_X2 U3828 ( .A(n4483), .ZN(n4727) );
  AND2_X2 U3829 ( .A1(n3339), .A2(n4589), .ZN(n3212) );
  AND2_X2 U3830 ( .A1(n3339), .A2(n4589), .ZN(n3213) );
  AND2_X1 U3831 ( .A1(n4589), .A2(n4588), .ZN(n3217) );
  AND2_X2 U3832 ( .A1(n4589), .A2(n4588), .ZN(n3218) );
  AND2_X2 U3833 ( .A1(n4593), .A2(n3223), .ZN(n3219) );
  INV_X1 U3835 ( .A(n3186), .ZN(n3229) );
  INV_X2 U3836 ( .A(n3460), .ZN(n3461) );
  NAND2_X2 U3837 ( .A1(n3345), .A2(n3344), .ZN(n3460) );
  BUF_X8 U3838 ( .A(n3492), .Z(n3226) );
  AND2_X1 U3839 ( .A1(n3633), .A2(n6426), .ZN(n5063) );
  NAND2_X2 U3840 ( .A1(n5655), .A2(n3735), .ZN(n5764) );
  NAND4_X4 U3841 ( .A1(n3375), .A2(n3374), .A3(n3373), .A4(n3372), .ZN(n3409)
         );
  AND3_X2 U3842 ( .A1(n3450), .A2(n4583), .A3(n3449), .ZN(n3328) );
  AND2_X2 U3843 ( .A1(n3786), .A2(n4688), .ZN(n3454) );
  BUF_X2 U3844 ( .A(n3376), .Z(n4688) );
  NAND2_X2 U3845 ( .A1(n3461), .A2(n3448), .ZN(n3467) );
  NAND2_X4 U3846 ( .A1(n3355), .A2(n3354), .ZN(n3448) );
  AND4_X2 U3847 ( .A1(n3417), .A2(n3416), .A3(n3415), .A4(n3414), .ZN(n3239)
         );
  NAND2_X2 U3848 ( .A1(n3491), .A2(n3490), .ZN(n3573) );
  AND2_X2 U3849 ( .A1(n3338), .A2(n3224), .ZN(n3233) );
  NOR2_X1 U3851 ( .A1(n3672), .A2(n3310), .ZN(n3309) );
  INV_X1 U3852 ( .A(n3658), .ZN(n3310) );
  OR2_X1 U3853 ( .A1(n3538), .A2(n3537), .ZN(n3718) );
  OR2_X1 U3854 ( .A1(n3502), .A2(n3501), .ZN(n3504) );
  INV_X1 U3855 ( .A(n3504), .ZN(n3601) );
  NAND2_X1 U3856 ( .A1(n4716), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3580) );
  OR2_X1 U3857 ( .A1(n3409), .A2(n6783), .ZN(n3579) );
  NAND2_X1 U3858 ( .A1(n3792), .A2(n3793), .ZN(n4308) );
  OR2_X1 U3859 ( .A1(n3794), .A2(n3791), .ZN(n3792) );
  AND2_X1 U3860 ( .A1(n6512), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3791)
         );
  INV_X1 U3861 ( .A(n5563), .ZN(n4150) );
  INV_X1 U3862 ( .A(n5571), .ZN(n4119) );
  NAND2_X1 U3863 ( .A1(n5585), .A2(n3295), .ZN(n3294) );
  INV_X1 U3864 ( .A(n5405), .ZN(n3295) );
  INV_X1 U3865 ( .A(n4290), .ZN(n4263) );
  NOR2_X1 U3866 ( .A1(n6630), .A2(n6783), .ZN(n4290) );
  OR2_X1 U3867 ( .A1(n5365), .A2(n5329), .ZN(n3307) );
  INV_X1 U3868 ( .A(n5177), .ZN(n3966) );
  NAND2_X1 U3869 ( .A1(n3461), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3987) );
  INV_X1 U3870 ( .A(n3298), .ZN(n3296) );
  NAND2_X1 U3871 ( .A1(n4456), .A2(n4455), .ZN(n4486) );
  AND2_X1 U3872 ( .A1(n5505), .A2(n5501), .ZN(n6777) );
  NAND2_X1 U3873 ( .A1(n3447), .A2(n4510), .ZN(n4445) );
  NAND2_X1 U3874 ( .A1(n3696), .A2(n3695), .ZN(n3704) );
  NAND2_X1 U3875 ( .A1(n3649), .A2(n3648), .ZN(n3658) );
  NAND2_X1 U3876 ( .A1(n3184), .A2(n3258), .ZN(n3320) );
  OAI211_X1 U3877 ( .C1(n3541), .C2(n3580), .A(n3540), .B(n3539), .ZN(n3614)
         );
  NAND2_X1 U3878 ( .A1(n3567), .A2(n3606), .ZN(n3616) );
  NOR2_X1 U3879 ( .A1(n4586), .A2(n4478), .ZN(n4481) );
  NOR2_X1 U3880 ( .A1(n4319), .A2(n4469), .ZN(n3290) );
  NOR2_X1 U3881 ( .A1(n4298), .A2(n3298), .ZN(n3297) );
  NAND2_X1 U3882 ( .A1(n3299), .A2(n5542), .ZN(n3298) );
  INV_X1 U3883 ( .A(n5536), .ZN(n3299) );
  XNOR2_X1 U3884 ( .A(n3657), .B(n3658), .ZN(n3933) );
  INV_X1 U3885 ( .A(n3320), .ZN(n3314) );
  NOR2_X1 U3886 ( .A1(n6103), .A2(n3317), .ZN(n3316) );
  INV_X1 U3887 ( .A(n3319), .ZN(n3317) );
  NOR2_X1 U3888 ( .A1(n5379), .A2(n3285), .ZN(n3284) );
  INV_X1 U3889 ( .A(n5373), .ZN(n3285) );
  INV_X1 U3890 ( .A(n4682), .ZN(n3282) );
  NAND2_X1 U3891 ( .A1(n4475), .A2(n3471), .ZN(n3543) );
  AND2_X1 U3892 ( .A1(n3470), .A2(n3469), .ZN(n3471) );
  AOI21_X1 U3893 ( .B1(n6782), .B2(n3465), .A(n3464), .ZN(n3470) );
  NOR2_X1 U3894 ( .A1(n4318), .A2(n3742), .ZN(n4302) );
  AND2_X1 U3895 ( .A1(n4301), .A2(n4302), .ZN(n4513) );
  AND2_X1 U3896 ( .A1(n3905), .A2(n5108), .ZN(n3950) );
  AND2_X1 U3897 ( .A1(n4457), .A2(n4509), .ZN(n4604) );
  INV_X1 U3898 ( .A(n4014), .ZN(n5414) );
  AND2_X1 U3899 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n3814), .ZN(n4225)
         );
  INV_X1 U3900 ( .A(n4205), .ZN(n3814) );
  AND2_X1 U3901 ( .A1(n6030), .A2(n4311), .ZN(n4206) );
  OR2_X1 U3902 ( .A1(n3303), .A2(n3301), .ZN(n3300) );
  INV_X1 U3903 ( .A(n5515), .ZN(n3301) );
  OR2_X1 U3904 ( .A1(n6050), .A2(n4269), .ZN(n4148) );
  AND2_X1 U3905 ( .A1(n5578), .A2(n3293), .ZN(n3292) );
  INV_X1 U3906 ( .A(n3294), .ZN(n3293) );
  NAND2_X1 U3907 ( .A1(n4032), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4048)
         );
  NAND2_X1 U3908 ( .A1(n3306), .A2(n5375), .ZN(n3305) );
  INV_X1 U3909 ( .A(n3307), .ZN(n3306) );
  NOR2_X1 U3910 ( .A1(n7149), .A2(n3981), .ZN(n3999) );
  NAND2_X1 U3911 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n3999), .ZN(n4013)
         );
  OR2_X1 U3912 ( .A1(n5182), .A2(n5329), .ZN(n5366) );
  AND2_X1 U3913 ( .A1(n4457), .A2(n3807), .ZN(n4515) );
  NAND2_X1 U3914 ( .A1(n3184), .A2(n5428), .ZN(n5429) );
  NAND2_X1 U3915 ( .A1(n3264), .A2(n3263), .ZN(n3727) );
  NAND2_X1 U3916 ( .A1(n3489), .A2(n3488), .ZN(n3490) );
  INV_X1 U3917 ( .A(n3487), .ZN(n3488) );
  NAND2_X1 U3918 ( .A1(n3205), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3489) );
  AOI21_X1 U3919 ( .B1(n4582), .B2(n6783), .A(n3592), .ZN(n4686) );
  INV_X1 U3920 ( .A(n3591), .ZN(n3592) );
  AND2_X1 U3921 ( .A1(n3799), .A2(n3798), .ZN(n3800) );
  OR2_X1 U3922 ( .A1(n3790), .A2(n3789), .ZN(n3802) );
  AND2_X1 U3923 ( .A1(n6749), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3803) );
  AND2_X1 U3924 ( .A1(n5456), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4417) );
  AND2_X1 U3925 ( .A1(n5593), .A2(n5370), .ZN(n6333) );
  INV_X1 U3926 ( .A(n5593), .ZN(n6332) );
  AND2_X1 U3927 ( .A1(n5593), .A2(n4559), .ZN(n5331) );
  AND2_X1 U3928 ( .A1(n3737), .A2(n3738), .ZN(n3739) );
  NOR2_X1 U3929 ( .A1(n4483), .A2(n4413), .ZN(n3476) );
  OR2_X1 U3930 ( .A1(n3694), .A2(n3693), .ZN(n3708) );
  OR2_X1 U3931 ( .A1(n3647), .A2(n3646), .ZN(n3675) );
  NOR2_X1 U3932 ( .A1(n3622), .A2(n3460), .ZN(n3472) );
  NAND2_X1 U3933 ( .A1(n3795), .A2(n3221), .ZN(n3796) );
  NAND2_X1 U3934 ( .A1(n3560), .A2(n3559), .ZN(n3604) );
  NAND2_X1 U3935 ( .A1(n3558), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3559) );
  AOI22_X1 U3936 ( .A1(n3428), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3516), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3398) );
  AOI22_X1 U3937 ( .A1(n3511), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3343) );
  OR2_X1 U3938 ( .A1(n3794), .A2(n3793), .ZN(n4303) );
  AOI22_X1 U3939 ( .A1(n3526), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3641), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3350) );
  NAND2_X1 U3940 ( .A1(n3304), .A2(n4150), .ZN(n3303) );
  INV_X1 U3941 ( .A(n5448), .ZN(n3304) );
  NOR2_X1 U3942 ( .A1(n3945), .A2(n3808), .ZN(n3900) );
  XNOR2_X1 U3943 ( .A(n3715), .B(n3706), .ZN(n3904) );
  OAI21_X1 U3944 ( .B1(n4656), .B2(n3269), .A(n3603), .ZN(n3630) );
  NOR3_X1 U3945 ( .A1(n3238), .A2(n3275), .A3(n3278), .ZN(n3277) );
  NAND2_X1 U3946 ( .A1(n4381), .A2(n5438), .ZN(n3275) );
  NAND2_X1 U3947 ( .A1(n5663), .A2(n3736), .ZN(n3319) );
  NAND2_X1 U3948 ( .A1(n5764), .A2(n3320), .ZN(n3318) );
  INV_X1 U3949 ( .A(n5564), .ZN(n3278) );
  INV_X1 U3950 ( .A(n5308), .ZN(n3311) );
  INV_X1 U3951 ( .A(n3267), .ZN(n3266) );
  INV_X1 U3952 ( .A(n5165), .ZN(n3268) );
  NOR2_X1 U3953 ( .A1(n5123), .A2(n3280), .ZN(n3279) );
  INV_X1 U3954 ( .A(n4809), .ZN(n3280) );
  AND4_X1 U3955 ( .A1(n4473), .A2(n4472), .A3(n4471), .A4(n4470), .ZN(n4474)
         );
  NAND2_X1 U3956 ( .A1(n3454), .A2(n4319), .ZN(n4583) );
  AND4_X1 U3957 ( .A1(n3461), .A2(n4716), .A3(n3409), .A4(n4576), .ZN(n3462)
         );
  AOI21_X1 U3958 ( .B1(n3778), .B2(n3777), .A(n3776), .ZN(n3790) );
  AND2_X1 U3959 ( .A1(n3775), .A2(n3774), .ZN(n3776) );
  OAI21_X1 U3960 ( .B1(n6787), .B2(n6669), .A(n5808), .ZN(n4687) );
  AND2_X1 U3961 ( .A1(n4582), .A2(n5853), .ZN(n4983) );
  XNOR2_X1 U3962 ( .A(n3615), .B(n3614), .ZN(n3618) );
  INV_X1 U3963 ( .A(n3616), .ZN(n3617) );
  INV_X1 U3964 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6643) );
  AND2_X1 U3965 ( .A1(n4632), .A2(n4631), .ZN(n6642) );
  AND2_X1 U3966 ( .A1(n4513), .A2(n4309), .ZN(n4508) );
  NOR2_X1 U3967 ( .A1(n4403), .A2(n4409), .ZN(n5461) );
  OR2_X1 U3968 ( .A1(n6109), .A2(n4269), .ZN(n4187) );
  AOI21_X1 U3969 ( .B1(n3936), .B2(n3996), .A(n3941), .ZN(n4799) );
  OR2_X1 U3970 ( .A1(n5626), .A2(n4269), .ZN(n4270) );
  AND2_X1 U3971 ( .A1(n4227), .A2(n4226), .ZN(n5542) );
  NAND2_X1 U3972 ( .A1(n5553), .A2(n5542), .ZN(n5543) );
  NAND2_X1 U3973 ( .A1(n4144), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4164)
         );
  INV_X1 U3974 ( .A(n5560), .ZN(n3302) );
  BUF_X1 U3975 ( .A(n5560), .Z(n5574) );
  AND2_X1 U3976 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n3812), .ZN(n4099)
         );
  INV_X1 U3977 ( .A(n4082), .ZN(n3812) );
  AND2_X1 U3978 ( .A1(n4084), .A2(n4083), .ZN(n5585) );
  NOR2_X1 U3979 ( .A1(n4048), .A2(n3811), .ZN(n4053) );
  NAND2_X1 U3980 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n4053), .ZN(n4082)
         );
  INV_X1 U3981 ( .A(n5391), .ZN(n4051) );
  INV_X1 U3982 ( .A(n5374), .ZN(n4052) );
  AND2_X1 U3983 ( .A1(n4034), .A2(n4033), .ZN(n5375) );
  NOR2_X1 U3984 ( .A1(n6943), .A2(n4013), .ZN(n4032) );
  AND2_X1 U3985 ( .A1(n4017), .A2(n4016), .ZN(n5365) );
  NOR2_X1 U3986 ( .A1(n5182), .A2(n3307), .ZN(n5376) );
  AND3_X1 U3987 ( .A1(n4002), .A2(n4001), .A3(n4000), .ZN(n5329) );
  INV_X1 U3988 ( .A(n5176), .ZN(n3965) );
  NAND2_X1 U3989 ( .A1(n3824), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3951)
         );
  INV_X1 U3990 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3952) );
  NOR2_X1 U3991 ( .A1(n3848), .A2(n3810), .ZN(n3824) );
  NAND2_X1 U3992 ( .A1(n3868), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3848)
         );
  AND2_X1 U3993 ( .A1(n5298), .A2(n5297), .ZN(n5295) );
  AND3_X1 U3994 ( .A1(n3865), .A2(n3864), .A3(n3863), .ZN(n5288) );
  OR2_X1 U3995 ( .A1(n5143), .A2(n5142), .ZN(n5287) );
  NAND2_X1 U3996 ( .A1(n3900), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3899)
         );
  NAND2_X1 U3997 ( .A1(n5116), .A2(n5115), .ZN(n5143) );
  AND2_X1 U3998 ( .A1(n5008), .A2(n5108), .ZN(n5116) );
  INV_X1 U3999 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6300) );
  NOR2_X1 U4000 ( .A1(n3929), .A2(n6300), .ZN(n3937) );
  NAND2_X1 U4001 ( .A1(n3935), .A2(n3934), .ZN(n4800) );
  INV_X1 U4002 ( .A(n4778), .ZN(n3935) );
  NAND2_X1 U4003 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3916) );
  NAND2_X1 U4004 ( .A1(n4579), .A2(n4580), .ZN(n4578) );
  NAND2_X1 U4005 ( .A1(n5547), .A2(n5538), .ZN(n4403) );
  AND2_X1 U4006 ( .A1(n5551), .A2(n5545), .ZN(n5547) );
  NOR2_X1 U4007 ( .A1(n5550), .A2(n5549), .ZN(n5551) );
  NAND2_X1 U4008 ( .A1(n3184), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5646) );
  AOI21_X1 U4009 ( .B1(n3316), .B2(n3314), .A(n3255), .ZN(n3313) );
  INV_X1 U4010 ( .A(n3316), .ZN(n3315) );
  NAND2_X1 U4011 ( .A1(n3277), .A2(n3276), .ZN(n5550) );
  INV_X1 U4012 ( .A(n5518), .ZN(n3276) );
  INV_X1 U4013 ( .A(n3277), .ZN(n5519) );
  NOR3_X1 U4014 ( .A1(n3238), .A2(n3278), .A3(n5568), .ZN(n5566) );
  NOR2_X1 U4015 ( .A1(n3238), .A2(n5568), .ZN(n5569) );
  NAND2_X1 U4016 ( .A1(n5663), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5427) );
  AND2_X1 U4017 ( .A1(n3284), .A2(n4368), .ZN(n3283) );
  OR2_X1 U4018 ( .A1(n6161), .A2(n4501), .ZN(n5441) );
  NAND2_X1 U4019 ( .A1(n5333), .A2(n3284), .ZN(n5401) );
  NAND2_X1 U4020 ( .A1(n5333), .A2(n5373), .ZN(n5378) );
  AND2_X1 U4021 ( .A1(n5683), .A2(n3734), .ZN(n3321) );
  NAND2_X1 U4022 ( .A1(n5242), .A2(n5243), .ZN(n5334) );
  NAND2_X1 U4023 ( .A1(n3262), .A2(n3266), .ZN(n3312) );
  OR2_X1 U4024 ( .A1(n3322), .A2(n3268), .ZN(n3262) );
  XNOR2_X1 U4025 ( .A(n3722), .B(n5095), .ZN(n5082) );
  AND2_X1 U4026 ( .A1(n4808), .A2(n3279), .ZN(n5121) );
  XNOR2_X1 U4027 ( .A(n3712), .B(n6470), .ZN(n5110) );
  NAND2_X1 U4028 ( .A1(n4808), .A2(n4809), .ZN(n5122) );
  XNOR2_X1 U4029 ( .A(n3700), .B(n5086), .ZN(n4805) );
  INV_X1 U4030 ( .A(n6501), .ZN(n5781) );
  XNOR2_X1 U4031 ( .A(n3654), .B(n3653), .ZN(n4669) );
  NAND2_X1 U4032 ( .A1(n4486), .A2(n4511), .ZN(n5089) );
  AND2_X1 U4033 ( .A1(n4327), .A2(n4326), .ZN(n4563) );
  INV_X1 U4034 ( .A(n4656), .ZN(n4816) );
  INV_X1 U4035 ( .A(n3599), .ZN(n3261) );
  OR2_X1 U4036 ( .A1(n3467), .A2(n3804), .ZN(n6630) );
  INV_X1 U4037 ( .A(n6635), .ZN(n5476) );
  OAI21_X1 U4038 ( .B1(n6519), .B2(n5852), .A(n6564), .ZN(n5861) );
  INV_X1 U4039 ( .A(n4782), .ZN(n4895) );
  AND2_X1 U4040 ( .A1(n5863), .A2(n4751), .ZN(n4821) );
  INV_X1 U4041 ( .A(n6566), .ZN(n5188) );
  OR2_X1 U4042 ( .A1(n3483), .A2(n4621), .ZN(n3578) );
  INV_X1 U4043 ( .A(n4319), .ZN(n4722) );
  NAND2_X1 U4044 ( .A1(n6783), .A2(n4687), .ZN(n4782) );
  INV_X1 U4045 ( .A(n5187), .ZN(n5903) );
  INV_X1 U4046 ( .A(n4757), .ZN(n4752) );
  INV_X1 U4047 ( .A(n4821), .ZN(n5129) );
  INV_X1 U4048 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n7152) );
  INV_X1 U4049 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6691) );
  AOI21_X1 U4050 ( .B1(n5512), .B2(n5513), .A(n3273), .ZN(n3272) );
  NAND2_X1 U4051 ( .A1(n5511), .A2(n5510), .ZN(n3273) );
  OR3_X1 U4052 ( .A1(n6777), .A2(n4453), .A3(n4419), .ZN(n6262) );
  INV_X1 U4053 ( .A(n6262), .ZN(n6307) );
  INV_X1 U4054 ( .A(n4582), .ZN(n6315) );
  AND2_X1 U4055 ( .A1(n6296), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6272) );
  NAND2_X1 U4056 ( .A1(n4683), .A2(n4682), .ZN(n4679) );
  INV_X1 U4057 ( .A(n5592), .ZN(n5557) );
  INV_X1 U4058 ( .A(n5591), .ZN(n5556) );
  NAND2_X2 U4059 ( .A1(n4575), .A2(n4574), .ZN(n5591) );
  INV_X1 U4060 ( .A(n6016), .ZN(n5604) );
  AOI21_X1 U4061 ( .B1(n4556), .B2(n4604), .A(n4555), .ZN(n4557) );
  INV_X1 U4062 ( .A(n5331), .ZN(n5338) );
  AND2_X1 U4063 ( .A1(n4556), .A2(n4535), .ZN(n6349) );
  INV_X1 U4064 ( .A(n6349), .ZN(n6360) );
  NAND2_X1 U4065 ( .A1(n4556), .A2(n4607), .ZN(n6421) );
  INV_X1 U4066 ( .A(n6421), .ZN(n6422) );
  OR2_X1 U4067 ( .A1(n4315), .A2(n4314), .ZN(n4316) );
  NAND2_X1 U4068 ( .A1(n5553), .A2(n3244), .ZN(n5418) );
  INV_X1 U4069 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6943) );
  INV_X1 U4070 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n7149) );
  INV_X1 U4071 ( .A(n6437), .ZN(n5709) );
  INV_X1 U4072 ( .A(n6438), .ZN(n6431) );
  NAND2_X1 U4073 ( .A1(n3322), .A2(n3242), .ZN(n3265) );
  INV_X1 U4074 ( .A(n6503), .ZN(n5783) );
  AND2_X1 U4075 ( .A1(n4486), .A2(n4461), .ZN(n6507) );
  AND2_X1 U4076 ( .A1(n4486), .A2(n4467), .ZN(n6503) );
  INV_X1 U4077 ( .A(n6564), .ZN(n6571) );
  INV_X1 U4078 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6765) );
  NOR2_X1 U4079 ( .A1(n6519), .A2(n6565), .ZN(n6758) );
  INV_X1 U4080 ( .A(n6763), .ZN(n6766) );
  INV_X1 U4081 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6512) );
  AND2_X1 U4082 ( .A1(n4944), .A2(n5187), .ZN(n5846) );
  NOR2_X1 U4083 ( .A1(n6519), .A2(n5903), .ZN(n6554) );
  NOR2_X1 U4084 ( .A1(n6519), .A2(n5129), .ZN(n6553) );
  INV_X1 U4085 ( .A(n5131), .ZN(n5276) );
  NAND2_X1 U4086 ( .A1(n5188), .A2(n5187), .ZN(n6628) );
  INV_X1 U4087 ( .A(n6535), .ZN(n6589) );
  NOR2_X1 U4088 ( .A1(n4757), .A2(n5903), .ZN(n5958) );
  NOR2_X2 U4089 ( .A1(n4757), .A2(n5129), .ZN(n5837) );
  INV_X1 U4090 ( .A(n6672), .ZN(n6787) );
  AND2_X1 U4091 ( .A1(n3803), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6664) );
  NOR2_X1 U4092 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6665) );
  NAND2_X1 U4093 ( .A1(n3274), .A2(n3270), .ZN(U2797) );
  OR2_X1 U4094 ( .A1(n5532), .A2(n6318), .ZN(n3274) );
  INV_X1 U4095 ( .A(n3271), .ZN(n3270) );
  OAI21_X1 U4096 ( .B1(n5506), .B2(n6278), .A(n3272), .ZN(n3271) );
  OR2_X1 U4097 ( .A1(n5506), .A2(n5714), .ZN(n4296) );
  AND2_X2 U4098 ( .A1(n4588), .A2(n4581), .ZN(n3516) );
  OR3_X1 U4099 ( .A1(n4757), .A2(n5863), .A3(n5862), .ZN(n3235) );
  INV_X1 U4100 ( .A(n3448), .ZN(n3474) );
  OR2_X1 U4101 ( .A1(n3184), .A2(n7009), .ZN(n3236) );
  AND2_X1 U4102 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n5472), .ZN(n3237)
         );
  OR2_X1 U4103 ( .A1(n5581), .A2(n5580), .ZN(n3238) );
  NAND2_X1 U4104 ( .A1(n3321), .A2(n3254), .ZN(n5682) );
  OR2_X1 U4105 ( .A1(n3481), .A2(n3329), .ZN(n3240) );
  NAND2_X1 U4106 ( .A1(n3318), .A2(n3316), .ZN(n4438) );
  NAND2_X1 U4107 ( .A1(n3318), .A2(n3319), .ZN(n5631) );
  NOR2_X1 U4108 ( .A1(n5560), .A2(n3303), .ZN(n5447) );
  NAND2_X1 U4109 ( .A1(n3448), .A2(n3376), .ZN(n3742) );
  AND4_X1 U4110 ( .A1(n3385), .A2(n3384), .A3(n3383), .A4(n3382), .ZN(n3241)
         );
  AND2_X1 U4111 ( .A1(n3253), .A2(n3726), .ZN(n3242) );
  INV_X1 U4112 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5499) );
  NOR2_X1 U4113 ( .A1(n5406), .A2(n5405), .ZN(n5407) );
  OAI21_X1 U4114 ( .B1(n5764), .B2(n3315), .A(n3313), .ZN(n3737) );
  NAND2_X1 U4115 ( .A1(n5553), .A2(n3296), .ZN(n3243) );
  INV_X1 U4116 ( .A(n3321), .ZN(n5692) );
  NOR2_X1 U4117 ( .A1(n3737), .A2(n5646), .ZN(n5640) );
  AND2_X1 U4118 ( .A1(n3297), .A2(n5412), .ZN(n3244) );
  AND2_X1 U4119 ( .A1(n3279), .A2(n5083), .ZN(n3245) );
  AND2_X1 U4120 ( .A1(n5640), .A2(n5472), .ZN(n3246) );
  AND2_X1 U4121 ( .A1(n3674), .A2(n3703), .ZN(n3936) );
  NAND2_X1 U4122 ( .A1(n3184), .A2(n4490), .ZN(n3247) );
  OR2_X1 U4123 ( .A1(n5352), .A2(n3311), .ZN(n3248) );
  AND2_X1 U4124 ( .A1(n3247), .A2(n3254), .ZN(n3249) );
  NOR2_X1 U4125 ( .A1(n5406), .A2(n3294), .ZN(n5577) );
  AND2_X1 U4126 ( .A1(n3249), .A2(n3734), .ZN(n3250) );
  NAND2_X1 U4127 ( .A1(n3288), .A2(n3286), .ZN(n4663) );
  AND2_X2 U4128 ( .A1(n5495), .A2(n3338), .ZN(n3641) );
  NOR2_X1 U4129 ( .A1(n4800), .A2(n4799), .ZN(n4801) );
  NAND2_X1 U4130 ( .A1(n3322), .A2(n3726), .ZN(n5164) );
  NAND2_X1 U4131 ( .A1(n3265), .A2(n5165), .ZN(n5306) );
  NAND2_X1 U4132 ( .A1(n3312), .A2(n5308), .ZN(n5349) );
  OR2_X1 U4133 ( .A1(n3866), .A2(n5288), .ZN(n3251) );
  NAND2_X1 U4134 ( .A1(n3323), .A2(n3458), .ZN(n4468) );
  OR2_X1 U4135 ( .A1(n5508), .A2(REIP_REG_29__SCAN_IN), .ZN(n3252) );
  NAND2_X1 U4136 ( .A1(n3184), .A2(n5168), .ZN(n3253) );
  NAND2_X1 U4137 ( .A1(n3184), .A2(n5785), .ZN(n3254) );
  AND2_X1 U4138 ( .A1(n3184), .A2(n6130), .ZN(n3255) );
  INV_X1 U4139 ( .A(n3308), .ZN(n4606) );
  NAND2_X1 U4140 ( .A1(n3473), .A2(n3472), .ZN(n3308) );
  OR2_X1 U4141 ( .A1(n4576), .A2(n6780), .ZN(n3256) );
  NAND2_X1 U4142 ( .A1(n3632), .A2(n3631), .ZN(n6426) );
  INV_X1 U4143 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6783) );
  INV_X1 U4144 ( .A(n3201), .ZN(n6757) );
  INV_X1 U4145 ( .A(n4329), .ZN(n4683) );
  AND2_X1 U4146 ( .A1(n4683), .A2(n3281), .ZN(n3257) );
  NAND2_X1 U4147 ( .A1(n5656), .A2(n4496), .ZN(n3258) );
  INV_X1 U4148 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5487) );
  NOR2_X1 U4149 ( .A1(n4743), .A2(n4727), .ZN(n3259) );
  NAND2_X1 U4150 ( .A1(n6745), .A2(n4687), .ZN(n4743) );
  INV_X1 U4151 ( .A(n3235), .ZN(n3260) );
  NOR3_X4 U4152 ( .A1(n6519), .A2(n5863), .A3(n5862), .ZN(n5938) );
  OAI21_X2 U4153 ( .B1(n3491), .B2(n3490), .A(n3573), .ZN(n4622) );
  NAND2_X2 U4154 ( .A1(n3597), .A2(n3598), .ZN(n3599) );
  NAND2_X1 U4155 ( .A1(n3322), .A2(n3266), .ZN(n3264) );
  NAND2_X2 U4156 ( .A1(n3448), .A2(n4483), .ZN(n3269) );
  NAND2_X4 U4157 ( .A1(n3239), .A2(n3181), .ZN(n4483) );
  NAND3_X1 U4158 ( .A1(n4683), .A2(n3281), .A3(n4673), .ZN(n4707) );
  AND2_X2 U4159 ( .A1(n5333), .A2(n3283), .ZN(n5586) );
  NAND2_X1 U4160 ( .A1(n3919), .A2(n3287), .ZN(n3286) );
  INV_X1 U4161 ( .A(n4578), .ZN(n3287) );
  NAND2_X1 U4162 ( .A1(n4665), .A2(n4664), .ZN(n3288) );
  INV_X1 U4163 ( .A(n3919), .ZN(n3289) );
  NAND2_X1 U4164 ( .A1(n3462), .A2(n3290), .ZN(n4625) );
  INV_X1 U4165 ( .A(n5406), .ZN(n3291) );
  NAND2_X1 U4166 ( .A1(n3291), .A2(n3292), .ZN(n5571) );
  NAND3_X1 U4167 ( .A1(n3473), .A2(n3472), .A3(n4318), .ZN(n4300) );
  NAND2_X1 U4168 ( .A1(n3659), .A2(n3309), .ZN(n3703) );
  NAND2_X1 U4169 ( .A1(n3659), .A2(n3658), .ZN(n3673) );
  NAND2_X2 U4170 ( .A1(n3725), .A2(n3236), .ZN(n3322) );
  NAND3_X1 U4171 ( .A1(n3323), .A2(n3458), .A3(n4319), .ZN(n3466) );
  OAI21_X1 U4172 ( .B1(n3920), .B2(n3269), .A(n3596), .ZN(n3634) );
  XNOR2_X1 U4173 ( .A(n3741), .B(n3740), .ZN(n5475) );
  INV_X1 U4174 ( .A(n5654), .ZN(n5670) );
  NAND2_X1 U4175 ( .A1(n5665), .A2(n7098), .ZN(n5435) );
  NAND2_X1 U4176 ( .A1(n5433), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U4177 ( .A1(n4301), .A2(n4727), .ZN(n3456) );
  AND2_X1 U4178 ( .A1(n3467), .A2(n4688), .ZN(n3459) );
  AND2_X1 U4179 ( .A1(n5863), .A2(n5862), .ZN(n5187) );
  INV_X1 U4180 ( .A(n5862), .ZN(n4751) );
  INV_X1 U4181 ( .A(n5339), .ZN(n6330) );
  OR2_X1 U4182 ( .A1(n6349), .A2(n6348), .ZN(n4536) );
  OR3_X1 U4183 ( .A1(n6777), .A2(n4349), .A3(n4412), .ZN(n6318) );
  INV_X1 U4184 ( .A(n6318), .ZN(n4435) );
  NOR2_X1 U4185 ( .A1(n5863), .A2(n4751), .ZN(n3324) );
  AND2_X1 U4186 ( .A1(n3456), .A2(n3455), .ZN(n3325) );
  INV_X1 U4187 ( .A(n4686), .ZN(n3593) );
  INV_X1 U4188 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4442) );
  INV_X1 U4189 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6165) );
  INV_X1 U4190 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5428) );
  OR3_X1 U4191 ( .A1(n5716), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n4503), 
        .ZN(n3327) );
  INV_X1 U4192 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3631) );
  NAND2_X1 U4193 ( .A1(n6780), .A2(n6781), .ZN(n4269) );
  BUF_X4 U4194 ( .A(n3551), .Z(n4280) );
  AND2_X1 U4195 ( .A1(n3480), .A2(n3207), .ZN(n3329) );
  AND2_X1 U4196 ( .A1(n6633), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3748)
         );
  AND2_X1 U4197 ( .A1(n3671), .A2(n3670), .ZN(n3672) );
  OR2_X1 U4198 ( .A1(n3522), .A2(n3521), .ZN(n3620) );
  NAND2_X1 U4199 ( .A1(n4318), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3743) );
  OR2_X1 U4200 ( .A1(n3669), .A2(n3668), .ZN(n3678) );
  OR2_X1 U4201 ( .A1(n3590), .A2(n3589), .ZN(n3595) );
  NAND2_X1 U4202 ( .A1(n3783), .A2(n3782), .ZN(n3794) );
  AOI22_X1 U4203 ( .A1(n3433), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3225), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3349) );
  INV_X1 U4204 ( .A(n3743), .ZN(n3503) );
  OR2_X1 U4205 ( .A1(n3563), .A2(n6783), .ZN(n3716) );
  AND2_X1 U4206 ( .A1(n3479), .A2(n3478), .ZN(n3480) );
  NAND2_X1 U4207 ( .A1(n4742), .A2(n4318), .ZN(n3457) );
  INV_X1 U4208 ( .A(n3899), .ZN(n3809) );
  NOR2_X1 U4209 ( .A1(n4243), .A2(n7068), .ZN(n4265) );
  NOR2_X1 U4210 ( .A1(n4115), .A2(n5666), .ZN(n4144) );
  OR2_X1 U4211 ( .A1(n3951), .A2(n3952), .ZN(n3981) );
  INV_X1 U4212 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3808) );
  INV_X1 U4213 ( .A(n4390), .ZN(n4394) );
  NAND2_X1 U4214 ( .A1(n3580), .A2(n3579), .ZN(n3799) );
  NAND2_X1 U4215 ( .A1(n3526), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3425) );
  NAND2_X1 U4216 ( .A1(n3809), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3867)
         );
  INV_X1 U4217 ( .A(n5572), .ZN(n4118) );
  INV_X1 U4218 ( .A(n4779), .ZN(n3934) );
  NAND2_X1 U4219 ( .A1(n4225), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4243)
         );
  AND2_X1 U4220 ( .A1(n4101), .A2(n4100), .ZN(n5578) );
  INV_X1 U4221 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3810) );
  INV_X1 U4222 ( .A(n3916), .ZN(n3921) );
  AND2_X1 U4223 ( .A1(n4486), .A2(n4479), .ZN(n4495) );
  NAND2_X1 U4224 ( .A1(n4322), .A2(n4406), .ZN(n4562) );
  AND2_X1 U4225 ( .A1(n3574), .A2(n4737), .ZN(n4894) );
  NOR2_X1 U4226 ( .A1(n6969), .A2(n3867), .ZN(n3868) );
  INV_X1 U4227 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6969) );
  NAND2_X1 U4228 ( .A1(n3921), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3929)
         );
  OR2_X1 U4229 ( .A1(n5395), .A2(n4349), .ZN(n4390) );
  AND2_X1 U4230 ( .A1(n4188), .A2(n4187), .ZN(n5515) );
  XNOR2_X1 U4231 ( .A(n4316), .B(n5421), .ZN(n5456) );
  NOR2_X1 U4232 ( .A1(n4164), .A2(n3813), .ZN(n4185) );
  NAND2_X1 U4233 ( .A1(n4099), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4115)
         );
  INV_X1 U4234 ( .A(n3987), .ZN(n3996) );
  INV_X1 U4235 ( .A(n6442), .ZN(n5707) );
  OR2_X1 U4236 ( .A1(n3184), .A2(n5428), .ZN(n5430) );
  NAND2_X1 U4237 ( .A1(n5299), .A2(n5253), .ZN(n5178) );
  AND2_X1 U4238 ( .A1(n4482), .A2(n5089), .ZN(n5799) );
  OR2_X1 U4239 ( .A1(n4582), .A2(n5126), .ZN(n5014) );
  AND2_X1 U4240 ( .A1(n3201), .A2(n4656), .ZN(n4944) );
  NAND2_X1 U4241 ( .A1(n4944), .A2(n4821), .ZN(n4924) );
  INV_X1 U4242 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6637) );
  AND2_X1 U4243 ( .A1(n6561), .A2(n3486), .ZN(n4787) );
  OR2_X1 U4244 ( .A1(n3201), .A2(n4816), .ZN(n6566) );
  NAND2_X1 U4245 ( .A1(n3578), .A2(n3577), .ZN(n6513) );
  INV_X1 U4246 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6633) );
  INV_X1 U4247 ( .A(n4269), .ZN(n4311) );
  NAND2_X1 U4248 ( .A1(n4433), .A2(n3252), .ZN(n4434) );
  OR2_X1 U4249 ( .A1(n6197), .A2(n4423), .ZN(n6085) );
  NAND2_X1 U4250 ( .A1(n6777), .A2(n4313), .ZN(n6296) );
  NAND2_X1 U4251 ( .A1(n3937), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3945)
         );
  INV_X1 U4252 ( .A(n6246), .ZN(n6325) );
  OAI21_X1 U4253 ( .B1(n6782), .B2(n6683), .A(n4526), .ZN(n6416) );
  INV_X1 U4254 ( .A(n6363), .ZN(n6792) );
  NAND2_X1 U4255 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n4185), .ZN(n4205)
         );
  NOR2_X1 U4256 ( .A1(n5287), .A2(n5288), .ZN(n5298) );
  AND2_X1 U4257 ( .A1(n4648), .A2(n6664), .ZN(n4556) );
  OR2_X1 U4258 ( .A1(n5761), .A2(n4494), .ZN(n5745) );
  NAND2_X1 U4259 ( .A1(n5799), .A2(n6499), .ZN(n6501) );
  INV_X1 U4260 ( .A(n5441), .ZN(n6141) );
  AND2_X1 U4261 ( .A1(n4709), .A2(n4500), .ZN(n5359) );
  INV_X1 U4262 ( .A(n5089), .ZN(n6488) );
  NAND2_X1 U4263 ( .A1(n4648), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5808) );
  NAND2_X1 U4264 ( .A1(n4944), .A2(n3324), .ZN(n5838) );
  AND2_X1 U4265 ( .A1(n4944), .A2(n4853), .ZN(n5847) );
  OAI21_X1 U4266 ( .B1(n4826), .B2(n4825), .A(n4824), .ZN(n4849) );
  INV_X1 U4267 ( .A(n5897), .ZN(n4930) );
  OAI21_X1 U4268 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n7152), .A(n4895), 
        .ZN(n6570) );
  INV_X1 U4269 ( .A(n5905), .ZN(n5934) );
  NOR2_X2 U4270 ( .A1(n6566), .A2(n4988), .ZN(n5952) );
  INV_X1 U4271 ( .A(n6628), .ZN(n6613) );
  INV_X1 U4272 ( .A(n6617), .ZN(n6622) );
  OAI211_X1 U4273 ( .C1(n5964), .C2(n7152), .A(n5963), .B(n5962), .ZN(n6002)
         );
  INV_X1 U4274 ( .A(n6551), .ZN(n6614) );
  NOR2_X1 U4275 ( .A1(n6749), .A2(n6780), .ZN(n6669) );
  INV_X1 U4276 ( .A(STATE_REG_0__SCAN_IN), .ZN(n7054) );
  CLKBUF_X1 U4277 ( .A(n6738), .Z(n6732) );
  NAND2_X1 U4278 ( .A1(n4556), .A2(n4514), .ZN(n5505) );
  INV_X1 U4279 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6781) );
  AOI21_X1 U4280 ( .B1(n4436), .B2(n4435), .A(n4434), .ZN(n4437) );
  INV_X1 U4281 ( .A(n6272), .ZN(n6314) );
  OR2_X1 U4282 ( .A1(n6777), .A2(n4416), .ZN(n6246) );
  NAND2_X1 U4283 ( .A1(n6296), .A2(n4317), .ZN(n6278) );
  INV_X1 U4284 ( .A(n6027), .ZN(n5607) );
  INV_X1 U4285 ( .A(n5702), .ZN(n5348) );
  NAND2_X1 U4286 ( .A1(n4557), .A2(n6421), .ZN(n5593) );
  INV_X2 U4287 ( .A(n4536), .ZN(n6358) );
  INV_X1 U4288 ( .A(n6416), .ZN(n6363) );
  NOR2_X1 U4290 ( .A1(n5745), .A2(n4497), .ZN(n6131) );
  NOR2_X1 U4291 ( .A1(n5791), .A2(n5359), .ZN(n6161) );
  INV_X1 U4292 ( .A(n6425), .ZN(n6498) );
  INV_X1 U4293 ( .A(n6507), .ZN(n6475) );
  INV_X1 U4294 ( .A(n5843), .ZN(n4887) );
  INV_X1 U4295 ( .A(n6554), .ZN(n5940) );
  INV_X1 U4296 ( .A(n6553), .ZN(n5278) );
  NAND2_X1 U4297 ( .A1(n5188), .A2(n3324), .ZN(n5131) );
  NAND2_X1 U4298 ( .A1(n5188), .A2(n4821), .ZN(n6617) );
  NAND2_X1 U4299 ( .A1(n4752), .A2(n3324), .ZN(n4977) );
  INV_X1 U4300 ( .A(n5958), .ZN(n6010) );
  INV_X1 U4301 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6749) );
  INV_X1 U4302 ( .A(n6743), .ZN(n6741) );
  INV_X1 U4303 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6682) );
  OAI21_X1 U4304 ( .B1(n5623), .B2(n6278), .A(n4437), .ZN(U2798) );
  INV_X1 U4305 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3331) );
  AND2_X2 U4306 ( .A1(n3331), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3339)
         );
  AOI22_X1 U4307 ( .A1(n3545), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3225), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3337) );
  NOR2_X4 U4308 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4589) );
  AOI22_X1 U4309 ( .A1(n3422), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3336) );
  AOI22_X1 U4310 ( .A1(n3526), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3213), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3335) );
  AND2_X2 U4311 ( .A1(n4592), .A2(n3333), .ZN(n3551) );
  AOI22_X1 U4312 ( .A1(n3214), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3551), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4313 ( .A1(n3233), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3210), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3342) );
  AOI22_X1 U4314 ( .A1(n3641), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3231), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3341) );
  AOI22_X1 U4315 ( .A1(n3546), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3528), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3340) );
  AOI22_X1 U4316 ( .A1(n3234), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3348) );
  AOI22_X1 U4317 ( .A1(n3545), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3210), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3347) );
  AOI22_X1 U4318 ( .A1(n3546), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3214), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3346) );
  AOI22_X1 U4319 ( .A1(n3422), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3511), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4320 ( .A1(n3528), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3516), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3352) );
  AOI22_X1 U4321 ( .A1(n3527), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3551), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3351) );
  INV_X1 U4322 ( .A(n3467), .ZN(n3377) );
  NAND2_X1 U4323 ( .A1(n3545), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3359)
         );
  NAND2_X1 U4324 ( .A1(n3225), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3358) );
  NAND2_X1 U4325 ( .A1(n3422), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3357) );
  NAND2_X1 U4326 ( .A1(n3183), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3356) );
  NAND2_X1 U4327 ( .A1(n3234), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3363) );
  NAND2_X1 U4328 ( .A1(n3641), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3362) );
  NAND2_X1 U4329 ( .A1(n4279), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3361)
         );
  NAND2_X1 U4330 ( .A1(n3516), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3360)
         );
  NAND2_X1 U4331 ( .A1(n3511), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3367) );
  NAND2_X1 U4332 ( .A1(n3546), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3366)
         );
  NAND2_X1 U4333 ( .A1(n3428), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3365)
         );
  NAND2_X1 U4334 ( .A1(n3528), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3364)
         );
  NAND2_X1 U4335 ( .A1(n3526), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3371) );
  NAND2_X1 U4336 ( .A1(n3433), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3370) );
  NAND2_X1 U4337 ( .A1(n3214), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3369) );
  NAND2_X1 U4338 ( .A1(n3551), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3368) );
  NAND2_X1 U4339 ( .A1(n3474), .A2(n3460), .ZN(n3387) );
  AOI22_X1 U4340 ( .A1(n3526), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3433), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3381) );
  AOI22_X1 U4341 ( .A1(n3545), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3380) );
  AOI22_X1 U4342 ( .A1(n3215), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3379) );
  AOI22_X1 U4343 ( .A1(n3211), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4344 ( .A1(n3234), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3385) );
  AOI22_X1 U4345 ( .A1(n3511), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3384) );
  AOI22_X1 U4346 ( .A1(n3641), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3516), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3383) );
  AOI22_X1 U4347 ( .A1(n3546), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3528), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4348 ( .A1(n3526), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3433), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3391) );
  AOI22_X1 U4349 ( .A1(n3545), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3390) );
  AOI22_X1 U4350 ( .A1(n3215), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3551), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3389) );
  AOI22_X1 U4351 ( .A1(n3422), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3388) );
  NAND4_X1 U4352 ( .A1(n3391), .A2(n3390), .A3(n3389), .A4(n3388), .ZN(n3397)
         );
  AOI22_X1 U4353 ( .A1(n3427), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4279), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3395) );
  AOI22_X1 U4354 ( .A1(n3511), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4355 ( .A1(n3641), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3516), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3393) );
  AOI22_X1 U4356 ( .A1(n3546), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3392) );
  NAND4_X1 U4357 ( .A1(n3395), .A2(n3394), .A3(n3393), .A4(n3392), .ZN(n3396)
         );
  AOI22_X1 U4358 ( .A1(n3545), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3641), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3401) );
  AOI22_X1 U4359 ( .A1(n3546), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3511), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3400) );
  AOI22_X1 U4360 ( .A1(n3427), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3215), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3399) );
  AOI22_X1 U4361 ( .A1(n3526), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3422), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3405) );
  AOI22_X1 U4362 ( .A1(n4279), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3404) );
  AOI22_X1 U4363 ( .A1(n3226), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3528), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3403) );
  AOI22_X1 U4364 ( .A1(n3433), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3551), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3402) );
  NOR2_X1 U4365 ( .A1(n3466), .A2(n4469), .ZN(n3806) );
  OAI21_X1 U4366 ( .B1(n3460), .B2(n3409), .A(n4576), .ZN(n3407) );
  INV_X1 U4367 ( .A(n3407), .ZN(n3413) );
  AND2_X1 U4368 ( .A1(n3460), .A2(n3448), .ZN(n3408) );
  NAND2_X1 U4369 ( .A1(n4742), .A2(n3408), .ZN(n3412) );
  NAND2_X1 U4370 ( .A1(n3742), .A2(n4469), .ZN(n3411) );
  NAND2_X1 U4371 ( .A1(n3467), .A2(n4319), .ZN(n3410) );
  AOI22_X1 U4372 ( .A1(n3526), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3417) );
  AOI22_X1 U4373 ( .A1(n3545), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3225), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3416) );
  AOI22_X1 U4374 ( .A1(n3214), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3551), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3415) );
  AOI22_X1 U4375 ( .A1(n3211), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3414) );
  AOI22_X1 U4376 ( .A1(n3427), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3209), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3421) );
  AOI22_X1 U4377 ( .A1(n3511), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3428), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3420) );
  AOI22_X1 U4378 ( .A1(n3641), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3419) );
  AOI22_X1 U4379 ( .A1(n3546), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3418) );
  NAND2_X1 U4380 ( .A1(n3641), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3426) );
  NAND2_X1 U4381 ( .A1(n4279), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3424)
         );
  NAND2_X1 U4382 ( .A1(n3422), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3423) );
  NAND2_X1 U4383 ( .A1(n3427), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3432) );
  NAND2_X1 U4384 ( .A1(n3545), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3431)
         );
  NAND2_X1 U4385 ( .A1(n3428), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3430)
         );
  NAND2_X1 U4386 ( .A1(n3182), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3429) );
  NAND2_X1 U4387 ( .A1(n3433), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3438) );
  NAND2_X1 U4388 ( .A1(n3225), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3437) );
  NAND2_X1 U4389 ( .A1(n3551), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3436) );
  NAND2_X1 U4390 ( .A1(n3214), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3435) );
  NAND2_X1 U4391 ( .A1(n3546), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3442)
         );
  NAND2_X1 U4392 ( .A1(n3511), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3441) );
  NAND2_X1 U4393 ( .A1(n3516), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3440)
         );
  NAND2_X1 U4394 ( .A1(n3528), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3439)
         );
  NAND2_X1 U4395 ( .A1(n3456), .A2(n4716), .ZN(n3451) );
  NAND2_X1 U4396 ( .A1(n3467), .A2(n4318), .ZN(n3447) );
  NAND2_X2 U4397 ( .A1(n4318), .A2(n4727), .ZN(n4510) );
  NAND2_X1 U4398 ( .A1(n4445), .A2(n3409), .ZN(n3450) );
  XNOR2_X1 U4399 ( .A(n6691), .B(STATE_REG_1__SCAN_IN), .ZN(n4413) );
  OR2_X1 U4400 ( .A1(n3476), .A2(n3448), .ZN(n3449) );
  NAND2_X1 U4401 ( .A1(n6665), .A2(n6783), .ZN(n3815) );
  MUX2_X1 U4402 ( .A(n3803), .B(n3815), .S(n6633), .Z(n3453) );
  INV_X1 U4403 ( .A(n3454), .ZN(n3455) );
  INV_X2 U4404 ( .A(n4510), .ZN(n6782) );
  NAND2_X1 U4405 ( .A1(n3459), .A2(n3458), .ZN(n4446) );
  NAND2_X1 U4406 ( .A1(n6665), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6169) );
  INV_X1 U4407 ( .A(n6169), .ZN(n3463) );
  NAND3_X1 U4408 ( .A1(n4583), .A2(n3463), .A3(n4625), .ZN(n3464) );
  AND2_X1 U4409 ( .A1(n3467), .A2(n3409), .ZN(n3468) );
  OAI21_X1 U4410 ( .B1(n3466), .B2(n3468), .A(n4483), .ZN(n3469) );
  INV_X1 U4411 ( .A(n4446), .ZN(n3473) );
  NAND2_X1 U4412 ( .A1(n4742), .A2(n4319), .ZN(n3622) );
  NAND2_X1 U4413 ( .A1(n4727), .A2(n4716), .ZN(n5216) );
  INV_X1 U4414 ( .A(n5216), .ZN(n4509) );
  AND2_X1 U4415 ( .A1(n3460), .A2(n4576), .ZN(n4452) );
  NAND2_X1 U4416 ( .A1(n4553), .A2(n4452), .ZN(n4458) );
  AND2_X1 U4417 ( .A1(n4302), .A2(n4727), .ZN(n3475) );
  OAI211_X1 U4418 ( .C1(n4300), .C2(n3476), .A(n4458), .B(n4636), .ZN(n3477)
         );
  NAND2_X1 U4419 ( .A1(n3477), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3481) );
  NAND2_X1 U4420 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3485) );
  OAI21_X1 U4421 ( .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n3485), .ZN(n4893) );
  OR2_X1 U4422 ( .A1(n3815), .A2(n4893), .ZN(n3479) );
  INV_X1 U4423 ( .A(n3803), .ZN(n3575) );
  NAND2_X1 U4424 ( .A1(n3575), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3478) );
  OAI211_X1 U4425 ( .C1(n3483), .C2(n3207), .A(n3481), .B(n3480), .ZN(n3508)
         );
  NAND2_X1 U4426 ( .A1(n3510), .A2(n3508), .ZN(n3482) );
  INV_X1 U4427 ( .A(n3485), .ZN(n3484) );
  NAND2_X1 U4428 ( .A1(n3484), .A2(n6643), .ZN(n6561) );
  NAND2_X1 U4429 ( .A1(n3485), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3486) );
  OAI22_X1 U4430 ( .A1(n4787), .A2(n3815), .B1(n3803), .B2(n6643), .ZN(n3487)
         );
  AOI22_X1 U4431 ( .A1(n4595), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3433), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3496) );
  AOI22_X1 U4432 ( .A1(n4274), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3495) );
  AOI22_X1 U4433 ( .A1(n3215), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3494) );
  AOI22_X1 U4434 ( .A1(n3219), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3493) );
  NAND4_X1 U4435 ( .A1(n3496), .A2(n3495), .A3(n3494), .A4(n3493), .ZN(n3502)
         );
  AOI22_X1 U4436 ( .A1(n3427), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3500) );
  AOI22_X1 U4437 ( .A1(n3229), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4281), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3499) );
  INV_X1 U4438 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n7080) );
  AOI22_X1 U4439 ( .A1(n3216), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3231), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3498) );
  AOI22_X1 U4440 ( .A1(n3222), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3497) );
  NAND4_X1 U4441 ( .A1(n3500), .A2(n3499), .A3(n3498), .A4(n3497), .ZN(n3501)
         );
  INV_X1 U4442 ( .A(n3580), .ZN(n3505) );
  AOI22_X1 U4443 ( .A1(n3795), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3505), 
        .B2(n3504), .ZN(n3506) );
  XNOR2_X2 U4444 ( .A(n3507), .B(n3506), .ZN(n3597) );
  NAND2_X1 U4445 ( .A1(n3240), .A2(n3508), .ZN(n3509) );
  XNOR2_X1 U4446 ( .A(n3510), .B(n3509), .ZN(n4652) );
  NAND2_X1 U4447 ( .A1(n4652), .A2(n6783), .ZN(n3525) );
  INV_X1 U4448 ( .A(n3579), .ZN(n3523) );
  AOI22_X1 U4449 ( .A1(n3526), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3222), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3515) );
  AOI22_X1 U4450 ( .A1(n3212), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3219), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3514) );
  AOI22_X1 U4451 ( .A1(n3226), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3513) );
  AOI22_X1 U4452 ( .A1(n3185), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4281), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3512) );
  NAND4_X1 U4453 ( .A1(n3515), .A2(n3514), .A3(n3513), .A4(n3512), .ZN(n3522)
         );
  AOI22_X1 U4454 ( .A1(n3234), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3215), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3520) );
  AOI22_X1 U4455 ( .A1(n3216), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3519) );
  AOI22_X1 U4456 ( .A1(n3182), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3518) );
  AOI22_X1 U4457 ( .A1(n4274), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3517) );
  NAND4_X1 U4458 ( .A1(n3520), .A2(n3519), .A3(n3518), .A4(n3517), .ZN(n3521)
         );
  NAND2_X1 U4459 ( .A1(n3523), .A2(n3620), .ZN(n3524) );
  INV_X1 U4460 ( .A(n3620), .ZN(n3541) );
  NAND2_X1 U4461 ( .A1(n3795), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3540) );
  AOI22_X1 U4462 ( .A1(n4274), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3216), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3532) );
  AOI22_X1 U4463 ( .A1(n3526), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4281), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3531) );
  AOI22_X1 U4464 ( .A1(n3213), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3530) );
  AOI22_X1 U4465 ( .A1(n3546), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3529) );
  NAND4_X1 U4466 ( .A1(n3532), .A2(n3531), .A3(n3530), .A4(n3529), .ZN(n3538)
         );
  AOI22_X1 U4467 ( .A1(n3427), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3536) );
  AOI22_X1 U4468 ( .A1(n4279), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3215), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3535) );
  AOI22_X1 U4469 ( .A1(n3219), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3534) );
  AOI22_X1 U4470 ( .A1(n3226), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3516), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3533) );
  NAND4_X1 U4471 ( .A1(n3536), .A2(n3535), .A3(n3534), .A4(n3533), .ZN(n3537)
         );
  NOR2_X1 U4472 ( .A1(n3579), .A2(n3718), .ZN(n3561) );
  INV_X1 U4473 ( .A(n3561), .ZN(n3539) );
  NAND2_X1 U4474 ( .A1(n3615), .A2(n3614), .ZN(n3568) );
  NAND2_X1 U4475 ( .A1(n3203), .A2(n3543), .ZN(n3542) );
  OAI21_X1 U4476 ( .B1(n3204), .B2(n3543), .A(n3542), .ZN(n3910) );
  NAND2_X1 U4477 ( .A1(n3910), .A2(n6783), .ZN(n3560) );
  NAND2_X1 U4478 ( .A1(n4688), .A2(n3718), .ZN(n3563) );
  AOI22_X1 U4479 ( .A1(n4595), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3433), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3550) );
  AOI22_X1 U4480 ( .A1(n4274), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3549) );
  AOI22_X1 U4481 ( .A1(n3234), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4281), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3548) );
  AOI22_X1 U4482 ( .A1(n3222), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3215), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3547) );
  NAND4_X1 U4483 ( .A1(n3550), .A2(n3549), .A3(n3548), .A4(n3547), .ZN(n3557)
         );
  AOI22_X1 U4484 ( .A1(n3226), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3185), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3555) );
  AOI22_X1 U4485 ( .A1(n3216), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4486 ( .A1(n3219), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3553) );
  AOI22_X1 U4487 ( .A1(n4251), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3552) );
  NAND4_X1 U4488 ( .A1(n3555), .A2(n3554), .A3(n3553), .A4(n3552), .ZN(n3556)
         );
  OR2_X1 U4489 ( .A1(n3563), .A2(n3621), .ZN(n3558) );
  NAND2_X1 U4490 ( .A1(n3561), .A2(n3621), .ZN(n3607) );
  AND2_X1 U4491 ( .A1(n3607), .A2(n3716), .ZN(n3562) );
  NAND2_X1 U4492 ( .A1(n3604), .A2(n3562), .ZN(n3567) );
  NAND2_X1 U4493 ( .A1(n3795), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3566) );
  AOI21_X1 U4494 ( .B1(n4716), .B2(n3621), .A(n6783), .ZN(n3564) );
  AND2_X1 U4495 ( .A1(n3564), .A2(n3563), .ZN(n3565) );
  NAND2_X1 U4496 ( .A1(n3566), .A2(n3565), .ZN(n3606) );
  NAND2_X1 U4497 ( .A1(n3568), .A2(n3616), .ZN(n3572) );
  INV_X1 U4498 ( .A(n3615), .ZN(n3570) );
  INV_X1 U4499 ( .A(n3614), .ZN(n3569) );
  NAND2_X1 U4500 ( .A1(n3570), .A2(n3569), .ZN(n3571) );
  INV_X1 U4501 ( .A(n3815), .ZN(n3576) );
  NOR3_X1 U4502 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6643), .A3(n6637), 
        .ZN(n6524) );
  NAND2_X1 U4503 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6524), .ZN(n6515) );
  NAND2_X1 U4504 ( .A1(n6765), .A2(n6515), .ZN(n3574) );
  NAND3_X1 U4505 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5957) );
  INV_X1 U4506 ( .A(n5957), .ZN(n4695) );
  NAND2_X1 U4507 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4695), .ZN(n4737) );
  AOI22_X1 U4508 ( .A1(n3576), .A2(n4894), .B1(n3575), .B2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3577) );
  XNOR2_X2 U4509 ( .A(n3573), .B(n6513), .ZN(n4582) );
  AOI22_X1 U4510 ( .A1(n4595), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3213), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3584) );
  AOI22_X1 U4511 ( .A1(n3233), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3216), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3583) );
  AOI22_X1 U4512 ( .A1(n3215), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3582) );
  AOI22_X1 U4513 ( .A1(n4281), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3581) );
  NAND4_X1 U4514 ( .A1(n3584), .A2(n3583), .A3(n3582), .A4(n3581), .ZN(n3590)
         );
  AOI22_X1 U4515 ( .A1(n4274), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3588) );
  AOI22_X1 U4516 ( .A1(n3222), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3185), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3587) );
  AOI22_X1 U4517 ( .A1(n3219), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4518 ( .A1(n3220), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3231), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3585) );
  NAND4_X1 U4519 ( .A1(n3588), .A2(n3587), .A3(n3586), .A4(n3585), .ZN(n3589)
         );
  AOI22_X1 U4520 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(n3795), .B1(n3799), 
        .B2(n3595), .ZN(n3591) );
  NAND2_X1 U4521 ( .A1(n3599), .A2(n4686), .ZN(n3594) );
  NAND2_X1 U4522 ( .A1(n3620), .A2(n3621), .ZN(n3619) );
  NAND2_X1 U4523 ( .A1(n3619), .A2(n3601), .ZN(n3600) );
  NAND2_X1 U4524 ( .A1(n3600), .A2(n3595), .ZN(n3677) );
  OAI211_X1 U4525 ( .C1(n3595), .C2(n3600), .A(n3677), .B(n6782), .ZN(n3596)
         );
  INV_X1 U4526 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6482) );
  XNOR2_X1 U4527 ( .A(n3634), .B(n6482), .ZN(n5064) );
  OAI21_X1 U4528 ( .B1(n3601), .B2(n3619), .A(n3600), .ZN(n3602) );
  AND2_X1 U4529 ( .A1(n4716), .A2(n4319), .ZN(n4476) );
  AOI21_X1 U4530 ( .B1(n3602), .B2(n6782), .A(n4476), .ZN(n3603) );
  NAND2_X1 U4531 ( .A1(n3630), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6427)
         );
  NAND2_X1 U4532 ( .A1(n3604), .A2(n3607), .ZN(n3605) );
  NAND2_X1 U4533 ( .A1(n3605), .A2(n3606), .ZN(n3610) );
  INV_X1 U4534 ( .A(n3606), .ZN(n3608) );
  NAND2_X1 U4535 ( .A1(n3608), .A2(n3607), .ZN(n3609) );
  INV_X1 U4536 ( .A(n4476), .ZN(n3611) );
  OAI21_X1 U4537 ( .B1(n4510), .B2(n3621), .A(n3611), .ZN(n3612) );
  INV_X1 U4538 ( .A(n3612), .ZN(n3613) );
  OAI21_X1 U4539 ( .B1(n5862), .B2(n3269), .A(n3613), .ZN(n4561) );
  NAND2_X1 U4540 ( .A1(n4561), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4560)
         );
  XNOR2_X1 U4541 ( .A(n4560), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5056)
         );
  NAND2_X1 U4542 ( .A1(n4650), .A2(n3221), .ZN(n3627) );
  OAI21_X1 U4543 ( .B1(n3621), .B2(n3620), .A(n3619), .ZN(n3624) );
  INV_X1 U4544 ( .A(n3622), .ZN(n3623) );
  OAI211_X1 U4545 ( .C1(n3624), .C2(n4510), .A(n3623), .B(n3448), .ZN(n3625)
         );
  INV_X1 U4546 ( .A(n3625), .ZN(n3626) );
  NAND2_X1 U4547 ( .A1(n3627), .A2(n3626), .ZN(n5055) );
  NAND2_X1 U4548 ( .A1(n5056), .A2(n5055), .ZN(n5057) );
  INV_X1 U4549 ( .A(n4560), .ZN(n3628) );
  NAND2_X1 U4550 ( .A1(n3628), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3629)
         );
  AND2_X1 U4551 ( .A1(n5057), .A2(n3629), .ZN(n6428) );
  NAND2_X1 U4552 ( .A1(n6427), .A2(n6428), .ZN(n3633) );
  INV_X1 U4553 ( .A(n3630), .ZN(n3632) );
  NAND2_X1 U4554 ( .A1(n5064), .A2(n5063), .ZN(n3636) );
  NAND2_X1 U4555 ( .A1(n3634), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3635)
         );
  NAND2_X1 U4556 ( .A1(n3636), .A2(n3635), .ZN(n4668) );
  NAND2_X1 U4557 ( .A1(n3795), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3649) );
  AOI22_X1 U4558 ( .A1(n4595), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3213), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4559 ( .A1(n4274), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4560 ( .A1(n3215), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3638) );
  AOI22_X1 U4561 ( .A1(n3219), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3637) );
  NAND4_X1 U4562 ( .A1(n3640), .A2(n3639), .A3(n3638), .A4(n3637), .ZN(n3647)
         );
  AOI22_X1 U4563 ( .A1(n3427), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4564 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n4281), .B1(n3185), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4565 ( .A1(n3216), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3516), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3643) );
  AOI22_X1 U4566 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3222), .B1(n4251), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3642) );
  NAND4_X1 U4567 ( .A1(n3645), .A2(n3644), .A3(n3643), .A4(n3642), .ZN(n3646)
         );
  NAND2_X1 U4568 ( .A1(n3799), .A2(n3675), .ZN(n3648) );
  NAND2_X1 U4569 ( .A1(n3933), .A2(n3221), .ZN(n3652) );
  XNOR2_X1 U4570 ( .A(n3677), .B(n3675), .ZN(n3650) );
  NAND2_X1 U4571 ( .A1(n3650), .A2(n6782), .ZN(n3651) );
  NAND2_X1 U4572 ( .A1(n3652), .A2(n3651), .ZN(n3654) );
  INV_X1 U4573 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3653) );
  NAND2_X1 U4574 ( .A1(n4668), .A2(n4669), .ZN(n3656) );
  NAND2_X1 U4575 ( .A1(n3654), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3655)
         );
  NAND2_X1 U4576 ( .A1(n3656), .A2(n3655), .ZN(n4703) );
  INV_X1 U4577 ( .A(n3657), .ZN(n3659) );
  NAND2_X1 U4578 ( .A1(n3795), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4579 ( .A1(n4274), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4580 ( .A1(n3222), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3662) );
  AOI22_X1 U4581 ( .A1(n3433), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3661) );
  AOI22_X1 U4582 ( .A1(n3234), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3660) );
  NAND4_X1 U4583 ( .A1(n3663), .A2(n3662), .A3(n3661), .A4(n3660), .ZN(n3669)
         );
  AOI22_X1 U4584 ( .A1(n3216), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4585 ( .A1(n4595), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3215), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3666) );
  AOI22_X1 U4586 ( .A1(n3219), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3665) );
  AOI22_X1 U4587 ( .A1(n4281), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3664) );
  NAND4_X1 U4588 ( .A1(n3667), .A2(n3666), .A3(n3665), .A4(n3664), .ZN(n3668)
         );
  NAND2_X1 U4589 ( .A1(n3799), .A2(n3678), .ZN(n3670) );
  NAND2_X1 U4590 ( .A1(n3673), .A2(n3672), .ZN(n3674) );
  NAND2_X1 U4591 ( .A1(n3936), .A2(n3221), .ZN(n3681) );
  INV_X1 U4592 ( .A(n3675), .ZN(n3676) );
  NOR2_X1 U4593 ( .A1(n3677), .A2(n3676), .ZN(n3679) );
  NAND2_X1 U4594 ( .A1(n3679), .A2(n3678), .ZN(n3707) );
  OAI211_X1 U4595 ( .C1(n3679), .C2(n3678), .A(n3707), .B(n6782), .ZN(n3680)
         );
  NAND2_X1 U4596 ( .A1(n3681), .A2(n3680), .ZN(n3682) );
  INV_X1 U4597 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4710) );
  XNOR2_X1 U4598 ( .A(n3682), .B(n4710), .ZN(n4702) );
  NAND2_X1 U4599 ( .A1(n4703), .A2(n4702), .ZN(n3684) );
  NAND2_X1 U4600 ( .A1(n3682), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3683)
         );
  NAND2_X1 U4601 ( .A1(n3684), .A2(n3683), .ZN(n4804) );
  AOI22_X1 U4602 ( .A1(n4595), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3213), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U4603 ( .A1(n4274), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4604 ( .A1(n3215), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U4605 ( .A1(n3219), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3685) );
  NAND4_X1 U4606 ( .A1(n3688), .A2(n3687), .A3(n3686), .A4(n3685), .ZN(n3694)
         );
  AOI22_X1 U4607 ( .A1(n3233), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3692) );
  AOI22_X1 U4608 ( .A1(n3185), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4281), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3691) );
  AOI22_X1 U4609 ( .A1(n3216), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3231), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3690) );
  INV_X1 U4610 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n7140) );
  AOI22_X1 U4611 ( .A1(n3222), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3689) );
  NAND4_X1 U4612 ( .A1(n3692), .A2(n3691), .A3(n3690), .A4(n3689), .ZN(n3693)
         );
  NAND2_X1 U4613 ( .A1(n3799), .A2(n3708), .ZN(n3696) );
  NAND2_X1 U4614 ( .A1(n3795), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3695) );
  XNOR2_X1 U4615 ( .A(n3703), .B(n3704), .ZN(n3942) );
  NAND2_X1 U4616 ( .A1(n3942), .A2(n3221), .ZN(n3699) );
  XNOR2_X1 U4617 ( .A(n3707), .B(n3708), .ZN(n3697) );
  NAND2_X1 U4618 ( .A1(n3697), .A2(n6782), .ZN(n3698) );
  NAND2_X1 U4619 ( .A1(n3699), .A2(n3698), .ZN(n3700) );
  INV_X1 U4620 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5086) );
  NAND2_X1 U4621 ( .A1(n4804), .A2(n4805), .ZN(n3702) );
  NAND2_X1 U4622 ( .A1(n3700), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3701)
         );
  INV_X1 U4623 ( .A(n3703), .ZN(n3705) );
  NAND2_X1 U4624 ( .A1(n3705), .A2(n3704), .ZN(n3715) );
  AOI22_X1 U4625 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n3795), .B1(n3799), 
        .B2(n3718), .ZN(n3706) );
  INV_X1 U4626 ( .A(n3707), .ZN(n3709) );
  NAND2_X1 U4627 ( .A1(n3709), .A2(n3708), .ZN(n3720) );
  XNOR2_X1 U4628 ( .A(n3720), .B(n3718), .ZN(n3710) );
  NAND2_X1 U4629 ( .A1(n3710), .A2(n6782), .ZN(n3711) );
  INV_X1 U4630 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6470) );
  NAND2_X1 U4631 ( .A1(n5109), .A2(n5110), .ZN(n3714) );
  NAND2_X1 U4632 ( .A1(n3712), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3713)
         );
  NAND2_X1 U4633 ( .A1(n3714), .A2(n3713), .ZN(n5081) );
  NOR2_X1 U4634 ( .A1(n3716), .A2(n3269), .ZN(n3717) );
  NAND2_X1 U4635 ( .A1(n6782), .A2(n3718), .ZN(n3719) );
  OR2_X1 U4636 ( .A1(n3720), .A2(n3719), .ZN(n3721) );
  NAND2_X1 U4637 ( .A1(n3728), .A2(n3721), .ZN(n3722) );
  INV_X1 U4638 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U4639 ( .A1(n3722), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3723)
         );
  NAND2_X1 U4640 ( .A1(n3724), .A2(n3723), .ZN(n5157) );
  INV_X1 U4641 ( .A(n5157), .ZN(n3725) );
  INV_X1 U4642 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n7009) );
  NAND2_X1 U4643 ( .A1(n3184), .A2(n7009), .ZN(n3726) );
  INV_X1 U4644 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5168) );
  OR2_X1 U4645 ( .A1(n3184), .A2(n5168), .ZN(n5165) );
  INV_X1 U4646 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n7122) );
  NAND2_X1 U4647 ( .A1(n3184), .A2(n7122), .ZN(n5307) );
  OR2_X1 U4648 ( .A1(n3184), .A2(n7122), .ZN(n5308) );
  INV_X1 U4649 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4352) );
  NOR2_X1 U4650 ( .A1(n3184), .A2(n4352), .ZN(n5352) );
  NAND2_X1 U4651 ( .A1(n3184), .A2(n4352), .ZN(n5350) );
  NAND2_X1 U4652 ( .A1(n3727), .A2(n5350), .ZN(n5383) );
  XNOR2_X1 U4653 ( .A(n3184), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5385)
         );
  NAND2_X1 U4654 ( .A1(n5383), .A2(n5385), .ZN(n5384) );
  INV_X1 U4655 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5792) );
  NAND2_X1 U4656 ( .A1(n3184), .A2(n5792), .ZN(n3729) );
  NAND2_X1 U4657 ( .A1(n5384), .A2(n3729), .ZN(n5705) );
  INV_X1 U4658 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4488) );
  OR2_X1 U4659 ( .A1(n3184), .A2(n4488), .ZN(n3730) );
  NAND2_X1 U4660 ( .A1(n3184), .A2(n4488), .ZN(n3731) );
  NAND2_X1 U4661 ( .A1(n3732), .A2(n3731), .ZN(n5697) );
  XNOR2_X1 U4662 ( .A(n3184), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5698)
         );
  NAND2_X1 U4663 ( .A1(n5697), .A2(n5698), .ZN(n5683) );
  INV_X1 U4664 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3733) );
  NAND2_X1 U4665 ( .A1(n3184), .A2(n3733), .ZN(n3734) );
  INV_X1 U4666 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U4667 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4490) );
  INV_X1 U4668 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U4669 ( .A1(n6145), .A2(n5785), .ZN(n5685) );
  OAI21_X1 U4670 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5685), .A(n5663), 
        .ZN(n3735) );
  NOR2_X1 U4671 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6133) );
  NOR2_X1 U4672 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5443) );
  NOR2_X1 U4673 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5748) );
  NAND3_X1 U4674 ( .A1(n6133), .A2(n5443), .A3(n5748), .ZN(n3736) );
  NAND2_X1 U4675 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U4676 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6134) );
  NOR2_X1 U4677 ( .A1(n5750), .A2(n6134), .ZN(n5656) );
  AND2_X1 U4678 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4496) );
  INV_X1 U4679 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6130) );
  XNOR2_X1 U4680 ( .A(n3184), .B(n6130), .ZN(n6103) );
  AND2_X1 U4681 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5472) );
  OR2_X1 U4682 ( .A1(n3184), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5647)
         );
  INV_X1 U4683 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5634) );
  INV_X1 U4684 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U4685 ( .A1(n5634), .A2(n5725), .ZN(n5718) );
  NOR2_X1 U4686 ( .A1(n5647), .A2(n5718), .ZN(n5484) );
  NAND2_X1 U4687 ( .A1(n5484), .A2(n5487), .ZN(n4439) );
  INV_X1 U4688 ( .A(n4439), .ZN(n3738) );
  INV_X1 U4689 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3740) );
  XNOR2_X1 U4690 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3752) );
  AOI21_X1 U4691 ( .B1(n3742), .B2(n3752), .A(n3743), .ZN(n3745) );
  NAND2_X1 U4692 ( .A1(n4727), .A2(n3448), .ZN(n3744) );
  NAND2_X1 U4693 ( .A1(n5216), .A2(n3744), .ZN(n3768) );
  OR2_X1 U4694 ( .A1(n3745), .A2(n3768), .ZN(n3757) );
  INV_X1 U4695 ( .A(n3748), .ZN(n3747) );
  XNOR2_X1 U4696 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3749) );
  INV_X1 U4697 ( .A(n3749), .ZN(n3746) );
  NAND2_X1 U4698 ( .A1(n3747), .A2(n3746), .ZN(n3750) );
  NAND2_X1 U4699 ( .A1(n3749), .A2(n3748), .ZN(n3762) );
  AND2_X1 U4700 ( .A1(n3750), .A2(n3762), .ZN(n4305) );
  INV_X1 U4701 ( .A(n4305), .ZN(n3756) );
  NAND2_X1 U4702 ( .A1(n3799), .A2(n4483), .ZN(n3751) );
  NAND2_X1 U4703 ( .A1(n3751), .A2(n3448), .ZN(n3758) );
  AND2_X1 U4704 ( .A1(n3799), .A2(n3752), .ZN(n3753) );
  OAI211_X1 U4705 ( .C1(n3758), .C2(n4305), .A(n3753), .B(n3757), .ZN(n3754)
         );
  NAND2_X1 U4706 ( .A1(n3754), .A2(n3796), .ZN(n3755) );
  OAI21_X1 U4707 ( .B1(n3757), .B2(n3756), .A(n3755), .ZN(n3760) );
  NAND3_X1 U4708 ( .A1(n3758), .A2(STATE2_REG_0__SCAN_IN), .A3(n4305), .ZN(
        n3759) );
  NAND2_X1 U4709 ( .A1(n3760), .A2(n3759), .ZN(n3766) );
  NAND2_X1 U4710 ( .A1(n6637), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3761) );
  NAND2_X1 U4711 ( .A1(n3762), .A2(n3761), .ZN(n3771) );
  XNOR2_X1 U4712 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3770) );
  INV_X1 U4713 ( .A(n3770), .ZN(n3763) );
  XNOR2_X1 U4714 ( .A(n3771), .B(n3763), .ZN(n4306) );
  INV_X1 U4715 ( .A(n3795), .ZN(n3775) );
  NAND2_X1 U4716 ( .A1(n3799), .A2(n4306), .ZN(n3767) );
  INV_X1 U4717 ( .A(n3768), .ZN(n3764) );
  OAI211_X1 U4718 ( .C1(n4306), .C2(n3775), .A(n3767), .B(n3764), .ZN(n3765)
         );
  NAND2_X1 U4719 ( .A1(n3766), .A2(n3765), .ZN(n3778) );
  INV_X1 U4720 ( .A(n3767), .ZN(n3769) );
  NAND2_X1 U4721 ( .A1(n3769), .A2(n3768), .ZN(n3777) );
  NAND2_X1 U4722 ( .A1(n3771), .A2(n3770), .ZN(n3773) );
  NAND2_X1 U4723 ( .A1(n6643), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3772) );
  NAND2_X1 U4724 ( .A1(n3773), .A2(n3772), .ZN(n3781) );
  XNOR2_X1 U4725 ( .A(n6765), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3779)
         );
  XNOR2_X1 U4726 ( .A(n3781), .B(n3779), .ZN(n4304) );
  INV_X1 U4727 ( .A(n4304), .ZN(n3774) );
  INV_X1 U4728 ( .A(n3779), .ZN(n3780) );
  NAND2_X1 U4729 ( .A1(n3781), .A2(n3780), .ZN(n3783) );
  NAND2_X1 U4730 ( .A1(n6765), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3782) );
  INV_X1 U4731 ( .A(n3794), .ZN(n3785) );
  NAND2_X1 U4732 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6165), .ZN(n3793) );
  INV_X1 U4733 ( .A(n3793), .ZN(n3784) );
  NAND3_X1 U4734 ( .A1(n3221), .A2(n3785), .A3(n3784), .ZN(n3788) );
  NAND2_X1 U4735 ( .A1(n6783), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3787) );
  OAI211_X1 U4736 ( .C1(n3796), .C2(n4304), .A(n3788), .B(n3787), .ZN(n3789)
         );
  OAI22_X1 U4737 ( .A1(n3796), .A2(n4308), .B1(n3795), .B2(n4303), .ZN(n3797)
         );
  INV_X1 U4738 ( .A(n3797), .ZN(n3801) );
  INV_X1 U4739 ( .A(n4308), .ZN(n3798) );
  NAND2_X1 U4740 ( .A1(n3409), .A2(n4576), .ZN(n3804) );
  NAND2_X1 U4741 ( .A1(n6630), .A2(n4716), .ZN(n3805) );
  AND2_X1 U4742 ( .A1(n3806), .A2(n3805), .ZN(n4457) );
  INV_X1 U4743 ( .A(n3742), .ZN(n3807) );
  INV_X1 U4744 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3811) );
  INV_X1 U4745 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5666) );
  INV_X1 U4746 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3813) );
  INV_X1 U4747 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n7068) );
  NAND2_X1 U4748 ( .A1(n4265), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4315)
         );
  XNOR2_X1 U4749 ( .A(n4315), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5509)
         );
  INV_X1 U4750 ( .A(n5509), .ZN(n3822) );
  AND2_X1 U4751 ( .A1(n6571), .A2(n3815), .ZN(n6778) );
  OR2_X1 U4752 ( .A1(n6778), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3816) );
  NAND2_X1 U4753 ( .A1(n6783), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3818) );
  NAND2_X1 U4754 ( .A1(n6781), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3817) );
  NAND2_X1 U4755 ( .A1(n3818), .A2(n3817), .ZN(n6441) );
  INV_X1 U4756 ( .A(n6441), .ZN(n3819) );
  OR2_X2 U4757 ( .A1(n6442), .A2(n3819), .ZN(n6437) );
  INV_X1 U4758 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4314) );
  AND2_X1 U4759 ( .A1(n6564), .A2(n6749), .ZN(n5502) );
  AND2_X2 U4760 ( .A1(n5502), .A2(n6783), .ZN(n6425) );
  NAND2_X1 U4761 ( .A1(n6425), .A2(REIP_REG_30__SCAN_IN), .ZN(n5467) );
  OAI21_X1 U4762 ( .B1(n5707), .B2(n4314), .A(n5467), .ZN(n3820) );
  INV_X1 U4763 ( .A(n3820), .ZN(n3821) );
  OAI21_X1 U4764 ( .B1(n3822), .B2(n6437), .A(n3821), .ZN(n3823) );
  INV_X1 U4765 ( .A(n3823), .ZN(n4297) );
  XOR2_X1 U4766 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3824), .Z(n6232) );
  AOI22_X1 U4767 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3427), .B1(n4595), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3828) );
  AOI22_X1 U4768 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n3216), .B1(n3222), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4769 ( .A1(n3215), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4770 ( .A1(n3226), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3825) );
  NAND4_X1 U4771 ( .A1(n3828), .A2(n3827), .A3(n3826), .A4(n3825), .ZN(n3834)
         );
  AOI22_X1 U4772 ( .A1(n3212), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4281), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4773 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n4274), .B1(n3220), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4774 ( .A1(n3219), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3830) );
  AOI22_X1 U4775 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n3185), .B1(n4251), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3829) );
  NAND4_X1 U4776 ( .A1(n3832), .A2(n3831), .A3(n3830), .A4(n3829), .ZN(n3833)
         );
  OR2_X1 U4777 ( .A1(n3834), .A2(n3833), .ZN(n3835) );
  NAND2_X1 U4778 ( .A1(n6780), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4014) );
  AOI22_X1 U4779 ( .A1(n3996), .A2(n3835), .B1(n5414), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3837) );
  INV_X2 U4780 ( .A(n3256), .ZN(n5415) );
  NAND2_X1 U4781 ( .A1(n5415), .A2(EAX_REG_12__SCAN_IN), .ZN(n3836) );
  OAI211_X1 U4782 ( .C1(n6232), .C2(n4269), .A(n3837), .B(n3836), .ZN(n5251)
         );
  AOI22_X1 U4783 ( .A1(n3213), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4784 ( .A1(n3216), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4785 ( .A1(n4595), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4786 ( .A1(n4281), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3838) );
  NAND4_X1 U4787 ( .A1(n3841), .A2(n3840), .A3(n3839), .A4(n3838), .ZN(n3847)
         );
  AOI22_X1 U4788 ( .A1(n4274), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3219), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4789 ( .A1(n3222), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4790 ( .A1(n3215), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3843) );
  AOI22_X1 U4791 ( .A1(n3234), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3516), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3842) );
  NAND4_X1 U4792 ( .A1(n3845), .A2(n3844), .A3(n3843), .A4(n3842), .ZN(n3846)
         );
  NOR2_X1 U4793 ( .A1(n3847), .A2(n3846), .ZN(n3852) );
  XNOR2_X1 U4794 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3848), .ZN(n6243)
         );
  OAI22_X1 U4795 ( .A1(n6243), .A2(n4269), .B1(n4014), .B2(n3810), .ZN(n3849)
         );
  INV_X1 U4796 ( .A(n3849), .ZN(n3851) );
  NAND2_X1 U4797 ( .A1(n5415), .A2(EAX_REG_11__SCAN_IN), .ZN(n3850) );
  OAI211_X1 U4798 ( .C1(n3987), .C2(n3852), .A(n3851), .B(n3850), .ZN(n5297)
         );
  NAND2_X1 U4799 ( .A1(n5251), .A2(n5297), .ZN(n3866) );
  AOI22_X1 U4800 ( .A1(n3234), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4801 ( .A1(n3216), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3185), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4802 ( .A1(n3219), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4803 ( .A1(n3222), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3853) );
  NAND4_X1 U4804 ( .A1(n3856), .A2(n3855), .A3(n3854), .A4(n3853), .ZN(n3862)
         );
  AOI22_X1 U4805 ( .A1(n4274), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4806 ( .A1(n4595), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3215), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4807 ( .A1(n3212), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4808 ( .A1(n4281), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3231), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3857) );
  NAND4_X1 U4809 ( .A1(n3860), .A2(n3859), .A3(n3858), .A4(n3857), .ZN(n3861)
         );
  OAI21_X1 U4810 ( .B1(n3862), .B2(n3861), .A(n3996), .ZN(n3865) );
  XOR2_X1 U4811 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3868), .Z(n6253) );
  INV_X1 U4812 ( .A(n6253), .ZN(n5291) );
  AOI22_X1 U4813 ( .A1(n5414), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n4311), 
        .B2(n5291), .ZN(n3864) );
  NAND2_X1 U4814 ( .A1(n5415), .A2(EAX_REG_10__SCAN_IN), .ZN(n3863) );
  NAND2_X1 U4815 ( .A1(n3867), .A2(n6969), .ZN(n3870) );
  INV_X1 U4816 ( .A(n3868), .ZN(n3869) );
  NAND2_X1 U4817 ( .A1(n3870), .A2(n3869), .ZN(n5160) );
  AOI22_X1 U4818 ( .A1(n3226), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3219), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4819 ( .A1(n3216), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4281), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4820 ( .A1(n3222), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3185), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4821 ( .A1(n3433), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3871) );
  NAND4_X1 U4822 ( .A1(n3874), .A2(n3873), .A3(n3872), .A4(n3871), .ZN(n3880)
         );
  AOI22_X1 U4823 ( .A1(n3233), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4824 ( .A1(n4595), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3215), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4825 ( .A1(n4274), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4826 ( .A1(n4251), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3875) );
  NAND4_X1 U4827 ( .A1(n3878), .A2(n3877), .A3(n3876), .A4(n3875), .ZN(n3879)
         );
  OAI21_X1 U4828 ( .B1(n3880), .B2(n3879), .A(n3996), .ZN(n3883) );
  NAND2_X1 U4829 ( .A1(n5415), .A2(EAX_REG_9__SCAN_IN), .ZN(n3882) );
  NAND2_X1 U4830 ( .A1(n5414), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3881)
         );
  NAND3_X1 U4831 ( .A1(n3883), .A2(n3882), .A3(n3881), .ZN(n3884) );
  AOI21_X1 U4832 ( .B1(n5160), .B2(n4311), .A(n3884), .ZN(n5142) );
  NOR2_X1 U4833 ( .A1(n3251), .A2(n5142), .ZN(n3898) );
  XNOR2_X1 U4834 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3899), .ZN(n5284) );
  AOI22_X1 U4835 ( .A1(n3427), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3216), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4836 ( .A1(n3219), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4837 ( .A1(n3182), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4838 ( .A1(n3229), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3885) );
  NAND4_X1 U4839 ( .A1(n3888), .A2(n3887), .A3(n3886), .A4(n3885), .ZN(n3894)
         );
  AOI22_X1 U4840 ( .A1(n3433), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4841 ( .A1(n3222), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4281), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4842 ( .A1(n4595), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3215), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4843 ( .A1(n4274), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3231), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3889) );
  NAND4_X1 U4844 ( .A1(n3892), .A2(n3891), .A3(n3890), .A4(n3889), .ZN(n3893)
         );
  OR2_X1 U4845 ( .A1(n3894), .A2(n3893), .ZN(n3895) );
  AOI22_X1 U4846 ( .A1(n3996), .A2(n3895), .B1(n5414), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3897) );
  NAND2_X1 U4847 ( .A1(n5415), .A2(EAX_REG_8__SCAN_IN), .ZN(n3896) );
  OAI211_X1 U4848 ( .C1(n5284), .C2(n4269), .A(n3897), .B(n3896), .ZN(n5115)
         );
  AND2_X1 U4849 ( .A1(n3898), .A2(n5115), .ZN(n3905) );
  OAI21_X1 U4850 ( .B1(n3900), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3899), 
        .ZN(n6264) );
  NAND2_X1 U4851 ( .A1(n6264), .A2(n4311), .ZN(n3902) );
  AOI22_X1 U4852 ( .A1(n5415), .A2(EAX_REG_7__SCAN_IN), .B1(n5414), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3901) );
  AND2_X1 U4853 ( .A1(n3902), .A2(n3901), .ZN(n3903) );
  OAI21_X2 U4854 ( .B1(n4656), .B2(n3987), .A(n4014), .ZN(n3919) );
  NAND2_X1 U4855 ( .A1(n4650), .A2(n3996), .ZN(n3909) );
  AOI22_X1 U4856 ( .A1(n5415), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6780), .ZN(n3907) );
  AND2_X1 U4857 ( .A1(n4452), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3915) );
  NAND2_X1 U4858 ( .A1(n3915), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3906) );
  AND2_X1 U4859 ( .A1(n3907), .A2(n3906), .ZN(n3908) );
  NAND2_X1 U4860 ( .A1(n3909), .A2(n3908), .ZN(n4579) );
  AOI21_X1 U4861 ( .B1(n5862), .B2(n3461), .A(n6780), .ZN(n4550) );
  AOI22_X1 U4862 ( .A1(n5415), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6780), .ZN(n3912) );
  NAND2_X1 U4863 ( .A1(n3915), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3911) );
  AND2_X1 U4864 ( .A1(n3912), .A2(n3911), .ZN(n3913) );
  OAI21_X1 U4865 ( .B1(n3230), .B2(n3987), .A(n3913), .ZN(n4549) );
  NAND2_X1 U4866 ( .A1(n4550), .A2(n4549), .ZN(n4552) );
  OR2_X1 U4867 ( .A1(n4549), .A2(n4269), .ZN(n3914) );
  NAND2_X1 U4868 ( .A1(n4552), .A2(n3914), .ZN(n4580) );
  INV_X1 U4869 ( .A(n3915), .ZN(n3928) );
  OAI21_X1 U4870 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3916), .ZN(n6436) );
  AOI22_X1 U4871 ( .A1(n4311), .A2(n6436), .B1(n5414), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3918) );
  NAND2_X1 U4872 ( .A1(n5415), .A2(EAX_REG_2__SCAN_IN), .ZN(n3917) );
  OAI211_X1 U4873 ( .C1(n3928), .C2(n3332), .A(n3918), .B(n3917), .ZN(n4664)
         );
  OAI21_X1 U4874 ( .B1(n3921), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n3929), 
        .ZN(n6320) );
  AOI22_X1 U4875 ( .A1(n6320), .A2(n4311), .B1(n5414), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3923) );
  NAND2_X1 U4876 ( .A1(n5415), .A2(EAX_REG_3__SCAN_IN), .ZN(n3922) );
  OAI211_X1 U4877 ( .C1(n3928), .C2(n4621), .A(n3923), .B(n3922), .ZN(n3924)
         );
  INV_X1 U4878 ( .A(n3924), .ZN(n3925) );
  OAI21_X1 U4879 ( .B1(n3201), .B2(n3987), .A(n3925), .ZN(n4678) );
  NAND2_X1 U4880 ( .A1(n4663), .A2(n4678), .ZN(n4778) );
  OAI21_X1 U4881 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n6781), .A(n6780), 
        .ZN(n3927) );
  NAND2_X1 U4882 ( .A1(n5415), .A2(EAX_REG_4__SCAN_IN), .ZN(n3926) );
  OAI211_X1 U4883 ( .C1(n3928), .C2(n6165), .A(n3927), .B(n3926), .ZN(n3931)
         );
  AOI21_X1 U4884 ( .B1(n3929), .B2(n6300), .A(n3937), .ZN(n6303) );
  NAND2_X1 U4885 ( .A1(n6303), .A2(n4311), .ZN(n3930) );
  AND2_X1 U4886 ( .A1(n3931), .A2(n3930), .ZN(n3932) );
  AOI21_X1 U4887 ( .B1(n3933), .B2(n3996), .A(n3932), .ZN(n4779) );
  INV_X1 U4888 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3940) );
  OAI21_X1 U4889 ( .B1(n3937), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3945), 
        .ZN(n6292) );
  NAND2_X1 U4890 ( .A1(n6292), .A2(n4311), .ZN(n3939) );
  NAND2_X1 U4891 ( .A1(n5414), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3938)
         );
  OAI211_X1 U4892 ( .C1(n3256), .C2(n3940), .A(n3939), .B(n3938), .ZN(n3941)
         );
  NAND2_X1 U4893 ( .A1(n3942), .A2(n3996), .ZN(n3949) );
  INV_X1 U4894 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3944) );
  OAI21_X1 U4895 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6781), .A(n6780), 
        .ZN(n3943) );
  OAI21_X1 U4896 ( .B1(n3256), .B2(n3944), .A(n3943), .ZN(n3947) );
  XNOR2_X1 U4897 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .B(n3945), .ZN(n5099) );
  NAND2_X1 U4898 ( .A1(n5099), .A2(n4311), .ZN(n3946) );
  NAND2_X1 U4899 ( .A1(n3947), .A2(n3946), .ZN(n3948) );
  NAND2_X1 U4900 ( .A1(n3949), .A2(n3948), .ZN(n5009) );
  XNOR2_X1 U4901 ( .A(n3951), .B(n3952), .ZN(n6219) );
  INV_X1 U4902 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6418) );
  OAI22_X1 U4903 ( .A1(n3256), .A2(n6418), .B1(n4014), .B2(n3952), .ZN(n3953)
         );
  AOI21_X1 U4904 ( .B1(n6219), .B2(n4311), .A(n3953), .ZN(n3968) );
  AOI22_X1 U4905 ( .A1(n4595), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3213), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4906 ( .A1(n4274), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4907 ( .A1(n3215), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4908 ( .A1(n3219), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3954) );
  NAND4_X1 U4909 ( .A1(n3957), .A2(n3956), .A3(n3955), .A4(n3954), .ZN(n3963)
         );
  AOI22_X1 U4910 ( .A1(n3427), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4911 ( .A1(n3229), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4281), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4912 ( .A1(n3216), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3516), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4913 ( .A1(n3222), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3958) );
  NAND4_X1 U4914 ( .A1(n3961), .A2(n3960), .A3(n3959), .A4(n3958), .ZN(n3962)
         );
  OR2_X1 U4915 ( .A1(n3963), .A2(n3962), .ZN(n3964) );
  NAND2_X1 U4916 ( .A1(n3996), .A2(n3964), .ZN(n5176) );
  NAND2_X1 U4917 ( .A1(n3966), .A2(n3965), .ZN(n3970) );
  AOI22_X1 U4918 ( .A1(n3226), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3219), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U4919 ( .A1(n4274), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4920 ( .A1(n3222), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3215), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4921 ( .A1(n4595), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3971) );
  NAND4_X1 U4922 ( .A1(n3974), .A2(n3973), .A3(n3972), .A4(n3971), .ZN(n3980)
         );
  AOI22_X1 U4923 ( .A1(n3216), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4924 ( .A1(n4281), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4925 ( .A1(n3234), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4926 ( .A1(n3213), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3975) );
  NAND4_X1 U4927 ( .A1(n3978), .A2(n3977), .A3(n3976), .A4(n3975), .ZN(n3979)
         );
  NOR2_X1 U4928 ( .A1(n3980), .A2(n3979), .ZN(n3986) );
  INV_X1 U4929 ( .A(n3981), .ZN(n3983) );
  INV_X1 U4930 ( .A(n3999), .ZN(n3982) );
  OAI21_X1 U4931 ( .B1(PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n3983), .A(n3982), 
        .ZN(n5241) );
  AOI22_X1 U4932 ( .A1(n4311), .A2(n5241), .B1(n5414), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3985) );
  NAND2_X1 U4933 ( .A1(n5415), .A2(EAX_REG_14__SCAN_IN), .ZN(n3984) );
  OAI211_X1 U4934 ( .C1(n3987), .C2(n3986), .A(n3985), .B(n3984), .ZN(n5183)
         );
  AOI22_X1 U4935 ( .A1(n3219), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4281), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U4936 ( .A1(n3220), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3215), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3990) );
  AOI22_X1 U4937 ( .A1(n3427), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3989) );
  AOI22_X1 U4938 ( .A1(n3183), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3988) );
  NAND4_X1 U4939 ( .A1(n3991), .A2(n3990), .A3(n3989), .A4(n3988), .ZN(n3998)
         );
  AOI22_X1 U4940 ( .A1(n4595), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3222), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U4941 ( .A1(n4274), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3216), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U4942 ( .A1(n3213), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U4943 ( .A1(n3229), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3516), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3992) );
  NAND4_X1 U4944 ( .A1(n3995), .A2(n3994), .A3(n3993), .A4(n3992), .ZN(n3997)
         );
  OAI21_X1 U4945 ( .B1(n3998), .B2(n3997), .A(n3996), .ZN(n4002) );
  OAI21_X1 U4946 ( .B1(PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n3999), .A(n4013), 
        .ZN(n5700) );
  AOI22_X1 U4947 ( .A1(n5414), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n4311), 
        .B2(n5700), .ZN(n4001) );
  NAND2_X1 U4948 ( .A1(n5415), .A2(EAX_REG_15__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4949 ( .A1(n4274), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U4950 ( .A1(n3216), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4281), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4005) );
  AOI22_X1 U4951 ( .A1(n3212), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U4952 ( .A1(n3219), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4003) );
  NAND4_X1 U4953 ( .A1(n4006), .A2(n4005), .A3(n4004), .A4(n4003), .ZN(n4012)
         );
  AOI22_X1 U4954 ( .A1(n3233), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U4955 ( .A1(n4595), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3215), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U4956 ( .A1(n3222), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4957 ( .A1(n3185), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4007) );
  NAND4_X1 U4958 ( .A1(n4010), .A2(n4009), .A3(n4008), .A4(n4007), .ZN(n4011)
         );
  OAI21_X1 U4959 ( .B1(n4012), .B2(n4011), .A(n4290), .ZN(n4017) );
  AOI21_X1 U4960 ( .B1(n6943), .B2(n4013), .A(n4032), .ZN(n6212) );
  OAI22_X1 U4961 ( .A1(n6212), .A2(n4269), .B1(n4014), .B2(n6943), .ZN(n4015)
         );
  AOI21_X1 U4962 ( .B1(n5415), .B2(EAX_REG_16__SCAN_IN), .A(n4015), .ZN(n4016)
         );
  AOI22_X1 U4963 ( .A1(n3427), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3216), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U4964 ( .A1(n4274), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3219), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4020) );
  AOI22_X1 U4965 ( .A1(n3222), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3215), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U4966 ( .A1(n3213), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4018) );
  NAND4_X1 U4967 ( .A1(n4021), .A2(n4020), .A3(n4019), .A4(n4018), .ZN(n4027)
         );
  AOI22_X1 U4968 ( .A1(n3220), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U4969 ( .A1(n4281), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U4970 ( .A1(n3226), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U4971 ( .A1(n4595), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4022) );
  NAND4_X1 U4972 ( .A1(n4025), .A2(n4024), .A3(n4023), .A4(n4022), .ZN(n4026)
         );
  NOR2_X1 U4973 ( .A1(n4027), .A2(n4026), .ZN(n4031) );
  NAND2_X1 U4974 ( .A1(n6780), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4028)
         );
  NAND2_X1 U4975 ( .A1(n4269), .A2(n4028), .ZN(n4029) );
  AOI21_X1 U4976 ( .B1(n5415), .B2(EAX_REG_17__SCAN_IN), .A(n4029), .ZN(n4030)
         );
  OAI21_X1 U4977 ( .B1(n4263), .B2(n4031), .A(n4030), .ZN(n4034) );
  OAI21_X1 U4978 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n4032), .A(n4048), 
        .ZN(n6204) );
  OR2_X1 U4979 ( .A1(n4269), .A2(n6204), .ZN(n4033) );
  AOI22_X1 U4980 ( .A1(n4595), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4038) );
  AOI22_X1 U4981 ( .A1(n4274), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4037) );
  AOI22_X1 U4982 ( .A1(n3215), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4036) );
  AOI22_X1 U4983 ( .A1(n3219), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4035) );
  NAND4_X1 U4984 ( .A1(n4038), .A2(n4037), .A3(n4036), .A4(n4035), .ZN(n4044)
         );
  AOI22_X1 U4985 ( .A1(n3233), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U4986 ( .A1(n3185), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4281), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U4987 ( .A1(n3216), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U4988 ( .A1(n3222), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4039) );
  NAND4_X1 U4989 ( .A1(n4042), .A2(n4041), .A3(n4040), .A4(n4039), .ZN(n4043)
         );
  NOR2_X1 U4990 ( .A1(n4044), .A2(n4043), .ZN(n4047) );
  AOI21_X1 U4991 ( .B1(n3811), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4045) );
  AOI21_X1 U4992 ( .B1(n5415), .B2(EAX_REG_18__SCAN_IN), .A(n4045), .ZN(n4046)
         );
  OAI21_X1 U4993 ( .B1(n4263), .B2(n4047), .A(n4046), .ZN(n4050) );
  XNOR2_X1 U4994 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n4048), .ZN(n6194)
         );
  NAND2_X1 U4995 ( .A1(n6194), .A2(n4311), .ZN(n4049) );
  NAND2_X1 U4996 ( .A1(n4050), .A2(n4049), .ZN(n5391) );
  OR2_X1 U4997 ( .A1(n4053), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4054)
         );
  NAND2_X1 U4998 ( .A1(n4054), .A2(n4082), .ZN(n6115) );
  AOI22_X1 U4999 ( .A1(n4595), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3219), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4058) );
  AOI22_X1 U5000 ( .A1(n3213), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4281), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U5001 ( .A1(n3215), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4056) );
  AOI22_X1 U5002 ( .A1(n3216), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4055) );
  NAND4_X1 U5003 ( .A1(n4058), .A2(n4057), .A3(n4056), .A4(n4055), .ZN(n4064)
         );
  AOI22_X1 U5004 ( .A1(n4274), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4062) );
  AOI22_X1 U5005 ( .A1(n3233), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U5006 ( .A1(n3185), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U5007 ( .A1(n3222), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3516), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4059) );
  NAND4_X1 U5008 ( .A1(n4062), .A2(n4061), .A3(n4060), .A4(n4059), .ZN(n4063)
         );
  NOR2_X1 U5009 ( .A1(n4064), .A2(n4063), .ZN(n4067) );
  OAI21_X1 U5010 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6994), .A(n4269), .ZN(
        n4065) );
  AOI21_X1 U5011 ( .B1(n5415), .B2(EAX_REG_19__SCAN_IN), .A(n4065), .ZN(n4066)
         );
  OAI21_X1 U5012 ( .B1(n4263), .B2(n4067), .A(n4066), .ZN(n4068) );
  OAI21_X1 U5013 ( .B1(n6115), .B2(n4269), .A(n4068), .ZN(n5405) );
  AOI22_X1 U5014 ( .A1(n3433), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3219), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4072) );
  AOI22_X1 U5015 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3216), .B1(n3220), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U5016 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3222), .B1(n3185), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4070) );
  AOI22_X1 U5017 ( .A1(n4595), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4069) );
  NAND4_X1 U5018 ( .A1(n4072), .A2(n4071), .A3(n4070), .A4(n4069), .ZN(n4078)
         );
  AOI22_X1 U5019 ( .A1(n4274), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U5020 ( .A1(n3215), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4075) );
  AOI22_X1 U5021 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n4281), .B1(n4251), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4074) );
  AOI22_X1 U5022 ( .A1(n3234), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3231), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4073) );
  NAND4_X1 U5023 ( .A1(n4076), .A2(n4075), .A3(n4074), .A4(n4073), .ZN(n4077)
         );
  NOR2_X1 U5024 ( .A1(n4078), .A2(n4077), .ZN(n4081) );
  INV_X1 U5025 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6088) );
  OAI21_X1 U5026 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6088), .A(n4269), .ZN(
        n4079) );
  AOI21_X1 U5027 ( .B1(n5415), .B2(EAX_REG_20__SCAN_IN), .A(n4079), .ZN(n4080)
         );
  OAI21_X1 U5028 ( .B1(n4263), .B2(n4081), .A(n4080), .ZN(n4084) );
  XNOR2_X1 U5029 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n4082), .ZN(n6080)
         );
  NAND2_X1 U5030 ( .A1(n6080), .A2(n4311), .ZN(n4083) );
  AOI22_X1 U5031 ( .A1(n4595), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3222), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4088) );
  AOI22_X1 U5032 ( .A1(n3226), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3219), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4087) );
  AOI22_X1 U5033 ( .A1(n3216), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4281), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4086) );
  AOI22_X1 U5034 ( .A1(n3212), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4085) );
  NAND4_X1 U5035 ( .A1(n4088), .A2(n4087), .A3(n4086), .A4(n4085), .ZN(n4094)
         );
  AOI22_X1 U5036 ( .A1(n3220), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4092) );
  AOI22_X1 U5037 ( .A1(n3233), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3215), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4091) );
  AOI22_X1 U5038 ( .A1(n4274), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4090) );
  AOI22_X1 U5039 ( .A1(n4251), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3516), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4089) );
  NAND4_X1 U5040 ( .A1(n4092), .A2(n4091), .A3(n4090), .A4(n4089), .ZN(n4093)
         );
  NOR2_X1 U5041 ( .A1(n4094), .A2(n4093), .ZN(n4098) );
  NAND2_X1 U5042 ( .A1(n6780), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4095)
         );
  NAND2_X1 U5043 ( .A1(n4269), .A2(n4095), .ZN(n4096) );
  AOI21_X1 U5044 ( .B1(n5415), .B2(EAX_REG_21__SCAN_IN), .A(n4096), .ZN(n4097)
         );
  OAI21_X1 U5045 ( .B1(n4263), .B2(n4098), .A(n4097), .ZN(n4101) );
  OAI21_X1 U5046 ( .B1(n4099), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n4115), 
        .ZN(n6070) );
  OR2_X1 U5047 ( .A1(n6070), .A2(n4269), .ZN(n4100) );
  AOI22_X1 U5048 ( .A1(n3212), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3222), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4105) );
  AOI22_X1 U5049 ( .A1(n4274), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U5050 ( .A1(n3216), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4281), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4103) );
  AOI22_X1 U5051 ( .A1(n3226), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4102) );
  NAND4_X1 U5052 ( .A1(n4105), .A2(n4104), .A3(n4103), .A4(n4102), .ZN(n4111)
         );
  AOI22_X1 U5053 ( .A1(n4595), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3427), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U5054 ( .A1(n3219), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U5055 ( .A1(n3215), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U5056 ( .A1(n4251), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3231), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4106) );
  NAND4_X1 U5057 ( .A1(n4109), .A2(n4108), .A3(n4107), .A4(n4106), .ZN(n4110)
         );
  NOR2_X1 U5058 ( .A1(n4111), .A2(n4110), .ZN(n4114) );
  OAI21_X1 U5059 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5666), .A(n4269), .ZN(
        n4112) );
  AOI21_X1 U5060 ( .B1(n5415), .B2(EAX_REG_22__SCAN_IN), .A(n4112), .ZN(n4113)
         );
  OAI21_X1 U5061 ( .B1(n4263), .B2(n4114), .A(n4113), .ZN(n4117) );
  XNOR2_X1 U5062 ( .A(n4115), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6061)
         );
  NAND2_X1 U5063 ( .A1(n6061), .A2(n4311), .ZN(n4116) );
  NAND2_X1 U5064 ( .A1(n4117), .A2(n4116), .ZN(n5572) );
  AOI22_X1 U5065 ( .A1(n4595), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4123) );
  AOI22_X1 U5066 ( .A1(n3234), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4122) );
  AOI22_X1 U5067 ( .A1(n3219), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4121) );
  AOI22_X1 U5068 ( .A1(n3222), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4120) );
  NAND4_X1 U5069 ( .A1(n4123), .A2(n4122), .A3(n4121), .A4(n4120), .ZN(n4129)
         );
  AOI22_X1 U5070 ( .A1(n4274), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4127) );
  AOI22_X1 U5071 ( .A1(n3185), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4281), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4126) );
  AOI22_X1 U5072 ( .A1(n3215), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U5073 ( .A1(n3216), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4124) );
  NAND4_X1 U5074 ( .A1(n4127), .A2(n4126), .A3(n4125), .A4(n4124), .ZN(n4128)
         );
  NOR2_X1 U5075 ( .A1(n4129), .A2(n4128), .ZN(n4151) );
  AOI22_X1 U5076 ( .A1(n4595), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3433), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4133) );
  AOI22_X1 U5077 ( .A1(n4274), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4132) );
  AOI22_X1 U5078 ( .A1(n3215), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U5079 ( .A1(n3219), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4130) );
  NAND4_X1 U5080 ( .A1(n4133), .A2(n4132), .A3(n4131), .A4(n4130), .ZN(n4139)
         );
  AOI22_X1 U5081 ( .A1(n3233), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4137) );
  AOI22_X1 U5082 ( .A1(n3229), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4281), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4136) );
  AOI22_X1 U5083 ( .A1(n3216), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3231), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4135) );
  AOI22_X1 U5084 ( .A1(n3222), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4134) );
  NAND4_X1 U5085 ( .A1(n4137), .A2(n4136), .A3(n4135), .A4(n4134), .ZN(n4138)
         );
  NOR2_X1 U5086 ( .A1(n4139), .A2(n4138), .ZN(n4152) );
  XNOR2_X1 U5087 ( .A(n4151), .B(n4152), .ZN(n4143) );
  NAND2_X1 U5088 ( .A1(n6780), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4140)
         );
  NAND2_X1 U5089 ( .A1(n4269), .A2(n4140), .ZN(n4141) );
  AOI21_X1 U5090 ( .B1(n5415), .B2(EAX_REG_23__SCAN_IN), .A(n4141), .ZN(n4142)
         );
  OAI21_X1 U5091 ( .B1(n4263), .B2(n4143), .A(n4142), .ZN(n4149) );
  INV_X1 U5092 ( .A(n4144), .ZN(n4146) );
  INV_X1 U5093 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4145) );
  NAND2_X1 U5094 ( .A1(n4146), .A2(n4145), .ZN(n4147) );
  NAND2_X1 U5095 ( .A1(n4164), .A2(n4147), .ZN(n6050) );
  NAND2_X1 U5096 ( .A1(n4149), .A2(n4148), .ZN(n5563) );
  NOR2_X1 U5097 ( .A1(n4152), .A2(n4151), .ZN(n4171) );
  AOI22_X1 U5098 ( .A1(n4595), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3213), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4156) );
  AOI22_X1 U5099 ( .A1(n4274), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4155) );
  AOI22_X1 U5100 ( .A1(n3215), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U5101 ( .A1(n3219), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3217), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4153) );
  NAND4_X1 U5102 ( .A1(n4156), .A2(n4155), .A3(n4154), .A4(n4153), .ZN(n4162)
         );
  AOI22_X1 U5103 ( .A1(n3234), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4160) );
  AOI22_X1 U5104 ( .A1(n3185), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4281), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4159) );
  AOI22_X1 U5105 ( .A1(n3216), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4158) );
  AOI22_X1 U5106 ( .A1(n3222), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4157) );
  NAND4_X1 U5107 ( .A1(n4160), .A2(n4159), .A3(n4158), .A4(n4157), .ZN(n4161)
         );
  OR2_X1 U5108 ( .A1(n4162), .A2(n4161), .ZN(n4170) );
  INV_X1 U5109 ( .A(n4170), .ZN(n4163) );
  XNOR2_X1 U5110 ( .A(n4171), .B(n4163), .ZN(n4169) );
  INV_X1 U5111 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4167) );
  XNOR2_X1 U5112 ( .A(n4164), .B(n3813), .ZN(n6040) );
  NAND2_X1 U5113 ( .A1(n6040), .A2(n4311), .ZN(n4166) );
  NAND2_X1 U5114 ( .A1(n5414), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4165)
         );
  OAI211_X1 U5115 ( .C1(n3256), .C2(n4167), .A(n4166), .B(n4165), .ZN(n4168)
         );
  AOI21_X1 U5116 ( .B1(n4169), .B2(n4290), .A(n4168), .ZN(n5448) );
  NAND2_X1 U5117 ( .A1(n4171), .A2(n4170), .ZN(n4189) );
  AOI22_X1 U5118 ( .A1(n4274), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4175) );
  AOI22_X1 U5119 ( .A1(n3427), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4174) );
  AOI22_X1 U5120 ( .A1(n3216), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4281), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4173) );
  AOI22_X1 U5121 ( .A1(n3212), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4172) );
  NAND4_X1 U5122 ( .A1(n4175), .A2(n4174), .A3(n4173), .A4(n4172), .ZN(n4181)
         );
  AOI22_X1 U5123 ( .A1(n4595), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3219), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4179) );
  AOI22_X1 U5124 ( .A1(n3222), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4178) );
  AOI22_X1 U5125 ( .A1(n3215), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4177) );
  AOI22_X1 U5126 ( .A1(n3229), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4176) );
  NAND4_X1 U5127 ( .A1(n4179), .A2(n4178), .A3(n4177), .A4(n4176), .ZN(n4180)
         );
  NOR2_X1 U5128 ( .A1(n4181), .A2(n4180), .ZN(n4190) );
  XNOR2_X1 U5129 ( .A(n4189), .B(n4190), .ZN(n4184) );
  OAI21_X1 U5130 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n7081), .A(n4269), .ZN(
        n4182) );
  AOI21_X1 U5131 ( .B1(n5415), .B2(EAX_REG_25__SCAN_IN), .A(n4182), .ZN(n4183)
         );
  OAI21_X1 U5132 ( .B1(n4184), .B2(n4263), .A(n4183), .ZN(n4188) );
  OR2_X1 U5133 ( .A1(n4185), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4186)
         );
  NAND2_X1 U5134 ( .A1(n4186), .A2(n4205), .ZN(n6109) );
  NOR2_X1 U5135 ( .A1(n4190), .A2(n4189), .ZN(n4220) );
  AOI22_X1 U5136 ( .A1(n4595), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3212), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4194) );
  AOI22_X1 U5137 ( .A1(n4274), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4193) );
  AOI22_X1 U5138 ( .A1(n3215), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4192) );
  AOI22_X1 U5139 ( .A1(n3219), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4191) );
  NAND4_X1 U5140 ( .A1(n4194), .A2(n4193), .A3(n4192), .A4(n4191), .ZN(n4200)
         );
  AOI22_X1 U5141 ( .A1(n3427), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4198) );
  AOI22_X1 U5142 ( .A1(n3229), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4281), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4197) );
  AOI22_X1 U5143 ( .A1(n3216), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3231), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4196) );
  AOI22_X1 U5144 ( .A1(n3222), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4195) );
  NAND4_X1 U5145 ( .A1(n4198), .A2(n4197), .A3(n4196), .A4(n4195), .ZN(n4199)
         );
  OR2_X1 U5146 ( .A1(n4200), .A2(n4199), .ZN(n4219) );
  INV_X1 U5147 ( .A(n4219), .ZN(n4201) );
  XNOR2_X1 U5148 ( .A(n4220), .B(n4201), .ZN(n4202) );
  NAND2_X1 U5149 ( .A1(n4202), .A2(n4290), .ZN(n4208) );
  NAND2_X1 U5150 ( .A1(n6780), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4203)
         );
  NAND2_X1 U5151 ( .A1(n4269), .A2(n4203), .ZN(n4204) );
  AOI21_X1 U5152 ( .B1(n5415), .B2(EAX_REG_26__SCAN_IN), .A(n4204), .ZN(n4207)
         );
  XNOR2_X1 U5153 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .B(n4205), .ZN(n6030)
         );
  AOI21_X1 U5154 ( .B1(n4208), .B2(n4207), .A(n4206), .ZN(n5555) );
  AND2_X2 U5155 ( .A1(n5514), .A2(n5555), .ZN(n5553) );
  AOI22_X1 U5156 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3212), .B1(n3219), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4212) );
  AOI22_X1 U5157 ( .A1(n3226), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4211) );
  AOI22_X1 U5158 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3234), .B1(n3185), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4210) );
  AOI22_X1 U5159 ( .A1(n4595), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4209) );
  NAND4_X1 U5160 ( .A1(n4212), .A2(n4211), .A3(n4210), .A4(n4209), .ZN(n4218)
         );
  AOI22_X1 U5161 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n4274), .B1(n3216), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4216) );
  AOI22_X1 U5162 ( .A1(n3215), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4215) );
  AOI22_X1 U5163 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n3222), .B1(n4251), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4214) );
  AOI22_X1 U5164 ( .A1(n4281), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3231), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4213) );
  NAND4_X1 U5165 ( .A1(n4216), .A2(n4215), .A3(n4214), .A4(n4213), .ZN(n4217)
         );
  NOR2_X1 U5166 ( .A1(n4218), .A2(n4217), .ZN(n4229) );
  NAND2_X1 U5167 ( .A1(n4220), .A2(n4219), .ZN(n4228) );
  XNOR2_X1 U5168 ( .A(n4229), .B(n4228), .ZN(n4224) );
  INV_X1 U5169 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4221) );
  AOI21_X1 U5170 ( .B1(n4221), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4222) );
  AOI21_X1 U5171 ( .B1(n5415), .B2(EAX_REG_27__SCAN_IN), .A(n4222), .ZN(n4223)
         );
  OAI21_X1 U5172 ( .B1(n4224), .B2(n4263), .A(n4223), .ZN(n4227) );
  OAI21_X1 U5173 ( .B1(n4225), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n4243), 
        .ZN(n6021) );
  OR2_X1 U5174 ( .A1(n6021), .A2(n4269), .ZN(n4226) );
  NOR2_X1 U5175 ( .A1(n4229), .A2(n4228), .ZN(n4259) );
  AOI22_X1 U5176 ( .A1(n4595), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3213), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4233) );
  AOI22_X1 U5177 ( .A1(n4274), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4232) );
  AOI22_X1 U5178 ( .A1(n3215), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4231) );
  AOI22_X1 U5179 ( .A1(n3219), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4230) );
  NAND4_X1 U5180 ( .A1(n4233), .A2(n4232), .A3(n4231), .A4(n4230), .ZN(n4239)
         );
  AOI22_X1 U5181 ( .A1(n3233), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4237) );
  AOI22_X1 U5182 ( .A1(n3185), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4281), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4236) );
  AOI22_X1 U5183 ( .A1(n3216), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4235) );
  AOI22_X1 U5184 ( .A1(n3222), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4234) );
  NAND4_X1 U5185 ( .A1(n4237), .A2(n4236), .A3(n4235), .A4(n4234), .ZN(n4238)
         );
  OR2_X1 U5186 ( .A1(n4239), .A2(n4238), .ZN(n4258) );
  XNOR2_X1 U5187 ( .A(n4259), .B(n4258), .ZN(n4242) );
  AOI21_X1 U5188 ( .B1(n7068), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4240) );
  AOI21_X1 U5189 ( .B1(n5415), .B2(EAX_REG_28__SCAN_IN), .A(n4240), .ZN(n4241)
         );
  OAI21_X1 U5190 ( .B1(n4242), .B2(n4263), .A(n4241), .ZN(n4246) );
  AND2_X1 U5191 ( .A1(n4243), .A2(n7068), .ZN(n4244) );
  NOR2_X1 U5192 ( .A1(n4265), .A2(n4244), .ZN(n6012) );
  NAND2_X1 U5193 ( .A1(n6012), .A2(n4311), .ZN(n4245) );
  NAND2_X1 U5194 ( .A1(n4246), .A2(n4245), .ZN(n5536) );
  AOI22_X1 U5195 ( .A1(n4274), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3219), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4250) );
  AOI22_X1 U5196 ( .A1(n3222), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4281), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4249) );
  AOI22_X1 U5197 ( .A1(n4595), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4248) );
  AOI22_X1 U5198 ( .A1(n3233), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3516), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4247) );
  NAND4_X1 U5199 ( .A1(n4250), .A2(n4249), .A3(n4248), .A4(n4247), .ZN(n4257)
         );
  AOI22_X1 U5200 ( .A1(n3433), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3226), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4255) );
  AOI22_X1 U5201 ( .A1(n3216), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4254) );
  AOI22_X1 U5202 ( .A1(n3215), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4253) );
  AOI22_X1 U5203 ( .A1(n3185), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4252) );
  NAND4_X1 U5204 ( .A1(n4255), .A2(n4254), .A3(n4253), .A4(n4252), .ZN(n4256)
         );
  NOR2_X1 U5205 ( .A1(n4257), .A2(n4256), .ZN(n4273) );
  NAND2_X1 U5206 ( .A1(n4259), .A2(n4258), .ZN(n4272) );
  XNOR2_X1 U5207 ( .A(n4273), .B(n4272), .ZN(n4264) );
  NAND2_X1 U5208 ( .A1(n6780), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4260)
         );
  NAND2_X1 U5209 ( .A1(n4269), .A2(n4260), .ZN(n4261) );
  AOI21_X1 U5210 ( .B1(n5415), .B2(EAX_REG_29__SCAN_IN), .A(n4261), .ZN(n4262)
         );
  OAI21_X1 U5211 ( .B1(n4264), .B2(n4263), .A(n4262), .ZN(n4271) );
  INV_X1 U5212 ( .A(n4265), .ZN(n4267) );
  INV_X1 U5213 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4266) );
  NAND2_X1 U5214 ( .A1(n4267), .A2(n4266), .ZN(n4268) );
  NAND2_X1 U5215 ( .A1(n4315), .A2(n4268), .ZN(n5626) );
  NAND2_X1 U5216 ( .A1(n4271), .A2(n4270), .ZN(n4298) );
  NOR2_X1 U5217 ( .A1(n4273), .A2(n4272), .ZN(n4289) );
  AOI22_X1 U5218 ( .A1(n4274), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3234), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4278) );
  AOI22_X1 U5219 ( .A1(n3212), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3219), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4277) );
  AOI22_X1 U5220 ( .A1(n4595), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3215), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4276) );
  AOI22_X1 U5221 ( .A1(n3216), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4251), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4275) );
  NAND4_X1 U5222 ( .A1(n4278), .A2(n4277), .A3(n4276), .A4(n4275), .ZN(n4287)
         );
  AOI22_X1 U5223 ( .A1(n3226), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3220), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4285) );
  AOI22_X1 U5224 ( .A1(n3222), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3185), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4284) );
  AOI22_X1 U5225 ( .A1(n3217), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4280), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4283) );
  AOI22_X1 U5226 ( .A1(n4281), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3232), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4282) );
  NAND4_X1 U5227 ( .A1(n4285), .A2(n4284), .A3(n4283), .A4(n4282), .ZN(n4286)
         );
  NOR2_X1 U5228 ( .A1(n4287), .A2(n4286), .ZN(n4288) );
  XNOR2_X1 U5229 ( .A(n4289), .B(n4288), .ZN(n4291) );
  NAND2_X1 U5230 ( .A1(n4291), .A2(n4290), .ZN(n4295) );
  AOI21_X1 U5231 ( .B1(n4314), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4292) );
  AOI21_X1 U5232 ( .B1(n5415), .B2(EAX_REG_30__SCAN_IN), .A(n4292), .ZN(n4294)
         );
  AND2_X1 U5233 ( .A1(n5509), .A2(n4311), .ZN(n4293) );
  AOI21_X1 U5234 ( .B1(n4295), .B2(n4294), .A(n4293), .ZN(n5412) );
  XNOR2_X1 U5235 ( .A(n5413), .B(n5412), .ZN(n5506) );
  AND2_X1 U5236 ( .A1(n6783), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4310) );
  NAND2_X1 U5237 ( .A1(n4310), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6676) );
  OAI211_X1 U5238 ( .C1(n5475), .C2(n6438), .A(n4297), .B(n4296), .ZN(U2956)
         );
  AND2_X1 U5239 ( .A1(n3243), .A2(n4298), .ZN(n4299) );
  INV_X1 U5240 ( .A(n4300), .ZN(n4514) );
  NAND4_X1 U5241 ( .A1(n4306), .A2(n4305), .A3(n4304), .A4(n4303), .ZN(n4307)
         );
  NAND2_X1 U5242 ( .A1(n4308), .A2(n4307), .ZN(n4512) );
  INV_X1 U5243 ( .A(n4512), .ZN(n4309) );
  NAND2_X1 U5244 ( .A1(n4508), .A2(n6664), .ZN(n5501) );
  NAND2_X1 U5245 ( .A1(n6749), .A2(n6780), .ZN(n6672) );
  NOR3_X1 U5246 ( .A1(n6783), .A2(n7152), .A3(n6672), .ZN(n6659) );
  AND2_X1 U5247 ( .A1(n4311), .A2(n4310), .ZN(n6668) );
  OR2_X1 U5248 ( .A1(n6425), .A2(n6668), .ZN(n4312) );
  NOR2_X1 U5249 ( .A1(n6659), .A2(n4312), .ZN(n4313) );
  INV_X1 U5250 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5421) );
  NOR2_X1 U5251 ( .A1(n5456), .A2(n6749), .ZN(n4317) );
  NAND2_X2 U5252 ( .A1(n4483), .A2(n4319), .ZN(n4406) );
  NAND2_X2 U5253 ( .A1(n4318), .A2(n4483), .ZN(n4349) );
  NAND2_X1 U5254 ( .A1(n5395), .A2(EBX_REG_9__SCAN_IN), .ZN(n4321) );
  NAND2_X1 U5255 ( .A1(n4387), .A2(n7009), .ZN(n4320) );
  OAI211_X1 U5256 ( .C1(n4390), .C2(EBX_REG_9__SCAN_IN), .A(n4321), .B(n4320), 
        .ZN(n5147) );
  OR2_X2 U5257 ( .A1(n4349), .A2(n4406), .ZN(n4401) );
  NAND2_X1 U5258 ( .A1(n4391), .A2(EBX_REG_1__SCAN_IN), .ZN(n4323) );
  NAND2_X1 U5259 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4349), .ZN(n4324)
         );
  OAI211_X2 U5260 ( .C1(n4401), .C2(EBX_REG_1__SCAN_IN), .A(n4325), .B(n4324), 
        .ZN(n4328) );
  NAND2_X1 U5261 ( .A1(n4322), .A2(EBX_REG_0__SCAN_IN), .ZN(n4327) );
  INV_X1 U5262 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5222) );
  NAND2_X1 U5263 ( .A1(n4406), .A2(n5222), .ZN(n4326) );
  XNOR2_X2 U5264 ( .A(n4328), .B(n4563), .ZN(n5313) );
  OAI21_X1 U5265 ( .B1(n5313), .B2(n4349), .A(n4328), .ZN(n4329) );
  NAND2_X1 U5266 ( .A1(n4391), .A2(EBX_REG_2__SCAN_IN), .ZN(n4330) );
  AND2_X1 U5267 ( .A1(n4378), .A2(n4330), .ZN(n4332) );
  NAND3_X1 U5268 ( .A1(n4349), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .A3(n4406), 
        .ZN(n4331) );
  OAI211_X1 U5269 ( .C1(n4401), .C2(EBX_REG_2__SCAN_IN), .A(n4332), .B(n4331), 
        .ZN(n4682) );
  NAND2_X1 U5270 ( .A1(n5395), .A2(EBX_REG_3__SCAN_IN), .ZN(n4334) );
  NAND2_X1 U5271 ( .A1(n4387), .A2(n6482), .ZN(n4333) );
  OAI211_X1 U5272 ( .C1(n4390), .C2(EBX_REG_3__SCAN_IN), .A(n4334), .B(n4333), 
        .ZN(n4680) );
  NAND2_X1 U5273 ( .A1(n4391), .A2(EBX_REG_4__SCAN_IN), .ZN(n4335) );
  AND2_X1 U5274 ( .A1(n4378), .A2(n4335), .ZN(n4337) );
  NAND2_X1 U5275 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n4349), .ZN(n4336)
         );
  OAI211_X1 U5276 ( .C1(n4401), .C2(EBX_REG_4__SCAN_IN), .A(n4337), .B(n4336), 
        .ZN(n4673) );
  NAND2_X1 U5277 ( .A1(n5395), .A2(EBX_REG_5__SCAN_IN), .ZN(n4339) );
  NAND2_X1 U5278 ( .A1(n4387), .A2(n4710), .ZN(n4338) );
  OAI211_X1 U5279 ( .C1(n4390), .C2(EBX_REG_5__SCAN_IN), .A(n4339), .B(n4338), 
        .ZN(n4708) );
  NOR2_X2 U5280 ( .A1(n4707), .A2(n4708), .ZN(n4808) );
  NAND2_X1 U5281 ( .A1(n4322), .A2(n5086), .ZN(n4340) );
  OAI211_X1 U5282 ( .C1(n4349), .C2(EBX_REG_6__SCAN_IN), .A(n4406), .B(n4340), 
        .ZN(n4341) );
  OAI21_X1 U5283 ( .B1(n4401), .B2(EBX_REG_6__SCAN_IN), .A(n4341), .ZN(n4809)
         );
  NAND2_X1 U5284 ( .A1(n5395), .A2(EBX_REG_7__SCAN_IN), .ZN(n4343) );
  NAND2_X1 U5285 ( .A1(n4387), .A2(n6470), .ZN(n4342) );
  OAI211_X1 U5286 ( .C1(n4390), .C2(EBX_REG_7__SCAN_IN), .A(n4343), .B(n4342), 
        .ZN(n5123) );
  NAND2_X1 U5287 ( .A1(n4322), .A2(n5095), .ZN(n4344) );
  OAI211_X1 U5288 ( .C1(n4349), .C2(EBX_REG_8__SCAN_IN), .A(n4406), .B(n4344), 
        .ZN(n4345) );
  OAI21_X1 U5289 ( .B1(n4401), .B2(EBX_REG_8__SCAN_IN), .A(n4345), .ZN(n5083)
         );
  NAND2_X1 U5290 ( .A1(n4391), .A2(EBX_REG_10__SCAN_IN), .ZN(n4346) );
  AND2_X1 U5291 ( .A1(n4378), .A2(n4346), .ZN(n4348) );
  NAND2_X1 U5292 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n4349), .ZN(n4347) );
  OAI211_X1 U5293 ( .C1(n4401), .C2(EBX_REG_10__SCAN_IN), .A(n4348), .B(n4347), 
        .ZN(n5170) );
  INV_X1 U5294 ( .A(n4349), .ZN(n4573) );
  INV_X1 U5295 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U5296 ( .A1(n4573), .A2(n6247), .ZN(n4350) );
  OAI211_X1 U5297 ( .C1(n5395), .C2(n7122), .A(n4350), .B(n4322), .ZN(n4351)
         );
  OAI21_X1 U5298 ( .B1(EBX_REG_11__SCAN_IN), .B2(n4390), .A(n4351), .ZN(n5301)
         );
  NAND2_X1 U5299 ( .A1(n4322), .A2(n4352), .ZN(n4353) );
  OAI211_X1 U5300 ( .C1(n4349), .C2(EBX_REG_12__SCAN_IN), .A(n4406), .B(n4353), 
        .ZN(n4354) );
  OAI21_X1 U5301 ( .B1(n4401), .B2(EBX_REG_12__SCAN_IN), .A(n4354), .ZN(n5253)
         );
  INV_X1 U5302 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5180) );
  AOI22_X1 U5303 ( .A1(n4394), .A2(n5180), .B1(n4387), .B2(n5792), .ZN(n4355)
         );
  OAI21_X1 U5304 ( .B1(n4406), .B2(n5180), .A(n4355), .ZN(n5179) );
  NOR2_X2 U5305 ( .A1(n5178), .A2(n5179), .ZN(n5242) );
  NAND2_X1 U5306 ( .A1(n4391), .A2(EBX_REG_14__SCAN_IN), .ZN(n4356) );
  AND2_X1 U5307 ( .A1(n4378), .A2(n4356), .ZN(n4358) );
  NAND2_X1 U5308 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n4349), .ZN(n4357) );
  OAI211_X1 U5309 ( .C1(n4401), .C2(EBX_REG_14__SCAN_IN), .A(n4358), .B(n4357), 
        .ZN(n5243) );
  INV_X1 U5310 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5340) );
  AOI22_X1 U5311 ( .A1(n4394), .A2(n5340), .B1(n4387), .B2(n3733), .ZN(n4359)
         );
  OAI21_X1 U5312 ( .B1(n4406), .B2(n5340), .A(n4359), .ZN(n5335) );
  NAND2_X1 U5313 ( .A1(n4391), .A2(EBX_REG_16__SCAN_IN), .ZN(n4360) );
  AND2_X1 U5314 ( .A1(n4378), .A2(n4360), .ZN(n4362) );
  NAND2_X1 U5315 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n4349), .ZN(n4361) );
  OAI211_X1 U5316 ( .C1(n4401), .C2(EBX_REG_16__SCAN_IN), .A(n4362), .B(n4361), 
        .ZN(n5373) );
  NAND2_X1 U5317 ( .A1(n4406), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4363) );
  OAI211_X1 U5318 ( .C1(n4349), .C2(EBX_REG_17__SCAN_IN), .A(n4322), .B(n4363), 
        .ZN(n4364) );
  OAI21_X1 U5319 ( .B1(n4390), .B2(EBX_REG_17__SCAN_IN), .A(n4364), .ZN(n5379)
         );
  NAND2_X1 U5320 ( .A1(n4391), .A2(EBX_REG_19__SCAN_IN), .ZN(n4365) );
  AND2_X1 U5321 ( .A1(n4378), .A2(n4365), .ZN(n4367) );
  NAND2_X1 U5322 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n4349), .ZN(n4366) );
  OAI211_X1 U5323 ( .C1(n4401), .C2(EBX_REG_19__SCAN_IN), .A(n4367), .B(n4366), 
        .ZN(n4368) );
  INV_X1 U5324 ( .A(n4368), .ZN(n5409) );
  OR2_X1 U5325 ( .A1(n4349), .A2(EBX_REG_20__SCAN_IN), .ZN(n4369) );
  OAI21_X1 U5326 ( .B1(n4562), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n4369), 
        .ZN(n4370) );
  INV_X1 U5327 ( .A(n4370), .ZN(n5588) );
  OR2_X1 U5328 ( .A1(n4349), .A2(EBX_REG_18__SCAN_IN), .ZN(n5394) );
  OAI21_X1 U5329 ( .B1(n4562), .B2(INSTADDRPOINTER_REG_18__SCAN_IN), .A(n5394), 
        .ZN(n5587) );
  NAND2_X1 U5330 ( .A1(n5395), .A2(EBX_REG_20__SCAN_IN), .ZN(n4372) );
  NAND2_X1 U5331 ( .A1(n5587), .A2(n4406), .ZN(n4371) );
  OAI211_X1 U5332 ( .C1(n5588), .C2(n5587), .A(n4372), .B(n4371), .ZN(n4373)
         );
  INV_X1 U5333 ( .A(n4373), .ZN(n4374) );
  NAND2_X1 U5334 ( .A1(n5586), .A2(n4374), .ZN(n5581) );
  NAND2_X1 U5335 ( .A1(n5395), .A2(EBX_REG_21__SCAN_IN), .ZN(n4376) );
  INV_X1 U5336 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U5337 ( .A1(n4387), .A2(n5756), .ZN(n4375) );
  OAI211_X1 U5338 ( .C1(n4390), .C2(EBX_REG_21__SCAN_IN), .A(n4376), .B(n4375), 
        .ZN(n5580) );
  NAND2_X1 U5339 ( .A1(n4391), .A2(EBX_REG_22__SCAN_IN), .ZN(n4377) );
  AND2_X1 U5340 ( .A1(n4378), .A2(n4377), .ZN(n4380) );
  NAND2_X1 U5341 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n4349), .ZN(n4379) );
  OAI211_X1 U5342 ( .C1(n4401), .C2(EBX_REG_22__SCAN_IN), .A(n4380), .B(n4379), 
        .ZN(n4381) );
  INV_X1 U5343 ( .A(n4381), .ZN(n5568) );
  INV_X1 U5344 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5567) );
  NAND2_X1 U5345 ( .A1(n4394), .A2(n5567), .ZN(n4384) );
  OAI22_X1 U5346 ( .A1(n4562), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5567), .B2(n4406), .ZN(n4382) );
  INV_X1 U5347 ( .A(n4382), .ZN(n4383) );
  AND2_X1 U5348 ( .A1(n4384), .A2(n4383), .ZN(n5564) );
  INV_X1 U5349 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U5350 ( .A1(n4322), .A2(n5444), .ZN(n4385) );
  OAI211_X1 U5351 ( .C1(n4349), .C2(EBX_REG_24__SCAN_IN), .A(n4406), .B(n4385), 
        .ZN(n4386) );
  OAI21_X1 U5352 ( .B1(n4401), .B2(EBX_REG_24__SCAN_IN), .A(n4386), .ZN(n5438)
         );
  NAND2_X1 U5353 ( .A1(n4387), .A2(n6130), .ZN(n4389) );
  NAND2_X1 U5354 ( .A1(n5395), .A2(EBX_REG_25__SCAN_IN), .ZN(n4388) );
  OAI211_X1 U5355 ( .C1(n4390), .C2(EBX_REG_25__SCAN_IN), .A(n4389), .B(n4388), 
        .ZN(n5518) );
  AOI22_X1 U5356 ( .A1(EBX_REG_26__SCAN_IN), .A2(n4391), .B1(n4349), .B2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4392) );
  OAI21_X1 U5357 ( .B1(n4401), .B2(EBX_REG_26__SCAN_IN), .A(n4392), .ZN(n4393)
         );
  INV_X1 U5358 ( .A(n4393), .ZN(n5549) );
  INV_X1 U5359 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U5360 ( .A1(n4394), .A2(n5548), .ZN(n4397) );
  OAI22_X1 U5361 ( .A1(n4562), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .B1(n4406), .B2(n5548), .ZN(n4395) );
  INV_X1 U5362 ( .A(n4395), .ZN(n4396) );
  AND2_X1 U5363 ( .A1(n4397), .A2(n4396), .ZN(n5545) );
  NAND2_X1 U5364 ( .A1(n4322), .A2(n5634), .ZN(n4398) );
  OAI211_X1 U5365 ( .C1(n4349), .C2(EBX_REG_28__SCAN_IN), .A(n4406), .B(n4398), 
        .ZN(n4399) );
  OAI21_X1 U5366 ( .B1(n4401), .B2(EBX_REG_28__SCAN_IN), .A(n4399), .ZN(n5538)
         );
  OR2_X1 U5367 ( .A1(n4349), .A2(EBX_REG_29__SCAN_IN), .ZN(n4400) );
  OAI21_X1 U5368 ( .B1(n4562), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n4400), 
        .ZN(n4409) );
  INV_X1 U5369 ( .A(n4401), .ZN(n4402) );
  INV_X1 U5370 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U5371 ( .A1(n4402), .A2(n5535), .ZN(n4408) );
  INV_X1 U5372 ( .A(n4408), .ZN(n4405) );
  INV_X1 U5373 ( .A(n4403), .ZN(n4404) );
  AOI22_X1 U5374 ( .A1(n5461), .A2(n4406), .B1(n4405), .B2(n4404), .ZN(n4407)
         );
  INV_X1 U5375 ( .A(n4407), .ZN(n4464) );
  OAI211_X1 U5376 ( .C1(n5395), .C2(n4409), .A(n4403), .B(n4408), .ZN(n4410)
         );
  INV_X1 U5377 ( .A(n4410), .ZN(n4411) );
  INV_X1 U5378 ( .A(n5534), .ZN(n4436) );
  INV_X1 U5379 ( .A(READY_N), .ZN(n6683) );
  NAND2_X1 U5380 ( .A1(n6683), .A2(n6781), .ZN(n4418) );
  NAND2_X1 U5381 ( .A1(n4418), .A2(EBX_REG_31__SCAN_IN), .ZN(n4412) );
  NAND2_X1 U5382 ( .A1(n4413), .A2(n7054), .ZN(n6681) );
  NOR3_X1 U5383 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .A3(n6681), .ZN(
        n6656) );
  INV_X1 U5384 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U5385 ( .A1(n4418), .A2(n5530), .ZN(n4414) );
  OAI22_X1 U5386 ( .A1(n4510), .A2(n6656), .B1(n4716), .B2(n4414), .ZN(n4415)
         );
  INV_X1 U5387 ( .A(n4415), .ZN(n4416) );
  NOR2_X1 U5388 ( .A1(n5626), .A2(n6319), .ZN(n4428) );
  INV_X1 U5389 ( .A(n6681), .ZN(n4605) );
  NOR2_X1 U5390 ( .A1(n4483), .A2(n4605), .ZN(n4453) );
  OR2_X1 U5391 ( .A1(n4716), .A2(n4418), .ZN(n4419) );
  NAND2_X1 U5392 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4426) );
  NAND2_X1 U5393 ( .A1(n6262), .A2(n6296), .ZN(n6297) );
  INV_X1 U5394 ( .A(n6297), .ZN(n4425) );
  NAND3_X1 U5395 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4432) );
  INV_X1 U5396 ( .A(n4432), .ZN(n4424) );
  INV_X1 U5397 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6722) );
  NAND2_X1 U5398 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n4431) );
  INV_X1 U5399 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6709) );
  INV_X1 U5400 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6702) );
  INV_X1 U5401 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6701) );
  INV_X1 U5402 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6698) );
  INV_X1 U5403 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6775) );
  INV_X1 U5404 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6695) );
  INV_X1 U5405 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6693) );
  NOR3_X1 U5406 ( .A1(n6775), .A2(n6695), .A3(n6693), .ZN(n6306) );
  NAND2_X1 U5407 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6306), .ZN(n6261) );
  NOR2_X1 U5408 ( .A1(n6698), .A2(n6261), .ZN(n6260) );
  NAND3_X1 U5409 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .A3(
        n6260), .ZN(n5234) );
  NOR2_X1 U5410 ( .A1(n6701), .A2(n5234), .ZN(n5150) );
  NAND3_X1 U5411 ( .A1(n5150), .A2(REIP_REG_9__SCAN_IN), .A3(
        REIP_REG_10__SCAN_IN), .ZN(n6236) );
  NOR2_X1 U5412 ( .A1(n6702), .A2(n6236), .ZN(n6222) );
  NAND4_X1 U5413 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6222), .A3(
        REIP_REG_13__SCAN_IN), .A4(REIP_REG_12__SCAN_IN), .ZN(n5341) );
  NOR2_X1 U5414 ( .A1(n6709), .A2(n5341), .ZN(n4429) );
  NAND3_X1 U5415 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        n4429), .ZN(n4420) );
  NAND2_X1 U5416 ( .A1(n6307), .A2(n4420), .ZN(n4421) );
  NAND2_X1 U5417 ( .A1(n4421), .A2(n6296), .ZN(n6197) );
  NAND2_X1 U5418 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n4430) );
  INV_X1 U5419 ( .A(n4430), .ZN(n4422) );
  AOI21_X1 U5420 ( .B1(REIP_REG_20__SCAN_IN), .B2(n4422), .A(n6262), .ZN(n4423) );
  AOI221_X1 U5421 ( .B1(n6722), .B2(n6297), .C1(n4431), .C2(n6297), .A(n6085), 
        .ZN(n6045) );
  OAI21_X1 U5422 ( .B1(n4425), .B2(n4424), .A(n6045), .ZN(n6036) );
  AOI21_X1 U5423 ( .B1(n6307), .B2(n4426), .A(n6036), .ZN(n6011) );
  INV_X1 U5424 ( .A(REIP_REG_29__SCAN_IN), .ZN(n7134) );
  OAI22_X1 U5425 ( .A1(n6011), .A2(n7134), .B1(n4266), .B2(n6314), .ZN(n4427)
         );
  AOI211_X1 U5426 ( .C1(n6325), .C2(EBX_REG_29__SCAN_IN), .A(n4428), .B(n4427), 
        .ZN(n4433) );
  INV_X1 U5427 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6712) );
  NAND2_X1 U5428 ( .A1(n6307), .A2(n4429), .ZN(n6206) );
  NOR2_X1 U5429 ( .A1(n6712), .A2(n6206), .ZN(n6198) );
  NAND2_X1 U5430 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6198), .ZN(n6093) );
  NOR2_X1 U5431 ( .A1(n6093), .A2(n4430), .ZN(n6084) );
  NAND2_X1 U5432 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6084), .ZN(n6060) );
  NOR2_X1 U5433 ( .A1(n6060), .A2(n4431), .ZN(n6056) );
  NAND2_X1 U5434 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6056), .ZN(n5521) );
  NOR2_X1 U5435 ( .A1(n5521), .A2(n4432), .ZN(n6024) );
  NAND3_X1 U5436 ( .A1(n6024), .A2(REIP_REG_28__SCAN_IN), .A3(
        REIP_REG_27__SCAN_IN), .ZN(n5508) );
  NOR3_X1 U5437 ( .A1(n4438), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n4439), 
        .ZN(n4440) );
  AOI21_X1 U5438 ( .B1(n4441), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n4440), 
        .ZN(n4443) );
  XNOR2_X1 U5439 ( .A(n4443), .B(n4442), .ZN(n5459) );
  NOR2_X1 U5440 ( .A1(n6630), .A2(n4727), .ZN(n4480) );
  INV_X1 U5441 ( .A(n4480), .ZN(n4450) );
  NAND2_X1 U5442 ( .A1(n4483), .A2(n6681), .ZN(n4444) );
  NOR2_X1 U5443 ( .A1(READY_N), .A2(n4512), .ZN(n4611) );
  NAND3_X1 U5444 ( .A1(n4444), .A2(n4611), .A3(n4469), .ZN(n4449) );
  NAND2_X1 U5445 ( .A1(n4446), .A2(n4445), .ZN(n4473) );
  NAND2_X1 U5446 ( .A1(n4457), .A2(n4473), .ZN(n4448) );
  INV_X1 U5447 ( .A(n4513), .ZN(n4447) );
  NAND2_X1 U5448 ( .A1(n4448), .A2(n4447), .ZN(n4614) );
  OAI211_X1 U5449 ( .C1(n4648), .C2(n4450), .A(n4449), .B(n4614), .ZN(n4451)
         );
  NAND2_X1 U5450 ( .A1(n4451), .A2(n6664), .ZN(n4456) );
  NAND2_X1 U5451 ( .A1(n4606), .A2(n6683), .ZN(n4527) );
  INV_X1 U5452 ( .A(n4452), .ZN(n5369) );
  OAI211_X1 U5453 ( .C1(n4527), .C2(n4453), .A(n4318), .B(n5369), .ZN(n4454)
         );
  NAND3_X1 U5454 ( .A1(n4556), .A2(n4742), .A3(n4454), .ZN(n4455) );
  INV_X1 U5455 ( .A(n4515), .ZN(n6647) );
  INV_X1 U5456 ( .A(n4604), .ZN(n4587) );
  INV_X1 U5457 ( .A(n4458), .ZN(n4459) );
  AOI22_X1 U5458 ( .A1(n4459), .A2(n3409), .B1(n4606), .B2(n4573), .ZN(n4460)
         );
  NAND4_X1 U5459 ( .A1(n6647), .A2(n4587), .A3(n4460), .A4(n4636), .ZN(n4461)
         );
  NAND2_X1 U5460 ( .A1(n4562), .A2(EBX_REG_30__SCAN_IN), .ZN(n4463) );
  NAND2_X1 U5461 ( .A1(n4349), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4462) );
  AND2_X1 U5462 ( .A1(n4463), .A2(n4462), .ZN(n5462) );
  NOR2_X1 U5463 ( .A1(n5461), .A2(n5395), .ZN(n5466) );
  AOI21_X1 U5464 ( .B1(n5462), .B2(n4464), .A(n5466), .ZN(n4466) );
  OAI22_X1 U5465 ( .A1(INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n4562), .B1(n4349), .B2(EBX_REG_31__SCAN_IN), .ZN(n4465) );
  XNOR2_X1 U5466 ( .A(n4466), .B(n4465), .ZN(n5529) );
  NAND2_X1 U5467 ( .A1(n4606), .A2(n6782), .ZN(n4533) );
  OAI21_X1 U5468 ( .B1(n4458), .B2(n3409), .A(n4533), .ZN(n4467) );
  NAND2_X1 U5469 ( .A1(n4716), .A2(n4483), .ZN(n5218) );
  NOR2_X1 U5470 ( .A1(n5218), .A2(n4469), .ZN(n4612) );
  OAI21_X1 U5471 ( .B1(n4612), .B2(n4562), .A(n3622), .ZN(n4472) );
  NAND2_X1 U5472 ( .A1(n4468), .A2(n5395), .ZN(n4471) );
  NAND2_X1 U5473 ( .A1(n5369), .A2(n4469), .ZN(n4470) );
  NAND2_X1 U5474 ( .A1(n4475), .A2(n4474), .ZN(n4586) );
  NAND2_X1 U5475 ( .A1(n3454), .A2(n4476), .ZN(n4477) );
  NAND2_X1 U5476 ( .A1(n4477), .A2(n4625), .ZN(n4478) );
  INV_X1 U5477 ( .A(n4481), .ZN(n4479) );
  INV_X1 U5478 ( .A(n4495), .ZN(n4482) );
  NAND2_X1 U5479 ( .A1(n4481), .A2(n4480), .ZN(n4603) );
  INV_X1 U5480 ( .A(n4603), .ZN(n4511) );
  AND2_X1 U5481 ( .A1(n4513), .A2(n4483), .ZN(n6632) );
  NAND2_X1 U5482 ( .A1(n4486), .A2(n6632), .ZN(n6499) );
  AND2_X1 U5483 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5732) );
  INV_X1 U5484 ( .A(n6499), .ZN(n5796) );
  NOR2_X1 U5485 ( .A1(n4495), .A2(n5796), .ZN(n4671) );
  NAND2_X1 U5486 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6486) );
  NAND2_X1 U5487 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4672) );
  NOR2_X1 U5488 ( .A1(n6486), .A2(n4672), .ZN(n4711) );
  NAND3_X1 U5489 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n4711), .ZN(n5093) );
  NOR2_X1 U5490 ( .A1(n6470), .A2(n5095), .ZN(n5167) );
  NAND3_X1 U5491 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n5167), .ZN(n4484) );
  NOR2_X1 U5492 ( .A1(n5093), .A2(n4484), .ZN(n4500) );
  INV_X1 U5493 ( .A(n4484), .ZN(n4485) );
  AOI21_X1 U5494 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n4670) );
  NOR2_X1 U5495 ( .A1(n4670), .A2(n4672), .ZN(n4704) );
  NAND2_X1 U5496 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4704), .ZN(n4705)
         );
  NOR2_X1 U5497 ( .A1(n5086), .A2(n4705), .ZN(n5090) );
  NAND2_X1 U5498 ( .A1(n4485), .A2(n5090), .ZN(n4499) );
  NOR2_X1 U5499 ( .A1(n4486), .A2(n6425), .ZN(n4567) );
  NOR2_X1 U5500 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5799), .ZN(n4566)
         );
  NOR2_X1 U5501 ( .A1(n4567), .A2(n4566), .ZN(n6511) );
  NOR2_X1 U5502 ( .A1(n6488), .A2(n6511), .ZN(n5092) );
  AOI21_X1 U5503 ( .B1(n6488), .B2(n4499), .A(n5092), .ZN(n4487) );
  OAI21_X1 U5504 ( .B1(n4671), .B2(n4500), .A(n4487), .ZN(n5795) );
  NOR2_X1 U5505 ( .A1(n7122), .A2(n4352), .ZN(n5798) );
  NAND2_X1 U5506 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5798), .ZN(n5803) );
  NOR2_X1 U5507 ( .A1(n4488), .A2(n5803), .ZN(n5784) );
  NAND3_X1 U5508 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5784), .ZN(n4501) );
  AND2_X1 U5509 ( .A1(n6501), .A2(n4501), .ZN(n4489) );
  NOR2_X1 U5510 ( .A1(n5795), .A2(n4489), .ZN(n6146) );
  INV_X1 U5511 ( .A(n4490), .ZN(n4492) );
  INV_X1 U5512 ( .A(n6134), .ZN(n4491) );
  NAND2_X1 U5513 ( .A1(n4492), .A2(n4491), .ZN(n5440) );
  NAND2_X1 U5514 ( .A1(n6501), .A2(n5440), .ZN(n4493) );
  NAND2_X1 U5515 ( .A1(n6146), .A2(n4493), .ZN(n5761) );
  AND2_X1 U5516 ( .A1(n6501), .A2(n5750), .ZN(n4494) );
  NAND2_X1 U5517 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n4495), .ZN(n5794)
         );
  NAND2_X1 U5518 ( .A1(n6499), .A2(n5794), .ZN(n4709) );
  INV_X1 U5519 ( .A(n4709), .ZN(n6490) );
  AOI21_X1 U5520 ( .B1(n6490), .B2(n5089), .A(n4496), .ZN(n4497) );
  OAI21_X1 U5521 ( .B1(n5781), .B2(n5732), .A(n6131), .ZN(n5729) );
  AND3_X1 U5522 ( .A1(n5472), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4502) );
  NOR2_X1 U5523 ( .A1(n5781), .A2(n4502), .ZN(n4498) );
  OAI21_X1 U5524 ( .B1(n5729), .B2(n4498), .A(INSTADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n4505) );
  AND2_X1 U5525 ( .A1(n6425), .A2(REIP_REG_31__SCAN_IN), .ZN(n5454) );
  INV_X1 U5526 ( .A(n5454), .ZN(n4504) );
  NOR2_X1 U5527 ( .A1(n5089), .A2(n4499), .ZN(n5791) );
  NAND3_X1 U5528 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n6141), .ZN(n6132) );
  NOR2_X1 U5529 ( .A1(n3258), .A2(n6132), .ZN(n6124) );
  NAND2_X1 U5530 ( .A1(n6124), .A2(n5732), .ZN(n5716) );
  INV_X1 U5531 ( .A(n4502), .ZN(n4503) );
  NAND3_X1 U5532 ( .A1(n4505), .A2(n4504), .A3(n3327), .ZN(n4506) );
  AOI21_X1 U5533 ( .B1(n5529), .B2(n6503), .A(n4506), .ZN(n4507) );
  OAI21_X1 U5534 ( .B1(n5459), .B2(n6475), .A(n4507), .ZN(U2987) );
  OAI22_X1 U5535 ( .A1(n4648), .A2(n4509), .B1(n4514), .B2(n4508), .ZN(n6167)
         );
  NAND2_X1 U5536 ( .A1(n4510), .A2(n5218), .ZN(n4525) );
  AOI21_X1 U5537 ( .B1(n4525), .B2(n6681), .A(READY_N), .ZN(n6785) );
  NOR2_X1 U5538 ( .A1(n6167), .A2(n6785), .ZN(n6646) );
  INV_X1 U5539 ( .A(n6664), .ZN(n6662) );
  NOR2_X1 U5540 ( .A1(n6646), .A2(n6662), .ZN(n6174) );
  INV_X1 U5541 ( .A(MORE_REG_SCAN_IN), .ZN(n4523) );
  NAND2_X1 U5542 ( .A1(n4511), .A2(n4648), .ZN(n4520) );
  NAND2_X1 U5543 ( .A1(n4513), .A2(n4512), .ZN(n4519) );
  OR2_X1 U5544 ( .A1(n4515), .A2(n4514), .ZN(n4516) );
  NOR2_X1 U5545 ( .A1(n4516), .A2(n4604), .ZN(n4517) );
  OR2_X1 U5546 ( .A1(n4648), .A2(n4517), .ZN(n4518) );
  AND3_X1 U5547 ( .A1(n4520), .A2(n4519), .A3(n4518), .ZN(n6648) );
  INV_X1 U5548 ( .A(n6648), .ZN(n4521) );
  NAND2_X1 U5549 ( .A1(n6174), .A2(n4521), .ZN(n4522) );
  OAI21_X1 U5550 ( .B1(n6174), .B2(n4523), .A(n4522), .ZN(U3471) );
  OAI21_X1 U5551 ( .B1(n5502), .B2(READREQUEST_REG_SCAN_IN), .A(n6777), .ZN(
        n4524) );
  OAI21_X1 U5552 ( .B1(n6777), .B2(n4525), .A(n4524), .ZN(U3474) );
  INV_X1 U5553 ( .A(n5505), .ZN(n4526) );
  INV_X1 U5554 ( .A(LWORD_REG_3__SCAN_IN), .ZN(n6815) );
  INV_X1 U5555 ( .A(n4533), .ZN(n6655) );
  INV_X1 U5556 ( .A(n6794), .ZN(n6419) );
  NOR2_X1 U5557 ( .A1(n4527), .A2(n4349), .ZN(n4607) );
  AND2_X1 U5558 ( .A1(n6422), .A2(DATAI_3_), .ZN(n6366) );
  AOI21_X1 U5559 ( .B1(n6419), .B2(EAX_REG_3__SCAN_IN), .A(n6366), .ZN(n4528)
         );
  OAI21_X1 U5560 ( .B1(n6363), .B2(n6815), .A(n4528), .ZN(U2942) );
  INV_X1 U5561 ( .A(UWORD_REG_2__SCAN_IN), .ZN(n7137) );
  AND2_X1 U5562 ( .A1(n6422), .A2(DATAI_2_), .ZN(n6395) );
  AOI21_X1 U5563 ( .B1(n6419), .B2(EAX_REG_18__SCAN_IN), .A(n6395), .ZN(n4529)
         );
  OAI21_X1 U5564 ( .B1(n6363), .B2(n7137), .A(n4529), .ZN(U2926) );
  INV_X1 U5565 ( .A(LWORD_REG_12__SCAN_IN), .ZN(n6344) );
  INV_X1 U5566 ( .A(DATAI_12_), .ZN(n5303) );
  NOR2_X1 U5567 ( .A1(n6421), .A2(n5303), .ZN(n4531) );
  AOI21_X1 U5568 ( .B1(n6419), .B2(EAX_REG_12__SCAN_IN), .A(n4531), .ZN(n4530)
         );
  OAI21_X1 U5569 ( .B1(n6363), .B2(n6344), .A(n4530), .ZN(U2951) );
  INV_X1 U5570 ( .A(UWORD_REG_12__SCAN_IN), .ZN(n7050) );
  AOI21_X1 U5571 ( .B1(n6419), .B2(EAX_REG_28__SCAN_IN), .A(n4531), .ZN(n4532)
         );
  OAI21_X1 U5572 ( .B1(n6363), .B2(n7050), .A(n4532), .ZN(U2936) );
  INV_X1 U5573 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6375) );
  INV_X1 U5574 ( .A(n6632), .ZN(n4534) );
  AOI21_X1 U5575 ( .B1(n4534), .B2(n4533), .A(n6681), .ZN(n4535) );
  NAND2_X1 U5576 ( .A1(n6349), .A2(n4318), .ZN(n6336) );
  NAND2_X1 U5577 ( .A1(n6783), .A2(n6669), .ZN(n6779) );
  INV_X2 U5578 ( .A(n6779), .ZN(n6348) );
  AOI22_X1 U5579 ( .A1(n6348), .A2(UWORD_REG_7__SCAN_IN), .B1(n6358), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4537) );
  OAI21_X1 U5580 ( .B1(n6375), .B2(n6336), .A(n4537), .ZN(U2900) );
  INV_X1 U5581 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6365) );
  AOI22_X1 U5582 ( .A1(n6348), .A2(UWORD_REG_1__SCAN_IN), .B1(n6358), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4538) );
  OAI21_X1 U5583 ( .B1(n6365), .B2(n6336), .A(n4538), .ZN(U2906) );
  INV_X1 U5584 ( .A(EAX_REG_19__SCAN_IN), .ZN(n6368) );
  AOI22_X1 U5585 ( .A1(n6348), .A2(UWORD_REG_3__SCAN_IN), .B1(n6358), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4539) );
  OAI21_X1 U5586 ( .B1(n6368), .B2(n6336), .A(n4539), .ZN(U2904) );
  INV_X1 U5587 ( .A(EAX_REG_20__SCAN_IN), .ZN(n6370) );
  AOI22_X1 U5588 ( .A1(n6348), .A2(UWORD_REG_4__SCAN_IN), .B1(n6358), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4540) );
  OAI21_X1 U5589 ( .B1(n6370), .B2(n6336), .A(n4540), .ZN(U2903) );
  INV_X1 U5590 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6372) );
  AOI22_X1 U5591 ( .A1(n6348), .A2(UWORD_REG_5__SCAN_IN), .B1(n6358), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4541) );
  OAI21_X1 U5592 ( .B1(n6372), .B2(n6336), .A(n4541), .ZN(U2902) );
  INV_X1 U5593 ( .A(EAX_REG_22__SCAN_IN), .ZN(n7095) );
  AOI22_X1 U5594 ( .A1(n6348), .A2(UWORD_REG_6__SCAN_IN), .B1(n6358), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4542) );
  OAI21_X1 U5595 ( .B1(n7095), .B2(n6336), .A(n4542), .ZN(U2901) );
  INV_X1 U5596 ( .A(EAX_REG_16__SCAN_IN), .ZN(n6362) );
  AOI22_X1 U5597 ( .A1(n6348), .A2(UWORD_REG_0__SCAN_IN), .B1(n6358), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4543) );
  OAI21_X1 U5598 ( .B1(n6362), .B2(n6336), .A(n4543), .ZN(U2907) );
  INV_X1 U5599 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6388) );
  AOI22_X1 U5600 ( .A1(n6348), .A2(UWORD_REG_14__SCAN_IN), .B1(n6358), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4544) );
  OAI21_X1 U5601 ( .B1(n6388), .B2(n6336), .A(n4544), .ZN(U2893) );
  INV_X1 U5602 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6386) );
  AOI22_X1 U5603 ( .A1(n6348), .A2(UWORD_REG_13__SCAN_IN), .B1(n6358), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4545) );
  OAI21_X1 U5604 ( .B1(n6386), .B2(n6336), .A(n4545), .ZN(U2894) );
  INV_X1 U5605 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6379) );
  AOI22_X1 U5606 ( .A1(n6348), .A2(UWORD_REG_9__SCAN_IN), .B1(n6358), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4546) );
  OAI21_X1 U5607 ( .B1(n6379), .B2(n6336), .A(n4546), .ZN(U2898) );
  INV_X1 U5608 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6382) );
  AOI22_X1 U5609 ( .A1(n6348), .A2(UWORD_REG_10__SCAN_IN), .B1(n6358), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4547) );
  OAI21_X1 U5610 ( .B1(n6382), .B2(n6336), .A(n4547), .ZN(U2897) );
  INV_X1 U5611 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6384) );
  AOI22_X1 U5612 ( .A1(n6348), .A2(UWORD_REG_11__SCAN_IN), .B1(
        DATAO_REG_27__SCAN_IN), .B2(n6358), .ZN(n4548) );
  OAI21_X1 U5613 ( .B1(n6384), .B2(n6336), .A(n4548), .ZN(U2896) );
  OR2_X1 U5614 ( .A1(n4550), .A2(n4549), .ZN(n4551) );
  NAND2_X1 U5615 ( .A1(n4552), .A2(n4551), .ZN(n6445) );
  NAND2_X1 U5616 ( .A1(n6664), .A2(n4611), .ZN(n4554) );
  INV_X1 U5617 ( .A(n4553), .ZN(n4584) );
  INV_X1 U5618 ( .A(n4576), .ZN(n5594) );
  NAND4_X1 U5619 ( .A1(n5594), .A2(n4688), .A3(n6664), .A4(n3460), .ZN(n4570)
         );
  OAI22_X1 U5620 ( .A1(n4636), .A2(n4554), .B1(n4584), .B2(n4570), .ZN(n4555)
         );
  NAND2_X1 U5621 ( .A1(n3467), .A2(n4576), .ZN(n4558) );
  NAND2_X2 U5622 ( .A1(n5593), .A2(n4558), .ZN(n5339) );
  INV_X1 U5623 ( .A(n4558), .ZN(n4559) );
  INV_X1 U5624 ( .A(DATAI_0_), .ZN(n4717) );
  INV_X1 U5625 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6391) );
  OAI222_X1 U5626 ( .A1(n6445), .A2(n5339), .B1(n5338), .B2(n4717), .C1(n5593), 
        .C2(n6391), .ZN(U2891) );
  OAI21_X1 U5627 ( .B1(n4561), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4560), 
        .ZN(n6439) );
  NOR2_X1 U5628 ( .A1(n4562), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4564)
         );
  NOR2_X1 U5629 ( .A1(n4564), .A2(n4563), .ZN(n5219) );
  INV_X1 U5630 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6769) );
  NOR2_X1 U5631 ( .A1(n6498), .A2(n6769), .ZN(n4565) );
  AOI211_X1 U5632 ( .C1(n6503), .C2(n5219), .A(n4566), .B(n4565), .ZN(n4569)
         );
  OAI21_X1 U5633 ( .B1(n4567), .B2(n5796), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4568) );
  OAI211_X1 U5634 ( .C1(n6439), .C2(n6475), .A(n4569), .B(n4568), .ZN(U3018)
         );
  INV_X1 U5635 ( .A(n5219), .ZN(n4577) );
  OR3_X1 U5636 ( .A1(n4603), .A2(n4648), .A3(n6662), .ZN(n4575) );
  INV_X1 U5637 ( .A(n4570), .ZN(n4571) );
  NAND3_X1 U5638 ( .A1(n4573), .A2(n4572), .A3(n4571), .ZN(n4574) );
  NAND2_X2 U5639 ( .A1(n5591), .A2(n4576), .ZN(n5575) );
  OAI222_X1 U5640 ( .A1(n4577), .A2(n5592), .B1(n5591), .B2(n5222), .C1(n5575), 
        .C2(n6445), .ZN(U2859) );
  OAI21_X1 U5641 ( .B1(n4580), .B2(n4579), .A(n4578), .ZN(n5320) );
  INV_X1 U5642 ( .A(DATAI_1_), .ZN(n7055) );
  INV_X1 U5643 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6394) );
  OAI222_X1 U5644 ( .A1(n5320), .A2(n5339), .B1(n5338), .B2(n7055), .C1(n5593), 
        .C2(n6394), .ZN(U2890) );
  INV_X1 U5645 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6173) );
  NAND2_X1 U5646 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6173), .ZN(n4643) );
  INV_X1 U5647 ( .A(n4581), .ZN(n4642) );
  NAND4_X1 U5648 ( .A1(n4636), .A2(n3308), .A3(n4584), .A4(n4583), .ZN(n4585)
         );
  NOR2_X1 U5649 ( .A1(n4586), .A2(n4585), .ZN(n6631) );
  INV_X1 U5650 ( .A(n6631), .ZN(n4602) );
  NAND2_X1 U5651 ( .A1(n4603), .A2(n4587), .ZN(n4628) );
  MUX2_X1 U5652 ( .A(n4589), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4588), 
        .Z(n4590) );
  NOR2_X1 U5653 ( .A1(n4590), .A2(n4581), .ZN(n4591) );
  NAND2_X1 U5654 ( .A1(n4628), .A2(n4591), .ZN(n4600) );
  XNOR2_X1 U5655 ( .A(n4592), .B(n4621), .ZN(n4598) );
  INV_X1 U5656 ( .A(n4593), .ZN(n4594) );
  OAI21_X1 U5657 ( .B1(n4588), .B2(n4621), .A(n4594), .ZN(n4596) );
  NOR2_X1 U5658 ( .A1(n4596), .A2(n4595), .ZN(n5809) );
  NOR2_X1 U5659 ( .A1(n4625), .A2(n5809), .ZN(n4597) );
  AOI21_X1 U5660 ( .B1(n6632), .B2(n4598), .A(n4597), .ZN(n4599) );
  NAND2_X1 U5661 ( .A1(n4600), .A2(n4599), .ZN(n4601) );
  AOI21_X1 U5662 ( .B1(n4582), .B2(n4602), .A(n4601), .ZN(n5810) );
  OR2_X1 U5663 ( .A1(n4603), .A2(n4648), .ZN(n4620) );
  NAND2_X1 U5664 ( .A1(n4648), .A2(n4604), .ZN(n4619) );
  OAI211_X1 U5665 ( .C1(n6632), .C2(n4606), .A(n4605), .B(n6683), .ZN(n4609)
         );
  INV_X1 U5666 ( .A(n4607), .ZN(n4608) );
  NAND2_X1 U5667 ( .A1(n4609), .A2(n4608), .ZN(n4610) );
  NAND2_X1 U5668 ( .A1(n4648), .A2(n4610), .ZN(n4618) );
  INV_X1 U5669 ( .A(n4611), .ZN(n4615) );
  INV_X1 U5670 ( .A(n4612), .ZN(n4613) );
  OAI211_X1 U5671 ( .C1(n4615), .C2(n4636), .A(n4614), .B(n4613), .ZN(n4616)
         );
  INV_X1 U5672 ( .A(n4616), .ZN(n4617) );
  NAND4_X1 U5673 ( .A1(n4620), .A2(n4619), .A3(n4618), .A4(n4617), .ZN(n6635)
         );
  MUX2_X1 U5674 ( .A(n4621), .B(n5810), .S(n6635), .Z(n6644) );
  INV_X1 U5675 ( .A(n6644), .ZN(n4633) );
  OR2_X1 U5676 ( .A1(n4622), .A2(n6631), .ZN(n4630) );
  XNOR2_X1 U5677 ( .A(n4588), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4627)
         );
  XNOR2_X1 U5678 ( .A(n3207), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4623)
         );
  NAND2_X1 U5679 ( .A1(n6632), .A2(n4623), .ZN(n4624) );
  OAI21_X1 U5680 ( .B1(n4627), .B2(n4625), .A(n4624), .ZN(n4626) );
  AOI21_X1 U5681 ( .B1(n4628), .B2(n4627), .A(n4626), .ZN(n4629) );
  AND2_X1 U5682 ( .A1(n4630), .A2(n4629), .ZN(n5477) );
  NAND2_X1 U5683 ( .A1(n5477), .A2(n6635), .ZN(n4632) );
  NAND2_X1 U5684 ( .A1(n5476), .A2(n3332), .ZN(n4631) );
  NAND3_X1 U5685 ( .A1(n4633), .A2(n6642), .A3(n6749), .ZN(n4641) );
  INV_X1 U5686 ( .A(n6513), .ZN(n4634) );
  OR2_X1 U5687 ( .A1(n3573), .A2(n4634), .ZN(n4635) );
  XNOR2_X1 U5688 ( .A(n4635), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6294)
         );
  INV_X1 U5689 ( .A(n4636), .ZN(n6162) );
  NAND2_X1 U5690 ( .A1(n6294), .A2(n6162), .ZN(n4638) );
  NAND2_X1 U5691 ( .A1(n5476), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4637) );
  NAND2_X1 U5692 ( .A1(n4638), .A2(n4637), .ZN(n4640) );
  NOR2_X1 U5693 ( .A1(n6165), .A2(n4643), .ZN(n4639) );
  AOI21_X1 U5694 ( .B1(n4640), .B2(n6749), .A(n4639), .ZN(n4645) );
  OAI211_X1 U5695 ( .C1(n4643), .C2(n4642), .A(n4641), .B(n4645), .ZN(n6651)
         );
  NAND2_X1 U5696 ( .A1(n4645), .A2(n3223), .ZN(n4646) );
  NAND2_X1 U5697 ( .A1(n6651), .A2(n4646), .ZN(n6660) );
  NAND2_X1 U5698 ( .A1(n6660), .A2(n6173), .ZN(n4647) );
  NAND2_X1 U5699 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6669), .ZN(n6673) );
  INV_X1 U5700 ( .A(n6673), .ZN(n6744) );
  NAND2_X1 U5701 ( .A1(n4647), .A2(n6744), .ZN(n4649) );
  NAND2_X1 U5702 ( .A1(n4649), .A2(n4782), .ZN(n6763) );
  INV_X1 U5703 ( .A(n5863), .ZN(n4651) );
  AOI21_X1 U5704 ( .B1(n4651), .B2(n6781), .A(n6571), .ZN(n4653) );
  NAND2_X1 U5705 ( .A1(n5863), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6565) );
  OR2_X1 U5706 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6749), .ZN(n6762) );
  AOI22_X1 U5707 ( .A1(n4653), .A2(n6565), .B1(n5317), .B2(n6762), .ZN(n4655)
         );
  NAND2_X1 U5708 ( .A1(n6766), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4654) );
  OAI21_X1 U5709 ( .B1(n6766), .B2(n4655), .A(n4654), .ZN(U3464) );
  XNOR2_X1 U5710 ( .A(n4816), .B(n6565), .ZN(n4658) );
  INV_X1 U5711 ( .A(n4622), .ZN(n4657) );
  AOI22_X1 U5712 ( .A1(n4658), .A2(n6564), .B1(n4657), .B2(n6762), .ZN(n4660)
         );
  NAND2_X1 U5713 ( .A1(n6766), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4659) );
  OAI21_X1 U5714 ( .B1(n6766), .B2(n4660), .A(n4659), .ZN(U3463) );
  INV_X1 U5715 ( .A(n3230), .ZN(n5853) );
  AOI222_X1 U5716 ( .A1(n6660), .A2(n6669), .B1(n4751), .B2(n6564), .C1(n5853), 
        .C2(n6762), .ZN(n4662) );
  NAND2_X1 U5717 ( .A1(n6766), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4661) );
  OAI21_X1 U5718 ( .B1(n6766), .B2(n4662), .A(n4661), .ZN(U3465) );
  NOR2_X1 U5719 ( .A1(n4665), .A2(n4664), .ZN(n4666) );
  NOR2_X1 U5720 ( .A1(n4663), .A2(n4666), .ZN(n6433) );
  INV_X1 U5721 ( .A(n6433), .ZN(n4684) );
  INV_X1 U5722 ( .A(DATAI_2_), .ZN(n4667) );
  INV_X1 U5723 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6397) );
  OAI222_X1 U5724 ( .A1(n4684), .A2(n5339), .B1(n5338), .B2(n4667), .C1(n5593), 
        .C2(n6397), .ZN(U2889) );
  XNOR2_X1 U5725 ( .A(n4668), .B(n4669), .ZN(n5080) );
  INV_X1 U5726 ( .A(n4670), .ZN(n6485) );
  INV_X1 U5727 ( .A(n4671), .ZN(n5094) );
  AOI21_X1 U5728 ( .B1(n5094), .B2(n6486), .A(n5092), .ZN(n6491) );
  OAI21_X1 U5729 ( .B1(n5089), .B2(n6485), .A(n6491), .ZN(n6472) );
  OAI21_X1 U5730 ( .B1(n6490), .B2(n6486), .A(n5089), .ZN(n4806) );
  NAND2_X1 U5731 ( .A1(n4806), .A2(n6485), .ZN(n6479) );
  OAI21_X1 U5732 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4672), .ZN(n4675) );
  OAI21_X1 U5733 ( .B1(n4673), .B2(n3257), .A(n4707), .ZN(n4890) );
  INV_X1 U5734 ( .A(n4890), .ZN(n6295) );
  AND2_X1 U5735 ( .A1(n6425), .A2(REIP_REG_4__SCAN_IN), .ZN(n5075) );
  AOI21_X1 U5736 ( .B1(n6503), .B2(n6295), .A(n5075), .ZN(n4674) );
  OAI21_X1 U5737 ( .B1(n6479), .B2(n4675), .A(n4674), .ZN(n4676) );
  AOI21_X1 U5738 ( .B1(n6472), .B2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4676), 
        .ZN(n4677) );
  OAI21_X1 U5739 ( .B1(n6475), .B2(n5080), .A(n4677), .ZN(U3014) );
  OAI21_X1 U5740 ( .B1(n4663), .B2(n4678), .A(n4778), .ZN(n6322) );
  INV_X1 U5741 ( .A(DATAI_3_), .ZN(n4723) );
  INV_X1 U5742 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6355) );
  OAI222_X1 U5743 ( .A1(n6322), .A2(n5339), .B1(n5338), .B2(n4723), .C1(n5593), 
        .C2(n6355), .ZN(U2888) );
  AOI21_X1 U5744 ( .B1(n4680), .B2(n4679), .A(n3257), .ZN(n6474) );
  AOI22_X1 U5745 ( .A1(n5557), .A2(n6474), .B1(n5556), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4681) );
  OAI21_X1 U5746 ( .B1(n6322), .B2(n5575), .A(n4681), .ZN(U2856) );
  XNOR2_X1 U5747 ( .A(n4683), .B(n4682), .ZN(n6484) );
  INV_X1 U5748 ( .A(EBX_REG_2__SCAN_IN), .ZN(n5324) );
  OAI222_X1 U5749 ( .A1(n4684), .A2(n5575), .B1(n5592), .B2(n6484), .C1(n5591), 
        .C2(n5324), .ZN(U2857) );
  XNOR2_X1 U5750 ( .A(n5313), .B(n4349), .ZN(n6502) );
  INV_X1 U5751 ( .A(n6502), .ZN(n4685) );
  INV_X1 U5752 ( .A(EBX_REG_1__SCAN_IN), .ZN(n6998) );
  OAI222_X1 U5753 ( .A1(n4685), .A2(n5592), .B1(n5591), .B2(n6998), .C1(n5575), 
        .C2(n5320), .ZN(U2858) );
  INV_X1 U5754 ( .A(DATAI_28_), .ZN(n7020) );
  NOR2_X1 U5755 ( .A1(n5714), .A2(n7020), .ZN(n6600) );
  INV_X1 U5756 ( .A(n6600), .ZN(n5882) );
  INV_X2 U5757 ( .A(n5714), .ZN(n6432) );
  NAND2_X1 U5758 ( .A1(n6432), .A2(DATAI_20_), .ZN(n6604) );
  INV_X1 U5759 ( .A(n6604), .ZN(n6540) );
  NOR2_X1 U5760 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n7152), .ZN(n6745) );
  NOR2_X1 U5761 ( .A1(n4743), .A2(n4688), .ZN(n6599) );
  INV_X1 U5762 ( .A(n6599), .ZN(n5988) );
  INV_X1 U5763 ( .A(n5317), .ZN(n5494) );
  OR2_X1 U5764 ( .A1(n5494), .A2(n4622), .ZN(n6514) );
  INV_X1 U5765 ( .A(n6514), .ZN(n5906) );
  NAND2_X1 U5766 ( .A1(n4983), .A2(n5906), .ZN(n4689) );
  NAND2_X1 U5767 ( .A1(n4689), .A2(n4737), .ZN(n4691) );
  AOI22_X1 U5768 ( .A1(n4691), .A2(n6564), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4695), .ZN(n4736) );
  INV_X1 U5769 ( .A(DATAI_4_), .ZN(n7086) );
  NOR2_X2 U5770 ( .A1(n7086), .A2(n4782), .ZN(n6601) );
  INV_X1 U5771 ( .A(n6601), .ZN(n6543) );
  OAI22_X1 U5772 ( .A1(n5988), .A2(n4737), .B1(n4736), .B2(n6543), .ZN(n4690)
         );
  AOI21_X1 U5773 ( .B1(n6540), .B2(n5837), .A(n4690), .ZN(n4697) );
  AOI21_X1 U5774 ( .B1(n4752), .B2(n5863), .A(n5714), .ZN(n4693) );
  NAND2_X1 U5775 ( .A1(n6564), .A2(n6781), .ZN(n4938) );
  INV_X1 U5776 ( .A(n4938), .ZN(n6761) );
  INV_X1 U5777 ( .A(n4691), .ZN(n4692) );
  OAI21_X1 U5778 ( .B1(n4693), .B2(n6761), .A(n4692), .ZN(n4694) );
  INV_X1 U5779 ( .A(n6570), .ZN(n6522) );
  OAI211_X1 U5780 ( .C1(n6564), .C2(n4695), .A(n4694), .B(n6522), .ZN(n4735)
         );
  NAND2_X1 U5781 ( .A1(n4735), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4696)
         );
  OAI211_X1 U5782 ( .C1(n6010), .C2(n5882), .A(n4697), .B(n4696), .ZN(U3144)
         );
  NAND2_X1 U5783 ( .A1(n6432), .A2(DATAI_29_), .ZN(n5887) );
  INV_X1 U5784 ( .A(DATAI_21_), .ZN(n4698) );
  NOR2_X1 U5785 ( .A1(n5714), .A2(n4698), .ZN(n6544) );
  INV_X1 U5786 ( .A(n6605), .ZN(n5992) );
  INV_X1 U5787 ( .A(DATAI_5_), .ZN(n7006) );
  NOR2_X2 U5788 ( .A1(n7006), .A2(n4782), .ZN(n6607) );
  INV_X1 U5789 ( .A(n6607), .ZN(n6547) );
  OAI22_X1 U5790 ( .A1(n5992), .A2(n4737), .B1(n4736), .B2(n6547), .ZN(n4699)
         );
  AOI21_X1 U5791 ( .B1(n6544), .B2(n5837), .A(n4699), .ZN(n4701) );
  NAND2_X1 U5792 ( .A1(n4735), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4700)
         );
  OAI211_X1 U5793 ( .C1(n6010), .C2(n5887), .A(n4701), .B(n4700), .ZN(U3145)
         );
  XNOR2_X1 U5794 ( .A(n4702), .B(n4703), .ZN(n5074) );
  AND2_X1 U5795 ( .A1(n6488), .A2(n4704), .ZN(n4706) );
  INV_X1 U5796 ( .A(n4705), .ZN(n4807) );
  OAI21_X1 U5797 ( .B1(n4807), .B2(n5781), .A(n6491), .ZN(n4813) );
  OAI21_X1 U5798 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4706), .A(n4813), 
        .ZN(n4714) );
  AOI21_X1 U5799 ( .B1(n4708), .B2(n4707), .A(n4808), .ZN(n6283) );
  AND2_X1 U5800 ( .A1(n6425), .A2(REIP_REG_5__SCAN_IN), .ZN(n5070) );
  AND3_X1 U5801 ( .A1(n4711), .A2(n4710), .A3(n4709), .ZN(n4712) );
  AOI211_X1 U5802 ( .C1(n6503), .C2(n6283), .A(n5070), .B(n4712), .ZN(n4713)
         );
  OAI211_X1 U5803 ( .C1(n5074), .C2(n6475), .A(n4714), .B(n4713), .ZN(U3013)
         );
  INV_X1 U5804 ( .A(DATAI_24_), .ZN(n4715) );
  NOR2_X1 U5805 ( .A1(n5714), .A2(n4715), .ZN(n6563) );
  INV_X1 U5806 ( .A(n6563), .ZN(n5865) );
  NAND2_X1 U5807 ( .A1(n6432), .A2(DATAI_16_), .ZN(n6580) );
  INV_X1 U5808 ( .A(n6580), .ZN(n6518) );
  INV_X1 U5809 ( .A(n6562), .ZN(n5969) );
  NOR2_X2 U5810 ( .A1(n4717), .A2(n4782), .ZN(n6577) );
  INV_X1 U5811 ( .A(n6577), .ZN(n6527) );
  OAI22_X1 U5812 ( .A1(n5969), .A2(n4737), .B1(n4736), .B2(n6527), .ZN(n4718)
         );
  AOI21_X1 U5813 ( .B1(n6518), .B2(n5837), .A(n4718), .ZN(n4720) );
  NAND2_X1 U5814 ( .A1(n4735), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4719)
         );
  OAI211_X1 U5815 ( .C1(n6010), .C2(n5865), .A(n4720), .B(n4719), .ZN(U3140)
         );
  NAND2_X1 U5816 ( .A1(n6432), .A2(DATAI_27_), .ZN(n6598) );
  INV_X1 U5817 ( .A(DATAI_19_), .ZN(n4721) );
  INV_X1 U5819 ( .A(n6593), .ZN(n5983) );
  NOR2_X2 U5820 ( .A1(n4723), .A2(n4782), .ZN(n6595) );
  INV_X1 U5821 ( .A(n6595), .ZN(n6539) );
  OAI22_X1 U5822 ( .A1(n5983), .A2(n4737), .B1(n4736), .B2(n6539), .ZN(n4724)
         );
  AOI21_X1 U5823 ( .B1(n6594), .B2(n5837), .A(n4724), .ZN(n4726) );
  NAND2_X1 U5824 ( .A1(n4735), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4725)
         );
  OAI211_X1 U5825 ( .C1(n6010), .C2(n6598), .A(n4726), .B(n4725), .ZN(U3143)
         );
  NAND2_X1 U5826 ( .A1(n6432), .A2(DATAI_25_), .ZN(n6586) );
  NOR2_X1 U5828 ( .A1(n4743), .A2(n4727), .ZN(n6581) );
  INV_X1 U5829 ( .A(n6581), .ZN(n5973) );
  NOR2_X2 U5830 ( .A1(n7055), .A2(n4782), .ZN(n6583) );
  INV_X1 U5831 ( .A(n6583), .ZN(n6531) );
  OAI22_X1 U5832 ( .A1(n5973), .A2(n4737), .B1(n4736), .B2(n6531), .ZN(n4728)
         );
  AOI21_X1 U5833 ( .B1(n6582), .B2(n5837), .A(n4728), .ZN(n4730) );
  NAND2_X1 U5834 ( .A1(n4735), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4729)
         );
  OAI211_X1 U5835 ( .C1(n6010), .C2(n6586), .A(n4730), .B(n4729), .ZN(U3141)
         );
  INV_X1 U5836 ( .A(DATAI_31_), .ZN(n6946) );
  NOR2_X1 U5837 ( .A1(n5714), .A2(n6946), .ZN(n6555) );
  INV_X1 U5838 ( .A(n6555), .ZN(n6629) );
  INV_X1 U5839 ( .A(DATAI_23_), .ZN(n4731) );
  INV_X1 U5841 ( .A(n6620), .ZN(n6005) );
  INV_X1 U5842 ( .A(DATAI_7_), .ZN(n5120) );
  NOR2_X2 U5843 ( .A1(n5120), .A2(n4782), .ZN(n6624) );
  INV_X1 U5844 ( .A(n6624), .ZN(n6559) );
  OAI22_X1 U5845 ( .A1(n6005), .A2(n4737), .B1(n4736), .B2(n6559), .ZN(n4732)
         );
  AOI21_X1 U5846 ( .B1(n6621), .B2(n5837), .A(n4732), .ZN(n4734) );
  NAND2_X1 U5847 ( .A1(n4735), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4733)
         );
  OAI211_X1 U5848 ( .C1(n6010), .C2(n6629), .A(n4734), .B(n4733), .ZN(U3147)
         );
  INV_X1 U5849 ( .A(n4735), .ZN(n4750) );
  INV_X1 U5850 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4741) );
  NAND2_X1 U5851 ( .A1(DATAI_6_), .A2(n4895), .ZN(n6551) );
  INV_X1 U5852 ( .A(n4736), .ZN(n4745) );
  INV_X1 U5853 ( .A(n4737), .ZN(n4744) );
  NOR2_X2 U5854 ( .A1(n4743), .A2(n3461), .ZN(n6611) );
  AOI22_X1 U5855 ( .A1(n6614), .A2(n4745), .B1(n4744), .B2(n6611), .ZN(n4740)
         );
  NAND2_X1 U5856 ( .A1(n6432), .A2(DATAI_30_), .ZN(n5997) );
  INV_X1 U5857 ( .A(n5997), .ZN(n6612) );
  INV_X1 U5858 ( .A(DATAI_22_), .ZN(n4738) );
  NOR2_X1 U5859 ( .A1(n5714), .A2(n4738), .ZN(n6548) );
  AOI22_X1 U5860 ( .A1(n6612), .A2(n5958), .B1(n5837), .B2(n6548), .ZN(n4739)
         );
  OAI211_X1 U5861 ( .C1(n4750), .C2(n4741), .A(n4740), .B(n4739), .ZN(U3146)
         );
  INV_X1 U5862 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4749) );
  NAND2_X1 U5863 ( .A1(DATAI_2_), .A2(n4895), .ZN(n6535) );
  NOR2_X2 U5864 ( .A1(n4743), .A2(n4742), .ZN(n6587) );
  AOI22_X1 U5865 ( .A1(n6589), .A2(n4745), .B1(n4744), .B2(n6587), .ZN(n4748)
         );
  NAND2_X1 U5866 ( .A1(n6432), .A2(DATAI_26_), .ZN(n5979) );
  INV_X1 U5867 ( .A(n5979), .ZN(n6588) );
  INV_X1 U5868 ( .A(DATAI_18_), .ZN(n4746) );
  NOR2_X1 U5869 ( .A1(n5714), .A2(n4746), .ZN(n6532) );
  AOI22_X1 U5870 ( .A1(n6588), .A2(n5958), .B1(n5837), .B2(n6532), .ZN(n4747)
         );
  OAI211_X1 U5871 ( .C1(n4750), .C2(n4749), .A(n4748), .B(n4747), .ZN(U3142)
         );
  NAND3_X1 U5872 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6637), .ZN(n4781) );
  INV_X1 U5873 ( .A(n4781), .ZN(n4754) );
  OR2_X1 U5874 ( .A1(n4622), .A2(n5317), .ZN(n4891) );
  INV_X1 U5875 ( .A(n4891), .ZN(n4786) );
  NOR2_X1 U5876 ( .A1(n6633), .A2(n4781), .ZN(n4774) );
  AOI21_X1 U5877 ( .B1(n4983), .B2(n4786), .A(n4774), .ZN(n4756) );
  OR2_X1 U5878 ( .A1(n5863), .A2(n6781), .ZN(n5852) );
  INV_X1 U5879 ( .A(n5852), .ZN(n4981) );
  NAND2_X1 U5880 ( .A1(n4752), .A2(n4981), .ZN(n4815) );
  NAND3_X1 U5881 ( .A1(n6564), .A2(n4756), .A3(n4815), .ZN(n4753) );
  OAI211_X1 U5882 ( .C1(n6564), .C2(n4754), .A(n6522), .B(n4753), .ZN(n4773)
         );
  NAND2_X1 U5883 ( .A1(n6564), .A2(n4815), .ZN(n4755) );
  OAI22_X1 U5884 ( .A1(n4756), .A2(n4755), .B1(n6780), .B2(n4781), .ZN(n4772)
         );
  AOI22_X1 U5885 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4773), .B1(n6589), 
        .B2(n4772), .ZN(n4759) );
  AOI22_X1 U5886 ( .A1(n3260), .A2(n6532), .B1(n4774), .B2(n6587), .ZN(n4758)
         );
  OAI211_X1 U5887 ( .C1(n4977), .C2(n5979), .A(n4759), .B(n4758), .ZN(U3126)
         );
  AOI22_X1 U5888 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4773), .B1(n6614), 
        .B2(n4772), .ZN(n4761) );
  AOI22_X1 U5889 ( .A1(n3260), .A2(n6548), .B1(n4774), .B2(n6611), .ZN(n4760)
         );
  OAI211_X1 U5890 ( .C1(n4977), .C2(n5997), .A(n4761), .B(n4760), .ZN(U3130)
         );
  AOI22_X1 U5891 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4773), .B1(n6583), 
        .B2(n4772), .ZN(n4763) );
  AOI22_X1 U5892 ( .A1(n3260), .A2(n6582), .B1(n4774), .B2(n3259), .ZN(n4762)
         );
  OAI211_X1 U5893 ( .C1(n4977), .C2(n6586), .A(n4763), .B(n4762), .ZN(U3125)
         );
  AOI22_X1 U5894 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4773), .B1(n6624), 
        .B2(n4772), .ZN(n4765) );
  AOI22_X1 U5895 ( .A1(n3260), .A2(n6621), .B1(n4774), .B2(n6620), .ZN(n4764)
         );
  OAI211_X1 U5896 ( .C1(n4977), .C2(n6629), .A(n4765), .B(n4764), .ZN(U3131)
         );
  AOI22_X1 U5897 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4773), .B1(n6595), 
        .B2(n4772), .ZN(n4767) );
  AOI22_X1 U5898 ( .A1(n3260), .A2(n6594), .B1(n4774), .B2(n6593), .ZN(n4766)
         );
  OAI211_X1 U5899 ( .C1(n4977), .C2(n6598), .A(n4767), .B(n4766), .ZN(U3127)
         );
  AOI22_X1 U5900 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4773), .B1(n6607), 
        .B2(n4772), .ZN(n4769) );
  AOI22_X1 U5901 ( .A1(n3260), .A2(n6544), .B1(n4774), .B2(n6605), .ZN(n4768)
         );
  OAI211_X1 U5902 ( .C1(n4977), .C2(n5887), .A(n4769), .B(n4768), .ZN(U3129)
         );
  AOI22_X1 U5903 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4773), .B1(n6601), 
        .B2(n4772), .ZN(n4771) );
  AOI22_X1 U5904 ( .A1(n3260), .A2(n6540), .B1(n4774), .B2(n6599), .ZN(n4770)
         );
  OAI211_X1 U5905 ( .C1(n4977), .C2(n5882), .A(n4771), .B(n4770), .ZN(U3128)
         );
  AOI22_X1 U5906 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4773), .B1(n6577), 
        .B2(n4772), .ZN(n4776) );
  AOI22_X1 U5907 ( .A1(n3260), .A2(n6518), .B1(n6562), .B2(n4774), .ZN(n4775)
         );
  OAI211_X1 U5908 ( .C1(n4977), .C2(n5865), .A(n4776), .B(n4775), .ZN(U3124)
         );
  INV_X1 U5909 ( .A(n4800), .ZN(n4777) );
  AOI21_X1 U5910 ( .B1(n4779), .B2(n4778), .A(n4777), .ZN(n6305) );
  INV_X1 U5911 ( .A(n6305), .ZN(n4888) );
  INV_X1 U5912 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6795) );
  OAI222_X1 U5913 ( .A1(n4888), .A2(n5339), .B1(n5338), .B2(n7086), .C1(n5593), 
        .C2(n6795), .ZN(U2887) );
  AOI21_X1 U5914 ( .B1(n6617), .B2(n4977), .A(n6781), .ZN(n4780) );
  AOI211_X1 U5915 ( .C1(n4786), .C2(n6513), .A(n6571), .B(n4780), .ZN(n4785)
         );
  NOR2_X1 U5916 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4781), .ZN(n4974)
         );
  AND2_X1 U5917 ( .A1(n4787), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5960) );
  INV_X1 U5918 ( .A(n5960), .ZN(n5194) );
  OAI21_X1 U5919 ( .B1(n7152), .B2(n4974), .A(n5194), .ZN(n4784) );
  NAND2_X1 U5920 ( .A1(n4894), .A2(n4893), .ZN(n4788) );
  AOI21_X1 U5921 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4788), .A(n4782), .ZN(
        n5136) );
  INV_X1 U5922 ( .A(n5136), .ZN(n4783) );
  NOR3_X1 U5923 ( .A1(n4785), .A2(n4784), .A3(n4783), .ZN(n4952) );
  INV_X1 U5924 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4794) );
  NAND2_X1 U5925 ( .A1(n4786), .A2(n6564), .ZN(n4900) );
  OR2_X1 U5926 ( .A1(n4900), .A2(n6315), .ZN(n4790) );
  NOR2_X1 U5927 ( .A1(n4787), .A2(n6780), .ZN(n5967) );
  INV_X1 U5928 ( .A(n4788), .ZN(n5127) );
  NAND2_X1 U5929 ( .A1(n5967), .A2(n5127), .ZN(n4789) );
  NAND2_X1 U5930 ( .A1(n4790), .A2(n4789), .ZN(n4973) );
  AOI22_X1 U5931 ( .A1(n6614), .A2(n4973), .B1(n6611), .B2(n4974), .ZN(n4793)
         );
  INV_X1 U5932 ( .A(n6548), .ZN(n6618) );
  OAI22_X1 U5933 ( .A1(n6617), .A2(n5997), .B1(n4977), .B2(n6618), .ZN(n4791)
         );
  INV_X1 U5934 ( .A(n4791), .ZN(n4792) );
  OAI211_X1 U5935 ( .C1(n4952), .C2(n4794), .A(n4793), .B(n4792), .ZN(U3122)
         );
  INV_X1 U5936 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4798) );
  AOI22_X1 U5937 ( .A1(n6589), .A2(n4973), .B1(n6587), .B2(n4974), .ZN(n4797)
         );
  INV_X1 U5938 ( .A(n6532), .ZN(n6592) );
  OAI22_X1 U5939 ( .A1(n6617), .A2(n5979), .B1(n4977), .B2(n6592), .ZN(n4795)
         );
  INV_X1 U5940 ( .A(n4795), .ZN(n4796) );
  OAI211_X1 U5941 ( .C1(n4952), .C2(n4798), .A(n4797), .B(n4796), .ZN(U3118)
         );
  AND2_X1 U5942 ( .A1(n4800), .A2(n4799), .ZN(n4802) );
  OR2_X1 U5943 ( .A1(n4802), .A2(n4801), .ZN(n5069) );
  AOI22_X1 U5944 ( .A1(n5557), .A2(n6283), .B1(n5556), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n4803) );
  OAI21_X1 U5945 ( .B1(n5069), .B2(n5575), .A(n4803), .ZN(U2854) );
  XNOR2_X1 U5946 ( .A(n4804), .B(n4805), .ZN(n5106) );
  NAND2_X1 U5947 ( .A1(n4807), .A2(n4806), .ZN(n5085) );
  NOR2_X1 U5948 ( .A1(n5085), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4812)
         );
  OR2_X1 U5949 ( .A1(n4809), .A2(n4808), .ZN(n4810) );
  NAND2_X1 U5950 ( .A1(n4810), .A2(n5122), .ZN(n6274) );
  NAND2_X1 U5951 ( .A1(n6425), .A2(REIP_REG_6__SCAN_IN), .ZN(n5100) );
  OAI21_X1 U5952 ( .B1(n5783), .B2(n6274), .A(n5100), .ZN(n4811) );
  AOI211_X1 U5953 ( .C1(n4813), .C2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n4812), 
        .B(n4811), .ZN(n4814) );
  OAI21_X1 U5954 ( .B1(n6475), .B2(n5106), .A(n4814), .ZN(U3012) );
  NAND2_X1 U5955 ( .A1(n4815), .A2(n6566), .ZN(n6759) );
  NOR3_X1 U5956 ( .A1(n6759), .A2(n4816), .A3(n6565), .ZN(n4817) );
  NOR2_X1 U5957 ( .A1(n4817), .A2(n6571), .ZN(n4823) );
  AND2_X1 U5958 ( .A1(n4622), .A2(n5317), .ZN(n5192) );
  NAND2_X1 U5959 ( .A1(n6315), .A2(n5192), .ZN(n4858) );
  OR2_X1 U5960 ( .A1(n4858), .A2(n3230), .ZN(n4819) );
  INV_X1 U5961 ( .A(n6561), .ZN(n4818) );
  NAND2_X1 U5962 ( .A1(n4818), .A2(n6765), .ZN(n4847) );
  NAND2_X1 U5963 ( .A1(n4819), .A2(n4847), .ZN(n4825) );
  NAND3_X1 U5964 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6765), .A3(n6643), .ZN(n4855) );
  INV_X1 U5965 ( .A(n4855), .ZN(n4820) );
  AOI22_X1 U5966 ( .A1(n4823), .A2(n4825), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4820), .ZN(n4852) );
  INV_X1 U5967 ( .A(n6621), .ZN(n6009) );
  OAI22_X1 U5968 ( .A1(n6005), .A2(n4847), .B1(n6009), .B2(n4924), .ZN(n4822)
         );
  AOI21_X1 U5969 ( .B1(n6555), .B2(n5846), .A(n4822), .ZN(n4828) );
  INV_X1 U5970 ( .A(n4823), .ZN(n4826) );
  AOI21_X1 U5971 ( .B1(n6571), .B2(n4855), .A(n6570), .ZN(n4824) );
  NAND2_X1 U5972 ( .A1(n4849), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4827) );
  OAI211_X1 U5973 ( .C1(n4852), .C2(n6559), .A(n4828), .B(n4827), .ZN(U3051)
         );
  INV_X1 U5974 ( .A(n6586), .ZN(n6528) );
  INV_X1 U5975 ( .A(n6582), .ZN(n5977) );
  OAI22_X1 U5976 ( .A1(n5973), .A2(n4847), .B1(n5977), .B2(n4924), .ZN(n4829)
         );
  AOI21_X1 U5977 ( .B1(n6528), .B2(n5846), .A(n4829), .ZN(n4831) );
  NAND2_X1 U5978 ( .A1(n4849), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4830) );
  OAI211_X1 U5979 ( .C1(n4852), .C2(n6531), .A(n4831), .B(n4830), .ZN(U3045)
         );
  OAI22_X1 U5980 ( .A1(n5988), .A2(n4847), .B1(n6604), .B2(n4924), .ZN(n4832)
         );
  AOI21_X1 U5981 ( .B1(n6600), .B2(n5846), .A(n4832), .ZN(n4834) );
  NAND2_X1 U5982 ( .A1(n4849), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4833) );
  OAI211_X1 U5983 ( .C1(n4852), .C2(n6543), .A(n4834), .B(n4833), .ZN(U3048)
         );
  INV_X1 U5984 ( .A(n6598), .ZN(n6536) );
  INV_X1 U5985 ( .A(n6594), .ZN(n5987) );
  OAI22_X1 U5986 ( .A1(n5983), .A2(n4847), .B1(n5987), .B2(n4924), .ZN(n4835)
         );
  AOI21_X1 U5987 ( .B1(n6536), .B2(n5846), .A(n4835), .ZN(n4837) );
  NAND2_X1 U5988 ( .A1(n4849), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4836) );
  OAI211_X1 U5989 ( .C1(n4852), .C2(n6539), .A(n4837), .B(n4836), .ZN(U3047)
         );
  INV_X1 U5990 ( .A(n5887), .ZN(n6606) );
  INV_X1 U5991 ( .A(n6544), .ZN(n6610) );
  OAI22_X1 U5992 ( .A1(n5992), .A2(n4847), .B1(n6610), .B2(n4924), .ZN(n4838)
         );
  AOI21_X1 U5993 ( .B1(n6606), .B2(n5846), .A(n4838), .ZN(n4840) );
  NAND2_X1 U5994 ( .A1(n4849), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4839) );
  OAI211_X1 U5995 ( .C1(n4852), .C2(n6547), .A(n4840), .B(n4839), .ZN(U3049)
         );
  INV_X1 U5996 ( .A(n6587), .ZN(n5978) );
  OAI22_X1 U5997 ( .A1(n5978), .A2(n4847), .B1(n6592), .B2(n4924), .ZN(n4841)
         );
  AOI21_X1 U5998 ( .B1(n6588), .B2(n5846), .A(n4841), .ZN(n4843) );
  NAND2_X1 U5999 ( .A1(n4849), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4842) );
  OAI211_X1 U6000 ( .C1(n4852), .C2(n6535), .A(n4843), .B(n4842), .ZN(U3046)
         );
  OAI22_X1 U6001 ( .A1(n5969), .A2(n4847), .B1(n6580), .B2(n4924), .ZN(n4844)
         );
  AOI21_X1 U6002 ( .B1(n6563), .B2(n5846), .A(n4844), .ZN(n4846) );
  NAND2_X1 U6003 ( .A1(n4849), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4845) );
  OAI211_X1 U6004 ( .C1(n4852), .C2(n6527), .A(n4846), .B(n4845), .ZN(U3044)
         );
  INV_X1 U6005 ( .A(n6611), .ZN(n5996) );
  OAI22_X1 U6006 ( .A1(n5996), .A2(n4847), .B1(n6618), .B2(n4924), .ZN(n4848)
         );
  AOI21_X1 U6007 ( .B1(n6612), .B2(n5846), .A(n4848), .ZN(n4851) );
  NAND2_X1 U6008 ( .A1(n4849), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4850) );
  OAI211_X1 U6009 ( .C1(n4852), .C2(n6551), .A(n4851), .B(n4850), .ZN(U3050)
         );
  OR2_X1 U6010 ( .A1(n5863), .A2(n5862), .ZN(n4988) );
  INV_X1 U6011 ( .A(n4988), .ZN(n4853) );
  OAI21_X1 U6012 ( .B1(n5846), .B2(n5847), .A(n4938), .ZN(n4854) );
  AOI21_X1 U6013 ( .B1(n4854), .B2(n4858), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4857) );
  NOR2_X1 U6014 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4855), .ZN(n5845)
         );
  NAND2_X1 U6015 ( .A1(n4893), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4856) );
  NAND2_X1 U6016 ( .A1(n4856), .A2(n4895), .ZN(n5961) );
  NOR2_X1 U6017 ( .A1(n5967), .A2(n5961), .ZN(n5199) );
  OAI21_X1 U6018 ( .B1(n4857), .B2(n5845), .A(n5199), .ZN(n5843) );
  INV_X1 U6019 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4864) );
  INV_X1 U6020 ( .A(n5847), .ZN(n4878) );
  OR2_X1 U6021 ( .A1(n4858), .A2(n6571), .ZN(n4860) );
  NOR2_X1 U6022 ( .A1(n4893), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5904)
         );
  NAND2_X1 U6023 ( .A1(n5960), .A2(n5904), .ZN(n4859) );
  NAND2_X1 U6024 ( .A1(n4860), .A2(n4859), .ZN(n5844) );
  AOI22_X1 U6025 ( .A1(n6593), .A2(n5845), .B1(n6595), .B2(n5844), .ZN(n4861)
         );
  OAI21_X1 U6026 ( .B1(n6598), .B2(n4878), .A(n4861), .ZN(n4862) );
  AOI21_X1 U6027 ( .B1(n6594), .B2(n5846), .A(n4862), .ZN(n4863) );
  OAI21_X1 U6028 ( .B1(n4887), .B2(n4864), .A(n4863), .ZN(U3039) );
  INV_X1 U6029 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4868) );
  AOI22_X1 U6030 ( .A1(n3259), .A2(n5845), .B1(n6583), .B2(n5844), .ZN(n4865)
         );
  OAI21_X1 U6031 ( .B1(n6586), .B2(n4878), .A(n4865), .ZN(n4866) );
  AOI21_X1 U6032 ( .B1(n6582), .B2(n5846), .A(n4866), .ZN(n4867) );
  OAI21_X1 U6033 ( .B1(n4887), .B2(n4868), .A(n4867), .ZN(U3037) );
  INV_X1 U6034 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4872) );
  AOI22_X1 U6035 ( .A1(n6620), .A2(n5845), .B1(n6624), .B2(n5844), .ZN(n4869)
         );
  OAI21_X1 U6036 ( .B1(n6629), .B2(n4878), .A(n4869), .ZN(n4870) );
  AOI21_X1 U6037 ( .B1(n6621), .B2(n5846), .A(n4870), .ZN(n4871) );
  OAI21_X1 U6038 ( .B1(n4887), .B2(n4872), .A(n4871), .ZN(U3043) );
  INV_X1 U6039 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4876) );
  AOI22_X1 U6040 ( .A1(n6605), .A2(n5845), .B1(n6607), .B2(n5844), .ZN(n4873)
         );
  OAI21_X1 U6041 ( .B1(n5887), .B2(n4878), .A(n4873), .ZN(n4874) );
  AOI21_X1 U6042 ( .B1(n6544), .B2(n5846), .A(n4874), .ZN(n4875) );
  OAI21_X1 U6043 ( .B1(n4887), .B2(n4876), .A(n4875), .ZN(U3041) );
  INV_X1 U6044 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4881) );
  AOI22_X1 U6045 ( .A1(n6599), .A2(n5845), .B1(n6601), .B2(n5844), .ZN(n4877)
         );
  OAI21_X1 U6046 ( .B1(n5882), .B2(n4878), .A(n4877), .ZN(n4879) );
  AOI21_X1 U6047 ( .B1(n6540), .B2(n5846), .A(n4879), .ZN(n4880) );
  OAI21_X1 U6048 ( .B1(n4887), .B2(n4881), .A(n4880), .ZN(U3040) );
  OAI222_X1 U6049 ( .A1(n5069), .A2(n5339), .B1(n5338), .B2(n7006), .C1(n5593), 
        .C2(n3940), .ZN(U2886) );
  AOI22_X1 U6050 ( .A1(n6589), .A2(n5844), .B1(n6587), .B2(n5845), .ZN(n4883)
         );
  AOI22_X1 U6051 ( .A1(n6588), .A2(n5847), .B1(n5846), .B2(n6532), .ZN(n4882)
         );
  OAI211_X1 U6052 ( .C1(n4887), .C2(n7138), .A(n4883), .B(n4882), .ZN(U3038)
         );
  INV_X1 U6053 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4886) );
  AOI22_X1 U6054 ( .A1(n6614), .A2(n5844), .B1(n6611), .B2(n5845), .ZN(n4885)
         );
  AOI22_X1 U6055 ( .A1(n6612), .A2(n5847), .B1(n5846), .B2(n6548), .ZN(n4884)
         );
  OAI211_X1 U6056 ( .C1(n4887), .C2(n4886), .A(n4885), .B(n4884), .ZN(U3042)
         );
  INV_X1 U6057 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4889) );
  OAI222_X1 U6058 ( .A1(n4890), .A2(n5592), .B1(n4889), .B2(n5591), .C1(n5575), 
        .C2(n4888), .ZN(U2855) );
  NOR2_X1 U6059 ( .A1(n4656), .A2(n3593), .ZN(n5128) );
  NAND2_X1 U6060 ( .A1(n5128), .A2(n3324), .ZN(n5897) );
  NAND3_X1 U6061 ( .A1(n4924), .A2(n6564), .A3(n5897), .ZN(n4892) );
  NOR2_X1 U6062 ( .A1(n4891), .A2(n6513), .ZN(n5854) );
  AOI21_X1 U6063 ( .B1(n4892), .B2(n4938), .A(n5854), .ZN(n4897) );
  INV_X1 U6064 ( .A(n4893), .ZN(n5193) );
  NOR2_X1 U6065 ( .A1(n5193), .A2(n4894), .ZN(n4942) );
  OAI21_X1 U6066 ( .B1(n4942), .B2(n6780), .A(n4895), .ZN(n4940) );
  NAND3_X1 U6067 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6765), .A3(n6637), .ZN(n5859) );
  NOR2_X1 U6068 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5859), .ZN(n4928)
         );
  NOR2_X1 U6069 ( .A1(n7152), .A2(n4928), .ZN(n4896) );
  NOR4_X2 U6070 ( .A1(n4897), .A2(n5960), .A3(n4940), .A4(n4896), .ZN(n4935)
         );
  INV_X1 U6071 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4904) );
  INV_X1 U6072 ( .A(n5967), .ZN(n4899) );
  INV_X1 U6073 ( .A(n4942), .ZN(n4898) );
  OAI22_X1 U6074 ( .A1(n4900), .A2(n4582), .B1(n4899), .B2(n4898), .ZN(n4929)
         );
  AOI22_X1 U6075 ( .A1(n6562), .A2(n4928), .B1(n6577), .B2(n4929), .ZN(n4901)
         );
  OAI21_X1 U6076 ( .B1(n5865), .B2(n4924), .A(n4901), .ZN(n4902) );
  AOI21_X1 U6077 ( .B1(n6518), .B2(n4930), .A(n4902), .ZN(n4903) );
  OAI21_X1 U6078 ( .B1(n4935), .B2(n4904), .A(n4903), .ZN(U3052) );
  INV_X1 U6079 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4908) );
  AOI22_X1 U6080 ( .A1(n6620), .A2(n4928), .B1(n6624), .B2(n4929), .ZN(n4905)
         );
  OAI21_X1 U6081 ( .B1(n6629), .B2(n4924), .A(n4905), .ZN(n4906) );
  AOI21_X1 U6082 ( .B1(n6621), .B2(n4930), .A(n4906), .ZN(n4907) );
  OAI21_X1 U6083 ( .B1(n4935), .B2(n4908), .A(n4907), .ZN(U3059) );
  INV_X1 U6084 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4912) );
  AOI22_X1 U6085 ( .A1(n6605), .A2(n4928), .B1(n6607), .B2(n4929), .ZN(n4909)
         );
  OAI21_X1 U6086 ( .B1(n5887), .B2(n4924), .A(n4909), .ZN(n4910) );
  AOI21_X1 U6087 ( .B1(n6544), .B2(n4930), .A(n4910), .ZN(n4911) );
  OAI21_X1 U6088 ( .B1(n4935), .B2(n4912), .A(n4911), .ZN(U3057) );
  INV_X1 U6089 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4916) );
  AOI22_X1 U6090 ( .A1(n6599), .A2(n4928), .B1(n6601), .B2(n4929), .ZN(n4913)
         );
  OAI21_X1 U6091 ( .B1(n5882), .B2(n4924), .A(n4913), .ZN(n4914) );
  AOI21_X1 U6092 ( .B1(n6540), .B2(n4930), .A(n4914), .ZN(n4915) );
  OAI21_X1 U6093 ( .B1(n4935), .B2(n4916), .A(n4915), .ZN(U3056) );
  AOI22_X1 U6094 ( .A1(n6581), .A2(n4928), .B1(n6583), .B2(n4929), .ZN(n4917)
         );
  OAI21_X1 U6095 ( .B1(n6586), .B2(n4924), .A(n4917), .ZN(n4918) );
  AOI21_X1 U6096 ( .B1(n6582), .B2(n4930), .A(n4918), .ZN(n4919) );
  OAI21_X1 U6097 ( .B1(n4935), .B2(n6981), .A(n4919), .ZN(U3053) );
  INV_X1 U6098 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4923) );
  AOI22_X1 U6099 ( .A1(n6593), .A2(n4928), .B1(n6595), .B2(n4929), .ZN(n4920)
         );
  OAI21_X1 U6100 ( .B1(n6598), .B2(n4924), .A(n4920), .ZN(n4921) );
  AOI21_X1 U6101 ( .B1(n6594), .B2(n4930), .A(n4921), .ZN(n4922) );
  OAI21_X1 U6102 ( .B1(n4935), .B2(n4923), .A(n4922), .ZN(U3055) );
  INV_X1 U6103 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4927) );
  AOI22_X1 U6104 ( .A1(n6614), .A2(n4929), .B1(n6611), .B2(n4928), .ZN(n4926)
         );
  INV_X1 U6105 ( .A(n4924), .ZN(n4931) );
  AOI22_X1 U6106 ( .A1(n4931), .A2(n6612), .B1(n4930), .B2(n6548), .ZN(n4925)
         );
  OAI211_X1 U6107 ( .C1(n4935), .C2(n4927), .A(n4926), .B(n4925), .ZN(U3058)
         );
  INV_X1 U6108 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4934) );
  AOI22_X1 U6109 ( .A1(n6589), .A2(n4929), .B1(n6587), .B2(n4928), .ZN(n4933)
         );
  AOI22_X1 U6110 ( .A1(n4931), .A2(n6588), .B1(n4930), .B2(n6532), .ZN(n4932)
         );
  OAI211_X1 U6111 ( .C1(n4935), .C2(n4934), .A(n4933), .B(n4932), .ZN(U3054)
         );
  NAND2_X1 U6112 ( .A1(n4622), .A2(n5494), .ZN(n5126) );
  INV_X1 U6113 ( .A(n5014), .ZN(n4937) );
  INV_X1 U6114 ( .A(n4944), .ZN(n4936) );
  OAI21_X1 U6115 ( .B1(n4936), .B2(n5852), .A(n6564), .ZN(n5019) );
  AOI211_X1 U6116 ( .C1(n5837), .C2(n4938), .A(n4937), .B(n5019), .ZN(n4941)
         );
  NAND3_X1 U6117 ( .A1(n6765), .A2(n6643), .A3(n6637), .ZN(n5017) );
  NOR2_X1 U6118 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5017), .ZN(n5836)
         );
  NOR2_X1 U6119 ( .A1(n7152), .A2(n5836), .ZN(n4939) );
  NOR4_X1 U6120 ( .A1(n4941), .A2(n4940), .A3(n5967), .A4(n4939), .ZN(n5813)
         );
  INV_X1 U6121 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4947) );
  NAND2_X1 U6122 ( .A1(n4942), .A2(n5960), .ZN(n4943) );
  OAI21_X1 U6123 ( .B1(n5014), .B2(n6571), .A(n4943), .ZN(n5835) );
  AOI22_X1 U6124 ( .A1(n6614), .A2(n5835), .B1(n6611), .B2(n5836), .ZN(n4946)
         );
  INV_X1 U6125 ( .A(n5838), .ZN(n4948) );
  AOI22_X1 U6126 ( .A1(n4948), .A2(n6548), .B1(n5837), .B2(n6612), .ZN(n4945)
         );
  OAI211_X1 U6127 ( .C1(n5813), .C2(n4947), .A(n4946), .B(n4945), .ZN(U3026)
         );
  INV_X1 U6128 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4951) );
  AOI22_X1 U6129 ( .A1(n6589), .A2(n5835), .B1(n6587), .B2(n5836), .ZN(n4950)
         );
  AOI22_X1 U6130 ( .A1(n4948), .A2(n6532), .B1(n5837), .B2(n6588), .ZN(n4949)
         );
  OAI211_X1 U6131 ( .C1(n5813), .C2(n4951), .A(n4950), .B(n4949), .ZN(U3022)
         );
  INV_X1 U6132 ( .A(n4952), .ZN(n4979) );
  NAND2_X1 U6133 ( .A1(n6622), .A2(n6600), .ZN(n4954) );
  AOI22_X1 U6134 ( .A1(n6599), .A2(n4974), .B1(n6601), .B2(n4973), .ZN(n4953)
         );
  OAI211_X1 U6135 ( .C1(n6604), .C2(n4977), .A(n4954), .B(n4953), .ZN(n4955)
         );
  AOI21_X1 U6136 ( .B1(n4979), .B2(INSTQUEUE_REG_12__4__SCAN_IN), .A(n4955), 
        .ZN(n4956) );
  INV_X1 U6137 ( .A(n4956), .ZN(U3120) );
  NAND2_X1 U6138 ( .A1(n6622), .A2(n6563), .ZN(n4958) );
  AOI22_X1 U6139 ( .A1(n6562), .A2(n4974), .B1(n6577), .B2(n4973), .ZN(n4957)
         );
  OAI211_X1 U6140 ( .C1(n6580), .C2(n4977), .A(n4958), .B(n4957), .ZN(n4959)
         );
  AOI21_X1 U6141 ( .B1(n4979), .B2(INSTQUEUE_REG_12__0__SCAN_IN), .A(n4959), 
        .ZN(n4960) );
  INV_X1 U6142 ( .A(n4960), .ZN(U3116) );
  NAND2_X1 U6143 ( .A1(n6622), .A2(n6536), .ZN(n4962) );
  AOI22_X1 U6144 ( .A1(n6593), .A2(n4974), .B1(n6595), .B2(n4973), .ZN(n4961)
         );
  OAI211_X1 U6145 ( .C1(n5987), .C2(n4977), .A(n4962), .B(n4961), .ZN(n4963)
         );
  AOI21_X1 U6146 ( .B1(n4979), .B2(INSTQUEUE_REG_12__3__SCAN_IN), .A(n4963), 
        .ZN(n4964) );
  INV_X1 U6147 ( .A(n4964), .ZN(U3119) );
  NAND2_X1 U6148 ( .A1(n6622), .A2(n6528), .ZN(n4966) );
  AOI22_X1 U6149 ( .A1(n6581), .A2(n4974), .B1(n6583), .B2(n4973), .ZN(n4965)
         );
  OAI211_X1 U6150 ( .C1(n5977), .C2(n4977), .A(n4966), .B(n4965), .ZN(n4967)
         );
  AOI21_X1 U6151 ( .B1(n4979), .B2(INSTQUEUE_REG_12__1__SCAN_IN), .A(n4967), 
        .ZN(n4968) );
  INV_X1 U6152 ( .A(n4968), .ZN(U3117) );
  NAND2_X1 U6153 ( .A1(n6622), .A2(n6606), .ZN(n4970) );
  AOI22_X1 U6154 ( .A1(n6605), .A2(n4974), .B1(n6607), .B2(n4973), .ZN(n4969)
         );
  OAI211_X1 U6155 ( .C1(n6610), .C2(n4977), .A(n4970), .B(n4969), .ZN(n4971)
         );
  AOI21_X1 U6156 ( .B1(n4979), .B2(INSTQUEUE_REG_12__5__SCAN_IN), .A(n4971), 
        .ZN(n4972) );
  INV_X1 U6157 ( .A(n4972), .ZN(U3121) );
  NAND2_X1 U6158 ( .A1(n6622), .A2(n6555), .ZN(n4976) );
  AOI22_X1 U6159 ( .A1(n6620), .A2(n4974), .B1(n6624), .B2(n4973), .ZN(n4975)
         );
  OAI211_X1 U6160 ( .C1(n6009), .C2(n4977), .A(n4976), .B(n4975), .ZN(n4978)
         );
  AOI21_X1 U6161 ( .B1(n4979), .B2(INSTQUEUE_REG_12__7__SCAN_IN), .A(n4978), 
        .ZN(n4980) );
  INV_X1 U6162 ( .A(n4980), .ZN(U3123) );
  AOI21_X1 U6163 ( .B1(n5188), .B2(n4981), .A(n6571), .ZN(n4985) );
  INV_X1 U6164 ( .A(n5126), .ZN(n4982) );
  NAND3_X1 U6165 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6643), .A3(n6637), .ZN(n5130) );
  NOR2_X1 U6166 ( .A1(n6633), .A2(n5130), .ZN(n5005) );
  AOI21_X1 U6167 ( .B1(n4983), .B2(n4982), .A(n5005), .ZN(n4987) );
  AOI22_X1 U6168 ( .A1(n4985), .A2(n4987), .B1(n6571), .B2(n5130), .ZN(n4984)
         );
  NAND2_X1 U6169 ( .A1(n6522), .A2(n4984), .ZN(n5004) );
  INV_X1 U6170 ( .A(n4985), .ZN(n4986) );
  OAI22_X1 U6171 ( .A1(n4987), .A2(n4986), .B1(n6780), .B2(n5130), .ZN(n5003)
         );
  AOI22_X1 U6172 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n5004), .B1(n6614), 
        .B2(n5003), .ZN(n4990) );
  AOI22_X1 U6173 ( .A1(n6548), .A2(n5952), .B1(n6611), .B2(n5005), .ZN(n4989)
         );
  OAI211_X1 U6174 ( .C1(n5997), .C2(n5131), .A(n4990), .B(n4989), .ZN(U3098)
         );
  AOI22_X1 U6175 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n5004), .B1(n6589), 
        .B2(n5003), .ZN(n4992) );
  AOI22_X1 U6176 ( .A1(n6532), .A2(n5952), .B1(n6587), .B2(n5005), .ZN(n4991)
         );
  OAI211_X1 U6177 ( .C1(n5979), .C2(n5131), .A(n4992), .B(n4991), .ZN(U3094)
         );
  AOI22_X1 U6178 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n5004), .B1(n6583), 
        .B2(n5003), .ZN(n4994) );
  AOI22_X1 U6179 ( .A1(n6582), .A2(n5952), .B1(n3259), .B2(n5005), .ZN(n4993)
         );
  OAI211_X1 U6180 ( .C1(n6586), .C2(n5131), .A(n4994), .B(n4993), .ZN(U3093)
         );
  AOI22_X1 U6181 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5004), .B1(n6624), 
        .B2(n5003), .ZN(n4996) );
  AOI22_X1 U6182 ( .A1(n6621), .A2(n5952), .B1(n6620), .B2(n5005), .ZN(n4995)
         );
  OAI211_X1 U6183 ( .C1(n6629), .C2(n5131), .A(n4996), .B(n4995), .ZN(U3099)
         );
  AOI22_X1 U6184 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n5004), .B1(n6595), 
        .B2(n5003), .ZN(n4998) );
  AOI22_X1 U6185 ( .A1(n6594), .A2(n5952), .B1(n6593), .B2(n5005), .ZN(n4997)
         );
  OAI211_X1 U6186 ( .C1(n6598), .C2(n5131), .A(n4998), .B(n4997), .ZN(U3095)
         );
  AOI22_X1 U6187 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5004), .B1(n6601), 
        .B2(n5003), .ZN(n5000) );
  AOI22_X1 U6188 ( .A1(n6540), .A2(n5952), .B1(n6599), .B2(n5005), .ZN(n4999)
         );
  OAI211_X1 U6189 ( .C1(n5882), .C2(n5131), .A(n5000), .B(n4999), .ZN(U3096)
         );
  AOI22_X1 U6190 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n5004), .B1(n6607), 
        .B2(n5003), .ZN(n5002) );
  AOI22_X1 U6191 ( .A1(n6544), .A2(n5952), .B1(n6605), .B2(n5005), .ZN(n5001)
         );
  OAI211_X1 U6192 ( .C1(n5887), .C2(n5131), .A(n5002), .B(n5001), .ZN(U3097)
         );
  AOI22_X1 U6193 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5004), .B1(n6577), 
        .B2(n5003), .ZN(n5007) );
  AOI22_X1 U6194 ( .A1(n6518), .A2(n5952), .B1(n6562), .B2(n5005), .ZN(n5006)
         );
  OAI211_X1 U6195 ( .C1(n5865), .C2(n5131), .A(n5007), .B(n5006), .ZN(U3092)
         );
  NOR2_X1 U6196 ( .A1(n4801), .A2(n5009), .ZN(n5010) );
  OR2_X1 U6197 ( .A1(n5008), .A2(n5010), .ZN(n6279) );
  INV_X1 U6198 ( .A(n6274), .ZN(n5011) );
  AOI22_X1 U6199 ( .A1(n5557), .A2(n5011), .B1(n5556), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n5012) );
  OAI21_X1 U6200 ( .B1(n6279), .B2(n5575), .A(n5012), .ZN(U2853) );
  NOR2_X1 U6201 ( .A1(n6633), .A2(n5017), .ZN(n5048) );
  INV_X1 U6202 ( .A(n5048), .ZN(n5013) );
  OAI21_X1 U6203 ( .B1(n5014), .B2(n3230), .A(n5013), .ZN(n5016) );
  NOR2_X1 U6204 ( .A1(n5019), .A2(n5016), .ZN(n5015) );
  INV_X1 U6205 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5023) );
  INV_X1 U6206 ( .A(n5016), .ZN(n5018) );
  OAI22_X1 U6207 ( .A1(n5019), .A2(n5018), .B1(n5017), .B2(n6780), .ZN(n5051)
         );
  AOI22_X1 U6208 ( .A1(n6548), .A2(n5847), .B1(n6611), .B2(n5048), .ZN(n5020)
         );
  OAI21_X1 U6209 ( .B1(n5997), .B2(n5838), .A(n5020), .ZN(n5021) );
  AOI21_X1 U6210 ( .B1(n5051), .B2(n6614), .A(n5021), .ZN(n5022) );
  OAI21_X1 U6211 ( .B1(n5054), .B2(n5023), .A(n5022), .ZN(U3034) );
  INV_X1 U6212 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5027) );
  AOI22_X1 U6213 ( .A1(n6621), .A2(n5847), .B1(n6620), .B2(n5048), .ZN(n5024)
         );
  OAI21_X1 U6214 ( .B1(n6629), .B2(n5838), .A(n5024), .ZN(n5025) );
  AOI21_X1 U6215 ( .B1(n5051), .B2(n6624), .A(n5025), .ZN(n5026) );
  OAI21_X1 U6216 ( .B1(n5054), .B2(n5027), .A(n5026), .ZN(U3035) );
  INV_X1 U6217 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n5031) );
  AOI22_X1 U6218 ( .A1(n6544), .A2(n5847), .B1(n6605), .B2(n5048), .ZN(n5028)
         );
  OAI21_X1 U6219 ( .B1(n5887), .B2(n5838), .A(n5028), .ZN(n5029) );
  AOI21_X1 U6220 ( .B1(n5051), .B2(n6607), .A(n5029), .ZN(n5030) );
  OAI21_X1 U6221 ( .B1(n5054), .B2(n5031), .A(n5030), .ZN(U3033) );
  INV_X1 U6222 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n5035) );
  AOI22_X1 U6223 ( .A1(n6582), .A2(n5847), .B1(n6581), .B2(n5048), .ZN(n5032)
         );
  OAI21_X1 U6224 ( .B1(n6586), .B2(n5838), .A(n5032), .ZN(n5033) );
  AOI21_X1 U6225 ( .B1(n5051), .B2(n6583), .A(n5033), .ZN(n5034) );
  OAI21_X1 U6226 ( .B1(n5054), .B2(n5035), .A(n5034), .ZN(U3029) );
  INV_X1 U6227 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n5039) );
  AOI22_X1 U6228 ( .A1(n6540), .A2(n5847), .B1(n6599), .B2(n5048), .ZN(n5036)
         );
  OAI21_X1 U6229 ( .B1(n5882), .B2(n5838), .A(n5036), .ZN(n5037) );
  AOI21_X1 U6230 ( .B1(n5051), .B2(n6601), .A(n5037), .ZN(n5038) );
  OAI21_X1 U6231 ( .B1(n5054), .B2(n5039), .A(n5038), .ZN(U3032) );
  INV_X1 U6232 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n5043) );
  AOI22_X1 U6233 ( .A1(n6594), .A2(n5847), .B1(n6593), .B2(n5048), .ZN(n5040)
         );
  OAI21_X1 U6234 ( .B1(n6598), .B2(n5838), .A(n5040), .ZN(n5041) );
  AOI21_X1 U6235 ( .B1(n5051), .B2(n6595), .A(n5041), .ZN(n5042) );
  OAI21_X1 U6236 ( .B1(n5054), .B2(n5043), .A(n5042), .ZN(U3031) );
  INV_X1 U6237 ( .A(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n5047) );
  AOI22_X1 U6238 ( .A1(n6518), .A2(n5847), .B1(n6562), .B2(n5048), .ZN(n5044)
         );
  OAI21_X1 U6239 ( .B1(n5865), .B2(n5838), .A(n5044), .ZN(n5045) );
  AOI21_X1 U6240 ( .B1(n5051), .B2(n6577), .A(n5045), .ZN(n5046) );
  OAI21_X1 U6241 ( .B1(n5054), .B2(n5047), .A(n5046), .ZN(U3028) );
  INV_X1 U6242 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n5053) );
  AOI22_X1 U6243 ( .A1(n6532), .A2(n5847), .B1(n6587), .B2(n5048), .ZN(n5049)
         );
  OAI21_X1 U6244 ( .B1(n5979), .B2(n5838), .A(n5049), .ZN(n5050) );
  AOI21_X1 U6245 ( .B1(n5051), .B2(n6589), .A(n5050), .ZN(n5052) );
  OAI21_X1 U6246 ( .B1(n5054), .B2(n5053), .A(n5052), .ZN(U3030) );
  OR2_X1 U6247 ( .A1(n5056), .A2(n5055), .ZN(n5058) );
  AND2_X1 U6248 ( .A1(n5058), .A2(n5057), .ZN(n6508) );
  AOI22_X1 U6249 ( .A1(n6442), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6425), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5059) );
  OAI21_X1 U6250 ( .B1(n6437), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n5059), 
        .ZN(n5060) );
  AOI21_X1 U6251 ( .B1(n6508), .B2(n6431), .A(n5060), .ZN(n5061) );
  OAI21_X1 U6252 ( .B1(n5320), .B2(n5714), .A(n5061), .ZN(U2985) );
  INV_X1 U6253 ( .A(DATAI_6_), .ZN(n5062) );
  OAI222_X1 U6254 ( .A1(n6279), .A2(n5339), .B1(n5338), .B2(n5062), .C1(n5593), 
        .C2(n3944), .ZN(U2885) );
  XNOR2_X1 U6255 ( .A(n5063), .B(n5064), .ZN(n6476) );
  INV_X1 U6256 ( .A(n6322), .ZN(n5067) );
  AND2_X1 U6257 ( .A1(n6425), .A2(REIP_REG_3__SCAN_IN), .ZN(n6473) );
  AOI21_X1 U6258 ( .B1(n6442), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n6473), 
        .ZN(n5065) );
  OAI21_X1 U6259 ( .B1(n6437), .B2(n6320), .A(n5065), .ZN(n5066) );
  AOI21_X1 U6260 ( .B1(n5067), .B2(n6432), .A(n5066), .ZN(n5068) );
  OAI21_X1 U6261 ( .B1(n6476), .B2(n6438), .A(n5068), .ZN(U2983) );
  INV_X1 U6262 ( .A(n5069), .ZN(n6287) );
  AOI21_X1 U6263 ( .B1(n6442), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n5070), 
        .ZN(n5071) );
  OAI21_X1 U6264 ( .B1(n6437), .B2(n6292), .A(n5071), .ZN(n5072) );
  AOI21_X1 U6265 ( .B1(n6287), .B2(n6432), .A(n5072), .ZN(n5073) );
  OAI21_X1 U6266 ( .B1(n6438), .B2(n5074), .A(n5073), .ZN(U2981) );
  INV_X1 U6267 ( .A(n6303), .ZN(n5077) );
  AOI21_X1 U6268 ( .B1(n6442), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n5075), 
        .ZN(n5076) );
  OAI21_X1 U6269 ( .B1(n6437), .B2(n5077), .A(n5076), .ZN(n5078) );
  AOI21_X1 U6270 ( .B1(n6305), .B2(n6432), .A(n5078), .ZN(n5079) );
  OAI21_X1 U6271 ( .B1(n6438), .B2(n5080), .A(n5079), .ZN(U2982) );
  XNOR2_X1 U6272 ( .A(n5081), .B(n5082), .ZN(n5286) );
  OR2_X1 U6273 ( .A1(n5083), .A2(n5121), .ZN(n5084) );
  NAND2_X1 U6274 ( .A1(n5084), .A2(n5146), .ZN(n5229) );
  INV_X1 U6275 ( .A(n5229), .ZN(n5118) );
  NAND2_X1 U6276 ( .A1(n6425), .A2(REIP_REG_8__SCAN_IN), .ZN(n5279) );
  AOI21_X1 U6277 ( .B1(n6470), .B2(n5095), .A(n5167), .ZN(n5087) );
  NOR2_X1 U6278 ( .A1(n5086), .A2(n5085), .ZN(n6462) );
  NAND2_X1 U6279 ( .A1(n5087), .A2(n6462), .ZN(n5088) );
  NAND2_X1 U6280 ( .A1(n5279), .A2(n5088), .ZN(n5097) );
  NOR2_X1 U6281 ( .A1(n5090), .A2(n5089), .ZN(n5091) );
  AOI211_X1 U6282 ( .C1(n5094), .C2(n5093), .A(n5092), .B(n5091), .ZN(n6471)
         );
  NOR2_X1 U6283 ( .A1(n6471), .A2(n5095), .ZN(n5096) );
  AOI211_X1 U6284 ( .C1(n6503), .C2(n5118), .A(n5097), .B(n5096), .ZN(n5098)
         );
  OAI21_X1 U6285 ( .B1(n6475), .B2(n5286), .A(n5098), .ZN(U3010) );
  INV_X1 U6286 ( .A(n6279), .ZN(n5104) );
  INV_X1 U6287 ( .A(n5099), .ZN(n6277) );
  INV_X1 U6288 ( .A(n5100), .ZN(n5101) );
  AOI21_X1 U6289 ( .B1(n6442), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n5101), 
        .ZN(n5102) );
  OAI21_X1 U6290 ( .B1(n6437), .B2(n6277), .A(n5102), .ZN(n5103) );
  AOI21_X1 U6291 ( .B1(n5104), .B2(n6432), .A(n5103), .ZN(n5105) );
  OAI21_X1 U6292 ( .B1(n6438), .B2(n5106), .A(n5105), .ZN(U2980) );
  INV_X1 U6293 ( .A(n5116), .ZN(n5107) );
  OAI21_X1 U6294 ( .B1(n5008), .B2(n5108), .A(n5107), .ZN(n6265) );
  XOR2_X1 U6295 ( .A(n5110), .B(n5109), .Z(n6468) );
  NAND2_X1 U6296 ( .A1(n6468), .A2(n6431), .ZN(n5114) );
  NAND2_X1 U6297 ( .A1(n6425), .A2(REIP_REG_7__SCAN_IN), .ZN(n6464) );
  INV_X1 U6298 ( .A(n6464), .ZN(n5112) );
  NOR2_X1 U6299 ( .A1(n6437), .A2(n6264), .ZN(n5111) );
  AOI211_X1 U6300 ( .C1(n6442), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n5112), 
        .B(n5111), .ZN(n5113) );
  OAI211_X1 U6301 ( .C1(n5714), .C2(n6265), .A(n5114), .B(n5113), .ZN(U2979)
         );
  OAI21_X1 U6302 ( .B1(n5116), .B2(n5115), .A(n5143), .ZN(n5281) );
  AOI22_X1 U6303 ( .A1(n5331), .A2(DATAI_8_), .B1(n6332), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n5117) );
  OAI21_X1 U6304 ( .B1(n5281), .B2(n5339), .A(n5117), .ZN(U2883) );
  AOI22_X1 U6305 ( .A1(n5557), .A2(n5118), .B1(n5556), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n5119) );
  OAI21_X1 U6306 ( .B1(n5281), .B2(n5575), .A(n5119), .ZN(U2851) );
  INV_X1 U6307 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6404) );
  OAI222_X1 U6308 ( .A1(n6265), .A2(n5339), .B1(n5338), .B2(n5120), .C1(n5593), 
        .C2(n6404), .ZN(U2884) );
  AOI21_X1 U6309 ( .B1(n5123), .B2(n5122), .A(n5121), .ZN(n6463) );
  INV_X1 U6310 ( .A(n6463), .ZN(n5125) );
  INV_X1 U6311 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5124) );
  OAI222_X1 U6312 ( .A1(n5125), .A2(n5592), .B1(n5124), .B2(n5591), .C1(n5575), 
        .C2(n6265), .ZN(U2852) );
  NOR2_X1 U6313 ( .A1(n6315), .A2(n5126), .ZN(n5132) );
  AOI22_X1 U6314 ( .A1(n5132), .A2(n6564), .B1(n5960), .B2(n5127), .ZN(n5255)
         );
  INV_X1 U6315 ( .A(n5128), .ZN(n6519) );
  AOI22_X1 U6316 ( .A1(n6588), .A2(n6553), .B1(n5276), .B2(n6532), .ZN(n5138)
         );
  NOR2_X1 U6317 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5130), .ZN(n5139)
         );
  INV_X1 U6318 ( .A(n5139), .ZN(n5274) );
  AOI21_X1 U6319 ( .B1(n5131), .B2(n5278), .A(n6781), .ZN(n5133) );
  NOR3_X1 U6320 ( .A1(n5133), .A2(n5132), .A3(n6571), .ZN(n5134) );
  AOI211_X1 U6321 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5274), .A(n5134), .B(
        n5967), .ZN(n5135) );
  NAND2_X1 U6322 ( .A1(n5136), .A2(n5135), .ZN(n5271) );
  AOI22_X1 U6323 ( .A1(n6587), .A2(n5139), .B1(INSTQUEUE_REG_8__2__SCAN_IN), 
        .B2(n5271), .ZN(n5137) );
  OAI211_X1 U6324 ( .C1(n6535), .C2(n5255), .A(n5138), .B(n5137), .ZN(U3086)
         );
  AOI22_X1 U6325 ( .A1(n6612), .A2(n6553), .B1(n5276), .B2(n6548), .ZN(n5141)
         );
  AOI22_X1 U6326 ( .A1(n6611), .A2(n5139), .B1(INSTQUEUE_REG_8__6__SCAN_IN), 
        .B2(n5271), .ZN(n5140) );
  OAI211_X1 U6327 ( .C1(n6551), .C2(n5255), .A(n5141), .B(n5140), .ZN(U3090)
         );
  NAND2_X1 U6328 ( .A1(n5143), .A2(n5142), .ZN(n5144) );
  NAND2_X1 U6329 ( .A1(n5287), .A2(n5144), .ZN(n5174) );
  AOI22_X1 U6330 ( .A1(n5331), .A2(DATAI_9_), .B1(n6332), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n5145) );
  OAI21_X1 U6331 ( .B1(n5174), .B2(n5339), .A(n5145), .ZN(U2882) );
  INV_X1 U6332 ( .A(n5160), .ZN(n5155) );
  NAND2_X1 U6333 ( .A1(n6307), .A2(n5150), .ZN(n6249) );
  NAND2_X1 U6334 ( .A1(n5147), .A2(n5146), .ZN(n5149) );
  INV_X1 U6335 ( .A(n5169), .ZN(n5148) );
  NAND2_X1 U6336 ( .A1(n5149), .A2(n5148), .ZN(n6454) );
  OAI22_X1 U6337 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6249), .B1(n6318), .B2(n6454), .ZN(n5154) );
  INV_X1 U6338 ( .A(n5150), .ZN(n5151) );
  NAND2_X1 U6339 ( .A1(n6307), .A2(n5151), .ZN(n5235) );
  NAND2_X1 U6340 ( .A1(n5235), .A2(n6296), .ZN(n6252) );
  AOI22_X1 U6341 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6325), .B1(
        REIP_REG_9__SCAN_IN), .B2(n6252), .ZN(n5152) );
  OAI211_X1 U6342 ( .C1(n6314), .C2(n6969), .A(n5152), .B(n6498), .ZN(n5153)
         );
  AOI211_X1 U6343 ( .C1(n6302), .C2(n5155), .A(n5154), .B(n5153), .ZN(n5156)
         );
  OAI21_X1 U6344 ( .B1(n6278), .B2(n5174), .A(n5156), .ZN(U2818) );
  XNOR2_X1 U6345 ( .A(n3184), .B(n7009), .ZN(n5158) );
  XNOR2_X1 U6346 ( .A(n5157), .B(n5158), .ZN(n6457) );
  NAND2_X1 U6347 ( .A1(n6457), .A2(n6431), .ZN(n5163) );
  INV_X1 U6348 ( .A(REIP_REG_9__SCAN_IN), .ZN(n5159) );
  NOR2_X1 U6349 ( .A1(n6498), .A2(n5159), .ZN(n6455) );
  NOR2_X1 U6350 ( .A1(n6437), .A2(n5160), .ZN(n5161) );
  AOI211_X1 U6351 ( .C1(n6442), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6455), 
        .B(n5161), .ZN(n5162) );
  OAI211_X1 U6352 ( .C1(n5714), .C2(n5174), .A(n5163), .B(n5162), .ZN(U2977)
         );
  NAND2_X1 U6353 ( .A1(n3253), .A2(n5165), .ZN(n5166) );
  XNOR2_X1 U6354 ( .A(n5164), .B(n5166), .ZN(n5294) );
  OAI21_X1 U6355 ( .B1(n5781), .B2(n5167), .A(n6471), .ZN(n6458) );
  NAND2_X1 U6356 ( .A1(n5167), .A2(n6462), .ZN(n6461) );
  AOI221_X1 U6357 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n7009), .C2(n5168), .A(n6461), 
        .ZN(n5172) );
  OAI21_X1 U6358 ( .B1(n5170), .B2(n5169), .A(n5300), .ZN(n6248) );
  INV_X1 U6359 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6703) );
  OAI22_X1 U6360 ( .A1(n5783), .A2(n6248), .B1(n6703), .B2(n6498), .ZN(n5171)
         );
  AOI211_X1 U6361 ( .C1(n6458), .C2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n5172), .B(n5171), .ZN(n5173) );
  OAI21_X1 U6362 ( .B1(n6475), .B2(n5294), .A(n5173), .ZN(U3008) );
  INV_X1 U6363 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5175) );
  OAI222_X1 U6364 ( .A1(n6454), .A2(n5592), .B1(n5591), .B2(n5175), .C1(n5575), 
        .C2(n5174), .ZN(U2850) );
  INV_X1 U6365 ( .A(DATAI_13_), .ZN(n7022) );
  XNOR2_X1 U6366 ( .A(n5177), .B(n5176), .ZN(n6218) );
  OAI222_X1 U6367 ( .A1(n5593), .A2(n6418), .B1(n5338), .B2(n7022), .C1(n5339), 
        .C2(n6218), .ZN(U2878) );
  AOI21_X1 U6368 ( .B1(n5179), .B2(n5178), .A(n5242), .ZN(n6216) );
  INV_X1 U6369 ( .A(n6216), .ZN(n5181) );
  OAI222_X1 U6370 ( .A1(n5181), .A2(n5592), .B1(n5575), .B2(n6218), .C1(n5591), 
        .C2(n5180), .ZN(U2846) );
  OR2_X1 U6371 ( .A1(n5184), .A2(n5183), .ZN(n5185) );
  NAND2_X1 U6372 ( .A1(n5182), .A2(n5185), .ZN(n5713) );
  AOI22_X1 U6373 ( .A1(n5331), .A2(DATAI_14_), .B1(n6332), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5186) );
  OAI21_X1 U6374 ( .B1(n5713), .B2(n5339), .A(n5186), .ZN(U2877) );
  INV_X1 U6375 ( .A(n5952), .ZN(n5189) );
  NAND2_X1 U6376 ( .A1(n5189), .A2(n6628), .ZN(n5190) );
  NAND2_X1 U6377 ( .A1(n5190), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5191) );
  NAND2_X1 U6378 ( .A1(n5191), .A2(n6564), .ZN(n5196) );
  NAND2_X1 U6379 ( .A1(n5192), .A2(n4582), .ZN(n6567) );
  NAND2_X1 U6380 ( .A1(n5193), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5965) );
  OAI22_X1 U6381 ( .A1(n5196), .A2(n6567), .B1(n5194), .B2(n5965), .ZN(n5949)
         );
  NAND3_X1 U6382 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6643), .ZN(n6574) );
  NOR2_X1 U6383 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6574), .ZN(n5951)
         );
  INV_X1 U6384 ( .A(n6567), .ZN(n5195) );
  OAI22_X1 U6385 ( .A1(n5196), .A2(n5195), .B1(n5951), .B2(n7152), .ZN(n5197)
         );
  INV_X1 U6386 ( .A(n5197), .ZN(n5198) );
  OAI211_X1 U6387 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6780), .A(n5199), .B(n5198), .ZN(n5950) );
  AOI22_X1 U6388 ( .A1(n6611), .A2(n5951), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5950), .ZN(n5201) );
  NAND2_X1 U6389 ( .A1(n5952), .A2(n6612), .ZN(n5200) );
  OAI211_X1 U6390 ( .C1(n6628), .C2(n6618), .A(n5201), .B(n5200), .ZN(n5202)
         );
  AOI21_X1 U6391 ( .B1(n5949), .B2(n6614), .A(n5202), .ZN(n5203) );
  INV_X1 U6392 ( .A(n5203), .ZN(U3106) );
  AOI22_X1 U6393 ( .A1(n6587), .A2(n5951), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5950), .ZN(n5205) );
  NAND2_X1 U6394 ( .A1(n5952), .A2(n6588), .ZN(n5204) );
  OAI211_X1 U6395 ( .C1(n6628), .C2(n6592), .A(n5205), .B(n5204), .ZN(n5206)
         );
  AOI21_X1 U6396 ( .B1(n5949), .B2(n6589), .A(n5206), .ZN(n5207) );
  INV_X1 U6397 ( .A(n5207), .ZN(U3102) );
  AOI22_X1 U6398 ( .A1(n6605), .A2(n5951), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5950), .ZN(n5209) );
  NAND2_X1 U6399 ( .A1(n5952), .A2(n6606), .ZN(n5208) );
  OAI211_X1 U6400 ( .C1(n6628), .C2(n6610), .A(n5209), .B(n5208), .ZN(n5210)
         );
  AOI21_X1 U6401 ( .B1(n5949), .B2(n6607), .A(n5210), .ZN(n5211) );
  INV_X1 U6402 ( .A(n5211), .ZN(U3105) );
  AOI22_X1 U6403 ( .A1(n6599), .A2(n5951), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5950), .ZN(n5213) );
  NAND2_X1 U6404 ( .A1(n5952), .A2(n6600), .ZN(n5212) );
  OAI211_X1 U6405 ( .C1(n6628), .C2(n6604), .A(n5213), .B(n5212), .ZN(n5214)
         );
  AOI21_X1 U6406 ( .B1(n5949), .B2(n6601), .A(n5214), .ZN(n5215) );
  INV_X1 U6407 ( .A(n5215), .ZN(U3104) );
  OR2_X1 U6408 ( .A1(n6777), .A2(n5216), .ZN(n5217) );
  NAND2_X1 U6409 ( .A1(n5217), .A2(n6278), .ZN(n6304) );
  INV_X1 U6410 ( .A(n6304), .ZN(n6321) );
  NOR2_X1 U6411 ( .A1(n6777), .A2(n5218), .ZN(n6293) );
  AOI22_X1 U6412 ( .A1(n6293), .A2(n5853), .B1(n4435), .B2(n5219), .ZN(n5221)
         );
  OAI21_X1 U6413 ( .B1(n6272), .B2(n6302), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5220) );
  OAI211_X1 U6414 ( .C1(n5222), .C2(n6246), .A(n5221), .B(n5220), .ZN(n5223)
         );
  AOI21_X1 U6415 ( .B1(REIP_REG_0__SCAN_IN), .B2(n6297), .A(n5223), .ZN(n5224)
         );
  OAI21_X1 U6416 ( .B1(n6321), .B2(n6445), .A(n5224), .ZN(U2827) );
  AOI22_X1 U6417 ( .A1(n6562), .A2(n5951), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5950), .ZN(n5226) );
  NAND2_X1 U6418 ( .A1(n5952), .A2(n6563), .ZN(n5225) );
  OAI211_X1 U6419 ( .C1(n6628), .C2(n6580), .A(n5226), .B(n5225), .ZN(n5227)
         );
  AOI21_X1 U6420 ( .B1(n5949), .B2(n6577), .A(n5227), .ZN(n5228) );
  INV_X1 U6421 ( .A(n5228), .ZN(U3100) );
  INV_X1 U6422 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5230) );
  OAI22_X1 U6423 ( .A1(n5230), .A2(n6246), .B1(n6318), .B2(n5229), .ZN(n5231)
         );
  NOR2_X1 U6424 ( .A1(n6425), .A2(n5231), .ZN(n5233) );
  AOI22_X1 U6425 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n6272), .B1(n6302), 
        .B2(n5284), .ZN(n5232) );
  OAI211_X1 U6426 ( .C1(n5235), .C2(n5234), .A(n5233), .B(n5232), .ZN(n5236)
         );
  AOI21_X1 U6427 ( .B1(REIP_REG_8__SCAN_IN), .B2(n6252), .A(n5236), .ZN(n5237)
         );
  OAI21_X1 U6428 ( .B1(n5281), .B2(n6278), .A(n5237), .ZN(U2819) );
  NAND2_X1 U6429 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n5239) );
  NAND2_X1 U6430 ( .A1(n6307), .A2(n6222), .ZN(n6223) );
  INV_X1 U6431 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5238) );
  OAI21_X1 U6432 ( .B1(n5239), .B2(n6223), .A(n5238), .ZN(n5249) );
  INV_X1 U6433 ( .A(n5341), .ZN(n5240) );
  NAND2_X1 U6434 ( .A1(n6296), .A2(n5240), .ZN(n6205) );
  NAND2_X1 U6435 ( .A1(n6297), .A2(n6205), .ZN(n5344) );
  INV_X1 U6436 ( .A(n5344), .ZN(n5248) );
  INV_X1 U6437 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5246) );
  INV_X1 U6438 ( .A(n5241), .ZN(n5710) );
  OAI21_X1 U6439 ( .B1(n5243), .B2(n5242), .A(n5334), .ZN(n5801) );
  OAI22_X1 U6440 ( .A1(n7149), .A2(n6314), .B1(n6318), .B2(n5801), .ZN(n5244)
         );
  AOI211_X1 U6441 ( .C1(n6302), .C2(n5710), .A(n5244), .B(n6425), .ZN(n5245)
         );
  OAI21_X1 U6442 ( .B1(n6246), .B2(n5246), .A(n5245), .ZN(n5247) );
  AOI21_X1 U6443 ( .B1(n5249), .B2(n5248), .A(n5247), .ZN(n5250) );
  OAI21_X1 U6444 ( .B1(n5713), .B2(n6278), .A(n5250), .ZN(U2813) );
  OAI21_X1 U6445 ( .B1(n5295), .B2(n5251), .A(n3967), .ZN(n5355) );
  INV_X1 U6446 ( .A(n5299), .ZN(n5252) );
  XNOR2_X1 U6447 ( .A(n5253), .B(n5252), .ZN(n6231) );
  AOI22_X1 U6448 ( .A1(n5557), .A2(n6231), .B1(n5556), .B2(EBX_REG_12__SCAN_IN), .ZN(n5254) );
  OAI21_X1 U6449 ( .B1(n5355), .B2(n5575), .A(n5254), .ZN(U2847) );
  INV_X1 U6450 ( .A(n5255), .ZN(n5272) );
  AOI22_X1 U6451 ( .A1(n5272), .A2(n6607), .B1(INSTQUEUE_REG_8__5__SCAN_IN), 
        .B2(n5271), .ZN(n5256) );
  OAI21_X1 U6452 ( .B1(n5992), .B2(n5274), .A(n5256), .ZN(n5257) );
  AOI21_X1 U6453 ( .B1(n6544), .B2(n5276), .A(n5257), .ZN(n5258) );
  OAI21_X1 U6454 ( .B1(n5887), .B2(n5278), .A(n5258), .ZN(U3089) );
  AOI22_X1 U6455 ( .A1(n5272), .A2(n6624), .B1(INSTQUEUE_REG_8__7__SCAN_IN), 
        .B2(n5271), .ZN(n5259) );
  OAI21_X1 U6456 ( .B1(n6005), .B2(n5274), .A(n5259), .ZN(n5260) );
  AOI21_X1 U6457 ( .B1(n6621), .B2(n5276), .A(n5260), .ZN(n5261) );
  OAI21_X1 U6458 ( .B1(n6629), .B2(n5278), .A(n5261), .ZN(U3091) );
  AOI22_X1 U6459 ( .A1(n5272), .A2(n6583), .B1(INSTQUEUE_REG_8__1__SCAN_IN), 
        .B2(n5271), .ZN(n5262) );
  OAI21_X1 U6460 ( .B1(n5973), .B2(n5274), .A(n5262), .ZN(n5263) );
  AOI21_X1 U6461 ( .B1(n6582), .B2(n5276), .A(n5263), .ZN(n5264) );
  OAI21_X1 U6462 ( .B1(n6586), .B2(n5278), .A(n5264), .ZN(U3085) );
  AOI22_X1 U6463 ( .A1(n5272), .A2(n6577), .B1(INSTQUEUE_REG_8__0__SCAN_IN), 
        .B2(n5271), .ZN(n5265) );
  OAI21_X1 U6464 ( .B1(n5969), .B2(n5274), .A(n5265), .ZN(n5266) );
  AOI21_X1 U6465 ( .B1(n6518), .B2(n5276), .A(n5266), .ZN(n5267) );
  OAI21_X1 U6466 ( .B1(n5865), .B2(n5278), .A(n5267), .ZN(U3084) );
  AOI22_X1 U6467 ( .A1(n5272), .A2(n6595), .B1(INSTQUEUE_REG_8__3__SCAN_IN), 
        .B2(n5271), .ZN(n5268) );
  OAI21_X1 U6468 ( .B1(n5983), .B2(n5274), .A(n5268), .ZN(n5269) );
  AOI21_X1 U6469 ( .B1(n6594), .B2(n5276), .A(n5269), .ZN(n5270) );
  OAI21_X1 U6470 ( .B1(n6598), .B2(n5278), .A(n5270), .ZN(U3087) );
  AOI22_X1 U6471 ( .A1(n5272), .A2(n6601), .B1(INSTQUEUE_REG_8__4__SCAN_IN), 
        .B2(n5271), .ZN(n5273) );
  OAI21_X1 U6472 ( .B1(n5988), .B2(n5274), .A(n5273), .ZN(n5275) );
  AOI21_X1 U6473 ( .B1(n6540), .B2(n5276), .A(n5275), .ZN(n5277) );
  OAI21_X1 U6474 ( .B1(n5882), .B2(n5278), .A(n5277), .ZN(U3088) );
  OAI222_X1 U6475 ( .A1(n5801), .A2(n5592), .B1(n5591), .B2(n5246), .C1(n5575), 
        .C2(n5713), .ZN(U2845) );
  INV_X1 U6476 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5280) );
  OAI21_X1 U6477 ( .B1(n5707), .B2(n5280), .A(n5279), .ZN(n5283) );
  NOR2_X1 U6478 ( .A1(n5281), .A2(n5714), .ZN(n5282) );
  AOI211_X1 U6479 ( .C1(n5709), .C2(n5284), .A(n5283), .B(n5282), .ZN(n5285)
         );
  OAI21_X1 U6480 ( .B1(n6438), .B2(n5286), .A(n5285), .ZN(U2978) );
  AOI21_X1 U6481 ( .B1(n5288), .B2(n5287), .A(n5298), .ZN(n6255) );
  INV_X1 U6482 ( .A(n6255), .ZN(n5304) );
  AOI22_X1 U6483 ( .A1(n5331), .A2(DATAI_10_), .B1(n6332), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5289) );
  OAI21_X1 U6484 ( .B1(n5304), .B2(n5339), .A(n5289), .ZN(U2881) );
  AOI22_X1 U6485 ( .A1(n6442), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6425), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5290) );
  OAI21_X1 U6486 ( .B1(n6437), .B2(n5291), .A(n5290), .ZN(n5292) );
  AOI21_X1 U6487 ( .B1(n6255), .B2(n6432), .A(n5292), .ZN(n5293) );
  OAI21_X1 U6488 ( .B1(n6438), .B2(n5294), .A(n5293), .ZN(U2976) );
  INV_X1 U6489 ( .A(n5295), .ZN(n5296) );
  OAI21_X1 U6490 ( .B1(n5298), .B2(n5297), .A(n5296), .ZN(n6241) );
  AOI21_X1 U6491 ( .B1(n5301), .B2(n5300), .A(n5299), .ZN(n6448) );
  AOI22_X1 U6492 ( .A1(n5557), .A2(n6448), .B1(n5556), .B2(EBX_REG_11__SCAN_IN), .ZN(n5302) );
  OAI21_X1 U6493 ( .B1(n6241), .B2(n5575), .A(n5302), .ZN(U2848) );
  INV_X1 U6494 ( .A(EAX_REG_12__SCAN_IN), .ZN(n7000) );
  OAI222_X1 U6495 ( .A1(n5338), .A2(n5303), .B1(n5593), .B2(n7000), .C1(n5339), 
        .C2(n5355), .ZN(U2879) );
  INV_X1 U6496 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5305) );
  OAI222_X1 U6497 ( .A1(n6248), .A2(n5592), .B1(n5305), .B2(n5591), .C1(n5575), 
        .C2(n5304), .ZN(U2849) );
  NAND2_X1 U6498 ( .A1(n5308), .A2(n5307), .ZN(n5309) );
  XNOR2_X1 U6499 ( .A(n5306), .B(n5309), .ZN(n6450) );
  NAND2_X1 U6500 ( .A1(n6450), .A2(n6431), .ZN(n5312) );
  NAND2_X1 U6501 ( .A1(n6425), .A2(REIP_REG_11__SCAN_IN), .ZN(n6446) );
  OAI21_X1 U6502 ( .B1(n5707), .B2(n3810), .A(n6446), .ZN(n5310) );
  AOI21_X1 U6503 ( .B1(n5709), .B2(n6243), .A(n5310), .ZN(n5311) );
  OAI211_X1 U6504 ( .C1(n5714), .C2(n6241), .A(n5312), .B(n5311), .ZN(U2975)
         );
  OAI22_X1 U6505 ( .A1(n6246), .A2(n6998), .B1(n6318), .B2(n5313), .ZN(n5315)
         );
  OAI22_X1 U6506 ( .A1(n6319), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6775), 
        .B2(n6296), .ZN(n5314) );
  AOI211_X1 U6507 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6272), .A(n5315), 
        .B(n5314), .ZN(n5319) );
  OR2_X1 U6508 ( .A1(n6262), .A2(REIP_REG_1__SCAN_IN), .ZN(n5321) );
  INV_X1 U6509 ( .A(n5321), .ZN(n5316) );
  AOI21_X1 U6510 ( .B1(n5317), .B2(n6293), .A(n5316), .ZN(n5318) );
  OAI211_X1 U6511 ( .C1(n6321), .C2(n5320), .A(n5319), .B(n5318), .ZN(U2826)
         );
  NAND2_X1 U6512 ( .A1(n6433), .A2(n6304), .ZN(n5328) );
  NAND2_X1 U6513 ( .A1(n5321), .A2(n6296), .ZN(n6312) );
  NAND3_X1 U6514 ( .A1(n6307), .A2(REIP_REG_1__SCAN_IN), .A3(n6693), .ZN(n5323) );
  NAND2_X1 U6515 ( .A1(n6272), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5322)
         );
  OAI211_X1 U6516 ( .C1(n6319), .C2(n6436), .A(n5323), .B(n5322), .ZN(n5326)
         );
  INV_X1 U6517 ( .A(n6293), .ZN(n6316) );
  OAI22_X1 U6518 ( .A1(n6316), .A2(n4622), .B1(n6246), .B2(n5324), .ZN(n5325)
         );
  AOI211_X1 U6519 ( .C1(REIP_REG_2__SCAN_IN), .C2(n6312), .A(n5326), .B(n5325), 
        .ZN(n5327) );
  OAI211_X1 U6520 ( .C1(n6484), .C2(n6318), .A(n5328), .B(n5327), .ZN(U2825)
         );
  NAND2_X1 U6521 ( .A1(n5182), .A2(n5329), .ZN(n5330) );
  AND2_X1 U6522 ( .A1(n5366), .A2(n5330), .ZN(n5702) );
  AOI22_X1 U6523 ( .A1(n5331), .A2(DATAI_15_), .B1(n6332), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5332) );
  OAI21_X1 U6524 ( .B1(n5348), .B2(n5339), .A(n5332), .ZN(U2876) );
  AOI21_X1 U6525 ( .B1(n5335), .B2(n5334), .A(n5333), .ZN(n6147) );
  AOI22_X1 U6526 ( .A1(n5557), .A2(n6147), .B1(n5556), .B2(EBX_REG_15__SCAN_IN), .ZN(n5336) );
  OAI21_X1 U6527 ( .B1(n5348), .B2(n5575), .A(n5336), .ZN(U2844) );
  INV_X1 U6528 ( .A(DATAI_11_), .ZN(n5337) );
  INV_X1 U6529 ( .A(EAX_REG_11__SCAN_IN), .ZN(n7157) );
  OAI222_X1 U6530 ( .A1(n6241), .A2(n5339), .B1(n5338), .B2(n5337), .C1(n5593), 
        .C2(n7157), .ZN(U2880) );
  OAI22_X1 U6531 ( .A1(n6319), .A2(n5700), .B1(n6246), .B2(n5340), .ZN(n5346)
         );
  NOR3_X1 U6532 ( .A1(n6262), .A2(REIP_REG_15__SCAN_IN), .A3(n5341), .ZN(n5342) );
  AOI211_X1 U6533 ( .C1(n6272), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6425), 
        .B(n5342), .ZN(n5343) );
  OAI21_X1 U6534 ( .B1(n6709), .B2(n5344), .A(n5343), .ZN(n5345) );
  AOI211_X1 U6535 ( .C1(n6147), .C2(n4435), .A(n5346), .B(n5345), .ZN(n5347)
         );
  OAI21_X1 U6536 ( .B1(n5348), .B2(n6278), .A(n5347), .ZN(U2812) );
  INV_X1 U6537 ( .A(n5350), .ZN(n5351) );
  NOR2_X1 U6538 ( .A1(n5352), .A2(n5351), .ZN(n5353) );
  XNOR2_X1 U6539 ( .A(n5349), .B(n5353), .ZN(n5364) );
  AND2_X1 U6540 ( .A1(n6425), .A2(REIP_REG_12__SCAN_IN), .ZN(n5358) );
  AND2_X1 U6541 ( .A1(n6442), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5354)
         );
  AOI211_X1 U6542 ( .C1(n5709), .C2(n6232), .A(n5358), .B(n5354), .ZN(n5357)
         );
  INV_X1 U6543 ( .A(n5355), .ZN(n6233) );
  NAND2_X1 U6544 ( .A1(n6233), .A2(n6432), .ZN(n5356) );
  OAI211_X1 U6545 ( .C1(n5364), .C2(n6438), .A(n5357), .B(n5356), .ZN(U2974)
         );
  AOI21_X1 U6546 ( .B1(n6503), .B2(n6231), .A(n5358), .ZN(n5363) );
  NOR2_X1 U6547 ( .A1(n6488), .A2(n5359), .ZN(n5767) );
  INV_X1 U6548 ( .A(n5795), .ZN(n6453) );
  OAI21_X1 U6549 ( .B1(n5798), .B2(n5767), .A(n6453), .ZN(n5361) );
  OAI21_X1 U6550 ( .B1(n6161), .B2(n7122), .A(n4352), .ZN(n5360) );
  NAND2_X1 U6551 ( .A1(n5361), .A2(n5360), .ZN(n5362) );
  OAI211_X1 U6552 ( .C1(n5364), .C2(n6475), .A(n5363), .B(n5362), .ZN(U3006)
         );
  INV_X1 U6553 ( .A(n5376), .ZN(n5368) );
  NAND2_X1 U6554 ( .A1(n5366), .A2(n5365), .ZN(n5367) );
  NAND2_X1 U6555 ( .A1(n5368), .A2(n5367), .ZN(n6210) );
  NOR2_X2 U6556 ( .A1(n6332), .A2(n5369), .ZN(n6329) );
  AOI22_X1 U6557 ( .A1(n6329), .A2(DATAI_16_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n6332), .ZN(n5372) );
  NOR2_X1 U6558 ( .A1(n5594), .A2(n3448), .ZN(n5370) );
  NAND2_X1 U6559 ( .A1(n6333), .A2(DATAI_0_), .ZN(n5371) );
  OAI211_X1 U6560 ( .C1(n6210), .C2(n5339), .A(n5372), .B(n5371), .ZN(U2875)
         );
  OAI21_X1 U6561 ( .B1(n5373), .B2(n5333), .A(n5378), .ZN(n6209) );
  INV_X1 U6562 ( .A(EBX_REG_16__SCAN_IN), .ZN(n6215) );
  OAI222_X1 U6563 ( .A1(n6209), .A2(n5592), .B1(n5591), .B2(n6215), .C1(n5575), 
        .C2(n6210), .ZN(U2843) );
  OR2_X1 U6564 ( .A1(n5376), .A2(n5375), .ZN(n5377) );
  AND2_X1 U6565 ( .A1(n5374), .A2(n5377), .ZN(n6331) );
  INV_X1 U6566 ( .A(n6331), .ZN(n5382) );
  NAND2_X1 U6567 ( .A1(n5379), .A2(n5378), .ZN(n5380) );
  AND2_X1 U6568 ( .A1(n5401), .A2(n5380), .ZN(n6201) );
  AOI22_X1 U6569 ( .A1(n5557), .A2(n6201), .B1(n5556), .B2(EBX_REG_17__SCAN_IN), .ZN(n5381) );
  OAI21_X1 U6570 ( .B1(n5382), .B2(n5575), .A(n5381), .ZN(U2842) );
  OAI21_X1 U6571 ( .B1(n5383), .B2(n5385), .A(n5384), .ZN(n6157) );
  NAND2_X1 U6572 ( .A1(n6157), .A2(n6431), .ZN(n5389) );
  INV_X1 U6573 ( .A(REIP_REG_13__SCAN_IN), .ZN(n5386) );
  NOR2_X1 U6574 ( .A1(n6498), .A2(n5386), .ZN(n6155) );
  NOR2_X1 U6575 ( .A1(n6437), .A2(n6219), .ZN(n5387) );
  AOI211_X1 U6576 ( .C1(n6442), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6155), 
        .B(n5387), .ZN(n5388) );
  OAI211_X1 U6577 ( .C1(n6218), .C2(n5714), .A(n5389), .B(n5388), .ZN(U2973)
         );
  INV_X1 U6578 ( .A(n5406), .ZN(n5390) );
  AOI21_X1 U6579 ( .B1(n5391), .B2(n5374), .A(n5390), .ZN(n5690) );
  INV_X1 U6580 ( .A(n5690), .ZN(n6192) );
  AOI22_X1 U6581 ( .A1(n6329), .A2(DATAI_18_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n6332), .ZN(n5393) );
  NAND2_X1 U6582 ( .A1(n6333), .A2(DATAI_2_), .ZN(n5392) );
  OAI211_X1 U6583 ( .C1(n6192), .C2(n5339), .A(n5393), .B(n5392), .ZN(U2873)
         );
  INV_X1 U6584 ( .A(n5401), .ZN(n5399) );
  OR2_X1 U6585 ( .A1(n5587), .A2(n5395), .ZN(n5398) );
  INV_X1 U6586 ( .A(n5394), .ZN(n5396) );
  NAND2_X1 U6587 ( .A1(n5396), .A2(n5395), .ZN(n5397) );
  NAND2_X1 U6588 ( .A1(n5398), .A2(n5397), .ZN(n5400) );
  NAND2_X1 U6589 ( .A1(n5399), .A2(n5400), .ZN(n5410) );
  INV_X1 U6590 ( .A(n5400), .ZN(n5402) );
  NAND2_X1 U6591 ( .A1(n5402), .A2(n5401), .ZN(n5403) );
  NAND2_X1 U6592 ( .A1(n5410), .A2(n5403), .ZN(n6196) );
  INV_X1 U6593 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5404) );
  OAI222_X1 U6594 ( .A1(n6196), .A2(n5592), .B1(n5591), .B2(n5404), .C1(n5575), 
        .C2(n6192), .ZN(U2841) );
  AND2_X1 U6595 ( .A1(n5406), .A2(n5405), .ZN(n5408) );
  OR2_X1 U6596 ( .A1(n5408), .A2(n5407), .ZN(n6110) );
  XNOR2_X1 U6597 ( .A(n5410), .B(n5409), .ZN(n6096) );
  INV_X1 U6598 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5411) );
  OAI222_X1 U6599 ( .A1(n6110), .A2(n5575), .B1(n5592), .B2(n6096), .C1(n5411), 
        .C2(n5591), .ZN(U2840) );
  AOI22_X1 U6600 ( .A1(n5415), .A2(EAX_REG_31__SCAN_IN), .B1(n5414), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5416) );
  INV_X1 U6601 ( .A(n5416), .ZN(n5417) );
  INV_X1 U6602 ( .A(n5595), .ZN(n5426) );
  INV_X1 U6603 ( .A(n6656), .ZN(n5419) );
  NAND3_X1 U6604 ( .A1(n6782), .A2(EBX_REG_31__SCAN_IN), .A3(n5419), .ZN(n5420) );
  OAI22_X1 U6605 ( .A1(n6314), .A2(n5421), .B1(n6777), .B2(n5420), .ZN(n5423)
         );
  INV_X1 U6606 ( .A(REIP_REG_30__SCAN_IN), .ZN(n5507) );
  NOR4_X1 U6607 ( .A1(n5508), .A2(REIP_REG_31__SCAN_IN), .A3(n5507), .A4(n7134), .ZN(n5422) );
  AOI211_X1 U6608 ( .C1(n5529), .C2(n4435), .A(n5423), .B(n5422), .ZN(n5425)
         );
  OAI211_X1 U6609 ( .C1(REIP_REG_29__SCAN_IN), .C2(n6262), .A(n6011), .B(
        REIP_REG_30__SCAN_IN), .ZN(n5513) );
  NAND3_X1 U6610 ( .A1(n5513), .A2(REIP_REG_31__SCAN_IN), .A3(n6297), .ZN(
        n5424) );
  OAI211_X1 U6611 ( .C1(n5426), .C2(n6278), .A(n5425), .B(n5424), .ZN(U2796)
         );
  XNOR2_X1 U6612 ( .A(n3184), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5766)
         );
  INV_X1 U6613 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5770) );
  NAND2_X1 U6614 ( .A1(n5765), .A2(n5427), .ZN(n5676) );
  NAND2_X1 U6615 ( .A1(n5431), .A2(n5430), .ZN(n5671) );
  XNOR2_X1 U6616 ( .A(n3184), .B(n5756), .ZN(n5672) );
  NAND2_X1 U6617 ( .A1(n3184), .A2(n5756), .ZN(n5432) );
  INV_X1 U6618 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n7098) );
  MUX2_X1 U6619 ( .A(n7098), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .S(n3184), 
        .Z(n5434) );
  NAND3_X1 U6620 ( .A1(n5436), .A2(n5435), .A3(n5434), .ZN(n5437) );
  XNOR2_X1 U6621 ( .A(n5437), .B(n5444), .ZN(n5453) );
  OR2_X1 U6622 ( .A1(n5566), .A2(n5438), .ZN(n5439) );
  NAND2_X1 U6623 ( .A1(n5519), .A2(n5439), .ZN(n6049) );
  INV_X1 U6624 ( .A(n6049), .ZN(n5558) );
  AND2_X1 U6625 ( .A1(n6425), .A2(REIP_REG_24__SCAN_IN), .ZN(n5449) );
  NOR2_X1 U6626 ( .A1(n5441), .A2(n5440), .ZN(n5757) );
  INV_X1 U6627 ( .A(n5750), .ZN(n5442) );
  NAND2_X1 U6628 ( .A1(n5757), .A2(n5442), .ZN(n5741) );
  AOI211_X1 U6629 ( .C1(n5444), .C2(n5741), .A(n5443), .B(n6131), .ZN(n5445)
         );
  AOI211_X1 U6630 ( .C1(n6503), .C2(n5558), .A(n5449), .B(n5445), .ZN(n5446)
         );
  OAI21_X1 U6631 ( .B1(n5453), .B2(n6475), .A(n5446), .ZN(U2994) );
  AOI21_X1 U6632 ( .B1(n5448), .B2(n5561), .A(n5447), .ZN(n6039) );
  AOI21_X1 U6633 ( .B1(n6442), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5449), 
        .ZN(n5450) );
  OAI21_X1 U6634 ( .B1(n6437), .B2(n6040), .A(n5450), .ZN(n5451) );
  AOI21_X1 U6635 ( .B1(n6039), .B2(n6432), .A(n5451), .ZN(n5452) );
  OAI21_X1 U6636 ( .B1(n5453), .B2(n6438), .A(n5452), .ZN(U2962) );
  AOI21_X1 U6637 ( .B1(n6442), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5454), 
        .ZN(n5455) );
  OAI21_X1 U6638 ( .B1(n6437), .B2(n5456), .A(n5455), .ZN(n5457) );
  AOI21_X1 U6639 ( .B1(n5595), .B2(n6432), .A(n5457), .ZN(n5458) );
  OAI21_X1 U6640 ( .B1(n5459), .B2(n6438), .A(n5458), .ZN(U2955) );
  INV_X1 U6641 ( .A(n5462), .ZN(n5460) );
  OAI21_X1 U6642 ( .B1(n5461), .B2(n4403), .A(n5460), .ZN(n5465) );
  INV_X1 U6643 ( .A(n5461), .ZN(n5463) );
  OAI211_X1 U6644 ( .C1(n4404), .C2(n4406), .A(n5463), .B(n5462), .ZN(n5464)
         );
  INV_X1 U6645 ( .A(n5532), .ZN(n5470) );
  INV_X1 U6646 ( .A(n5467), .ZN(n5469) );
  INV_X1 U6647 ( .A(n5472), .ZN(n5717) );
  NOR4_X1 U6648 ( .A1(n5716), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5487), 
        .A4(n5717), .ZN(n5468) );
  AOI211_X1 U6649 ( .C1(n5470), .C2(n6503), .A(n5469), .B(n5468), .ZN(n5474)
         );
  INV_X1 U6650 ( .A(n6131), .ZN(n5738) );
  INV_X1 U6651 ( .A(n5729), .ZN(n5471) );
  OAI211_X1 U6652 ( .C1(n5781), .C2(n5472), .A(n5471), .B(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5490) );
  OAI211_X1 U6653 ( .C1(n5738), .C2(n6501), .A(n5490), .B(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5473) );
  OAI211_X1 U6654 ( .C1(n5475), .C2(n6475), .A(n5474), .B(n5473), .ZN(U2988)
         );
  INV_X1 U6655 ( .A(n5808), .ZN(n6657) );
  INV_X1 U6656 ( .A(n4588), .ZN(n5478) );
  OAI22_X1 U6657 ( .A1(n5476), .A2(n6662), .B1(n6673), .B2(n6173), .ZN(n6163)
         );
  NOR2_X1 U6658 ( .A1(n6163), .A2(n6745), .ZN(n5811) );
  AOI21_X1 U6659 ( .B1(n6657), .B2(n5478), .A(n5811), .ZN(n5483) );
  INV_X1 U6660 ( .A(n5477), .ZN(n5481) );
  INV_X1 U6661 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n7025) );
  INV_X1 U6662 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6510) );
  AOI22_X1 U6663 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4442), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6510), .ZN(n5497) );
  NOR3_X1 U6664 ( .A1(n6749), .A2(n7025), .A3(n5497), .ZN(n5480) );
  NOR3_X1 U6665 ( .A1(n5808), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n5478), 
        .ZN(n5479) );
  AOI211_X1 U6666 ( .C1(n5481), .C2(n6665), .A(n5480), .B(n5479), .ZN(n5482)
         );
  OAI22_X1 U6667 ( .A1(n5483), .A2(n3332), .B1(n5811), .B2(n5482), .ZN(U3459)
         );
  AND2_X1 U6668 ( .A1(n3737), .A2(n5484), .ZN(n5485) );
  XNOR2_X1 U6669 ( .A(n5486), .B(n5487), .ZN(n5630) );
  OAI21_X1 U6670 ( .B1(n5716), .B2(n5717), .A(n5487), .ZN(n5489) );
  NOR2_X1 U6671 ( .A1(n5534), .A2(n5783), .ZN(n5488) );
  AND2_X1 U6672 ( .A1(n6425), .A2(REIP_REG_29__SCAN_IN), .ZN(n5624) );
  OAI21_X1 U6673 ( .B1(n5630), .B2(n6475), .A(n5491), .ZN(U2989) );
  NOR3_X1 U6674 ( .A1(n6630), .A2(n3224), .A3(n4588), .ZN(n5492) );
  AOI21_X1 U6675 ( .B1(n6632), .B2(n3207), .A(n5492), .ZN(n5493) );
  OAI21_X1 U6676 ( .B1(n5494), .B2(n6631), .A(n5493), .ZN(n6636) );
  NOR2_X1 U6677 ( .A1(n6749), .A2(n7025), .ZN(n5496) );
  AOI222_X1 U6678 ( .A1(n6636), .A2(n6665), .B1(n5497), .B2(n5496), .C1(n5495), 
        .C2(n6657), .ZN(n5500) );
  INV_X1 U6679 ( .A(n5811), .ZN(n6753) );
  OAI21_X1 U6680 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5808), .A(n6753), 
        .ZN(n6751) );
  INV_X1 U6681 ( .A(n6751), .ZN(n5498) );
  OAI22_X1 U6682 ( .A1(n5811), .A2(n5500), .B1(n3207), .B2(n5498), .ZN(U3460)
         );
  NAND2_X1 U6683 ( .A1(MEMORYFETCH_REG_SCAN_IN), .A2(n5501), .ZN(n5504) );
  INV_X1 U6684 ( .A(n5502), .ZN(n5503) );
  NAND3_X1 U6685 ( .A1(n5505), .A2(n5504), .A3(n5503), .ZN(U2788) );
  OAI21_X1 U6686 ( .B1(n5508), .B2(n7134), .A(n5507), .ZN(n5512) );
  AOI22_X1 U6687 ( .A1(n5509), .A2(n6302), .B1(n6272), .B2(
        PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5511) );
  NAND2_X1 U6688 ( .A1(n6325), .A2(EBX_REG_30__SCAN_IN), .ZN(n5510) );
  NOR2_X1 U6689 ( .A1(n5447), .A2(n5515), .ZN(n5516) );
  OR2_X1 U6690 ( .A1(n5514), .A2(n5516), .ZN(n5612) );
  INV_X1 U6691 ( .A(n5612), .ZN(n6106) );
  INV_X1 U6692 ( .A(n5521), .ZN(n5517) );
  NAND2_X1 U6693 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5517), .ZN(n6031) );
  OAI22_X1 U6694 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6031), .B1(n6109), .B2(
        n6319), .ZN(n5527) );
  NAND2_X1 U6695 ( .A1(n5519), .A2(n5518), .ZN(n5520) );
  NAND2_X1 U6696 ( .A1(n5550), .A2(n5520), .ZN(n6125) );
  NOR2_X1 U6697 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5521), .ZN(n6046) );
  INV_X1 U6698 ( .A(n6045), .ZN(n6055) );
  OAI21_X1 U6699 ( .B1(n6046), .B2(n6055), .A(REIP_REG_25__SCAN_IN), .ZN(n5525) );
  INV_X1 U6700 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5522) );
  INV_X1 U6701 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n7081) );
  OAI22_X1 U6702 ( .A1(n5522), .A2(n6246), .B1(n7081), .B2(n6314), .ZN(n5523)
         );
  INV_X1 U6703 ( .A(n5523), .ZN(n5524) );
  OAI211_X1 U6704 ( .C1(n6125), .C2(n6318), .A(n5525), .B(n5524), .ZN(n5526)
         );
  AOI211_X1 U6705 ( .C1(n6106), .C2(n6254), .A(n5527), .B(n5526), .ZN(n5528)
         );
  INV_X1 U6706 ( .A(n5528), .ZN(U2802) );
  INV_X1 U6707 ( .A(n5529), .ZN(n5531) );
  OAI22_X1 U6708 ( .A1(n5531), .A2(n5592), .B1(n5530), .B2(n5591), .ZN(U2828)
         );
  INV_X1 U6709 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5533) );
  OAI222_X1 U6710 ( .A1(n5575), .A2(n5506), .B1(n5591), .B2(n5533), .C1(n5532), 
        .C2(n5592), .ZN(U2829) );
  OAI222_X1 U6711 ( .A1(n5575), .A2(n5623), .B1(n5591), .B2(n5535), .C1(n5534), 
        .C2(n5592), .ZN(U2830) );
  NAND2_X1 U6712 ( .A1(n5543), .A2(n5536), .ZN(n5537) );
  OR2_X1 U6713 ( .A1(n5547), .A2(n5538), .ZN(n5539) );
  NAND2_X1 U6714 ( .A1(n4403), .A2(n5539), .ZN(n6019) );
  INV_X1 U6715 ( .A(EBX_REG_28__SCAN_IN), .ZN(n7058) );
  OAI22_X1 U6716 ( .A1(n6019), .A2(n5592), .B1(n7058), .B2(n5591), .ZN(n5540)
         );
  INV_X1 U6717 ( .A(n5540), .ZN(n5541) );
  OAI21_X1 U6718 ( .B1(n5604), .B2(n5575), .A(n5541), .ZN(U2831) );
  OR2_X1 U6719 ( .A1(n5553), .A2(n5542), .ZN(n5544) );
  NOR2_X1 U6720 ( .A1(n5551), .A2(n5545), .ZN(n5546) );
  OR2_X1 U6721 ( .A1(n5547), .A2(n5546), .ZN(n6025) );
  OAI222_X1 U6722 ( .A1(n5575), .A2(n5607), .B1(n5591), .B2(n5548), .C1(n6025), 
        .C2(n5592), .ZN(U2832) );
  AND2_X1 U6723 ( .A1(n5550), .A2(n5549), .ZN(n5552) );
  OR2_X1 U6724 ( .A1(n5552), .A2(n5551), .ZN(n6032) );
  INV_X1 U6725 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6945) );
  INV_X1 U6726 ( .A(n5553), .ZN(n5554) );
  OAI21_X1 U6727 ( .B1(n5555), .B2(n5514), .A(n5554), .ZN(n6033) );
  OAI222_X1 U6728 ( .A1(n6032), .A2(n5592), .B1(n5591), .B2(n6945), .C1(n5575), 
        .C2(n6033), .ZN(U2833) );
  OAI222_X1 U6729 ( .A1(n5612), .A2(n5575), .B1(n5591), .B2(n5522), .C1(n6125), 
        .C2(n5592), .ZN(U2834) );
  INV_X1 U6730 ( .A(n6039), .ZN(n5615) );
  AOI22_X1 U6731 ( .A1(n5558), .A2(n5557), .B1(n5556), .B2(EBX_REG_24__SCAN_IN), .ZN(n5559) );
  OAI21_X1 U6732 ( .B1(n5615), .B2(n5575), .A(n5559), .ZN(U2835) );
  INV_X1 U6733 ( .A(n5561), .ZN(n5562) );
  AOI21_X1 U6734 ( .B1(n5563), .B2(n5574), .A(n5562), .ZN(n6054) );
  INV_X1 U6735 ( .A(n6054), .ZN(n5618) );
  NOR2_X1 U6736 ( .A1(n5569), .A2(n5564), .ZN(n5565) );
  OR2_X1 U6737 ( .A1(n5566), .A2(n5565), .ZN(n6052) );
  OAI222_X1 U6738 ( .A1(n5575), .A2(n5618), .B1(n5591), .B2(n5567), .C1(n6052), 
        .C2(n5592), .ZN(U2836) );
  AND2_X1 U6739 ( .A1(n3238), .A2(n5568), .ZN(n5570) );
  OR2_X1 U6740 ( .A1(n5570), .A2(n5569), .ZN(n6069) );
  INV_X1 U6741 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U6742 ( .A1(n5571), .A2(n5572), .ZN(n5573) );
  NAND2_X1 U6743 ( .A1(n5574), .A2(n5573), .ZN(n6066) );
  OAI222_X1 U6744 ( .A1(n6069), .A2(n5592), .B1(n5591), .B2(n5576), .C1(n5575), 
        .C2(n6066), .ZN(U2837) );
  OR2_X1 U6745 ( .A1(n5577), .A2(n5578), .ZN(n5579) );
  AND2_X1 U6746 ( .A1(n5571), .A2(n5579), .ZN(n6097) );
  INV_X1 U6747 ( .A(n6097), .ZN(n5583) );
  INV_X1 U6748 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5582) );
  XNOR2_X1 U6749 ( .A(n5581), .B(n5580), .ZN(n6079) );
  OAI222_X1 U6750 ( .A1(n5583), .A2(n5575), .B1(n5591), .B2(n5582), .C1(n6079), 
        .C2(n5592), .ZN(U2838) );
  INV_X1 U6751 ( .A(n5577), .ZN(n5584) );
  OAI21_X1 U6752 ( .B1(n5585), .B2(n5407), .A(n5584), .ZN(n6082) );
  MUX2_X1 U6753 ( .A(n4406), .B(n5587), .S(n5586), .Z(n5589) );
  XNOR2_X1 U6754 ( .A(n5589), .B(n5588), .ZN(n6136) );
  INV_X1 U6755 ( .A(n6136), .ZN(n6081) );
  INV_X1 U6756 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5590) );
  OAI222_X1 U6757 ( .A1(n6082), .A2(n5575), .B1(n5592), .B2(n6081), .C1(n5591), 
        .C2(n5590), .ZN(U2839) );
  NAND3_X1 U6758 ( .A1(n5595), .A2(n5594), .A3(n5593), .ZN(n5597) );
  AOI22_X1 U6759 ( .A1(n6329), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6332), .ZN(n5596) );
  NAND2_X1 U6760 ( .A1(n5597), .A2(n5596), .ZN(U2860) );
  AOI22_X1 U6761 ( .A1(n6329), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6332), .ZN(n5599) );
  NAND2_X1 U6762 ( .A1(n6333), .A2(DATAI_14_), .ZN(n5598) );
  OAI211_X1 U6763 ( .C1(n5506), .C2(n5339), .A(n5599), .B(n5598), .ZN(U2861)
         );
  AOI22_X1 U6764 ( .A1(n6333), .A2(DATAI_13_), .B1(n6332), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5601) );
  NAND2_X1 U6765 ( .A1(n6329), .A2(DATAI_29_), .ZN(n5600) );
  OAI211_X1 U6766 ( .C1(n5623), .C2(n5339), .A(n5601), .B(n5600), .ZN(U2862)
         );
  AOI22_X1 U6767 ( .A1(n6333), .A2(DATAI_12_), .B1(n6332), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U6768 ( .A1(n6329), .A2(DATAI_28_), .ZN(n5602) );
  OAI211_X1 U6769 ( .C1(n5604), .C2(n5339), .A(n5603), .B(n5602), .ZN(U2863)
         );
  AOI22_X1 U6770 ( .A1(n6333), .A2(DATAI_11_), .B1(n6332), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U6771 ( .A1(n6329), .A2(DATAI_27_), .ZN(n5605) );
  OAI211_X1 U6772 ( .C1(n5607), .C2(n5339), .A(n5606), .B(n5605), .ZN(U2864)
         );
  AOI22_X1 U6773 ( .A1(n6333), .A2(DATAI_10_), .B1(n6332), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U6774 ( .A1(n6329), .A2(DATAI_26_), .ZN(n5608) );
  OAI211_X1 U6775 ( .C1(n6033), .C2(n5339), .A(n5609), .B(n5608), .ZN(U2865)
         );
  AOI22_X1 U6776 ( .A1(n6329), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n6332), .ZN(n5611) );
  NAND2_X1 U6777 ( .A1(n6333), .A2(DATAI_9_), .ZN(n5610) );
  OAI211_X1 U6778 ( .C1(n5612), .C2(n5339), .A(n5611), .B(n5610), .ZN(U2866)
         );
  AOI22_X1 U6779 ( .A1(n6333), .A2(DATAI_8_), .B1(n6332), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5614) );
  NAND2_X1 U6780 ( .A1(n6329), .A2(DATAI_24_), .ZN(n5613) );
  OAI211_X1 U6781 ( .C1(n5615), .C2(n5339), .A(n5614), .B(n5613), .ZN(U2867)
         );
  AOI22_X1 U6782 ( .A1(n6333), .A2(DATAI_7_), .B1(n6332), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U6783 ( .A1(n6329), .A2(DATAI_23_), .ZN(n5616) );
  OAI211_X1 U6784 ( .C1(n5618), .C2(n5339), .A(n5617), .B(n5616), .ZN(U2868)
         );
  AOI22_X1 U6785 ( .A1(n6333), .A2(DATAI_6_), .B1(n6332), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5620) );
  NAND2_X1 U6786 ( .A1(n6329), .A2(DATAI_22_), .ZN(n5619) );
  OAI211_X1 U6787 ( .C1(n6066), .C2(n5339), .A(n5620), .B(n5619), .ZN(U2869)
         );
  AOI22_X1 U6788 ( .A1(n6333), .A2(DATAI_4_), .B1(n6332), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5622) );
  NAND2_X1 U6789 ( .A1(n6329), .A2(DATAI_20_), .ZN(n5621) );
  OAI211_X1 U6790 ( .C1(n6082), .C2(n5339), .A(n5622), .B(n5621), .ZN(U2871)
         );
  INV_X1 U6791 ( .A(n5623), .ZN(n5628) );
  AOI21_X1 U6792 ( .B1(n6442), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5624), 
        .ZN(n5625) );
  OAI21_X1 U6793 ( .B1(n6437), .B2(n5626), .A(n5625), .ZN(n5627) );
  AOI21_X1 U6794 ( .B1(n5628), .B2(n6432), .A(n5627), .ZN(n5629) );
  OAI21_X1 U6795 ( .B1(n5630), .B2(n6438), .A(n5629), .ZN(U2957) );
  NOR3_X1 U6796 ( .A1(n3737), .A2(n5663), .A3(n5725), .ZN(n5633) );
  OR2_X1 U6797 ( .A1(n5647), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5632)
         );
  NOR2_X1 U6798 ( .A1(n5631), .A2(n5632), .ZN(n5641) );
  OAI22_X1 U6799 ( .A1(n5633), .A2(n5641), .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n5725), .ZN(n5635) );
  XNOR2_X1 U6800 ( .A(n5635), .B(n5634), .ZN(n5723) );
  INV_X1 U6801 ( .A(n6012), .ZN(n5637) );
  AND2_X1 U6802 ( .A1(n6425), .A2(REIP_REG_28__SCAN_IN), .ZN(n5715) );
  AOI21_X1 U6803 ( .B1(n6442), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5715), 
        .ZN(n5636) );
  OAI21_X1 U6804 ( .B1(n6437), .B2(n5637), .A(n5636), .ZN(n5638) );
  AOI21_X1 U6805 ( .B1(n6016), .B2(n6432), .A(n5638), .ZN(n5639) );
  OAI21_X1 U6806 ( .B1(n6438), .B2(n5723), .A(n5639), .ZN(U2958) );
  NOR2_X1 U6807 ( .A1(n5640), .A2(n5641), .ZN(n5642) );
  XNOR2_X1 U6808 ( .A(n5642), .B(n5725), .ZN(n5731) );
  AND2_X1 U6809 ( .A1(n6425), .A2(REIP_REG_27__SCAN_IN), .ZN(n5724) );
  AOI21_X1 U6810 ( .B1(n6442), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5724), 
        .ZN(n5643) );
  OAI21_X1 U6811 ( .B1(n6437), .B2(n6021), .A(n5643), .ZN(n5644) );
  AOI21_X1 U6812 ( .B1(n6027), .B2(n6432), .A(n5644), .ZN(n5645) );
  OAI21_X1 U6813 ( .B1(n5731), .B2(n6438), .A(n5645), .ZN(U2959) );
  NAND2_X1 U6814 ( .A1(n5647), .A2(n5646), .ZN(n5648) );
  XOR2_X1 U6815 ( .A(n5648), .B(n3737), .Z(n5740) );
  INV_X1 U6816 ( .A(n6033), .ZN(n5652) );
  INV_X1 U6817 ( .A(n6030), .ZN(n5650) );
  AND2_X1 U6818 ( .A1(n6425), .A2(REIP_REG_26__SCAN_IN), .ZN(n5734) );
  AOI21_X1 U6819 ( .B1(n6442), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5734), 
        .ZN(n5649) );
  OAI21_X1 U6820 ( .B1(n6437), .B2(n5650), .A(n5649), .ZN(n5651) );
  AOI21_X1 U6821 ( .B1(n5652), .B2(n6432), .A(n5651), .ZN(n5653) );
  OAI21_X1 U6822 ( .B1(n5740), .B2(n6438), .A(n5653), .ZN(U2960) );
  NAND2_X1 U6823 ( .A1(n5663), .A2(n7098), .ZN(n5662) );
  NAND2_X1 U6824 ( .A1(n3184), .A2(n5656), .ZN(n5657) );
  OAI22_X1 U6825 ( .A1(n5654), .A2(n5662), .B1(n5655), .B2(n5657), .ZN(n5658)
         );
  XNOR2_X1 U6826 ( .A(n5658), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5747)
         );
  NAND2_X1 U6827 ( .A1(n6425), .A2(REIP_REG_23__SCAN_IN), .ZN(n5742) );
  NAND2_X1 U6828 ( .A1(n6442), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5659)
         );
  OAI211_X1 U6829 ( .C1(n6437), .C2(n6050), .A(n5742), .B(n5659), .ZN(n5660)
         );
  AOI21_X1 U6830 ( .B1(n6054), .B2(n6432), .A(n5660), .ZN(n5661) );
  OAI21_X1 U6831 ( .B1(n5747), .B2(n6438), .A(n5661), .ZN(U2963) );
  OAI21_X1 U6832 ( .B1(n5663), .B2(n7098), .A(n5662), .ZN(n5664) );
  XNOR2_X1 U6833 ( .A(n5665), .B(n5664), .ZN(n5755) );
  NAND2_X1 U6834 ( .A1(n6425), .A2(REIP_REG_22__SCAN_IN), .ZN(n5751) );
  OAI21_X1 U6835 ( .B1(n5707), .B2(n5666), .A(n5751), .ZN(n5668) );
  NOR2_X1 U6836 ( .A1(n6066), .A2(n5714), .ZN(n5667) );
  AOI211_X1 U6837 ( .C1(n5709), .C2(n6061), .A(n5668), .B(n5667), .ZN(n5669)
         );
  OAI21_X1 U6838 ( .B1(n5755), .B2(n6438), .A(n5669), .ZN(U2964) );
  AOI21_X1 U6839 ( .B1(n5672), .B2(n5671), .A(n5670), .ZN(n5763) );
  NAND2_X1 U6840 ( .A1(n6425), .A2(REIP_REG_21__SCAN_IN), .ZN(n5758) );
  NAND2_X1 U6841 ( .A1(n6442), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5673)
         );
  OAI211_X1 U6842 ( .C1(n6437), .C2(n6070), .A(n5758), .B(n5673), .ZN(n5674)
         );
  AOI21_X1 U6843 ( .B1(n6097), .B2(n6432), .A(n5674), .ZN(n5675) );
  OAI21_X1 U6844 ( .B1(n5763), .B2(n6438), .A(n5675), .ZN(U2965) );
  XNOR2_X1 U6845 ( .A(n5663), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5677)
         );
  XNOR2_X1 U6846 ( .A(n5676), .B(n5677), .ZN(n6137) );
  NAND2_X1 U6847 ( .A1(n6137), .A2(n6431), .ZN(n5681) );
  INV_X1 U6848 ( .A(REIP_REG_20__SCAN_IN), .ZN(n5678) );
  OAI22_X1 U6849 ( .A1(n5707), .A2(n6088), .B1(n6498), .B2(n5678), .ZN(n5679)
         );
  AOI21_X1 U6850 ( .B1(n5709), .B2(n6080), .A(n5679), .ZN(n5680) );
  OAI211_X1 U6851 ( .C1(n5714), .C2(n6082), .A(n5681), .B(n5680), .ZN(U2966)
         );
  NAND2_X1 U6852 ( .A1(n3184), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6120) );
  OR3_X1 U6853 ( .A1(n5684), .A2(n3184), .A3(n5685), .ZN(n6118) );
  OAI21_X1 U6854 ( .B1(n5682), .B2(n6120), .A(n6118), .ZN(n5686) );
  XNOR2_X1 U6855 ( .A(n5686), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5780)
         );
  INV_X1 U6856 ( .A(n6194), .ZN(n5688) );
  NAND2_X1 U6857 ( .A1(n6442), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5687)
         );
  NAND2_X1 U6858 ( .A1(n6425), .A2(REIP_REG_18__SCAN_IN), .ZN(n5775) );
  OAI211_X1 U6859 ( .C1(n6437), .C2(n5688), .A(n5687), .B(n5775), .ZN(n5689)
         );
  AOI21_X1 U6860 ( .B1(n5690), .B2(n6432), .A(n5689), .ZN(n5691) );
  OAI21_X1 U6861 ( .B1(n6438), .B2(n5780), .A(n5691), .ZN(U2968) );
  OR2_X1 U6862 ( .A1(n3184), .A2(n5785), .ZN(n6116) );
  NAND2_X1 U6863 ( .A1(n3254), .A2(n6116), .ZN(n5693) );
  XNOR2_X1 U6864 ( .A(n5692), .B(n5693), .ZN(n5789) );
  NAND2_X1 U6865 ( .A1(n6425), .A2(REIP_REG_16__SCAN_IN), .ZN(n5782) );
  NOR2_X1 U6866 ( .A1(n6210), .A2(n5714), .ZN(n5694) );
  AOI211_X1 U6867 ( .C1(n5709), .C2(n6212), .A(n5695), .B(n5694), .ZN(n5696)
         );
  OAI21_X1 U6868 ( .B1(n6438), .B2(n5789), .A(n5696), .ZN(U2970) );
  OAI21_X1 U6869 ( .B1(n5697), .B2(n5698), .A(n5684), .ZN(n6148) );
  INV_X1 U6870 ( .A(n6148), .ZN(n5704) );
  AOI22_X1 U6871 ( .A1(n6442), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n6425), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5699) );
  OAI21_X1 U6872 ( .B1(n6437), .B2(n5700), .A(n5699), .ZN(n5701) );
  AOI21_X1 U6873 ( .B1(n5702), .B2(n6432), .A(n5701), .ZN(n5703) );
  OAI21_X1 U6874 ( .B1(n5704), .B2(n6438), .A(n5703), .ZN(U2971) );
  XNOR2_X1 U6875 ( .A(n3184), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5706)
         );
  XNOR2_X1 U6876 ( .A(n5705), .B(n5706), .ZN(n5790) );
  NAND2_X1 U6877 ( .A1(n5790), .A2(n6431), .ZN(n5712) );
  AOI21_X1 U6878 ( .B1(n5710), .B2(n5709), .A(n5708), .ZN(n5711) );
  OAI211_X1 U6879 ( .C1(n5714), .C2(n5713), .A(n5712), .B(n5711), .ZN(U2972)
         );
  INV_X1 U6880 ( .A(n5715), .ZN(n5720) );
  INV_X1 U6881 ( .A(n5716), .ZN(n5726) );
  NAND3_X1 U6882 ( .A1(n5726), .A2(n5718), .A3(n5717), .ZN(n5719) );
  OAI211_X1 U6883 ( .C1(n6019), .C2(n5783), .A(n5720), .B(n5719), .ZN(n5721)
         );
  AOI21_X1 U6884 ( .B1(n5729), .B2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n5721), 
        .ZN(n5722) );
  OAI21_X1 U6885 ( .B1(n5723), .B2(n6475), .A(n5722), .ZN(U2990) );
  AOI21_X1 U6886 ( .B1(n5726), .B2(n5725), .A(n5724), .ZN(n5727) );
  OAI21_X1 U6887 ( .B1(n6025), .B2(n5783), .A(n5727), .ZN(n5728) );
  AOI21_X1 U6888 ( .B1(n5729), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5728), 
        .ZN(n5730) );
  OAI21_X1 U6889 ( .B1(n5731), .B2(n6475), .A(n5730), .ZN(U2991) );
  INV_X1 U6890 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5733) );
  AOI21_X1 U6891 ( .B1(n5733), .B2(n6130), .A(n5732), .ZN(n5735) );
  AOI21_X1 U6892 ( .B1(n6124), .B2(n5735), .A(n5734), .ZN(n5736) );
  OAI21_X1 U6893 ( .B1(n6032), .B2(n5783), .A(n5736), .ZN(n5737) );
  AOI21_X1 U6894 ( .B1(n5738), .B2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5737), 
        .ZN(n5739) );
  OAI21_X1 U6895 ( .B1(n5740), .B2(n6475), .A(n5739), .ZN(U2992) );
  NOR2_X1 U6896 ( .A1(n5741), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5744)
         );
  OAI21_X1 U6897 ( .B1(n5783), .B2(n6052), .A(n5742), .ZN(n5743) );
  AOI211_X1 U6898 ( .C1(n5745), .C2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n5744), .B(n5743), .ZN(n5746) );
  OAI21_X1 U6899 ( .B1(n5747), .B2(n6475), .A(n5746), .ZN(U2995) );
  INV_X1 U6900 ( .A(n5748), .ZN(n5749) );
  NAND3_X1 U6901 ( .A1(n5757), .A2(n5750), .A3(n5749), .ZN(n5752) );
  OAI211_X1 U6902 ( .C1(n5783), .C2(n6069), .A(n5752), .B(n5751), .ZN(n5753)
         );
  AOI21_X1 U6903 ( .B1(n5761), .B2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5753), 
        .ZN(n5754) );
  OAI21_X1 U6904 ( .B1(n5755), .B2(n6475), .A(n5754), .ZN(U2996) );
  NAND2_X1 U6905 ( .A1(n5757), .A2(n5756), .ZN(n5759) );
  OAI211_X1 U6906 ( .C1(n5783), .C2(n6079), .A(n5759), .B(n5758), .ZN(n5760)
         );
  AOI21_X1 U6907 ( .B1(n5761), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5760), 
        .ZN(n5762) );
  OAI21_X1 U6908 ( .B1(n5763), .B2(n6475), .A(n5762), .ZN(U2997) );
  OAI21_X1 U6909 ( .B1(n5764), .B2(n5766), .A(n5765), .ZN(n6111) );
  INV_X1 U6910 ( .A(n6096), .ZN(n5772) );
  INV_X1 U6911 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5768) );
  OAI21_X1 U6912 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5767), .A(n6146), 
        .ZN(n5778) );
  AOI21_X1 U6913 ( .B1(n5768), .B2(n6501), .A(n5778), .ZN(n6140) );
  NAND2_X1 U6914 ( .A1(n6425), .A2(REIP_REG_19__SCAN_IN), .ZN(n5769) );
  OAI221_X1 U6915 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n6132), .C1(
        n5770), .C2(n6140), .A(n5769), .ZN(n5771) );
  AOI21_X1 U6916 ( .B1(n6503), .B2(n5772), .A(n5771), .ZN(n5773) );
  OAI21_X1 U6917 ( .B1(n6111), .B2(n6475), .A(n5773), .ZN(U2999) );
  NOR2_X1 U6918 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n6145), .ZN(n5774)
         );
  NAND2_X1 U6919 ( .A1(n6141), .A2(n5774), .ZN(n5776) );
  OAI211_X1 U6920 ( .C1(n5783), .C2(n6196), .A(n5776), .B(n5775), .ZN(n5777)
         );
  AOI21_X1 U6921 ( .B1(n5778), .B2(INSTADDRPOINTER_REG_18__SCAN_IN), .A(n5777), 
        .ZN(n5779) );
  OAI21_X1 U6922 ( .B1(n5780), .B2(n6475), .A(n5779), .ZN(U3000) );
  OAI21_X1 U6923 ( .B1(n5781), .B2(n5784), .A(n6453), .ZN(n6151) );
  OAI21_X1 U6924 ( .B1(n5783), .B2(n6209), .A(n5782), .ZN(n5787) );
  INV_X1 U6925 ( .A(n6161), .ZN(n6449) );
  NAND2_X1 U6926 ( .A1(n5784), .A2(n6449), .ZN(n6149) );
  AOI221_X1 U6927 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .C1(n3733), .C2(n5785), .A(n6149), 
        .ZN(n5786) );
  AOI211_X1 U6928 ( .C1(INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n6151), .A(n5787), .B(n5786), .ZN(n5788) );
  OAI21_X1 U6929 ( .B1(n5789), .B2(n6475), .A(n5788), .ZN(U3002) );
  NAND2_X1 U6930 ( .A1(n5790), .A2(n6507), .ZN(n5807) );
  INV_X1 U6931 ( .A(n5791), .ZN(n5793) );
  NAND2_X1 U6932 ( .A1(n5798), .A2(n5792), .ZN(n6160) );
  AOI21_X1 U6933 ( .B1(n5794), .B2(n5793), .A(n6160), .ZN(n5800) );
  AOI21_X1 U6934 ( .B1(n5796), .B2(n5803), .A(n5795), .ZN(n5797) );
  OAI21_X1 U6935 ( .B1(n5799), .B2(n5798), .A(n5797), .ZN(n6156) );
  OAI21_X1 U6936 ( .B1(n5800), .B2(n6156), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5806) );
  INV_X1 U6937 ( .A(n5801), .ZN(n5802) );
  AOI22_X1 U6938 ( .A1(n6503), .A2(n5802), .B1(n6425), .B2(
        REIP_REG_14__SCAN_IN), .ZN(n5805) );
  OR3_X1 U6939 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6161), .A3(n5803), 
        .ZN(n5804) );
  NAND4_X1 U6940 ( .A1(n5807), .A2(n5806), .A3(n5805), .A4(n5804), .ZN(U3004)
         );
  INV_X1 U6941 ( .A(n6665), .ZN(n6755) );
  OAI22_X1 U6942 ( .A1(n5810), .A2(n6755), .B1(n5809), .B2(n5808), .ZN(n5812)
         );
  MUX2_X1 U6943 ( .A(n5812), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n5811), 
        .Z(U3456) );
  INV_X1 U6944 ( .A(n5813), .ZN(n5834) );
  NAND2_X1 U6945 ( .A1(n5834), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5817) );
  AOI22_X1 U6946 ( .A1(n6562), .A2(n5836), .B1(n6577), .B2(n5835), .ZN(n5816)
         );
  NAND2_X1 U6947 ( .A1(n5837), .A2(n6563), .ZN(n5815) );
  OR2_X1 U6948 ( .A1(n5838), .A2(n6580), .ZN(n5814) );
  NAND4_X1 U6949 ( .A1(n5817), .A2(n5816), .A3(n5815), .A4(n5814), .ZN(U3020)
         );
  NAND2_X1 U6950 ( .A1(n5834), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5821) );
  AOI22_X1 U6951 ( .A1(n3259), .A2(n5836), .B1(n6583), .B2(n5835), .ZN(n5820)
         );
  NAND2_X1 U6952 ( .A1(n5837), .A2(n6528), .ZN(n5819) );
  OR2_X1 U6953 ( .A1(n5838), .A2(n5977), .ZN(n5818) );
  NAND4_X1 U6954 ( .A1(n5821), .A2(n5820), .A3(n5819), .A4(n5818), .ZN(U3021)
         );
  NAND2_X1 U6955 ( .A1(n5834), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5825) );
  AOI22_X1 U6956 ( .A1(n6593), .A2(n5836), .B1(n6595), .B2(n5835), .ZN(n5824)
         );
  NAND2_X1 U6957 ( .A1(n5837), .A2(n6536), .ZN(n5823) );
  OR2_X1 U6958 ( .A1(n5838), .A2(n5987), .ZN(n5822) );
  NAND4_X1 U6959 ( .A1(n5825), .A2(n5824), .A3(n5823), .A4(n5822), .ZN(U3023)
         );
  NAND2_X1 U6960 ( .A1(n5834), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5829) );
  AOI22_X1 U6961 ( .A1(n6599), .A2(n5836), .B1(n6601), .B2(n5835), .ZN(n5828)
         );
  NAND2_X1 U6962 ( .A1(n5837), .A2(n6600), .ZN(n5827) );
  OR2_X1 U6963 ( .A1(n5838), .A2(n6604), .ZN(n5826) );
  NAND4_X1 U6964 ( .A1(n5829), .A2(n5828), .A3(n5827), .A4(n5826), .ZN(U3024)
         );
  NAND2_X1 U6965 ( .A1(n5834), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5833) );
  AOI22_X1 U6966 ( .A1(n6605), .A2(n5836), .B1(n6607), .B2(n5835), .ZN(n5832)
         );
  NAND2_X1 U6967 ( .A1(n5837), .A2(n6606), .ZN(n5831) );
  OR2_X1 U6968 ( .A1(n5838), .A2(n6610), .ZN(n5830) );
  NAND4_X1 U6969 ( .A1(n5833), .A2(n5832), .A3(n5831), .A4(n5830), .ZN(U3025)
         );
  NAND2_X1 U6970 ( .A1(n5834), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5842) );
  AOI22_X1 U6971 ( .A1(n6620), .A2(n5836), .B1(n6624), .B2(n5835), .ZN(n5841)
         );
  NAND2_X1 U6972 ( .A1(n5837), .A2(n6555), .ZN(n5840) );
  OR2_X1 U6973 ( .A1(n5838), .A2(n6009), .ZN(n5839) );
  NAND4_X1 U6974 ( .A1(n5842), .A2(n5841), .A3(n5840), .A4(n5839), .ZN(U3027)
         );
  NAND2_X1 U6975 ( .A1(n5843), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5851) );
  AOI22_X1 U6976 ( .A1(n6562), .A2(n5845), .B1(n6577), .B2(n5844), .ZN(n5850)
         );
  NAND2_X1 U6977 ( .A1(n5846), .A2(n6518), .ZN(n5849) );
  NAND2_X1 U6978 ( .A1(n5847), .A2(n6563), .ZN(n5848) );
  NAND4_X1 U6979 ( .A1(n5851), .A2(n5850), .A3(n5849), .A4(n5848), .ZN(U3036)
         );
  NAND2_X1 U6980 ( .A1(n5854), .A2(n5853), .ZN(n5856) );
  NOR2_X1 U6981 ( .A1(n6633), .A2(n5859), .ZN(n5895) );
  INV_X1 U6982 ( .A(n5895), .ZN(n5855) );
  NAND2_X1 U6983 ( .A1(n5856), .A2(n5855), .ZN(n5858) );
  NOR2_X1 U6984 ( .A1(n5861), .A2(n5858), .ZN(n5857) );
  INV_X1 U6985 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n5868) );
  INV_X1 U6986 ( .A(n5858), .ZN(n5860) );
  OAI22_X1 U6987 ( .A1(n5861), .A2(n5860), .B1(n5859), .B2(n6780), .ZN(n5899)
         );
  AOI22_X1 U6988 ( .A1(n5938), .A2(n6518), .B1(n6562), .B2(n5895), .ZN(n5864)
         );
  OAI21_X1 U6989 ( .B1(n5865), .B2(n5897), .A(n5864), .ZN(n5866) );
  AOI21_X1 U6990 ( .B1(n6577), .B2(n5899), .A(n5866), .ZN(n5867) );
  OAI21_X1 U6991 ( .B1(n5902), .B2(n5868), .A(n5867), .ZN(U3060) );
  INV_X1 U6992 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n5872) );
  AOI22_X1 U6993 ( .A1(n5938), .A2(n6582), .B1(n6581), .B2(n5895), .ZN(n5869)
         );
  OAI21_X1 U6994 ( .B1(n6586), .B2(n5897), .A(n5869), .ZN(n5870) );
  AOI21_X1 U6995 ( .B1(n6583), .B2(n5899), .A(n5870), .ZN(n5871) );
  OAI21_X1 U6996 ( .B1(n5902), .B2(n5872), .A(n5871), .ZN(U3061) );
  INV_X1 U6997 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n5876) );
  AOI22_X1 U6998 ( .A1(n5938), .A2(n6532), .B1(n6587), .B2(n5895), .ZN(n5873)
         );
  OAI21_X1 U6999 ( .B1(n5979), .B2(n5897), .A(n5873), .ZN(n5874) );
  AOI21_X1 U7000 ( .B1(n6589), .B2(n5899), .A(n5874), .ZN(n5875) );
  OAI21_X1 U7001 ( .B1(n5902), .B2(n5876), .A(n5875), .ZN(U3062) );
  INV_X1 U7002 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n5880) );
  AOI22_X1 U7003 ( .A1(n5938), .A2(n6594), .B1(n6593), .B2(n5895), .ZN(n5877)
         );
  OAI21_X1 U7004 ( .B1(n6598), .B2(n5897), .A(n5877), .ZN(n5878) );
  AOI21_X1 U7005 ( .B1(n6595), .B2(n5899), .A(n5878), .ZN(n5879) );
  OAI21_X1 U7006 ( .B1(n5902), .B2(n5880), .A(n5879), .ZN(U3063) );
  INV_X1 U7007 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n5885) );
  AOI22_X1 U7008 ( .A1(n5938), .A2(n6540), .B1(n6599), .B2(n5895), .ZN(n5881)
         );
  OAI21_X1 U7009 ( .B1(n5882), .B2(n5897), .A(n5881), .ZN(n5883) );
  AOI21_X1 U7010 ( .B1(n6601), .B2(n5899), .A(n5883), .ZN(n5884) );
  OAI21_X1 U7011 ( .B1(n5902), .B2(n5885), .A(n5884), .ZN(U3064) );
  INV_X1 U7012 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n5890) );
  AOI22_X1 U7013 ( .A1(n5938), .A2(n6544), .B1(n6605), .B2(n5895), .ZN(n5886)
         );
  OAI21_X1 U7014 ( .B1(n5887), .B2(n5897), .A(n5886), .ZN(n5888) );
  AOI21_X1 U7015 ( .B1(n6607), .B2(n5899), .A(n5888), .ZN(n5889) );
  OAI21_X1 U7016 ( .B1(n5902), .B2(n5890), .A(n5889), .ZN(U3065) );
  INV_X1 U7017 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5894) );
  AOI22_X1 U7018 ( .A1(n5938), .A2(n6548), .B1(n6611), .B2(n5895), .ZN(n5891)
         );
  OAI21_X1 U7019 ( .B1(n5997), .B2(n5897), .A(n5891), .ZN(n5892) );
  AOI21_X1 U7020 ( .B1(n6614), .B2(n5899), .A(n5892), .ZN(n5893) );
  OAI21_X1 U7021 ( .B1(n5902), .B2(n5894), .A(n5893), .ZN(U3066) );
  INV_X1 U7022 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5901) );
  AOI22_X1 U7023 ( .A1(n5938), .A2(n6621), .B1(n6620), .B2(n5895), .ZN(n5896)
         );
  OAI21_X1 U7024 ( .B1(n6629), .B2(n5897), .A(n5896), .ZN(n5898) );
  AOI21_X1 U7025 ( .B1(n6624), .B2(n5899), .A(n5898), .ZN(n5900) );
  OAI21_X1 U7026 ( .B1(n5902), .B2(n5901), .A(n5900), .ZN(U3067) );
  AND2_X1 U7027 ( .A1(n6633), .A2(n6524), .ZN(n5928) );
  INV_X1 U7028 ( .A(n5928), .ZN(n5936) );
  NOR2_X1 U7029 ( .A1(n6514), .A2(n6571), .ZN(n5968) );
  AOI22_X1 U7030 ( .A1(n5968), .A2(n6315), .B1(n5904), .B2(n5967), .ZN(n5905)
         );
  NOR2_X1 U7031 ( .A1(n5906), .A2(n6571), .ZN(n5908) );
  OAI21_X1 U7032 ( .B1(n5938), .B2(n6554), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5907) );
  AOI211_X1 U7033 ( .C1(n5908), .C2(n5907), .A(n5960), .B(n5961), .ZN(n5909)
         );
  OAI211_X1 U7034 ( .C1(n5928), .C2(n7152), .A(n5909), .B(n6765), .ZN(n5933)
         );
  AOI22_X1 U7035 ( .A1(n5934), .A2(n6577), .B1(INSTQUEUE_REG_6__0__SCAN_IN), 
        .B2(n5933), .ZN(n5910) );
  OAI21_X1 U7036 ( .B1(n5969), .B2(n5936), .A(n5910), .ZN(n5911) );
  AOI21_X1 U7037 ( .B1(n6563), .B2(n5938), .A(n5911), .ZN(n5912) );
  OAI21_X1 U7038 ( .B1(n6580), .B2(n5940), .A(n5912), .ZN(U3068) );
  AOI22_X1 U7039 ( .A1(n5934), .A2(n6583), .B1(INSTQUEUE_REG_6__1__SCAN_IN), 
        .B2(n5933), .ZN(n5913) );
  OAI21_X1 U7040 ( .B1(n5973), .B2(n5936), .A(n5913), .ZN(n5914) );
  AOI21_X1 U7041 ( .B1(n6528), .B2(n5938), .A(n5914), .ZN(n5915) );
  OAI21_X1 U7042 ( .B1(n5977), .B2(n5940), .A(n5915), .ZN(U3069) );
  INV_X1 U7043 ( .A(n5938), .ZN(n5930) );
  AOI22_X1 U7044 ( .A1(n6587), .A2(n5928), .B1(INSTQUEUE_REG_6__2__SCAN_IN), 
        .B2(n5933), .ZN(n5916) );
  OAI21_X1 U7045 ( .B1(n5930), .B2(n5979), .A(n5916), .ZN(n5917) );
  AOI21_X1 U7046 ( .B1(n6589), .B2(n5934), .A(n5917), .ZN(n5918) );
  OAI21_X1 U7047 ( .B1(n6592), .B2(n5940), .A(n5918), .ZN(U3070) );
  AOI22_X1 U7048 ( .A1(n5934), .A2(n6595), .B1(INSTQUEUE_REG_6__3__SCAN_IN), 
        .B2(n5933), .ZN(n5919) );
  OAI21_X1 U7049 ( .B1(n5983), .B2(n5936), .A(n5919), .ZN(n5920) );
  AOI21_X1 U7050 ( .B1(n6536), .B2(n5938), .A(n5920), .ZN(n5921) );
  OAI21_X1 U7051 ( .B1(n5987), .B2(n5940), .A(n5921), .ZN(U3071) );
  AOI22_X1 U7052 ( .A1(n5934), .A2(n6601), .B1(INSTQUEUE_REG_6__4__SCAN_IN), 
        .B2(n5933), .ZN(n5922) );
  OAI21_X1 U7053 ( .B1(n5988), .B2(n5936), .A(n5922), .ZN(n5923) );
  AOI21_X1 U7054 ( .B1(n6600), .B2(n5938), .A(n5923), .ZN(n5924) );
  OAI21_X1 U7055 ( .B1(n6604), .B2(n5940), .A(n5924), .ZN(U3072) );
  AOI22_X1 U7056 ( .A1(n5934), .A2(n6607), .B1(INSTQUEUE_REG_6__5__SCAN_IN), 
        .B2(n5933), .ZN(n5925) );
  OAI21_X1 U7057 ( .B1(n5992), .B2(n5936), .A(n5925), .ZN(n5926) );
  AOI21_X1 U7058 ( .B1(n6606), .B2(n5938), .A(n5926), .ZN(n5927) );
  OAI21_X1 U7059 ( .B1(n6610), .B2(n5940), .A(n5927), .ZN(U3073) );
  AOI22_X1 U7060 ( .A1(n6611), .A2(n5928), .B1(INSTQUEUE_REG_6__6__SCAN_IN), 
        .B2(n5933), .ZN(n5929) );
  OAI21_X1 U7061 ( .B1(n5930), .B2(n5997), .A(n5929), .ZN(n5931) );
  AOI21_X1 U7062 ( .B1(n6614), .B2(n5934), .A(n5931), .ZN(n5932) );
  OAI21_X1 U7063 ( .B1(n6618), .B2(n5940), .A(n5932), .ZN(U3074) );
  AOI22_X1 U7064 ( .A1(n5934), .A2(n6624), .B1(INSTQUEUE_REG_6__7__SCAN_IN), 
        .B2(n5933), .ZN(n5935) );
  OAI21_X1 U7065 ( .B1(n6005), .B2(n5936), .A(n5935), .ZN(n5937) );
  AOI21_X1 U7066 ( .B1(n6555), .B2(n5938), .A(n5937), .ZN(n5939) );
  OAI21_X1 U7067 ( .B1(n6009), .B2(n5940), .A(n5939), .ZN(U3075) );
  NAND2_X1 U7068 ( .A1(n5949), .A2(n6583), .ZN(n5944) );
  AOI22_X1 U7069 ( .A1(n3259), .A2(n5951), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5950), .ZN(n5943) );
  NAND2_X1 U7070 ( .A1(n6613), .A2(n6582), .ZN(n5942) );
  NAND2_X1 U7071 ( .A1(n5952), .A2(n6528), .ZN(n5941) );
  NAND4_X1 U7072 ( .A1(n5944), .A2(n5943), .A3(n5942), .A4(n5941), .ZN(U3101)
         );
  NAND2_X1 U7073 ( .A1(n5949), .A2(n6595), .ZN(n5948) );
  AOI22_X1 U7074 ( .A1(n6593), .A2(n5951), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5950), .ZN(n5947) );
  NAND2_X1 U7075 ( .A1(n6613), .A2(n6594), .ZN(n5946) );
  NAND2_X1 U7076 ( .A1(n5952), .A2(n6536), .ZN(n5945) );
  NAND4_X1 U7077 ( .A1(n5948), .A2(n5947), .A3(n5946), .A4(n5945), .ZN(U3103)
         );
  NAND2_X1 U7078 ( .A1(n5949), .A2(n6624), .ZN(n5956) );
  AOI22_X1 U7079 ( .A1(n6620), .A2(n5951), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5950), .ZN(n5955) );
  NAND2_X1 U7080 ( .A1(n6613), .A2(n6621), .ZN(n5954) );
  NAND2_X1 U7081 ( .A1(n5952), .A2(n6555), .ZN(n5953) );
  NAND4_X1 U7082 ( .A1(n5956), .A2(n5955), .A3(n5954), .A4(n5953), .ZN(U3107)
         );
  NOR2_X1 U7083 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5957), .ZN(n5964)
         );
  OAI21_X1 U7084 ( .B1(n3260), .B2(n5958), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5959) );
  NAND3_X1 U7085 ( .A1(n6514), .A2(n6564), .A3(n5959), .ZN(n5963) );
  NOR3_X1 U7086 ( .A1(n5961), .A2(n6765), .A3(n5960), .ZN(n5962) );
  NAND2_X1 U7087 ( .A1(n6002), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5972)
         );
  INV_X1 U7088 ( .A(n5964), .ZN(n6004) );
  INV_X1 U7089 ( .A(n5965), .ZN(n5966) );
  AOI22_X1 U7090 ( .A1(n5968), .A2(n4582), .B1(n5967), .B2(n5966), .ZN(n6003)
         );
  OAI22_X1 U7091 ( .A1(n5969), .A2(n6004), .B1(n6003), .B2(n6527), .ZN(n5970)
         );
  AOI21_X1 U7092 ( .B1(n6563), .B2(n3260), .A(n5970), .ZN(n5971) );
  OAI211_X1 U7093 ( .C1(n6010), .C2(n6580), .A(n5972), .B(n5971), .ZN(U3132)
         );
  NAND2_X1 U7094 ( .A1(n6002), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5976)
         );
  OAI22_X1 U7095 ( .A1(n5973), .A2(n6004), .B1(n6003), .B2(n6531), .ZN(n5974)
         );
  AOI21_X1 U7096 ( .B1(n3260), .B2(n6528), .A(n5974), .ZN(n5975) );
  OAI211_X1 U7097 ( .C1(n6010), .C2(n5977), .A(n5976), .B(n5975), .ZN(U3133)
         );
  INV_X1 U7098 ( .A(n6003), .ZN(n5999) );
  OAI22_X1 U7099 ( .A1(n3235), .A2(n5979), .B1(n5978), .B2(n6004), .ZN(n5980)
         );
  AOI21_X1 U7100 ( .B1(n6589), .B2(n5999), .A(n5980), .ZN(n5982) );
  NAND2_X1 U7101 ( .A1(n6002), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5981)
         );
  OAI211_X1 U7102 ( .C1(n6010), .C2(n6592), .A(n5982), .B(n5981), .ZN(U3134)
         );
  NAND2_X1 U7103 ( .A1(n6002), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5986)
         );
  OAI22_X1 U7104 ( .A1(n5983), .A2(n6004), .B1(n6003), .B2(n6539), .ZN(n5984)
         );
  AOI21_X1 U7105 ( .B1(n3260), .B2(n6536), .A(n5984), .ZN(n5985) );
  OAI211_X1 U7106 ( .C1(n6010), .C2(n5987), .A(n5986), .B(n5985), .ZN(U3135)
         );
  NAND2_X1 U7107 ( .A1(n6002), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5991)
         );
  OAI22_X1 U7108 ( .A1(n5988), .A2(n6004), .B1(n6003), .B2(n6543), .ZN(n5989)
         );
  AOI21_X1 U7109 ( .B1(n3260), .B2(n6600), .A(n5989), .ZN(n5990) );
  OAI211_X1 U7110 ( .C1(n6010), .C2(n6604), .A(n5991), .B(n5990), .ZN(U3136)
         );
  NAND2_X1 U7111 ( .A1(n6002), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5995)
         );
  OAI22_X1 U7112 ( .A1(n5992), .A2(n6004), .B1(n6003), .B2(n6547), .ZN(n5993)
         );
  AOI21_X1 U7113 ( .B1(n3260), .B2(n6606), .A(n5993), .ZN(n5994) );
  OAI211_X1 U7114 ( .C1(n6010), .C2(n6610), .A(n5995), .B(n5994), .ZN(U3137)
         );
  OAI22_X1 U7115 ( .A1(n3235), .A2(n5997), .B1(n5996), .B2(n6004), .ZN(n5998)
         );
  AOI21_X1 U7116 ( .B1(n6614), .B2(n5999), .A(n5998), .ZN(n6001) );
  NAND2_X1 U7117 ( .A1(n6002), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n6000)
         );
  OAI211_X1 U7118 ( .C1(n6010), .C2(n6618), .A(n6001), .B(n6000), .ZN(U3138)
         );
  NAND2_X1 U7119 ( .A1(n6002), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n6008)
         );
  OAI22_X1 U7120 ( .A1(n6005), .A2(n6004), .B1(n6003), .B2(n6559), .ZN(n6006)
         );
  AOI21_X1 U7121 ( .B1(n3260), .B2(n6555), .A(n6006), .ZN(n6007) );
  OAI211_X1 U7122 ( .C1(n6010), .C2(n6009), .A(n6008), .B(n6007), .ZN(U3139)
         );
  AND2_X1 U7123 ( .A1(n6358), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U7124 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6731) );
  NOR2_X1 U7125 ( .A1(n6011), .A2(n6731), .ZN(n6015) );
  AOI22_X1 U7126 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n6272), .B1(n6302), 
        .B2(n6012), .ZN(n6013) );
  OAI21_X1 U7127 ( .B1(n7058), .B2(n6246), .A(n6013), .ZN(n6014) );
  AOI211_X1 U7128 ( .C1(n6016), .C2(n6254), .A(n6015), .B(n6014), .ZN(n6018)
         );
  NAND3_X1 U7129 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6024), .A3(n6731), .ZN(
        n6017) );
  OAI211_X1 U7130 ( .C1(n6318), .C2(n6019), .A(n6018), .B(n6017), .ZN(U2799)
         );
  INV_X1 U7131 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6023) );
  AOI22_X1 U7132 ( .A1(EBX_REG_27__SCAN_IN), .A2(n6325), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6272), .ZN(n6020) );
  OAI21_X1 U7133 ( .B1(n6021), .B2(n6319), .A(n6020), .ZN(n6022) );
  AOI221_X1 U7134 ( .B1(n6024), .B2(n6023), .C1(n6036), .C2(
        REIP_REG_27__SCAN_IN), .A(n6022), .ZN(n6029) );
  NOR2_X1 U7135 ( .A1(n6025), .A2(n6318), .ZN(n6026) );
  AOI21_X1 U7136 ( .B1(n6027), .B2(n6254), .A(n6026), .ZN(n6028) );
  NAND2_X1 U7137 ( .A1(n6029), .A2(n6028), .ZN(U2800) );
  AOI22_X1 U7138 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n6272), .B1(n6030), 
        .B2(n6302), .ZN(n6038) );
  INV_X1 U7139 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6724) );
  INV_X1 U7140 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6727) );
  OAI21_X1 U7141 ( .B1(n6724), .B2(n6031), .A(n6727), .ZN(n6035) );
  OAI22_X1 U7142 ( .A1(n6033), .A2(n6278), .B1(n6318), .B2(n6032), .ZN(n6034)
         );
  OAI211_X1 U7143 ( .C1(n6945), .C2(n6246), .A(n6038), .B(n6037), .ZN(U2801)
         );
  INV_X1 U7144 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6044) );
  NAND2_X1 U7145 ( .A1(n6039), .A2(n6254), .ZN(n6043) );
  OAI22_X1 U7146 ( .A1(n6040), .A2(n6319), .B1(n6314), .B2(n3813), .ZN(n6041)
         );
  AOI21_X1 U7147 ( .B1(n6325), .B2(EBX_REG_24__SCAN_IN), .A(n6041), .ZN(n6042)
         );
  OAI211_X1 U7148 ( .C1(n6045), .C2(n6044), .A(n6043), .B(n6042), .ZN(n6047)
         );
  NOR2_X1 U7149 ( .A1(n6047), .A2(n6046), .ZN(n6048) );
  OAI21_X1 U7150 ( .B1(n6049), .B2(n6318), .A(n6048), .ZN(U2803) );
  OAI22_X1 U7151 ( .A1(n4145), .A2(n6314), .B1(n6050), .B2(n6319), .ZN(n6051)
         );
  AOI21_X1 U7152 ( .B1(EBX_REG_23__SCAN_IN), .B2(n6325), .A(n6051), .ZN(n6059)
         );
  INV_X1 U7153 ( .A(n6052), .ZN(n6053) );
  AOI22_X1 U7154 ( .A1(n6054), .A2(n6254), .B1(n4435), .B2(n6053), .ZN(n6058)
         );
  OAI21_X1 U7155 ( .B1(REIP_REG_23__SCAN_IN), .B2(n6056), .A(n6055), .ZN(n6057) );
  NAND3_X1 U7156 ( .A1(n6059), .A2(n6058), .A3(n6057), .ZN(U2804) );
  NOR2_X1 U7157 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6060), .ZN(n6076) );
  NOR2_X1 U7158 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6060), .ZN(n6064) );
  AOI22_X1 U7159 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n6272), .B1(n6302), 
        .B2(n6061), .ZN(n6062) );
  OAI21_X1 U7160 ( .B1(n5576), .B2(n6246), .A(n6062), .ZN(n6063) );
  AOI21_X1 U7161 ( .B1(n6064), .B2(REIP_REG_21__SCAN_IN), .A(n6063), .ZN(n6065) );
  OAI21_X1 U7162 ( .B1(n6066), .B2(n6278), .A(n6065), .ZN(n6067) );
  AOI221_X1 U7163 ( .B1(n6076), .B2(REIP_REG_22__SCAN_IN), .C1(n6085), .C2(
        REIP_REG_22__SCAN_IN), .A(n6067), .ZN(n6068) );
  OAI21_X1 U7164 ( .B1(n6069), .B2(n6318), .A(n6068), .ZN(U2805) );
  INV_X1 U7165 ( .A(n6070), .ZN(n6071) );
  NAND2_X1 U7166 ( .A1(n6302), .A2(n6071), .ZN(n6074) );
  NAND2_X1 U7167 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6085), .ZN(n6073) );
  AOI22_X1 U7168 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6325), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6272), .ZN(n6072) );
  NAND3_X1 U7169 ( .A1(n6074), .A2(n6073), .A3(n6072), .ZN(n6075) );
  OR2_X1 U7170 ( .A1(n6076), .A2(n6075), .ZN(n6077) );
  AOI21_X1 U7171 ( .B1(n6097), .B2(n6254), .A(n6077), .ZN(n6078) );
  OAI21_X1 U7172 ( .B1(n6079), .B2(n6318), .A(n6078), .ZN(U2806) );
  AOI22_X1 U7173 ( .A1(EBX_REG_20__SCAN_IN), .A2(n6325), .B1(n6080), .B2(n6302), .ZN(n6087) );
  OAI22_X1 U7174 ( .A1(n6082), .A2(n6278), .B1(n6081), .B2(n6318), .ZN(n6083)
         );
  AOI221_X1 U7175 ( .B1(REIP_REG_20__SCAN_IN), .B2(n6085), .C1(n6084), .C2(
        n6085), .A(n6083), .ZN(n6086) );
  OAI211_X1 U7176 ( .C1(n6088), .C2(n6314), .A(n6087), .B(n6086), .ZN(U2807)
         );
  INV_X1 U7177 ( .A(n6110), .ZN(n6100) );
  INV_X1 U7178 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6714) );
  NOR3_X1 U7179 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6093), .A3(n6714), .ZN(n6092) );
  INV_X1 U7180 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6994) );
  INV_X1 U7181 ( .A(n6115), .ZN(n6089) );
  AOI22_X1 U7182 ( .A1(EBX_REG_19__SCAN_IN), .A2(n6325), .B1(n6089), .B2(n6302), .ZN(n6090) );
  OAI211_X1 U7183 ( .C1(n6314), .C2(n6994), .A(n6090), .B(n6498), .ZN(n6091)
         );
  AOI211_X1 U7184 ( .C1(n6100), .C2(n6254), .A(n6092), .B(n6091), .ZN(n6095)
         );
  NOR2_X1 U7185 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6093), .ZN(n6189) );
  OAI21_X1 U7186 ( .B1(n6197), .B2(n6189), .A(REIP_REG_19__SCAN_IN), .ZN(n6094) );
  OAI211_X1 U7187 ( .C1(n6096), .C2(n6318), .A(n6095), .B(n6094), .ZN(U2808)
         );
  AOI22_X1 U7188 ( .A1(n6097), .A2(n6330), .B1(n6329), .B2(DATAI_21_), .ZN(
        n6099) );
  AOI22_X1 U7189 ( .A1(n6333), .A2(DATAI_5_), .B1(n6332), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7190 ( .A1(n6099), .A2(n6098), .ZN(U2870) );
  AOI22_X1 U7191 ( .A1(n6100), .A2(n6330), .B1(n6329), .B2(DATAI_19_), .ZN(
        n6102) );
  AOI22_X1 U7192 ( .A1(n6333), .A2(DATAI_3_), .B1(n6332), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U7193 ( .A1(n6102), .A2(n6101), .ZN(U2872) );
  AOI22_X1 U7194 ( .A1(n6425), .A2(REIP_REG_25__SCAN_IN), .B1(n6442), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6108) );
  INV_X1 U7195 ( .A(n5631), .ZN(n6105) );
  INV_X1 U7196 ( .A(n6103), .ZN(n6104) );
  OAI21_X1 U7197 ( .B1(n6105), .B2(n6104), .A(n4438), .ZN(n6127) );
  AOI22_X1 U7198 ( .A1(n6106), .A2(n6432), .B1(n6431), .B2(n6127), .ZN(n6107)
         );
  OAI211_X1 U7199 ( .C1(n6437), .C2(n6109), .A(n6108), .B(n6107), .ZN(U2961)
         );
  AOI22_X1 U7200 ( .A1(n6425), .A2(REIP_REG_19__SCAN_IN), .B1(n6442), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6114) );
  OAI22_X1 U7201 ( .A1(n6111), .A2(n6438), .B1(n5714), .B2(n6110), .ZN(n6112)
         );
  INV_X1 U7202 ( .A(n6112), .ZN(n6113) );
  OAI211_X1 U7203 ( .C1(n6437), .C2(n6115), .A(n6114), .B(n6113), .ZN(U2967)
         );
  AOI22_X1 U7204 ( .A1(n6425), .A2(REIP_REG_17__SCAN_IN), .B1(n6442), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6123) );
  INV_X1 U7205 ( .A(n5682), .ZN(n6121) );
  NAND2_X1 U7206 ( .A1(n5682), .A2(n6116), .ZN(n6117) );
  OAI211_X1 U7207 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n3184), .A(n6117), .B(n6120), .ZN(n6119) );
  OAI211_X1 U7208 ( .C1(n6121), .C2(n6120), .A(n6119), .B(n6118), .ZN(n6142)
         );
  AOI22_X1 U7209 ( .A1(n6142), .A2(n6431), .B1(n6432), .B2(n6331), .ZN(n6122)
         );
  OAI211_X1 U7210 ( .C1(n6437), .C2(n6204), .A(n6123), .B(n6122), .ZN(U2969)
         );
  AOI22_X1 U7211 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6425), .B1(n6124), .B2(
        n6130), .ZN(n6129) );
  INV_X1 U7212 ( .A(n6125), .ZN(n6126) );
  AOI22_X1 U7213 ( .A1(n6127), .A2(n6507), .B1(n6503), .B2(n6126), .ZN(n6128)
         );
  OAI211_X1 U7214 ( .C1(n6131), .C2(n6130), .A(n6129), .B(n6128), .ZN(U2993)
         );
  NOR2_X1 U7215 ( .A1(n6133), .A2(n6132), .ZN(n6135) );
  AOI22_X1 U7216 ( .A1(n6425), .A2(REIP_REG_20__SCAN_IN), .B1(n6135), .B2(
        n6134), .ZN(n6139) );
  AOI22_X1 U7217 ( .A1(n6137), .A2(n6507), .B1(n6503), .B2(n6136), .ZN(n6138)
         );
  OAI211_X1 U7218 ( .C1(n6140), .C2(n5428), .A(n6139), .B(n6138), .ZN(U2998)
         );
  AOI22_X1 U7219 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6425), .B1(n6141), .B2(
        n6145), .ZN(n6144) );
  AOI22_X1 U7220 ( .A1(n6142), .A2(n6507), .B1(n6503), .B2(n6201), .ZN(n6143)
         );
  OAI211_X1 U7221 ( .C1(n6146), .C2(n6145), .A(n6144), .B(n6143), .ZN(U3001)
         );
  AOI22_X1 U7222 ( .A1(n6148), .A2(n6507), .B1(n6503), .B2(n6147), .ZN(n6154)
         );
  INV_X1 U7223 ( .A(n6149), .ZN(n6152) );
  NOR2_X1 U7224 ( .A1(n6498), .A2(n6709), .ZN(n6150) );
  AOI221_X1 U7225 ( .B1(n6152), .B2(n3733), .C1(n6151), .C2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A(n6150), .ZN(n6153) );
  NAND2_X1 U7226 ( .A1(n6154), .A2(n6153), .ZN(U3003) );
  AOI21_X1 U7227 ( .B1(n6503), .B2(n6216), .A(n6155), .ZN(n6159) );
  AOI22_X1 U7228 ( .A1(n6157), .A2(n6507), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n6156), .ZN(n6158) );
  OAI211_X1 U7229 ( .C1(n6161), .C2(n6160), .A(n6159), .B(n6158), .ZN(U3005)
         );
  NAND4_X1 U7230 ( .A1(n6163), .A2(n6665), .A3(n6162), .A4(n6294), .ZN(n6164)
         );
  OAI21_X1 U7231 ( .B1(n6753), .B2(n6165), .A(n6164), .ZN(U3455) );
  AOI21_X1 U7232 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6691), .A(n7054), .ZN(n6171) );
  INV_X1 U7233 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6166) );
  NOR2_X2 U7234 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6682), .ZN(n6790) );
  AOI21_X1 U7235 ( .B1(n6171), .B2(n6166), .A(n6790), .ZN(U2789) );
  OAI21_X1 U7236 ( .B1(n6167), .B2(n6662), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6168) );
  OAI21_X1 U7237 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6169), .A(n6168), .ZN(
        U2790) );
  INV_X1 U7238 ( .A(n6790), .ZN(n6738) );
  NOR2_X1 U7239 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6172) );
  OAI21_X1 U7240 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6172), .A(n6732), .ZN(n6170)
         );
  OAI21_X1 U7241 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6738), .A(n6170), .ZN(
        U2791) );
  NOR2_X1 U7242 ( .A1(n6790), .A2(n6171), .ZN(n6743) );
  OAI21_X1 U7243 ( .B1(n6172), .B2(BS16_N), .A(n6743), .ZN(n6742) );
  OAI21_X1 U7244 ( .B1(n6743), .B2(n6781), .A(n6742), .ZN(U2792) );
  OAI21_X1 U7245 ( .B1(n6174), .B2(n6173), .A(n6438), .ZN(U2793) );
  NOR4_X1 U7246 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(
        DATAWIDTH_REG_4__SCAN_IN), .ZN(n6184) );
  AOI211_X1 U7247 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_30__SCAN_IN), .B(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6183) );
  NOR4_X1 U7248 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(
        n6175) );
  INV_X1 U7249 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n7151) );
  INV_X1 U7250 ( .A(DATAWIDTH_REG_29__SCAN_IN), .ZN(n7173) );
  NAND3_X1 U7251 ( .A1(n6175), .A2(n7151), .A3(n7173), .ZN(n6181) );
  NOR4_X1 U7252 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n6179) );
  NOR4_X1 U7253 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_12__SCAN_IN), .A4(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6178)
         );
  NOR4_X1 U7254 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(
        DATAWIDTH_REG_26__SCAN_IN), .A3(DATAWIDTH_REG_27__SCAN_IN), .A4(
        DATAWIDTH_REG_28__SCAN_IN), .ZN(n6177) );
  NOR4_X1 U7255 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n6176) );
  NAND4_X1 U7256 ( .A1(n6179), .A2(n6178), .A3(n6177), .A4(n6176), .ZN(n6180)
         );
  NOR4_X1 U7257 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(n6181), .A4(n6180), .ZN(n6182) );
  NAND3_X1 U7258 ( .A1(n6184), .A2(n6183), .A3(n6182), .ZN(n6776) );
  INV_X1 U7259 ( .A(n6776), .ZN(n6773) );
  NAND2_X1 U7260 ( .A1(n6773), .A2(n6769), .ZN(n6772) );
  NOR3_X1 U7261 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(n6772), .ZN(n6186) );
  AOI21_X1 U7262 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(n6776), .A(n6186), .ZN(
        n6185) );
  OAI21_X1 U7263 ( .B1(n6775), .B2(n6776), .A(n6185), .ZN(U2794) );
  NAND2_X1 U7264 ( .A1(n6773), .A2(n6775), .ZN(n6767) );
  AOI21_X1 U7265 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(n6776), .A(n6186), .ZN(
        n6187) );
  OAI21_X1 U7266 ( .B1(DATAWIDTH_REG_1__SCAN_IN), .B2(n6767), .A(n6187), .ZN(
        U2795) );
  AOI21_X1 U7267 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6272), .A(n6425), 
        .ZN(n6188) );
  OAI21_X1 U7268 ( .B1(n5404), .B2(n6246), .A(n6188), .ZN(n6190) );
  AOI211_X1 U7269 ( .C1(REIP_REG_18__SCAN_IN), .C2(n6197), .A(n6190), .B(n6189), .ZN(n6191) );
  OAI21_X1 U7270 ( .B1(n6192), .B2(n6278), .A(n6191), .ZN(n6193) );
  AOI21_X1 U7271 ( .B1(n6194), .B2(n6302), .A(n6193), .ZN(n6195) );
  OAI21_X1 U7272 ( .B1(n6318), .B2(n6196), .A(n6195), .ZN(U2809) );
  INV_X1 U7273 ( .A(EBX_REG_17__SCAN_IN), .ZN(n7073) );
  OAI21_X1 U7274 ( .B1(REIP_REG_17__SCAN_IN), .B2(n6198), .A(n6197), .ZN(n6199) );
  OAI211_X1 U7275 ( .C1(n6246), .C2(n7073), .A(n6498), .B(n6199), .ZN(n6200)
         );
  AOI21_X1 U7276 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6272), .A(n6200), 
        .ZN(n6203) );
  AOI22_X1 U7277 ( .A1(n6331), .A2(n6254), .B1(n4435), .B2(n6201), .ZN(n6202)
         );
  OAI211_X1 U7278 ( .C1(n6204), .C2(n6319), .A(n6203), .B(n6202), .ZN(U2810)
         );
  OAI21_X1 U7279 ( .B1(n6709), .B2(n6205), .A(n6297), .ZN(n6207) );
  AOI22_X1 U7280 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6207), .B1(n6206), .B2(
        n6712), .ZN(n6208) );
  AOI211_X1 U7281 ( .C1(n6272), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6425), 
        .B(n6208), .ZN(n6214) );
  OAI22_X1 U7282 ( .A1(n6210), .A2(n6278), .B1(n6318), .B2(n6209), .ZN(n6211)
         );
  AOI21_X1 U7283 ( .B1(n6212), .B2(n6302), .A(n6211), .ZN(n6213) );
  OAI211_X1 U7284 ( .C1(n6215), .C2(n6246), .A(n6214), .B(n6213), .ZN(U2811)
         );
  AOI22_X1 U7285 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6325), .B1(n4435), .B2(n6216), .ZN(n6227) );
  INV_X1 U7286 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6706) );
  NOR3_X1 U7287 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6706), .A3(n6223), .ZN(n6217) );
  AOI211_X1 U7288 ( .C1(n6272), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6425), 
        .B(n6217), .ZN(n6226) );
  INV_X1 U7289 ( .A(n6218), .ZN(n6221) );
  INV_X1 U7290 ( .A(n6219), .ZN(n6220) );
  AOI22_X1 U7291 ( .A1(n6221), .A2(n6254), .B1(n6302), .B2(n6220), .ZN(n6225)
         );
  OAI21_X1 U7292 ( .B1(n6262), .B2(n6222), .A(n6296), .ZN(n6237) );
  NOR2_X1 U7293 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6223), .ZN(n6230) );
  OAI21_X1 U7294 ( .B1(n6237), .B2(n6230), .A(REIP_REG_13__SCAN_IN), .ZN(n6224) );
  NAND4_X1 U7295 ( .A1(n6227), .A2(n6226), .A3(n6225), .A4(n6224), .ZN(U2814)
         );
  INV_X1 U7296 ( .A(EBX_REG_12__SCAN_IN), .ZN(n7074) );
  AOI22_X1 U7297 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n6272), .B1(
        REIP_REG_12__SCAN_IN), .B2(n6237), .ZN(n6228) );
  OAI211_X1 U7298 ( .C1(n6246), .C2(n7074), .A(n6228), .B(n6498), .ZN(n6229)
         );
  AOI211_X1 U7299 ( .C1(n6231), .C2(n4435), .A(n6230), .B(n6229), .ZN(n6235)
         );
  AOI22_X1 U7300 ( .A1(n6233), .A2(n6254), .B1(n6302), .B2(n6232), .ZN(n6234)
         );
  NAND2_X1 U7301 ( .A1(n6235), .A2(n6234), .ZN(U2815) );
  OAI21_X1 U7302 ( .B1(n6262), .B2(n6236), .A(n6702), .ZN(n6238) );
  NAND2_X1 U7303 ( .A1(n6238), .A2(n6237), .ZN(n6245) );
  OAI21_X1 U7304 ( .B1(n6314), .B2(n3810), .A(n6498), .ZN(n6239) );
  AOI21_X1 U7305 ( .B1(n4435), .B2(n6448), .A(n6239), .ZN(n6240) );
  OAI21_X1 U7306 ( .B1(n6241), .B2(n6278), .A(n6240), .ZN(n6242) );
  AOI21_X1 U7307 ( .B1(n6243), .B2(n6302), .A(n6242), .ZN(n6244) );
  OAI211_X1 U7308 ( .C1(n6247), .C2(n6246), .A(n6245), .B(n6244), .ZN(U2816)
         );
  INV_X1 U7309 ( .A(n6248), .ZN(n6251) );
  AOI221_X1 U7310 ( .B1(REIP_REG_9__SCAN_IN), .B2(REIP_REG_10__SCAN_IN), .C1(
        n5159), .C2(n6703), .A(n6249), .ZN(n6250) );
  AOI21_X1 U7311 ( .B1(n6251), .B2(n4435), .A(n6250), .ZN(n6259) );
  AOI22_X1 U7312 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6325), .B1(
        PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n6272), .ZN(n6258) );
  AOI21_X1 U7313 ( .B1(REIP_REG_10__SCAN_IN), .B2(n6252), .A(n6425), .ZN(n6257) );
  AOI22_X1 U7314 ( .A1(n6255), .A2(n6254), .B1(n6302), .B2(n6253), .ZN(n6256)
         );
  NAND4_X1 U7315 ( .A1(n6259), .A2(n6258), .A3(n6257), .A4(n6256), .ZN(U2817)
         );
  AOI21_X1 U7316 ( .B1(n6272), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6425), 
        .ZN(n6271) );
  AOI22_X1 U7317 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6325), .B1(n4435), .B2(n6463), 
        .ZN(n6270) );
  OAI21_X1 U7318 ( .B1(n6262), .B2(n6260), .A(n6296), .ZN(n6288) );
  NOR2_X1 U7319 ( .A1(n6262), .A2(n6261), .ZN(n6289) );
  AND2_X1 U7320 ( .A1(n6289), .A2(REIP_REG_5__SCAN_IN), .ZN(n6267) );
  INV_X1 U7321 ( .A(n6267), .ZN(n6263) );
  NOR2_X1 U7322 ( .A1(n6263), .A2(REIP_REG_6__SCAN_IN), .ZN(n6276) );
  OAI22_X1 U7323 ( .A1(n6265), .A2(n6278), .B1(n6264), .B2(n6319), .ZN(n6266)
         );
  AOI221_X1 U7324 ( .B1(n6288), .B2(REIP_REG_7__SCAN_IN), .C1(n6276), .C2(
        REIP_REG_7__SCAN_IN), .A(n6266), .ZN(n6269) );
  INV_X1 U7325 ( .A(REIP_REG_7__SCAN_IN), .ZN(n7170) );
  NAND3_X1 U7326 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6267), .A3(n7170), .ZN(n6268) );
  NAND4_X1 U7327 ( .A1(n6271), .A2(n6270), .A3(n6269), .A4(n6268), .ZN(U2820)
         );
  AOI22_X1 U7328 ( .A1(EBX_REG_6__SCAN_IN), .A2(n6325), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6272), .ZN(n6273) );
  OAI211_X1 U7329 ( .C1(n6318), .C2(n6274), .A(n6273), .B(n6498), .ZN(n6275)
         );
  AOI211_X1 U7330 ( .C1(n6288), .C2(REIP_REG_6__SCAN_IN), .A(n6276), .B(n6275), 
        .ZN(n6282) );
  OAI22_X1 U7331 ( .A1(n6279), .A2(n6278), .B1(n6277), .B2(n6319), .ZN(n6280)
         );
  INV_X1 U7332 ( .A(n6280), .ZN(n6281) );
  NAND2_X1 U7333 ( .A1(n6282), .A2(n6281), .ZN(U2821) );
  INV_X1 U7334 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6285) );
  AOI22_X1 U7335 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6325), .B1(n4435), .B2(n6283), 
        .ZN(n6284) );
  OAI211_X1 U7336 ( .C1(n6314), .C2(n6285), .A(n6284), .B(n6498), .ZN(n6286)
         );
  AOI21_X1 U7337 ( .B1(n6287), .B2(n6304), .A(n6286), .ZN(n6291) );
  OAI21_X1 U7338 ( .B1(REIP_REG_5__SCAN_IN), .B2(n6289), .A(n6288), .ZN(n6290)
         );
  OAI211_X1 U7339 ( .C1(n6319), .C2(n6292), .A(n6291), .B(n6290), .ZN(U2822)
         );
  AOI22_X1 U7340 ( .A1(n4435), .A2(n6295), .B1(n6294), .B2(n6293), .ZN(n6311)
         );
  INV_X1 U7341 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6696) );
  INV_X1 U7342 ( .A(n6296), .ZN(n6299) );
  INV_X1 U7343 ( .A(n6306), .ZN(n6298) );
  OAI21_X1 U7344 ( .B1(n6299), .B2(n6298), .A(n6297), .ZN(n6328) );
  OAI22_X1 U7345 ( .A1(n6300), .A2(n6314), .B1(n6696), .B2(n6328), .ZN(n6301)
         );
  AOI211_X1 U7346 ( .C1(n6325), .C2(EBX_REG_4__SCAN_IN), .A(n6425), .B(n6301), 
        .ZN(n6310) );
  AOI22_X1 U7347 ( .A1(n6305), .A2(n6304), .B1(n6303), .B2(n6302), .ZN(n6309)
         );
  NAND3_X1 U7348 ( .A1(n6307), .A2(n6306), .A3(n6696), .ZN(n6308) );
  NAND4_X1 U7349 ( .A1(n6311), .A2(n6310), .A3(n6309), .A4(n6308), .ZN(U2823)
         );
  OR2_X1 U7350 ( .A1(n6312), .A2(n6693), .ZN(n6327) );
  INV_X1 U7351 ( .A(n6474), .ZN(n6317) );
  INV_X1 U7352 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6313) );
  OAI222_X1 U7353 ( .A1(n6318), .A2(n6317), .B1(n6316), .B2(n6315), .C1(n6314), 
        .C2(n6313), .ZN(n6324) );
  OAI22_X1 U7354 ( .A1(n6322), .A2(n6321), .B1(n6320), .B2(n6319), .ZN(n6323)
         );
  AOI211_X1 U7355 ( .C1(EBX_REG_3__SCAN_IN), .C2(n6325), .A(n6324), .B(n6323), 
        .ZN(n6326) );
  OAI221_X1 U7356 ( .B1(n6328), .B2(n6695), .C1(n6328), .C2(n6327), .A(n6326), 
        .ZN(U2824) );
  AOI22_X1 U7357 ( .A1(n6331), .A2(n6330), .B1(n6329), .B2(DATAI_17_), .ZN(
        n6335) );
  AOI22_X1 U7358 ( .A1(n6333), .A2(DATAI_1_), .B1(n6332), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6334) );
  NAND2_X1 U7359 ( .A1(n6335), .A2(n6334), .ZN(U2874) );
  INV_X1 U7360 ( .A(n6336), .ZN(n6339) );
  AOI22_X1 U7361 ( .A1(n6358), .A2(DATAO_REG_28__SCAN_IN), .B1(n6339), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n6337) );
  OAI21_X1 U7362 ( .B1(n6779), .B2(n7050), .A(n6337), .ZN(U2895) );
  INV_X1 U7363 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n7067) );
  AOI22_X1 U7364 ( .A1(n6339), .A2(EAX_REG_24__SCAN_IN), .B1(n6348), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n6338) );
  OAI21_X1 U7365 ( .B1(n7067), .B2(n4536), .A(n6338), .ZN(U2899) );
  AOI22_X1 U7366 ( .A1(n6358), .A2(DATAO_REG_18__SCAN_IN), .B1(n6339), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6340) );
  OAI21_X1 U7367 ( .B1(n6779), .B2(n7137), .A(n6340), .ZN(U2905) );
  INV_X1 U7368 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6424) );
  AOI22_X1 U7369 ( .A1(n6348), .A2(LWORD_REG_15__SCAN_IN), .B1(n6358), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6341) );
  OAI21_X1 U7370 ( .B1(n6424), .B2(n6360), .A(n6341), .ZN(U2908) );
  INV_X1 U7371 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n7096) );
  AOI22_X1 U7372 ( .A1(EAX_REG_14__SCAN_IN), .A2(n6349), .B1(n6348), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n6342) );
  OAI21_X1 U7373 ( .B1(n7096), .B2(n4536), .A(n6342), .ZN(U2909) );
  AOI22_X1 U7374 ( .A1(n6348), .A2(LWORD_REG_13__SCAN_IN), .B1(n6358), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6343) );
  OAI21_X1 U7375 ( .B1(n6418), .B2(n6360), .A(n6343), .ZN(U2910) );
  INV_X1 U7376 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n7064) );
  OAI222_X1 U7377 ( .A1(n6779), .A2(n6344), .B1(n6360), .B2(n7000), .C1(n7064), 
        .C2(n4536), .ZN(U2911) );
  AOI22_X1 U7378 ( .A1(n6348), .A2(LWORD_REG_11__SCAN_IN), .B1(n6358), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6345) );
  OAI21_X1 U7379 ( .B1(n7157), .B2(n6360), .A(n6345), .ZN(U2912) );
  INV_X1 U7380 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6412) );
  AOI22_X1 U7381 ( .A1(n6348), .A2(LWORD_REG_10__SCAN_IN), .B1(n6358), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6346) );
  OAI21_X1 U7382 ( .B1(n6412), .B2(n6360), .A(n6346), .ZN(U2913) );
  INV_X1 U7383 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6409) );
  AOI22_X1 U7384 ( .A1(n6348), .A2(LWORD_REG_9__SCAN_IN), .B1(
        DATAO_REG_9__SCAN_IN), .B2(n6358), .ZN(n6347) );
  OAI21_X1 U7385 ( .B1(n6409), .B2(n6360), .A(n6347), .ZN(U2914) );
  INV_X1 U7386 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n7101) );
  AOI22_X1 U7387 ( .A1(EAX_REG_8__SCAN_IN), .A2(n6349), .B1(n6348), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n6350) );
  OAI21_X1 U7388 ( .B1(n7101), .B2(n4536), .A(n6350), .ZN(U2915) );
  AOI22_X1 U7389 ( .A1(n6348), .A2(LWORD_REG_7__SCAN_IN), .B1(n6358), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6351) );
  OAI21_X1 U7390 ( .B1(n6404), .B2(n6360), .A(n6351), .ZN(U2916) );
  AOI22_X1 U7391 ( .A1(n6348), .A2(LWORD_REG_6__SCAN_IN), .B1(
        DATAO_REG_6__SCAN_IN), .B2(n6358), .ZN(n6352) );
  OAI21_X1 U7392 ( .B1(n3944), .B2(n6360), .A(n6352), .ZN(U2917) );
  AOI22_X1 U7393 ( .A1(n6348), .A2(LWORD_REG_5__SCAN_IN), .B1(n6358), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6353) );
  OAI21_X1 U7394 ( .B1(n3940), .B2(n6360), .A(n6353), .ZN(U2918) );
  INV_X1 U7395 ( .A(LWORD_REG_4__SCAN_IN), .ZN(n6354) );
  INV_X1 U7396 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n6972) );
  OAI222_X1 U7397 ( .A1(n6779), .A2(n6354), .B1(n6360), .B2(n6795), .C1(n6972), 
        .C2(n4536), .ZN(U2919) );
  INV_X1 U7398 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n7100) );
  OAI222_X1 U7399 ( .A1(n6779), .A2(n6815), .B1(n6360), .B2(n6355), .C1(n7100), 
        .C2(n4536), .ZN(U2920) );
  AOI22_X1 U7400 ( .A1(n6348), .A2(LWORD_REG_2__SCAN_IN), .B1(n6358), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6356) );
  OAI21_X1 U7401 ( .B1(n6397), .B2(n6360), .A(n6356), .ZN(U2921) );
  AOI22_X1 U7402 ( .A1(n6348), .A2(LWORD_REG_1__SCAN_IN), .B1(n6358), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6357) );
  OAI21_X1 U7403 ( .B1(n6394), .B2(n6360), .A(n6357), .ZN(U2922) );
  AOI22_X1 U7404 ( .A1(n6348), .A2(LWORD_REG_0__SCAN_IN), .B1(n6358), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6359) );
  OAI21_X1 U7405 ( .B1(n6391), .B2(n6360), .A(n6359), .ZN(U2923) );
  AND2_X1 U7406 ( .A1(n6422), .A2(DATAI_0_), .ZN(n6389) );
  AOI21_X1 U7407 ( .B1(UWORD_REG_0__SCAN_IN), .B2(n6416), .A(n6389), .ZN(n6361) );
  OAI21_X1 U7408 ( .B1(n6362), .B2(n6794), .A(n6361), .ZN(U2924) );
  AND2_X1 U7409 ( .A1(n6422), .A2(DATAI_1_), .ZN(n6392) );
  AOI21_X1 U7410 ( .B1(UWORD_REG_1__SCAN_IN), .B2(n6792), .A(n6392), .ZN(n6364) );
  OAI21_X1 U7411 ( .B1(n6365), .B2(n6794), .A(n6364), .ZN(U2925) );
  AOI21_X1 U7412 ( .B1(UWORD_REG_3__SCAN_IN), .B2(n6792), .A(n6366), .ZN(n6367) );
  OAI21_X1 U7413 ( .B1(n6368), .B2(n6794), .A(n6367), .ZN(U2927) );
  AND2_X1 U7414 ( .A1(n6422), .A2(DATAI_4_), .ZN(n6791) );
  AOI21_X1 U7415 ( .B1(UWORD_REG_4__SCAN_IN), .B2(n6792), .A(n6791), .ZN(n6369) );
  OAI21_X1 U7416 ( .B1(n6370), .B2(n6794), .A(n6369), .ZN(U2928) );
  AND2_X1 U7417 ( .A1(n6422), .A2(DATAI_5_), .ZN(n6398) );
  AOI21_X1 U7418 ( .B1(UWORD_REG_5__SCAN_IN), .B2(n6792), .A(n6398), .ZN(n6371) );
  OAI21_X1 U7419 ( .B1(n6372), .B2(n6794), .A(n6371), .ZN(U2929) );
  AND2_X1 U7420 ( .A1(n6422), .A2(DATAI_6_), .ZN(n6400) );
  AOI21_X1 U7421 ( .B1(UWORD_REG_6__SCAN_IN), .B2(n6792), .A(n6400), .ZN(n6373) );
  OAI21_X1 U7422 ( .B1(n7095), .B2(n6794), .A(n6373), .ZN(U2930) );
  AND2_X1 U7423 ( .A1(n6422), .A2(DATAI_7_), .ZN(n6402) );
  AOI21_X1 U7424 ( .B1(UWORD_REG_7__SCAN_IN), .B2(n6792), .A(n6402), .ZN(n6374) );
  OAI21_X1 U7425 ( .B1(n6375), .B2(n6794), .A(n6374), .ZN(U2931) );
  AOI22_X1 U7426 ( .A1(n6792), .A2(UWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_24__SCAN_IN), .B2(n6419), .ZN(n6376) );
  NAND2_X1 U7427 ( .A1(n6422), .A2(DATAI_8_), .ZN(n6405) );
  NAND2_X1 U7428 ( .A1(n6376), .A2(n6405), .ZN(U2932) );
  INV_X1 U7429 ( .A(DATAI_9_), .ZN(n6377) );
  NOR2_X1 U7430 ( .A1(n6421), .A2(n6377), .ZN(n6407) );
  AOI21_X1 U7431 ( .B1(UWORD_REG_9__SCAN_IN), .B2(n6792), .A(n6407), .ZN(n6378) );
  OAI21_X1 U7432 ( .B1(n6379), .B2(n6794), .A(n6378), .ZN(U2933) );
  INV_X1 U7433 ( .A(DATAI_10_), .ZN(n6380) );
  NOR2_X1 U7434 ( .A1(n6421), .A2(n6380), .ZN(n6410) );
  AOI21_X1 U7435 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n6792), .A(n6410), .ZN(
        n6381) );
  OAI21_X1 U7436 ( .B1(n6382), .B2(n6794), .A(n6381), .ZN(U2934) );
  AND2_X1 U7437 ( .A1(n6422), .A2(DATAI_11_), .ZN(n6413) );
  AOI21_X1 U7438 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n6792), .A(n6413), .ZN(
        n6383) );
  OAI21_X1 U7439 ( .B1(n6384), .B2(n6794), .A(n6383), .ZN(U2935) );
  AND2_X1 U7440 ( .A1(n6422), .A2(DATAI_13_), .ZN(n6415) );
  AOI21_X1 U7441 ( .B1(UWORD_REG_13__SCAN_IN), .B2(n6792), .A(n6415), .ZN(
        n6385) );
  OAI21_X1 U7442 ( .B1(n6386), .B2(n6794), .A(n6385), .ZN(U2937) );
  AOI22_X1 U7443 ( .A1(n6792), .A2(UWORD_REG_14__SCAN_IN), .B1(n6422), .B2(
        DATAI_14_), .ZN(n6387) );
  OAI21_X1 U7444 ( .B1(n6388), .B2(n6794), .A(n6387), .ZN(U2938) );
  AOI21_X1 U7445 ( .B1(LWORD_REG_0__SCAN_IN), .B2(n6792), .A(n6389), .ZN(n6390) );
  OAI21_X1 U7446 ( .B1(n6391), .B2(n6794), .A(n6390), .ZN(U2939) );
  AOI21_X1 U7447 ( .B1(LWORD_REG_1__SCAN_IN), .B2(n6792), .A(n6392), .ZN(n6393) );
  OAI21_X1 U7448 ( .B1(n6394), .B2(n6794), .A(n6393), .ZN(U2940) );
  AOI21_X1 U7449 ( .B1(LWORD_REG_2__SCAN_IN), .B2(n6792), .A(n6395), .ZN(n6396) );
  OAI21_X1 U7450 ( .B1(n6397), .B2(n6794), .A(n6396), .ZN(U2941) );
  AOI21_X1 U7451 ( .B1(LWORD_REG_5__SCAN_IN), .B2(n6792), .A(n6398), .ZN(n6399) );
  OAI21_X1 U7452 ( .B1(n3940), .B2(n6794), .A(n6399), .ZN(U2944) );
  AOI21_X1 U7453 ( .B1(LWORD_REG_6__SCAN_IN), .B2(n6792), .A(n6400), .ZN(n6401) );
  OAI21_X1 U7454 ( .B1(n3944), .B2(n6794), .A(n6401), .ZN(U2945) );
  AOI21_X1 U7455 ( .B1(LWORD_REG_7__SCAN_IN), .B2(n6416), .A(n6402), .ZN(n6403) );
  OAI21_X1 U7456 ( .B1(n6404), .B2(n6794), .A(n6403), .ZN(U2946) );
  AOI22_X1 U7457 ( .A1(n6792), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n6419), .ZN(n6406) );
  NAND2_X1 U7458 ( .A1(n6406), .A2(n6405), .ZN(U2947) );
  AOI21_X1 U7459 ( .B1(LWORD_REG_9__SCAN_IN), .B2(n6416), .A(n6407), .ZN(n6408) );
  OAI21_X1 U7460 ( .B1(n6409), .B2(n6794), .A(n6408), .ZN(U2948) );
  AOI21_X1 U7461 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n6416), .A(n6410), .ZN(
        n6411) );
  OAI21_X1 U7462 ( .B1(n6412), .B2(n6794), .A(n6411), .ZN(U2949) );
  AOI21_X1 U7463 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n6416), .A(n6413), .ZN(
        n6414) );
  OAI21_X1 U7464 ( .B1(n7157), .B2(n6794), .A(n6414), .ZN(U2950) );
  AOI21_X1 U7465 ( .B1(LWORD_REG_13__SCAN_IN), .B2(n6416), .A(n6415), .ZN(
        n6417) );
  OAI21_X1 U7466 ( .B1(n6418), .B2(n6794), .A(n6417), .ZN(U2952) );
  INV_X1 U7467 ( .A(DATAI_14_), .ZN(n7119) );
  AOI22_X1 U7468 ( .A1(n6792), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n6419), .ZN(n6420) );
  OAI21_X1 U7469 ( .B1(n6421), .B2(n7119), .A(n6420), .ZN(U2953) );
  AOI22_X1 U7470 ( .A1(n6792), .A2(LWORD_REG_15__SCAN_IN), .B1(n6422), .B2(
        DATAI_15_), .ZN(n6423) );
  OAI21_X1 U7471 ( .B1(n6424), .B2(n6794), .A(n6423), .ZN(U2954) );
  AOI22_X1 U7472 ( .A1(n6425), .A2(REIP_REG_2__SCAN_IN), .B1(n6442), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6435) );
  NAND2_X1 U7473 ( .A1(n6426), .A2(n6427), .ZN(n6430) );
  INV_X1 U7474 ( .A(n6428), .ZN(n6429) );
  XNOR2_X1 U7475 ( .A(n6430), .B(n6429), .ZN(n6493) );
  AOI22_X1 U7476 ( .A1(n6433), .A2(n6432), .B1(n6493), .B2(n6431), .ZN(n6434)
         );
  OAI211_X1 U7477 ( .C1(n6437), .C2(n6436), .A(n6435), .B(n6434), .ZN(U2984)
         );
  OAI22_X1 U7478 ( .A1(n6439), .A2(n6438), .B1(n6498), .B2(n6769), .ZN(n6440)
         );
  INV_X1 U7479 ( .A(n6440), .ZN(n6444) );
  OAI21_X1 U7480 ( .B1(n6442), .B2(n6441), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n6443) );
  OAI211_X1 U7481 ( .C1(n6445), .C2(n5714), .A(n6444), .B(n6443), .ZN(U2986)
         );
  INV_X1 U7482 ( .A(n6446), .ZN(n6447) );
  AOI21_X1 U7483 ( .B1(n6503), .B2(n6448), .A(n6447), .ZN(n6452) );
  AOI22_X1 U7484 ( .A1(n6507), .A2(n6450), .B1(n7122), .B2(n6449), .ZN(n6451)
         );
  OAI211_X1 U7485 ( .C1(n6453), .C2(n7122), .A(n6452), .B(n6451), .ZN(U3007)
         );
  INV_X1 U7486 ( .A(n6454), .ZN(n6456) );
  AOI21_X1 U7487 ( .B1(n6503), .B2(n6456), .A(n6455), .ZN(n6460) );
  AOI22_X1 U7488 ( .A1(n6458), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .B1(n6507), 
        .B2(n6457), .ZN(n6459) );
  OAI211_X1 U7489 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6461), .A(n6460), 
        .B(n6459), .ZN(U3009) );
  INV_X1 U7490 ( .A(n6462), .ZN(n6466) );
  NAND2_X1 U7491 ( .A1(n6503), .A2(n6463), .ZN(n6465) );
  OAI211_X1 U7492 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n6466), .A(n6465), 
        .B(n6464), .ZN(n6467) );
  AOI21_X1 U7493 ( .B1(n6468), .B2(n6507), .A(n6467), .ZN(n6469) );
  OAI21_X1 U7494 ( .B1(n6471), .B2(n6470), .A(n6469), .ZN(U3011) );
  INV_X1 U7495 ( .A(n6472), .ZN(n6483) );
  AOI21_X1 U7496 ( .B1(n6503), .B2(n6474), .A(n6473), .ZN(n6478) );
  OR2_X1 U7497 ( .A1(n6476), .A2(n6475), .ZN(n6477) );
  OAI211_X1 U7498 ( .C1(n6479), .C2(INSTADDRPOINTER_REG_3__SCAN_IN), .A(n6478), 
        .B(n6477), .ZN(n6480) );
  INV_X1 U7499 ( .A(n6480), .ZN(n6481) );
  OAI21_X1 U7500 ( .B1(n6483), .B2(n6482), .A(n6481), .ZN(U3015) );
  INV_X1 U7501 ( .A(n6484), .ZN(n6489) );
  OAI21_X1 U7502 ( .B1(n6486), .B2(n7025), .A(n6485), .ZN(n6487) );
  AOI22_X1 U7503 ( .A1(n6489), .A2(n6503), .B1(n6488), .B2(n6487), .ZN(n6497)
         );
  OAI33_X1 U7505 ( .A1(1'b0), .A2(n6491), .A3(n3631), .B1(
        INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6490), .B3(n6510), .ZN(n6495) );
  AND2_X1 U7506 ( .A1(n6493), .A2(n6507), .ZN(n6494) );
  NOR2_X1 U7507 ( .A1(n6495), .A2(n6494), .ZN(n6496) );
  OAI211_X1 U7508 ( .C1(n6498), .C2(n6693), .A(n6497), .B(n6496), .ZN(U3016)
         );
  AOI21_X1 U7509 ( .B1(n6499), .B2(n7025), .A(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .ZN(n6500) );
  NAND2_X1 U7510 ( .A1(n6501), .A2(n6500), .ZN(n6505) );
  AOI22_X1 U7511 ( .A1(n6503), .A2(n6502), .B1(n6425), .B2(REIP_REG_1__SCAN_IN), .ZN(n6504) );
  NAND2_X1 U7512 ( .A1(n6505), .A2(n6504), .ZN(n6506) );
  AOI21_X1 U7513 ( .B1(n6508), .B2(n6507), .A(n6506), .ZN(n6509) );
  OAI21_X1 U7514 ( .B1(n6511), .B2(n6510), .A(n6509), .ZN(U3017) );
  NOR2_X1 U7515 ( .A1(n6512), .A2(n6763), .ZN(U3019) );
  NOR3_X1 U7516 ( .A1(n6514), .A2(n6513), .A3(n3230), .ZN(n6516) );
  INV_X1 U7517 ( .A(n6515), .ZN(n6552) );
  NOR2_X1 U7518 ( .A1(n6516), .A2(n6552), .ZN(n6520) );
  NOR2_X1 U7519 ( .A1(n6520), .A2(n6571), .ZN(n6517) );
  AOI21_X1 U7520 ( .B1(n6524), .B2(STATE2_REG_2__SCAN_IN), .A(n6517), .ZN(
        n6560) );
  AOI22_X1 U7521 ( .A1(n6553), .A2(n6518), .B1(n6552), .B2(n6562), .ZN(n6526)
         );
  INV_X1 U7522 ( .A(n6758), .ZN(n6521) );
  NAND3_X1 U7523 ( .A1(n6521), .A2(n6564), .A3(n6520), .ZN(n6523) );
  OAI211_X1 U7524 ( .C1(n6524), .C2(n6564), .A(n6523), .B(n6522), .ZN(n6556)
         );
  AOI22_X1 U7525 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6556), .B1(n6563), 
        .B2(n6554), .ZN(n6525) );
  OAI211_X1 U7526 ( .C1(n6560), .C2(n6527), .A(n6526), .B(n6525), .ZN(U3076)
         );
  AOI22_X1 U7527 ( .A1(n6554), .A2(n6528), .B1(n6552), .B2(n3259), .ZN(n6530)
         );
  AOI22_X1 U7528 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6556), .B1(n6582), 
        .B2(n6553), .ZN(n6529) );
  OAI211_X1 U7529 ( .C1(n6560), .C2(n6531), .A(n6530), .B(n6529), .ZN(U3077)
         );
  AOI22_X1 U7530 ( .A1(n6554), .A2(n6588), .B1(n6552), .B2(n6587), .ZN(n6534)
         );
  AOI22_X1 U7531 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6556), .B1(n6532), 
        .B2(n6553), .ZN(n6533) );
  OAI211_X1 U7532 ( .C1(n6560), .C2(n6535), .A(n6534), .B(n6533), .ZN(U3078)
         );
  AOI22_X1 U7533 ( .A1(n6554), .A2(n6536), .B1(n6552), .B2(n6593), .ZN(n6538)
         );
  AOI22_X1 U7534 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6556), .B1(n6594), 
        .B2(n6553), .ZN(n6537) );
  OAI211_X1 U7535 ( .C1(n6560), .C2(n6539), .A(n6538), .B(n6537), .ZN(U3079)
         );
  AOI22_X1 U7536 ( .A1(n6553), .A2(n6540), .B1(n6552), .B2(n6599), .ZN(n6542)
         );
  AOI22_X1 U7537 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6556), .B1(n6600), 
        .B2(n6554), .ZN(n6541) );
  OAI211_X1 U7538 ( .C1(n6560), .C2(n6543), .A(n6542), .B(n6541), .ZN(U3080)
         );
  AOI22_X1 U7539 ( .A1(n6554), .A2(n6606), .B1(n6552), .B2(n6605), .ZN(n6546)
         );
  AOI22_X1 U7540 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6556), .B1(n6544), 
        .B2(n6553), .ZN(n6545) );
  OAI211_X1 U7541 ( .C1(n6560), .C2(n6547), .A(n6546), .B(n6545), .ZN(U3081)
         );
  AOI22_X1 U7542 ( .A1(n6554), .A2(n6612), .B1(n6552), .B2(n6611), .ZN(n6550)
         );
  AOI22_X1 U7543 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6556), .B1(n6548), 
        .B2(n6553), .ZN(n6549) );
  OAI211_X1 U7544 ( .C1(n6560), .C2(n6551), .A(n6550), .B(n6549), .ZN(U3082)
         );
  AOI22_X1 U7545 ( .A1(n6553), .A2(n6621), .B1(n6552), .B2(n6620), .ZN(n6558)
         );
  AOI22_X1 U7546 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6556), .B1(n6555), 
        .B2(n6554), .ZN(n6557) );
  OAI211_X1 U7547 ( .C1(n6560), .C2(n6559), .A(n6558), .B(n6557), .ZN(U3083)
         );
  NOR2_X1 U7548 ( .A1(n6561), .A2(n6765), .ZN(n6619) );
  AOI22_X1 U7549 ( .A1(n6613), .A2(n6563), .B1(n6562), .B2(n6619), .ZN(n6579)
         );
  OAI21_X1 U7550 ( .B1(n6566), .B2(n6565), .A(n6564), .ZN(n6576) );
  OR2_X1 U7551 ( .A1(n6567), .A2(n3230), .ZN(n6569) );
  INV_X1 U7552 ( .A(n6619), .ZN(n6568) );
  AND2_X1 U7553 ( .A1(n6569), .A2(n6568), .ZN(n6575) );
  INV_X1 U7554 ( .A(n6575), .ZN(n6573) );
  AOI21_X1 U7555 ( .B1(n6571), .B2(n6574), .A(n6570), .ZN(n6572) );
  OAI21_X1 U7556 ( .B1(n6576), .B2(n6573), .A(n6572), .ZN(n6625) );
  OAI22_X1 U7557 ( .A1(n6576), .A2(n6575), .B1(n6574), .B2(n6780), .ZN(n6623)
         );
  AOI22_X1 U7558 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6625), .B1(n6577), 
        .B2(n6623), .ZN(n6578) );
  OAI211_X1 U7559 ( .C1(n6580), .C2(n6617), .A(n6579), .B(n6578), .ZN(U3108)
         );
  AOI22_X1 U7560 ( .A1(n6622), .A2(n6582), .B1(n3259), .B2(n6619), .ZN(n6585)
         );
  AOI22_X1 U7561 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6625), .B1(n6583), 
        .B2(n6623), .ZN(n6584) );
  OAI211_X1 U7562 ( .C1(n6586), .C2(n6628), .A(n6585), .B(n6584), .ZN(U3109)
         );
  AOI22_X1 U7563 ( .A1(n6613), .A2(n6588), .B1(n6587), .B2(n6619), .ZN(n6591)
         );
  AOI22_X1 U7564 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6625), .B1(n6589), 
        .B2(n6623), .ZN(n6590) );
  OAI211_X1 U7565 ( .C1(n6592), .C2(n6617), .A(n6591), .B(n6590), .ZN(U3110)
         );
  AOI22_X1 U7566 ( .A1(n6622), .A2(n6594), .B1(n6593), .B2(n6619), .ZN(n6597)
         );
  AOI22_X1 U7567 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6625), .B1(n6595), 
        .B2(n6623), .ZN(n6596) );
  OAI211_X1 U7568 ( .C1(n6598), .C2(n6628), .A(n6597), .B(n6596), .ZN(U3111)
         );
  AOI22_X1 U7569 ( .A1(n6613), .A2(n6600), .B1(n6599), .B2(n6619), .ZN(n6603)
         );
  AOI22_X1 U7570 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6625), .B1(n6601), 
        .B2(n6623), .ZN(n6602) );
  OAI211_X1 U7571 ( .C1(n6604), .C2(n6617), .A(n6603), .B(n6602), .ZN(U3112)
         );
  AOI22_X1 U7572 ( .A1(n6613), .A2(n6606), .B1(n6605), .B2(n6619), .ZN(n6609)
         );
  AOI22_X1 U7573 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6625), .B1(n6607), 
        .B2(n6623), .ZN(n6608) );
  OAI211_X1 U7574 ( .C1(n6610), .C2(n6617), .A(n6609), .B(n6608), .ZN(U3113)
         );
  AOI22_X1 U7575 ( .A1(n6613), .A2(n6612), .B1(n6611), .B2(n6619), .ZN(n6616)
         );
  AOI22_X1 U7576 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6625), .B1(n6614), 
        .B2(n6623), .ZN(n6615) );
  OAI211_X1 U7577 ( .C1(n6618), .C2(n6617), .A(n6616), .B(n6615), .ZN(U3114)
         );
  AOI22_X1 U7578 ( .A1(n6622), .A2(n6621), .B1(n6620), .B2(n6619), .ZN(n6627)
         );
  AOI22_X1 U7579 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6625), .B1(n6624), 
        .B2(n6623), .ZN(n6626) );
  OAI211_X1 U7580 ( .C1(n6629), .C2(n6628), .A(n6627), .B(n6626), .ZN(U3115)
         );
  OAI22_X1 U7581 ( .A1(n3230), .A2(n6631), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6630), .ZN(n6748) );
  NAND2_X1 U7582 ( .A1(n6632), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6756) );
  INV_X1 U7583 ( .A(n6756), .ZN(n6634) );
  NOR3_X1 U7584 ( .A1(n6748), .A2(n6634), .A3(n6633), .ZN(n6640) );
  INV_X1 U7585 ( .A(n6640), .ZN(n6638) );
  OAI211_X1 U7586 ( .C1(n6638), .C2(n6637), .A(n6636), .B(n6635), .ZN(n6639)
         );
  OAI21_X1 U7587 ( .B1(n6640), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n6639), 
        .ZN(n6641) );
  AOI222_X1 U7588 ( .A1(n6643), .A2(n6642), .B1(n6643), .B2(n6641), .C1(n6642), 
        .C2(n6641), .ZN(n6645) );
  OAI21_X1 U7589 ( .B1(n6645), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n6644), 
        .ZN(n6653) );
  AOI21_X1 U7590 ( .B1(n6645), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6652) );
  OAI21_X1 U7591 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6646), 
        .ZN(n6649) );
  NAND3_X1 U7592 ( .A1(n6649), .A2(n6648), .A3(n6647), .ZN(n6650) );
  AOI211_X1 U7593 ( .C1(n6653), .C2(n6652), .A(n6651), .B(n6650), .ZN(n6663)
         );
  AOI22_X1 U7594 ( .A1(n6663), .A2(n6664), .B1(READY_N), .B2(n6348), .ZN(n6654) );
  AOI21_X1 U7595 ( .B1(n6656), .B2(n6655), .A(n6654), .ZN(n6746) );
  AOI211_X1 U7596 ( .C1(n6657), .C2(n6787), .A(STATE2_REG_0__SCAN_IN), .B(
        n6746), .ZN(n6658) );
  AOI211_X1 U7597 ( .C1(n6744), .C2(n6660), .A(n6659), .B(n6658), .ZN(n6661)
         );
  OAI221_X1 U7598 ( .B1(n6746), .B2(READY_N), .C1(n6746), .C2(n6780), .A(
        STATE2_REG_0__SCAN_IN), .ZN(n6671) );
  OAI211_X1 U7599 ( .C1(n6663), .C2(n6662), .A(n6661), .B(n6671), .ZN(U3148)
         );
  NOR2_X1 U7600 ( .A1(READY_N), .A2(n6783), .ZN(n6674) );
  AOI21_X1 U7601 ( .B1(n6665), .B2(n6674), .A(n6664), .ZN(n6666) );
  NOR2_X1 U7602 ( .A1(n6666), .A2(n6746), .ZN(n6667) );
  AOI211_X1 U7603 ( .C1(n6746), .C2(n6669), .A(n6668), .B(n6667), .ZN(n6670)
         );
  OAI21_X1 U7604 ( .B1(n6749), .B2(n6671), .A(n6670), .ZN(U3149) );
  OAI211_X1 U7605 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6674), .A(n6673), .B(
        n6672), .ZN(n6675) );
  NAND2_X1 U7606 ( .A1(n6676), .A2(n6675), .ZN(U3150) );
  AND2_X1 U7607 ( .A1(n6741), .A2(DATAWIDTH_REG_31__SCAN_IN), .ZN(U3151) );
  AND2_X1 U7608 ( .A1(n6741), .A2(DATAWIDTH_REG_30__SCAN_IN), .ZN(U3152) );
  NOR2_X1 U7609 ( .A1(n6743), .A2(n7173), .ZN(U3153) );
  AND2_X1 U7610 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6741), .ZN(U3154) );
  AND2_X1 U7611 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6741), .ZN(U3155) );
  AND2_X1 U7612 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6741), .ZN(U3156) );
  AND2_X1 U7613 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6741), .ZN(U3157) );
  INV_X1 U7614 ( .A(DATAWIDTH_REG_24__SCAN_IN), .ZN(n6963) );
  NOR2_X1 U7615 ( .A1(n6743), .A2(n6963), .ZN(U3158) );
  AND2_X1 U7616 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6741), .ZN(U3159) );
  AND2_X1 U7617 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6741), .ZN(U3160) );
  AND2_X1 U7618 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6741), .ZN(U3161) );
  AND2_X1 U7619 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6741), .ZN(U3162) );
  AND2_X1 U7620 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6741), .ZN(U3163) );
  AND2_X1 U7621 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6741), .ZN(U3164) );
  AND2_X1 U7622 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6741), .ZN(U3165) );
  AND2_X1 U7623 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6741), .ZN(U3166) );
  AND2_X1 U7624 ( .A1(n6741), .A2(DATAWIDTH_REG_15__SCAN_IN), .ZN(U3167) );
  AND2_X1 U7625 ( .A1(n6741), .A2(DATAWIDTH_REG_14__SCAN_IN), .ZN(U3168) );
  AND2_X1 U7626 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6741), .ZN(U3169) );
  AND2_X1 U7627 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6741), .ZN(U3170) );
  AND2_X1 U7628 ( .A1(n6741), .A2(DATAWIDTH_REG_11__SCAN_IN), .ZN(U3171) );
  AND2_X1 U7629 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6741), .ZN(U3172) );
  AND2_X1 U7630 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6741), .ZN(U3173) );
  AND2_X1 U7631 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6741), .ZN(U3174) );
  NOR2_X1 U7632 ( .A1(n6743), .A2(n7151), .ZN(U3175) );
  AND2_X1 U7633 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6741), .ZN(U3176) );
  AND2_X1 U7634 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6741), .ZN(U3177) );
  INV_X1 U7635 ( .A(DATAWIDTH_REG_4__SCAN_IN), .ZN(n7034) );
  NOR2_X1 U7636 ( .A1(n6743), .A2(n7034), .ZN(U3178) );
  AND2_X1 U7637 ( .A1(n6741), .A2(DATAWIDTH_REG_3__SCAN_IN), .ZN(U3179) );
  AND2_X1 U7638 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6741), .ZN(U3180) );
  NOR2_X1 U7639 ( .A1(n6682), .A2(n6691), .ZN(n6685) );
  AOI22_X1 U7640 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6688) );
  AND2_X1 U7641 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6679) );
  INV_X1 U7642 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6984) );
  INV_X1 U7643 ( .A(NA_N), .ZN(n6960) );
  AOI211_X1 U7644 ( .C1(STATE_REG_2__SCAN_IN), .C2(n6960), .A(
        STATE_REG_0__SCAN_IN), .B(n6685), .ZN(n6690) );
  AOI221_X1 U7645 ( .B1(n6679), .B2(n6732), .C1(n6984), .C2(n6732), .A(n6690), 
        .ZN(n6677) );
  OAI21_X1 U7646 ( .B1(n6685), .B2(n6688), .A(n6677), .ZN(U3181) );
  NOR2_X1 U7647 ( .A1(n7054), .A2(n6984), .ZN(n6686) );
  NAND2_X1 U7648 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6678) );
  OAI21_X1 U7649 ( .B1(n6686), .B2(n6679), .A(n6678), .ZN(n6680) );
  OAI211_X1 U7650 ( .C1(n6682), .C2(n6683), .A(n6681), .B(n6680), .ZN(U3182)
         );
  AOI221_X1 U7651 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6683), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6684) );
  AOI221_X1 U7652 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6684), .C2(HOLD), .A(n7054), .ZN(n6689) );
  AOI21_X1 U7653 ( .B1(n6686), .B2(n6960), .A(n6685), .ZN(n6687) );
  OAI22_X1 U7654 ( .A1(n6690), .A2(n6689), .B1(n6688), .B2(n6687), .ZN(U3183)
         );
  NAND2_X1 U7655 ( .A1(n6790), .A2(n6691), .ZN(n6737) );
  INV_X1 U7656 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n7163) );
  NAND2_X1 U7657 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6790), .ZN(n6735) );
  OAI222_X1 U7658 ( .A1(n6737), .A2(n6693), .B1(n7163), .B2(n6790), .C1(n6775), 
        .C2(n6735), .ZN(U3184) );
  INV_X1 U7659 ( .A(n6737), .ZN(n6729) );
  AOI22_X1 U7660 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6729), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6732), .ZN(n6692) );
  OAI21_X1 U7661 ( .B1(n6693), .B2(n6735), .A(n6692), .ZN(U3185) );
  AOI22_X1 U7662 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6729), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6732), .ZN(n6694) );
  OAI21_X1 U7663 ( .B1(n6695), .B2(n6735), .A(n6694), .ZN(U3186) );
  INV_X1 U7664 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n7052) );
  OAI222_X1 U7665 ( .A1(n6735), .A2(n6696), .B1(n7052), .B2(n6790), .C1(n6698), 
        .C2(n6737), .ZN(U3187) );
  AOI22_X1 U7666 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6729), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6732), .ZN(n6697) );
  OAI21_X1 U7667 ( .B1(n6698), .B2(n6735), .A(n6697), .ZN(U3188) );
  INV_X1 U7668 ( .A(n6735), .ZN(n6733) );
  AOI22_X1 U7669 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6738), .ZN(n6699) );
  OAI21_X1 U7670 ( .B1(n7170), .B2(n6737), .A(n6699), .ZN(U3189) );
  AOI22_X1 U7671 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6738), .ZN(n6700) );
  OAI21_X1 U7672 ( .B1(n6701), .B2(n6737), .A(n6700), .ZN(U3190) );
  INV_X1 U7673 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n7142) );
  OAI222_X1 U7674 ( .A1(n6737), .A2(n5159), .B1(n7142), .B2(n6790), .C1(n6701), 
        .C2(n6735), .ZN(U3191) );
  INV_X1 U7675 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n7070) );
  OAI222_X1 U7676 ( .A1(n6737), .A2(n6703), .B1(n7070), .B2(n6790), .C1(n5159), 
        .C2(n6735), .ZN(U3192) );
  INV_X1 U7677 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n7118) );
  OAI222_X1 U7678 ( .A1(n6735), .A2(n6703), .B1(n7118), .B2(n6790), .C1(n6702), 
        .C2(n6737), .ZN(U3193) );
  AOI22_X1 U7679 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6738), .ZN(n6704) );
  OAI21_X1 U7680 ( .B1(n6706), .B2(n6737), .A(n6704), .ZN(U3194) );
  INV_X1 U7681 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n6705) );
  OAI222_X1 U7682 ( .A1(n6735), .A2(n6706), .B1(n6705), .B2(n6790), .C1(n5386), 
        .C2(n6737), .ZN(U3195) );
  AOI22_X1 U7683 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6729), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6738), .ZN(n6707) );
  OAI21_X1 U7684 ( .B1(n5386), .B2(n6735), .A(n6707), .ZN(U3196) );
  AOI22_X1 U7685 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6732), .ZN(n6708) );
  OAI21_X1 U7686 ( .B1(n6709), .B2(n6737), .A(n6708), .ZN(U3197) );
  AOI22_X1 U7687 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6732), .ZN(n6710) );
  OAI21_X1 U7688 ( .B1(n6712), .B2(n6737), .A(n6710), .ZN(U3198) );
  AOI22_X1 U7689 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6729), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6738), .ZN(n6711) );
  OAI21_X1 U7690 ( .B1(n6712), .B2(n6735), .A(n6711), .ZN(U3199) );
  AOI22_X1 U7691 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6732), .ZN(n6713) );
  OAI21_X1 U7692 ( .B1(n6714), .B2(n6737), .A(n6713), .ZN(U3200) );
  INV_X1 U7693 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n7135) );
  INV_X1 U7694 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6716) );
  OAI222_X1 U7695 ( .A1(n6735), .A2(n6714), .B1(n7135), .B2(n6790), .C1(n6716), 
        .C2(n6737), .ZN(U3201) );
  AOI22_X1 U7696 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6729), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6738), .ZN(n6715) );
  OAI21_X1 U7697 ( .B1(n6716), .B2(n6735), .A(n6715), .ZN(U3202) );
  INV_X1 U7698 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6719) );
  AOI22_X1 U7699 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6732), .ZN(n6717) );
  OAI21_X1 U7700 ( .B1(n6719), .B2(n6737), .A(n6717), .ZN(U3203) );
  AOI22_X1 U7701 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6729), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6732), .ZN(n6718) );
  OAI21_X1 U7702 ( .B1(n6719), .B2(n6735), .A(n6718), .ZN(U3204) );
  AOI22_X1 U7703 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6732), .ZN(n6720) );
  OAI21_X1 U7704 ( .B1(n6722), .B2(n6737), .A(n6720), .ZN(U3205) );
  AOI22_X1 U7705 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6729), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6732), .ZN(n6721) );
  OAI21_X1 U7706 ( .B1(n6722), .B2(n6735), .A(n6721), .ZN(U3206) );
  AOI22_X1 U7707 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6732), .ZN(n6723) );
  OAI21_X1 U7708 ( .B1(n6724), .B2(n6737), .A(n6723), .ZN(U3207) );
  AOI22_X1 U7709 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6732), .ZN(n6725) );
  OAI21_X1 U7710 ( .B1(n6727), .B2(n6737), .A(n6725), .ZN(U3208) );
  AOI22_X1 U7711 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6729), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6732), .ZN(n6726) );
  OAI21_X1 U7712 ( .B1(n6727), .B2(n6735), .A(n6726), .ZN(U3209) );
  AOI22_X1 U7713 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6732), .ZN(n6728) );
  OAI21_X1 U7714 ( .B1(n6731), .B2(n6737), .A(n6728), .ZN(U3210) );
  AOI22_X1 U7715 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6729), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6732), .ZN(n6730) );
  OAI21_X1 U7716 ( .B1(n6731), .B2(n6735), .A(n6730), .ZN(U3211) );
  AOI22_X1 U7717 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6733), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6732), .ZN(n6734) );
  OAI21_X1 U7718 ( .B1(n5507), .B2(n6737), .A(n6734), .ZN(U3212) );
  INV_X1 U7719 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6736) );
  INV_X1 U7720 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n7103) );
  OAI222_X1 U7721 ( .A1(n6737), .A2(n6736), .B1(n7103), .B2(n6790), .C1(n5507), 
        .C2(n6735), .ZN(U3213) );
  MUX2_X1 U7722 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6790), .Z(U3445) );
  MUX2_X1 U7723 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6790), .Z(U3446) );
  MUX2_X1 U7724 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6790), .Z(U3447) );
  INV_X1 U7725 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6739) );
  INV_X1 U7726 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n7128) );
  AOI22_X1 U7727 ( .A1(n6790), .A2(n6739), .B1(n7128), .B2(n6738), .ZN(U3448)
         );
  INV_X1 U7728 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n7155) );
  INV_X1 U7729 ( .A(n6742), .ZN(n6740) );
  AOI21_X1 U7730 ( .B1(n7155), .B2(n6741), .A(n6740), .ZN(U3451) );
  INV_X1 U7731 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6768) );
  OAI21_X1 U7732 ( .B1(n6743), .B2(n6768), .A(n6742), .ZN(U3452) );
  AOI211_X1 U7733 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6746), .A(n6745), .B(
        n6744), .ZN(n6747) );
  INV_X1 U7734 ( .A(n6747), .ZN(U3453) );
  INV_X1 U7735 ( .A(n6748), .ZN(n6750) );
  OAI22_X1 U7736 ( .A1(n6750), .A2(n6755), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6749), .ZN(n6752) );
  OAI22_X1 U7737 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6753), .B1(n6752), .B2(n6751), .ZN(n6754) );
  OAI21_X1 U7738 ( .B1(n6756), .B2(n6755), .A(n6754), .ZN(U3461) );
  OR2_X1 U7739 ( .A1(n6759), .A2(n6758), .ZN(n6760) );
  AOI222_X1 U7740 ( .A1(n6762), .A2(n4582), .B1(n6757), .B2(n6761), .C1(n6760), 
        .C2(n6564), .ZN(n6764) );
  AOI22_X1 U7741 ( .A1(n6766), .A2(n6765), .B1(n6764), .B2(n6763), .ZN(U3462)
         );
  AOI221_X1 U7742 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6769), .C1(n7155), 
        .C2(n6768), .A(n6767), .ZN(n6771) );
  OAI22_X1 U7743 ( .A1(n6773), .A2(BYTEENABLE_REG_2__SCAN_IN), .B1(n6775), 
        .B2(n6772), .ZN(n6770) );
  NOR2_X1 U7744 ( .A1(n6771), .A2(n6770), .ZN(U3468) );
  OAI21_X1 U7745 ( .B1(n6773), .B2(BYTEENABLE_REG_0__SCAN_IN), .A(n6772), .ZN(
        n6774) );
  OAI21_X1 U7746 ( .B1(n6776), .B2(n6775), .A(n6774), .ZN(U3469) );
  INV_X1 U7747 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n7169) );
  MUX2_X1 U7748 ( .A(W_R_N_REG_SCAN_IN), .B(n7169), .S(n6790), .Z(U3470) );
  OAI211_X1 U7749 ( .C1(READY_N), .C2(n6779), .A(n6778), .B(n6777), .ZN(n6789)
         );
  AOI21_X1 U7750 ( .B1(n6782), .B2(n6781), .A(n6780), .ZN(n6784) );
  AOI21_X1 U7751 ( .B1(n6785), .B2(n6784), .A(n6783), .ZN(n6786) );
  OAI21_X1 U7752 ( .B1(n6787), .B2(n6786), .A(n6789), .ZN(n6788) );
  OAI21_X1 U7753 ( .B1(n6789), .B2(n6984), .A(n6788), .ZN(U3472) );
  MUX2_X1 U7754 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6790), .Z(U3473) );
  AOI21_X1 U7755 ( .B1(LWORD_REG_4__SCAN_IN), .B2(n6792), .A(n6791), .ZN(n6793) );
  OAI21_X1 U7756 ( .B1(n6795), .B2(n6794), .A(n6793), .ZN(n7189) );
  OAI22_X1 U7757 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(keyinput102), .B1(
        keyinput85), .B2(DATAI_28_), .ZN(n6796) );
  AOI221_X1 U7758 ( .B1(INSTQUEUE_REG_7__0__SCAN_IN), .B2(keyinput102), .C1(
        DATAI_28_), .C2(keyinput85), .A(n6796), .ZN(n6803) );
  OAI22_X1 U7759 ( .A1(REIP_REG_13__SCAN_IN), .A2(keyinput83), .B1(DATAI_13_), 
        .B2(keyinput80), .ZN(n6797) );
  AOI221_X1 U7760 ( .B1(REIP_REG_13__SCAN_IN), .B2(keyinput83), .C1(keyinput80), .C2(DATAI_13_), .A(n6797), .ZN(n6802) );
  OAI22_X1 U7761 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(keyinput78), .B1(
        keyinput101), .B2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6798) );
  AOI221_X1 U7762 ( .B1(INSTQUEUE_REG_11__0__SCAN_IN), .B2(keyinput78), .C1(
        INSTADDRPOINTER_REG_7__SCAN_IN), .C2(keyinput101), .A(n6798), .ZN(
        n6801) );
  OAI22_X1 U7763 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(keyinput116), 
        .B1(keyinput30), .B2(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6799) );
  AOI221_X1 U7764 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(keyinput116), 
        .C1(DATAWIDTH_REG_14__SCAN_IN), .C2(keyinput30), .A(n6799), .ZN(n6800)
         );
  NAND4_X1 U7765 ( .A1(n6803), .A2(n6802), .A3(n6801), .A4(n6800), .ZN(n6833)
         );
  OAI22_X1 U7766 ( .A1(DATAI_5_), .A2(keyinput86), .B1(keyinput126), .B2(
        DATAWIDTH_REG_11__SCAN_IN), .ZN(n6804) );
  AOI221_X1 U7767 ( .B1(DATAI_5_), .B2(keyinput86), .C1(
        DATAWIDTH_REG_11__SCAN_IN), .C2(keyinput126), .A(n6804), .ZN(n6811) );
  OAI22_X1 U7768 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(keyinput71), .B1(
        DATAO_REG_6__SCAN_IN), .B2(keyinput7), .ZN(n6805) );
  AOI221_X1 U7769 ( .B1(INSTQUEUE_REG_3__4__SCAN_IN), .B2(keyinput71), .C1(
        keyinput7), .C2(DATAO_REG_6__SCAN_IN), .A(n6805), .ZN(n6810) );
  OAI22_X1 U7770 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(keyinput51), .B1(
        keyinput18), .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n6806) );
  AOI221_X1 U7771 ( .B1(INSTQUEUE_REG_15__1__SCAN_IN), .B2(keyinput51), .C1(
        INSTQUEUE_REG_11__5__SCAN_IN), .C2(keyinput18), .A(n6806), .ZN(n6809)
         );
  OAI22_X1 U7772 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(keyinput39), .B1(
        PHYADDRPOINTER_REG_16__SCAN_IN), .B2(keyinput54), .ZN(n6807) );
  AOI221_X1 U7773 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(keyinput39), .C1(
        keyinput54), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6807), .ZN(n6808) );
  NAND4_X1 U7774 ( .A1(n6811), .A2(n6810), .A3(n6809), .A4(n6808), .ZN(n6832)
         );
  OAI22_X1 U7775 ( .A1(n7000), .A2(keyinput64), .B1(keyinput24), .B2(
        REIP_REG_21__SCAN_IN), .ZN(n6812) );
  AOI221_X1 U7776 ( .B1(n7000), .B2(keyinput64), .C1(REIP_REG_21__SCAN_IN), 
        .C2(keyinput24), .A(n6812), .ZN(n6821) );
  OAI22_X1 U7777 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(keyinput123), .B1(
        DATAWIDTH_REG_24__SCAN_IN), .B2(keyinput32), .ZN(n6813) );
  AOI221_X1 U7778 ( .B1(INSTQUEUE_REG_11__1__SCAN_IN), .B2(keyinput123), .C1(
        keyinput32), .C2(DATAWIDTH_REG_24__SCAN_IN), .A(n6813), .ZN(n6820) );
  OAI22_X1 U7779 ( .A1(n6945), .A2(keyinput9), .B1(n6815), .B2(keyinput46), 
        .ZN(n6814) );
  AOI221_X1 U7780 ( .B1(n6945), .B2(keyinput9), .C1(keyinput46), .C2(n6815), 
        .A(n6814), .ZN(n6819) );
  INV_X1 U7781 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n6817) );
  OAI22_X1 U7782 ( .A1(n6817), .A2(keyinput108), .B1(n3940), .B2(keyinput97), 
        .ZN(n6816) );
  AOI221_X1 U7783 ( .B1(n6817), .B2(keyinput108), .C1(keyinput97), .C2(n3940), 
        .A(n6816), .ZN(n6818) );
  NAND4_X1 U7784 ( .A1(n6821), .A2(n6820), .A3(n6819), .A4(n6818), .ZN(n6831)
         );
  OAI22_X1 U7785 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(keyinput41), .B1(
        DATAO_REG_9__SCAN_IN), .B2(keyinput11), .ZN(n6822) );
  AOI221_X1 U7786 ( .B1(INSTQUEUE_REG_1__6__SCAN_IN), .B2(keyinput41), .C1(
        keyinput11), .C2(DATAO_REG_9__SCAN_IN), .A(n6822), .ZN(n6829) );
  OAI22_X1 U7787 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(keyinput104), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(keyinput5), .ZN(n6823) );
  AOI221_X1 U7788 ( .B1(INSTQUEUE_REG_1__2__SCAN_IN), .B2(keyinput104), .C1(
        keyinput5), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6823), .ZN(n6828)
         );
  OAI22_X1 U7789 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(keyinput89), .B1(
        REIP_REG_9__SCAN_IN), .B2(keyinput106), .ZN(n6824) );
  AOI221_X1 U7790 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(keyinput89), 
        .C1(keyinput106), .C2(REIP_REG_9__SCAN_IN), .A(n6824), .ZN(n6827) );
  OAI22_X1 U7791 ( .A1(INSTQUEUE_REG_4__1__SCAN_IN), .A2(keyinput67), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(keyinput66), .ZN(n6825) );
  AOI221_X1 U7792 ( .B1(INSTQUEUE_REG_4__1__SCAN_IN), .B2(keyinput67), .C1(
        keyinput66), .C2(ADDRESS_REG_11__SCAN_IN), .A(n6825), .ZN(n6826) );
  NAND4_X1 U7793 ( .A1(n6829), .A2(n6828), .A3(n6827), .A4(n6826), .ZN(n6830)
         );
  NOR4_X1 U7794 ( .A1(n6833), .A2(n6832), .A3(n6831), .A4(n6830), .ZN(n7187)
         );
  OAI22_X1 U7795 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(keyinput82), .B1(
        INSTQUEUE_REG_6__0__SCAN_IN), .B2(keyinput15), .ZN(n6834) );
  AOI221_X1 U7796 ( .B1(INSTQUEUE_REG_9__1__SCAN_IN), .B2(keyinput82), .C1(
        keyinput15), .C2(INSTQUEUE_REG_6__0__SCAN_IN), .A(n6834), .ZN(n6841)
         );
  OAI22_X1 U7797 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(keyinput59), .B1(
        REQUESTPENDING_REG_SCAN_IN), .B2(keyinput111), .ZN(n6835) );
  AOI221_X1 U7798 ( .B1(INSTQUEUE_REG_10__5__SCAN_IN), .B2(keyinput59), .C1(
        keyinput111), .C2(REQUESTPENDING_REG_SCAN_IN), .A(n6835), .ZN(n6840)
         );
  OAI22_X1 U7799 ( .A1(LWORD_REG_7__SCAN_IN), .A2(keyinput91), .B1(keyinput73), 
        .B2(DATAO_REG_4__SCAN_IN), .ZN(n6836) );
  AOI221_X1 U7800 ( .B1(LWORD_REG_7__SCAN_IN), .B2(keyinput91), .C1(
        DATAO_REG_4__SCAN_IN), .C2(keyinput73), .A(n6836), .ZN(n6839) );
  OAI22_X1 U7801 ( .A1(EBX_REG_16__SCAN_IN), .A2(keyinput48), .B1(keyinput29), 
        .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6837) );
  AOI221_X1 U7802 ( .B1(EBX_REG_16__SCAN_IN), .B2(keyinput48), .C1(
        INSTADDRPOINTER_REG_0__SCAN_IN), .C2(keyinput29), .A(n6837), .ZN(n6838) );
  NAND4_X1 U7803 ( .A1(n6841), .A2(n6840), .A3(n6839), .A4(n6838), .ZN(n6869)
         );
  OAI22_X1 U7804 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(keyinput37), .B1(
        EAX_REG_16__SCAN_IN), .B2(keyinput81), .ZN(n6842) );
  AOI221_X1 U7805 ( .B1(INSTQUEUE_REG_1__5__SCAN_IN), .B2(keyinput37), .C1(
        keyinput81), .C2(EAX_REG_16__SCAN_IN), .A(n6842), .ZN(n6849) );
  OAI22_X1 U7806 ( .A1(REIP_REG_8__SCAN_IN), .A2(keyinput90), .B1(keyinput68), 
        .B2(LWORD_REG_12__SCAN_IN), .ZN(n6843) );
  AOI221_X1 U7807 ( .B1(REIP_REG_8__SCAN_IN), .B2(keyinput90), .C1(
        LWORD_REG_12__SCAN_IN), .C2(keyinput68), .A(n6843), .ZN(n6848) );
  OAI22_X1 U7808 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(keyinput113), .B1(
        keyinput114), .B2(DATAWIDTH_REG_30__SCAN_IN), .ZN(n6844) );
  AOI221_X1 U7809 ( .B1(INSTQUEUE_REG_14__0__SCAN_IN), .B2(keyinput113), .C1(
        DATAWIDTH_REG_30__SCAN_IN), .C2(keyinput114), .A(n6844), .ZN(n6847) );
  OAI22_X1 U7810 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(keyinput84), .B1(
        UWORD_REG_9__SCAN_IN), .B2(keyinput28), .ZN(n6845) );
  AOI221_X1 U7811 ( .B1(PHYADDRPOINTER_REG_9__SCAN_IN), .B2(keyinput84), .C1(
        keyinput28), .C2(UWORD_REG_9__SCAN_IN), .A(n6845), .ZN(n6846) );
  NAND4_X1 U7812 ( .A1(n6849), .A2(n6848), .A3(n6847), .A4(n6846), .ZN(n6868)
         );
  OAI22_X1 U7813 ( .A1(EBX_REG_1__SCAN_IN), .A2(keyinput87), .B1(keyinput47), 
        .B2(DATAI_31_), .ZN(n6850) );
  AOI221_X1 U7814 ( .B1(EBX_REG_1__SCAN_IN), .B2(keyinput87), .C1(DATAI_31_), 
        .C2(keyinput47), .A(n6850), .ZN(n6857) );
  OAI22_X1 U7815 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(keyinput14), .B1(
        DATAWIDTH_REG_3__SCAN_IN), .B2(keyinput95), .ZN(n6851) );
  AOI221_X1 U7816 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(keyinput14), .C1(
        keyinput95), .C2(DATAWIDTH_REG_3__SCAN_IN), .A(n6851), .ZN(n6856) );
  OAI22_X1 U7817 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(keyinput117), .B1(
        keyinput17), .B2(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6852) );
  AOI221_X1 U7818 ( .B1(INSTQUEUE_REG_5__1__SCAN_IN), .B2(keyinput117), .C1(
        DATAWIDTH_REG_4__SCAN_IN), .C2(keyinput17), .A(n6852), .ZN(n6855) );
  OAI22_X1 U7819 ( .A1(EBX_REG_8__SCAN_IN), .A2(keyinput49), .B1(keyinput57), 
        .B2(NA_N), .ZN(n6853) );
  AOI221_X1 U7820 ( .B1(EBX_REG_8__SCAN_IN), .B2(keyinput49), .C1(NA_N), .C2(
        keyinput57), .A(n6853), .ZN(n6854) );
  NAND4_X1 U7821 ( .A1(n6857), .A2(n6856), .A3(n6855), .A4(n6854), .ZN(n6867)
         );
  OAI22_X1 U7822 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(keyinput35), .B1(
        DATAWIDTH_REG_31__SCAN_IN), .B2(keyinput42), .ZN(n6858) );
  AOI221_X1 U7823 ( .B1(INSTQUEUE_REG_7__2__SCAN_IN), .B2(keyinput35), .C1(
        keyinput42), .C2(DATAWIDTH_REG_31__SCAN_IN), .A(n6858), .ZN(n6865) );
  OAI22_X1 U7824 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(keyinput20), .B1(
        keyinput50), .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n6859) );
  AOI221_X1 U7825 ( .B1(INSTQUEUE_REG_13__1__SCAN_IN), .B2(keyinput20), .C1(
        INSTQUEUE_REG_8__4__SCAN_IN), .C2(keyinput50), .A(n6859), .ZN(n6864)
         );
  OAI22_X1 U7826 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(keyinput105), .B1(
        DATAWIDTH_REG_15__SCAN_IN), .B2(keyinput4), .ZN(n6860) );
  AOI221_X1 U7827 ( .B1(INSTQUEUE_REG_13__0__SCAN_IN), .B2(keyinput105), .C1(
        keyinput4), .C2(DATAWIDTH_REG_15__SCAN_IN), .A(n6860), .ZN(n6863) );
  OAI22_X1 U7828 ( .A1(REIP_REG_20__SCAN_IN), .A2(keyinput19), .B1(keyinput36), 
        .B2(LWORD_REG_5__SCAN_IN), .ZN(n6861) );
  AOI221_X1 U7829 ( .B1(REIP_REG_20__SCAN_IN), .B2(keyinput19), .C1(
        LWORD_REG_5__SCAN_IN), .C2(keyinput36), .A(n6861), .ZN(n6862) );
  NAND4_X1 U7830 ( .A1(n6865), .A2(n6864), .A3(n6863), .A4(n6862), .ZN(n6866)
         );
  NOR4_X1 U7831 ( .A1(n6869), .A2(n6868), .A3(n6867), .A4(n6866), .ZN(n7186)
         );
  AOI22_X1 U7832 ( .A1(INSTQUEUE_REG_6__2__SCAN_IN), .A2(keyinput161), .B1(
        INSTQUEUE_REG_0__0__SCAN_IN), .B2(keyinput138), .ZN(n6870) );
  OAI221_X1 U7833 ( .B1(INSTQUEUE_REG_6__2__SCAN_IN), .B2(keyinput161), .C1(
        INSTQUEUE_REG_0__0__SCAN_IN), .C2(keyinput138), .A(n6870), .ZN(n6877)
         );
  AOI22_X1 U7834 ( .A1(ADDRESS_REG_0__SCAN_IN), .A2(keyinput227), .B1(
        LWORD_REG_5__SCAN_IN), .B2(keyinput164), .ZN(n6871) );
  OAI221_X1 U7835 ( .B1(ADDRESS_REG_0__SCAN_IN), .B2(keyinput227), .C1(
        LWORD_REG_5__SCAN_IN), .C2(keyinput164), .A(n6871), .ZN(n6876) );
  AOI22_X1 U7836 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(keyinput254), .B1(
        INSTQUEUE_REG_9__7__SCAN_IN), .B2(keyinput198), .ZN(n6872) );
  OAI221_X1 U7837 ( .B1(DATAWIDTH_REG_11__SCAN_IN), .B2(keyinput254), .C1(
        INSTQUEUE_REG_9__7__SCAN_IN), .C2(keyinput198), .A(n6872), .ZN(n6875)
         );
  AOI22_X1 U7838 ( .A1(UWORD_REG_9__SCAN_IN), .A2(keyinput156), .B1(
        REIP_REG_20__SCAN_IN), .B2(keyinput147), .ZN(n6873) );
  OAI221_X1 U7839 ( .B1(UWORD_REG_9__SCAN_IN), .B2(keyinput156), .C1(
        REIP_REG_20__SCAN_IN), .C2(keyinput147), .A(n6873), .ZN(n6874) );
  NOR4_X1 U7840 ( .A1(n6877), .A2(n6876), .A3(n6875), .A4(n6874), .ZN(n6905)
         );
  AOI22_X1 U7841 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(keyinput132), .B1(
        LWORD_REG_7__SCAN_IN), .B2(keyinput219), .ZN(n6878) );
  OAI221_X1 U7842 ( .B1(DATAWIDTH_REG_15__SCAN_IN), .B2(keyinput132), .C1(
        LWORD_REG_7__SCAN_IN), .C2(keyinput219), .A(n6878), .ZN(n6885) );
  AOI22_X1 U7843 ( .A1(REIP_REG_9__SCAN_IN), .A2(keyinput234), .B1(
        EBX_REG_7__SCAN_IN), .B2(keyinput173), .ZN(n6879) );
  OAI221_X1 U7844 ( .B1(REIP_REG_9__SCAN_IN), .B2(keyinput234), .C1(
        EBX_REG_7__SCAN_IN), .C2(keyinput173), .A(n6879), .ZN(n6884) );
  AOI22_X1 U7845 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(keyinput131), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(keyinput128), .ZN(n6880) );
  OAI221_X1 U7846 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(keyinput131), .C1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .C2(keyinput128), .A(n6880), .ZN(
        n6883) );
  AOI22_X1 U7847 ( .A1(DATAO_REG_8__SCAN_IN), .A2(keyinput190), .B1(
        INSTQUEUE_REG_10__6__SCAN_IN), .B2(keyinput231), .ZN(n6881) );
  OAI221_X1 U7848 ( .B1(DATAO_REG_8__SCAN_IN), .B2(keyinput190), .C1(
        INSTQUEUE_REG_10__6__SCAN_IN), .C2(keyinput231), .A(n6881), .ZN(n6882)
         );
  NOR4_X1 U7849 ( .A1(n6885), .A2(n6884), .A3(n6883), .A4(n6882), .ZN(n6904)
         );
  AOI22_X1 U7850 ( .A1(ADDRESS_REG_8__SCAN_IN), .A2(keyinput235), .B1(
        EBX_REG_8__SCAN_IN), .B2(keyinput177), .ZN(n6886) );
  OAI221_X1 U7851 ( .B1(ADDRESS_REG_8__SCAN_IN), .B2(keyinput235), .C1(
        EBX_REG_8__SCAN_IN), .C2(keyinput177), .A(n6886), .ZN(n6893) );
  AOI22_X1 U7852 ( .A1(DATAO_REG_9__SCAN_IN), .A2(keyinput139), .B1(
        INSTADDRPOINTER_REG_7__SCAN_IN), .B2(keyinput229), .ZN(n6887) );
  OAI221_X1 U7853 ( .B1(DATAO_REG_9__SCAN_IN), .B2(keyinput139), .C1(
        INSTADDRPOINTER_REG_7__SCAN_IN), .C2(keyinput229), .A(n6887), .ZN(
        n6892) );
  AOI22_X1 U7854 ( .A1(STATE_REG_0__SCAN_IN), .A2(keyinput237), .B1(
        INSTQUEUE_REG_6__1__SCAN_IN), .B2(keyinput250), .ZN(n6888) );
  OAI221_X1 U7855 ( .B1(STATE_REG_0__SCAN_IN), .B2(keyinput237), .C1(
        INSTQUEUE_REG_6__1__SCAN_IN), .C2(keyinput250), .A(n6888), .ZN(n6891)
         );
  AOI22_X1 U7856 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(keyinput226), .B1(
        EAX_REG_22__SCAN_IN), .B2(keyinput166), .ZN(n6889) );
  OAI221_X1 U7857 ( .B1(DATAWIDTH_REG_7__SCAN_IN), .B2(keyinput226), .C1(
        EAX_REG_22__SCAN_IN), .C2(keyinput166), .A(n6889), .ZN(n6890) );
  NOR4_X1 U7858 ( .A1(n6893), .A2(n6892), .A3(n6891), .A4(n6890), .ZN(n6903)
         );
  AOI22_X1 U7859 ( .A1(REIP_REG_8__SCAN_IN), .A2(keyinput218), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(keyinput151), .ZN(n6894) );
  OAI221_X1 U7860 ( .B1(REIP_REG_8__SCAN_IN), .B2(keyinput218), .C1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .C2(keyinput151), .A(n6894), .ZN(
        n6901) );
  AOI22_X1 U7861 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(keyinput205), 
        .B1(INSTQUEUE_REG_5__1__SCAN_IN), .B2(keyinput245), .ZN(n6895) );
  OAI221_X1 U7862 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(keyinput205), 
        .C1(INSTQUEUE_REG_5__1__SCAN_IN), .C2(keyinput245), .A(n6895), .ZN(
        n6900) );
  AOI22_X1 U7863 ( .A1(ADDRESS_REG_9__SCAN_IN), .A2(keyinput130), .B1(
        INSTQUEUE_REG_8__3__SCAN_IN), .B2(keyinput134), .ZN(n6896) );
  OAI221_X1 U7864 ( .B1(ADDRESS_REG_9__SCAN_IN), .B2(keyinput130), .C1(
        INSTQUEUE_REG_8__3__SCAN_IN), .C2(keyinput134), .A(n6896), .ZN(n6899)
         );
  AOI22_X1 U7865 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(keyinput170), .B1(
        INSTQUEUE_REG_1__5__SCAN_IN), .B2(keyinput165), .ZN(n6897) );
  OAI221_X1 U7866 ( .B1(DATAWIDTH_REG_31__SCAN_IN), .B2(keyinput170), .C1(
        INSTQUEUE_REG_1__5__SCAN_IN), .C2(keyinput165), .A(n6897), .ZN(n6898)
         );
  NOR4_X1 U7867 ( .A1(n6901), .A2(n6900), .A3(n6899), .A4(n6898), .ZN(n6902)
         );
  NAND4_X1 U7868 ( .A1(n6905), .A2(n6904), .A3(n6903), .A4(n6902), .ZN(n7047)
         );
  AOI22_X1 U7869 ( .A1(ADDRESS_REG_3__SCAN_IN), .A2(keyinput248), .B1(
        REIP_REG_13__SCAN_IN), .B2(keyinput211), .ZN(n6906) );
  OAI221_X1 U7870 ( .B1(ADDRESS_REG_3__SCAN_IN), .B2(keyinput248), .C1(
        REIP_REG_13__SCAN_IN), .C2(keyinput211), .A(n6906), .ZN(n6913) );
  AOI22_X1 U7871 ( .A1(LWORD_REG_12__SCAN_IN), .A2(keyinput196), .B1(
        INSTADDRPOINTER_REG_13__SCAN_IN), .B2(keyinput244), .ZN(n6907) );
  OAI221_X1 U7872 ( .B1(LWORD_REG_12__SCAN_IN), .B2(keyinput196), .C1(
        INSTADDRPOINTER_REG_13__SCAN_IN), .C2(keyinput244), .A(n6907), .ZN(
        n6912) );
  AOI22_X1 U7873 ( .A1(REIP_REG_21__SCAN_IN), .A2(keyinput152), .B1(
        EBX_REG_16__SCAN_IN), .B2(keyinput176), .ZN(n6908) );
  OAI221_X1 U7874 ( .B1(REIP_REG_21__SCAN_IN), .B2(keyinput152), .C1(
        EBX_REG_16__SCAN_IN), .C2(keyinput176), .A(n6908), .ZN(n6911) );
  AOI22_X1 U7875 ( .A1(LWORD_REG_3__SCAN_IN), .A2(keyinput174), .B1(
        INSTADDRPOINTER_REG_2__SCAN_IN), .B2(keyinput142), .ZN(n6909) );
  OAI221_X1 U7876 ( .B1(LWORD_REG_3__SCAN_IN), .B2(keyinput174), .C1(
        INSTADDRPOINTER_REG_2__SCAN_IN), .C2(keyinput142), .A(n6909), .ZN(
        n6910) );
  NOR4_X1 U7877 ( .A1(n6913), .A2(n6912), .A3(n6911), .A4(n6910), .ZN(n6941)
         );
  AOI22_X1 U7878 ( .A1(ADDRESS_REG_11__SCAN_IN), .A2(keyinput194), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(keyinput189), .ZN(n6914) );
  OAI221_X1 U7879 ( .B1(ADDRESS_REG_11__SCAN_IN), .B2(keyinput194), .C1(
        ADDRESS_REG_7__SCAN_IN), .C2(keyinput189), .A(n6914), .ZN(n6921) );
  AOI22_X1 U7880 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(keyinput223), .B1(
        DATAWIDTH_REG_30__SCAN_IN), .B2(keyinput242), .ZN(n6915) );
  OAI221_X1 U7881 ( .B1(DATAWIDTH_REG_3__SCAN_IN), .B2(keyinput223), .C1(
        DATAWIDTH_REG_30__SCAN_IN), .C2(keyinput242), .A(n6915), .ZN(n6920) );
  AOI22_X1 U7882 ( .A1(ADDRESS_REG_29__SCAN_IN), .A2(keyinput144), .B1(
        INSTQUEUE_REG_13__5__SCAN_IN), .B2(keyinput155), .ZN(n6916) );
  OAI221_X1 U7883 ( .B1(ADDRESS_REG_29__SCAN_IN), .B2(keyinput144), .C1(
        INSTQUEUE_REG_13__5__SCAN_IN), .C2(keyinput155), .A(n6916), .ZN(n6919)
         );
  AOI22_X1 U7884 ( .A1(UWORD_REG_12__SCAN_IN), .A2(keyinput255), .B1(
        EBX_REG_17__SCAN_IN), .B2(keyinput184), .ZN(n6917) );
  OAI221_X1 U7885 ( .B1(UWORD_REG_12__SCAN_IN), .B2(keyinput255), .C1(
        EBX_REG_17__SCAN_IN), .C2(keyinput184), .A(n6917), .ZN(n6918) );
  NOR4_X1 U7886 ( .A1(n6921), .A2(n6920), .A3(n6919), .A4(n6918), .ZN(n6940)
         );
  AOI22_X1 U7887 ( .A1(UWORD_REG_2__SCAN_IN), .A2(keyinput183), .B1(
        BE_N_REG_0__SCAN_IN), .B2(keyinput193), .ZN(n6922) );
  OAI221_X1 U7888 ( .B1(UWORD_REG_2__SCAN_IN), .B2(keyinput183), .C1(
        BE_N_REG_0__SCAN_IN), .C2(keyinput193), .A(n6922), .ZN(n6929) );
  AOI22_X1 U7889 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(keyinput243), .B1(
        INSTQUEUE_REG_11__5__SCAN_IN), .B2(keyinput146), .ZN(n6923) );
  OAI221_X1 U7890 ( .B1(PHYADDRPOINTER_REG_15__SCAN_IN), .B2(keyinput243), 
        .C1(INSTQUEUE_REG_11__5__SCAN_IN), .C2(keyinput146), .A(n6923), .ZN(
        n6928) );
  AOI22_X1 U7891 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(keyinput232), .B1(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(keyinput222), .ZN(n6924) );
  OAI221_X1 U7892 ( .B1(INSTQUEUE_REG_1__2__SCAN_IN), .B2(keyinput232), .C1(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(keyinput222), .A(n6924), .ZN(
        n6927) );
  AOI22_X1 U7893 ( .A1(EAX_REG_16__SCAN_IN), .A2(keyinput209), .B1(
        INSTQUEUE_REG_2__4__SCAN_IN), .B2(keyinput204), .ZN(n6925) );
  OAI221_X1 U7894 ( .B1(EAX_REG_16__SCAN_IN), .B2(keyinput209), .C1(
        INSTQUEUE_REG_2__4__SCAN_IN), .C2(keyinput204), .A(n6925), .ZN(n6926)
         );
  NOR4_X1 U7895 ( .A1(n6929), .A2(n6928), .A3(n6927), .A4(n6926), .ZN(n6939)
         );
  AOI22_X1 U7896 ( .A1(DATAI_17_), .A2(keyinput181), .B1(
        INSTQUEUE_REG_12__7__SCAN_IN), .B2(keyinput236), .ZN(n6930) );
  OAI221_X1 U7897 ( .B1(DATAI_17_), .B2(keyinput181), .C1(
        INSTQUEUE_REG_12__7__SCAN_IN), .C2(keyinput236), .A(n6930), .ZN(n6937)
         );
  AOI22_X1 U7898 ( .A1(REIP_REG_7__SCAN_IN), .A2(keyinput240), .B1(
        INSTQUEUE_REG_6__7__SCAN_IN), .B2(keyinput168), .ZN(n6931) );
  OAI221_X1 U7899 ( .B1(REIP_REG_7__SCAN_IN), .B2(keyinput240), .C1(
        INSTQUEUE_REG_6__7__SCAN_IN), .C2(keyinput168), .A(n6931), .ZN(n6936)
         );
  AOI22_X1 U7900 ( .A1(DATAO_REG_6__SCAN_IN), .A2(keyinput135), .B1(
        INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(keyinput217), .ZN(n6932) );
  OAI221_X1 U7901 ( .B1(DATAO_REG_6__SCAN_IN), .B2(keyinput135), .C1(
        INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(keyinput217), .A(n6932), .ZN(
        n6935) );
  AOI22_X1 U7902 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(keyinput158), .B1(
        INSTQUEUE_REG_8__4__SCAN_IN), .B2(keyinput178), .ZN(n6933) );
  OAI221_X1 U7903 ( .B1(DATAWIDTH_REG_14__SCAN_IN), .B2(keyinput158), .C1(
        INSTQUEUE_REG_8__4__SCAN_IN), .C2(keyinput178), .A(n6933), .ZN(n6934)
         );
  NOR4_X1 U7904 ( .A1(n6937), .A2(n6936), .A3(n6935), .A4(n6934), .ZN(n6938)
         );
  NAND4_X1 U7905 ( .A1(n6941), .A2(n6940), .A3(n6939), .A4(n6938), .ZN(n7046)
         );
  AOI22_X1 U7906 ( .A1(n6946), .A2(keyinput175), .B1(n6945), .B2(keyinput137), 
        .ZN(n6944) );
  OAI221_X1 U7907 ( .B1(n6946), .B2(keyinput175), .C1(n6945), .C2(keyinput137), 
        .A(n6944), .ZN(n6954) );
  INV_X1 U7908 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n6948) );
  AOI22_X1 U7909 ( .A1(n7055), .A2(keyinput246), .B1(n6948), .B2(keyinput148), 
        .ZN(n6947) );
  OAI221_X1 U7910 ( .B1(n7055), .B2(keyinput246), .C1(n6948), .C2(keyinput148), 
        .A(n6947), .ZN(n6953) );
  INV_X1 U7911 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n6951) );
  INV_X1 U7912 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n6950) );
  AOI22_X1 U7913 ( .A1(n6951), .A2(keyinput143), .B1(n6950), .B2(keyinput199), 
        .ZN(n6949) );
  OAI221_X1 U7914 ( .B1(n6951), .B2(keyinput143), .C1(n6950), .C2(keyinput199), 
        .A(n6949), .ZN(n6952) );
  NOR4_X1 U7915 ( .A1(n6955), .A2(n6954), .A3(n6953), .A4(n6952), .ZN(n6992)
         );
  INV_X1 U7916 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n7083) );
  AOI22_X1 U7917 ( .A1(n7083), .A2(keyinput129), .B1(keyinput154), .B2(n7173), 
        .ZN(n6956) );
  OAI221_X1 U7918 ( .B1(n7083), .B2(keyinput129), .C1(n7173), .C2(keyinput154), 
        .A(n6956), .ZN(n6967) );
  INV_X1 U7919 ( .A(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n6958) );
  AOI22_X1 U7920 ( .A1(n6958), .A2(keyinput230), .B1(keyinput207), .B2(n3944), 
        .ZN(n6957) );
  OAI221_X1 U7921 ( .B1(n6958), .B2(keyinput230), .C1(n3944), .C2(keyinput207), 
        .A(n6957), .ZN(n6966) );
  INV_X1 U7922 ( .A(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n6961) );
  AOI22_X1 U7923 ( .A1(n6961), .A2(keyinput206), .B1(keyinput185), .B2(n6960), 
        .ZN(n6959) );
  OAI221_X1 U7924 ( .B1(n6961), .B2(keyinput206), .C1(n6960), .C2(keyinput185), 
        .A(n6959), .ZN(n6965) );
  AOI22_X1 U7925 ( .A1(n7134), .A2(keyinput186), .B1(keyinput160), .B2(n6963), 
        .ZN(n6962) );
  OAI221_X1 U7926 ( .B1(n7134), .B2(keyinput186), .C1(n6963), .C2(keyinput160), 
        .A(n6962), .ZN(n6964) );
  NOR4_X1 U7927 ( .A1(n6967), .A2(n6966), .A3(n6965), .A4(n6964), .ZN(n6991)
         );
  INV_X1 U7928 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n7089) );
  AOI22_X1 U7929 ( .A1(n7140), .A2(keyinput252), .B1(keyinput197), .B2(n7096), 
        .ZN(n6970) );
  OAI221_X1 U7930 ( .B1(n7140), .B2(keyinput252), .C1(n7096), .C2(keyinput197), 
        .A(n6970), .ZN(n6977) );
  AOI22_X1 U7931 ( .A1(n6972), .A2(keyinput201), .B1(keyinput216), .B2(n7100), 
        .ZN(n6971) );
  OAI221_X1 U7932 ( .B1(n6972), .B2(keyinput201), .C1(n7100), .C2(keyinput216), 
        .A(n6971), .ZN(n6976) );
  INV_X1 U7933 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n7104) );
  INV_X1 U7934 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n6974) );
  AOI22_X1 U7935 ( .A1(n7104), .A2(keyinput247), .B1(n6974), .B2(keyinput233), 
        .ZN(n6973) );
  OAI221_X1 U7936 ( .B1(n7104), .B2(keyinput247), .C1(n6974), .C2(keyinput233), 
        .A(n6973), .ZN(n6975) );
  NOR4_X1 U7937 ( .A1(n6978), .A2(n6977), .A3(n6976), .A4(n6975), .ZN(n6990)
         );
  AOI22_X1 U7938 ( .A1(n7058), .A2(keyinput136), .B1(keyinput202), .B2(n7135), 
        .ZN(n6979) );
  OAI221_X1 U7939 ( .B1(n7058), .B2(keyinput136), .C1(n7135), .C2(keyinput202), 
        .A(n6979), .ZN(n6988) );
  INV_X1 U7940 ( .A(DATAI_27_), .ZN(n7143) );
  INV_X1 U7941 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n6981) );
  AOI22_X1 U7942 ( .A1(n7143), .A2(keyinput200), .B1(n6981), .B2(keyinput195), 
        .ZN(n6980) );
  OAI221_X1 U7943 ( .B1(n7143), .B2(keyinput200), .C1(n6981), .C2(keyinput195), 
        .A(n6980), .ZN(n6987) );
  AOI22_X1 U7944 ( .A1(n7157), .A2(keyinput150), .B1(n7152), .B2(keyinput228), 
        .ZN(n6982) );
  OAI221_X1 U7945 ( .B1(n7157), .B2(keyinput150), .C1(n7152), .C2(keyinput228), 
        .A(n6982), .ZN(n6986) );
  INV_X1 U7946 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n7138) );
  AOI22_X1 U7947 ( .A1(n6984), .A2(keyinput239), .B1(n7138), .B2(keyinput220), 
        .ZN(n6983) );
  OAI221_X1 U7948 ( .B1(n6984), .B2(keyinput239), .C1(n7138), .C2(keyinput220), 
        .A(n6983), .ZN(n6985) );
  NOR4_X1 U7949 ( .A1(n6988), .A2(n6987), .A3(n6986), .A4(n6985), .ZN(n6989)
         );
  NAND4_X1 U7950 ( .A1(n6992), .A2(n6991), .A3(n6990), .A4(n6989), .ZN(n7045)
         );
  AOI22_X1 U7951 ( .A1(n7067), .A2(keyinput188), .B1(n7074), .B2(keyinput221), 
        .ZN(n6995) );
  OAI221_X1 U7952 ( .B1(n7067), .B2(keyinput188), .C1(n7074), .C2(keyinput221), 
        .A(n6995), .ZN(n7003) );
  INV_X1 U7953 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n6997) );
  AOI22_X1 U7954 ( .A1(n6998), .A2(keyinput215), .B1(n6997), .B2(keyinput179), 
        .ZN(n6996) );
  OAI221_X1 U7955 ( .B1(n6998), .B2(keyinput215), .C1(n6997), .C2(keyinput179), 
        .A(n6996), .ZN(n7002) );
  AOI22_X1 U7956 ( .A1(n7000), .A2(keyinput192), .B1(keyinput162), .B2(n7086), 
        .ZN(n6999) );
  OAI221_X1 U7957 ( .B1(n7000), .B2(keyinput192), .C1(n7086), .C2(keyinput162), 
        .A(n6999), .ZN(n7001) );
  NOR4_X1 U7958 ( .A1(n7004), .A2(n7003), .A3(n7002), .A4(n7001), .ZN(n7043)
         );
  INV_X1 U7959 ( .A(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n7007) );
  AOI22_X1 U7960 ( .A1(n7007), .A2(keyinput163), .B1(keyinput214), .B2(n7006), 
        .ZN(n7005) );
  OAI221_X1 U7961 ( .B1(n7007), .B2(keyinput163), .C1(n7006), .C2(keyinput214), 
        .A(n7005), .ZN(n7018) );
  INV_X1 U7962 ( .A(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n7057) );
  AOI22_X1 U7963 ( .A1(n7009), .A2(keyinput167), .B1(n7057), .B2(keyinput171), 
        .ZN(n7008) );
  OAI221_X1 U7964 ( .B1(n7009), .B2(keyinput167), .C1(n7057), .C2(keyinput171), 
        .A(n7008), .ZN(n7017) );
  INV_X1 U7965 ( .A(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n7012) );
  INV_X1 U7966 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n7011) );
  AOI22_X1 U7967 ( .A1(n7012), .A2(keyinput210), .B1(keyinput241), .B2(n7011), 
        .ZN(n7010) );
  OAI221_X1 U7968 ( .B1(n7012), .B2(keyinput210), .C1(n7011), .C2(keyinput241), 
        .A(n7010), .ZN(n7016) );
  INV_X1 U7969 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n7014) );
  AOI22_X1 U7970 ( .A1(n7014), .A2(keyinput187), .B1(keyinput203), .B2(n5507), 
        .ZN(n7013) );
  OAI221_X1 U7971 ( .B1(n7014), .B2(keyinput187), .C1(n5507), .C2(keyinput203), 
        .A(n7013), .ZN(n7015) );
  NOR4_X1 U7972 ( .A1(n7018), .A2(n7017), .A3(n7016), .A4(n7015), .ZN(n7042)
         );
  AOI22_X1 U7973 ( .A1(n4904), .A2(keyinput153), .B1(keyinput213), .B2(n7020), 
        .ZN(n7019) );
  OAI221_X1 U7974 ( .B1(n4904), .B2(keyinput153), .C1(n7020), .C2(keyinput213), 
        .A(n7019), .ZN(n7029) );
  AOI22_X1 U7975 ( .A1(n4442), .A2(keyinput249), .B1(keyinput208), .B2(n7022), 
        .ZN(n7021) );
  OAI221_X1 U7976 ( .B1(n4442), .B2(keyinput249), .C1(n7022), .C2(keyinput208), 
        .A(n7021), .ZN(n7028) );
  INV_X1 U7977 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n7065) );
  INV_X1 U7978 ( .A(EBX_REG_3__SCAN_IN), .ZN(n7071) );
  AOI22_X1 U7979 ( .A1(n7065), .A2(keyinput141), .B1(keyinput149), .B2(n7071), 
        .ZN(n7023) );
  OAI221_X1 U7980 ( .B1(n7065), .B2(keyinput141), .C1(n7071), .C2(keyinput149), 
        .A(n7023), .ZN(n7027) );
  AOI22_X1 U7981 ( .A1(n3940), .A2(keyinput225), .B1(n7025), .B2(keyinput157), 
        .ZN(n7024) );
  OAI221_X1 U7982 ( .B1(n3940), .B2(keyinput225), .C1(n7025), .C2(keyinput157), 
        .A(n7024), .ZN(n7026) );
  NOR4_X1 U7983 ( .A1(n7029), .A2(n7028), .A3(n7027), .A4(n7026), .ZN(n7041)
         );
  INV_X1 U7984 ( .A(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n7031) );
  AOI22_X1 U7985 ( .A1(n5023), .A2(keyinput169), .B1(n7031), .B2(keyinput251), 
        .ZN(n7030) );
  OAI221_X1 U7986 ( .B1(n5023), .B2(keyinput169), .C1(n7031), .C2(keyinput251), 
        .A(n7030), .ZN(n7039) );
  INV_X1 U7987 ( .A(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n7049) );
  AOI22_X1 U7988 ( .A1(n7049), .A2(keyinput253), .B1(keyinput224), .B2(n7064), 
        .ZN(n7032) );
  OAI221_X1 U7989 ( .B1(n7049), .B2(keyinput253), .C1(n7064), .C2(keyinput224), 
        .A(n7032), .ZN(n7038) );
  AOI22_X1 U7990 ( .A1(n7034), .A2(keyinput145), .B1(n7119), .B2(keyinput191), 
        .ZN(n7033) );
  OAI221_X1 U7991 ( .B1(n7034), .B2(keyinput145), .C1(n7119), .C2(keyinput191), 
        .A(n7033), .ZN(n7037) );
  INV_X1 U7992 ( .A(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n7114) );
  AOI22_X1 U7993 ( .A1(n7169), .A2(keyinput172), .B1(n7114), .B2(keyinput180), 
        .ZN(n7035) );
  OAI221_X1 U7994 ( .B1(n7169), .B2(keyinput172), .C1(n7114), .C2(keyinput180), 
        .A(n7035), .ZN(n7036) );
  NOR4_X1 U7995 ( .A1(n7039), .A2(n7038), .A3(n7037), .A4(n7036), .ZN(n7040)
         );
  NAND4_X1 U7996 ( .A1(n7043), .A2(n7042), .A3(n7041), .A4(n7040), .ZN(n7044)
         );
  NOR4_X1 U7997 ( .A1(n7047), .A2(n7046), .A3(n7045), .A4(n7044), .ZN(n7184)
         );
  AOI22_X1 U7998 ( .A1(n7050), .A2(keyinput127), .B1(n7049), .B2(keyinput125), 
        .ZN(n7048) );
  OAI221_X1 U7999 ( .B1(n7050), .B2(keyinput127), .C1(n7049), .C2(keyinput125), 
        .A(n7048), .ZN(n7062) );
  AOI22_X1 U8000 ( .A1(n4881), .A2(keyinput76), .B1(keyinput120), .B2(n7052), 
        .ZN(n7051) );
  OAI221_X1 U8001 ( .B1(n4881), .B2(keyinput76), .C1(n7052), .C2(keyinput120), 
        .A(n7051), .ZN(n7061) );
  AOI22_X1 U8002 ( .A1(n7055), .A2(keyinput118), .B1(n7054), .B2(keyinput109), 
        .ZN(n7053) );
  OAI221_X1 U8003 ( .B1(n7055), .B2(keyinput118), .C1(n7054), .C2(keyinput109), 
        .A(n7053), .ZN(n7060) );
  AOI22_X1 U8004 ( .A1(n7058), .A2(keyinput8), .B1(n7057), .B2(keyinput43), 
        .ZN(n7056) );
  OAI221_X1 U8005 ( .B1(n7058), .B2(keyinput8), .C1(n7057), .C2(keyinput43), 
        .A(n7056), .ZN(n7059) );
  NOR4_X1 U8006 ( .A1(n7062), .A2(n7061), .A3(n7060), .A4(n7059), .ZN(n7112)
         );
  AOI22_X1 U8007 ( .A1(n7065), .A2(keyinput13), .B1(keyinput96), .B2(n7064), 
        .ZN(n7063) );
  OAI221_X1 U8008 ( .B1(n7065), .B2(keyinput13), .C1(n7064), .C2(keyinput96), 
        .A(n7063), .ZN(n7078) );
  AOI22_X1 U8009 ( .A1(n7068), .A2(keyinput0), .B1(keyinput60), .B2(n7067), 
        .ZN(n7066) );
  OAI221_X1 U8010 ( .B1(n7068), .B2(keyinput0), .C1(n7067), .C2(keyinput60), 
        .A(n7066), .ZN(n7077) );
  AOI22_X1 U8011 ( .A1(n7071), .A2(keyinput21), .B1(keyinput107), .B2(n7070), 
        .ZN(n7069) );
  OAI221_X1 U8012 ( .B1(n7071), .B2(keyinput21), .C1(n7070), .C2(keyinput107), 
        .A(n7069), .ZN(n7076) );
  AOI22_X1 U8013 ( .A1(n7074), .A2(keyinput93), .B1(keyinput56), .B2(n7073), 
        .ZN(n7072) );
  OAI221_X1 U8014 ( .B1(n7074), .B2(keyinput93), .C1(n7073), .C2(keyinput56), 
        .A(n7072), .ZN(n7075) );
  NOR4_X1 U8015 ( .A1(n7078), .A2(n7077), .A3(n7076), .A4(n7075), .ZN(n7111)
         );
  AOI22_X1 U8016 ( .A1(n7081), .A2(keyinput23), .B1(n7080), .B2(keyinput33), 
        .ZN(n7079) );
  OAI221_X1 U8017 ( .B1(n7081), .B2(keyinput23), .C1(n7080), .C2(keyinput33), 
        .A(n7079), .ZN(n7093) );
  AOI22_X1 U8018 ( .A1(n7083), .A2(keyinput1), .B1(keyinput45), .B2(n5124), 
        .ZN(n7082) );
  OAI221_X1 U8019 ( .B1(n7083), .B2(keyinput1), .C1(n5124), .C2(keyinput45), 
        .A(n7082), .ZN(n7092) );
  INV_X1 U8020 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n7085) );
  AOI22_X1 U8021 ( .A1(n7086), .A2(keyinput34), .B1(n7085), .B2(keyinput10), 
        .ZN(n7084) );
  OAI221_X1 U8022 ( .B1(n7086), .B2(keyinput34), .C1(n7085), .C2(keyinput10), 
        .A(n7084), .ZN(n7091) );
  INV_X1 U8023 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n7088) );
  AOI22_X1 U8024 ( .A1(n7089), .A2(keyinput110), .B1(n7088), .B2(keyinput40), 
        .ZN(n7087) );
  OAI221_X1 U8025 ( .B1(n7089), .B2(keyinput110), .C1(n7088), .C2(keyinput40), 
        .A(n7087), .ZN(n7090) );
  NOR4_X1 U8026 ( .A1(n7093), .A2(n7092), .A3(n7091), .A4(n7090), .ZN(n7110)
         );
  AOI22_X1 U8027 ( .A1(n7096), .A2(keyinput69), .B1(n7095), .B2(keyinput38), 
        .ZN(n7094) );
  OAI221_X1 U8028 ( .B1(n7096), .B2(keyinput69), .C1(n7095), .C2(keyinput38), 
        .A(n7094), .ZN(n7108) );
  AOI22_X1 U8029 ( .A1(n4442), .A2(keyinput121), .B1(n7098), .B2(keyinput12), 
        .ZN(n7097) );
  OAI221_X1 U8030 ( .B1(n4442), .B2(keyinput121), .C1(n7098), .C2(keyinput12), 
        .A(n7097), .ZN(n7107) );
  AOI22_X1 U8031 ( .A1(n7101), .A2(keyinput62), .B1(keyinput88), .B2(n7100), 
        .ZN(n7099) );
  OAI221_X1 U8032 ( .B1(n7101), .B2(keyinput62), .C1(n7100), .C2(keyinput88), 
        .A(n7099), .ZN(n7106) );
  AOI22_X1 U8033 ( .A1(n7104), .A2(keyinput119), .B1(keyinput16), .B2(n7103), 
        .ZN(n7102) );
  OAI221_X1 U8034 ( .B1(n7104), .B2(keyinput119), .C1(n7103), .C2(keyinput16), 
        .A(n7102), .ZN(n7105) );
  NOR4_X1 U8035 ( .A1(n7108), .A2(n7107), .A3(n7106), .A4(n7105), .ZN(n7109)
         );
  NAND4_X1 U8036 ( .A1(n7112), .A2(n7111), .A3(n7110), .A4(n7109), .ZN(n7183)
         );
  INV_X1 U8037 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n7115) );
  AOI22_X1 U8038 ( .A1(n7115), .A2(keyinput6), .B1(n7114), .B2(keyinput52), 
        .ZN(n7113) );
  OAI221_X1 U8039 ( .B1(n7115), .B2(keyinput6), .C1(n7114), .C2(keyinput52), 
        .A(n7113), .ZN(n7116) );
  INV_X1 U8040 ( .A(n7116), .ZN(n7132) );
  AOI22_X1 U8041 ( .A1(n7119), .A2(keyinput63), .B1(keyinput2), .B2(n7118), 
        .ZN(n7117) );
  OAI221_X1 U8042 ( .B1(n7119), .B2(keyinput63), .C1(n7118), .C2(keyinput2), 
        .A(n7117), .ZN(n7120) );
  INV_X1 U8043 ( .A(n7120), .ZN(n7131) );
  INV_X1 U8044 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n7123) );
  AOI22_X1 U8045 ( .A1(n7123), .A2(keyinput103), .B1(keyinput77), .B2(n7122), 
        .ZN(n7121) );
  OAI221_X1 U8046 ( .B1(n7123), .B2(keyinput103), .C1(n7122), .C2(keyinput77), 
        .A(n7121), .ZN(n7126) );
  INV_X1 U8047 ( .A(keyinput94), .ZN(n7124) );
  XNOR2_X1 U8048 ( .A(n7124), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n7125)
         );
  NOR2_X1 U8049 ( .A1(n7126), .A2(n7125), .ZN(n7130) );
  INV_X1 U8050 ( .A(keyinput65), .ZN(n7127) );
  XNOR2_X1 U8051 ( .A(n7128), .B(n7127), .ZN(n7129) );
  AND4_X1 U8052 ( .A1(n7132), .A2(n7131), .A3(n7130), .A4(n7129), .ZN(n7181)
         );
  AOI22_X1 U8053 ( .A1(n7135), .A2(keyinput74), .B1(n7134), .B2(keyinput58), 
        .ZN(n7133) );
  OAI221_X1 U8054 ( .B1(n7135), .B2(keyinput74), .C1(n7134), .C2(keyinput58), 
        .A(n7133), .ZN(n7147) );
  AOI22_X1 U8055 ( .A1(n7138), .A2(keyinput92), .B1(keyinput55), .B2(n7137), 
        .ZN(n7136) );
  OAI221_X1 U8056 ( .B1(n7138), .B2(keyinput92), .C1(n7137), .C2(keyinput55), 
        .A(n7136), .ZN(n7146) );
  AOI22_X1 U8057 ( .A1(n7140), .A2(keyinput124), .B1(keyinput75), .B2(n5507), 
        .ZN(n7139) );
  OAI221_X1 U8058 ( .B1(n7140), .B2(keyinput124), .C1(n5507), .C2(keyinput75), 
        .A(n7139), .ZN(n7145) );
  AOI22_X1 U8059 ( .A1(n7143), .A2(keyinput72), .B1(keyinput61), .B2(n7142), 
        .ZN(n7141) );
  OAI221_X1 U8060 ( .B1(n7143), .B2(keyinput72), .C1(n7142), .C2(keyinput61), 
        .A(n7141), .ZN(n7144) );
  NOR4_X1 U8061 ( .A1(n7147), .A2(n7146), .A3(n7145), .A4(n7144), .ZN(n7180)
         );
  AOI22_X1 U8062 ( .A1(n7152), .A2(keyinput100), .B1(keyinput98), .B2(n7151), 
        .ZN(n7150) );
  OAI221_X1 U8063 ( .B1(n7152), .B2(keyinput100), .C1(n7151), .C2(keyinput98), 
        .A(n7150), .ZN(n7160) );
  INV_X1 U8064 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n7154) );
  AOI22_X1 U8065 ( .A1(n7155), .A2(keyinput3), .B1(n7154), .B2(keyinput27), 
        .ZN(n7153) );
  OAI221_X1 U8066 ( .B1(n7155), .B2(keyinput3), .C1(n7154), .C2(keyinput27), 
        .A(n7153), .ZN(n7159) );
  AOI22_X1 U8067 ( .A1(n3944), .A2(keyinput79), .B1(keyinput22), .B2(n7157), 
        .ZN(n7156) );
  OAI221_X1 U8068 ( .B1(n3944), .B2(keyinput79), .C1(n7157), .C2(keyinput22), 
        .A(n7156), .ZN(n7158) );
  NOR4_X1 U8069 ( .A1(n7161), .A2(n7160), .A3(n7159), .A4(n7158), .ZN(n7179)
         );
  INV_X1 U8070 ( .A(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n7164) );
  AOI22_X1 U8071 ( .A1(n7164), .A2(keyinput70), .B1(keyinput99), .B2(n7163), 
        .ZN(n7162) );
  OAI221_X1 U8072 ( .B1(n7164), .B2(keyinput70), .C1(n7163), .C2(keyinput99), 
        .A(n7162), .ZN(n7177) );
  INV_X1 U8073 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n7167) );
  INV_X1 U8074 ( .A(DATAI_17_), .ZN(n7166) );
  AOI22_X1 U8075 ( .A1(n7167), .A2(keyinput115), .B1(keyinput53), .B2(n7166), 
        .ZN(n7165) );
  OAI221_X1 U8076 ( .B1(n7167), .B2(keyinput115), .C1(n7166), .C2(keyinput53), 
        .A(n7165), .ZN(n7176) );
  AOI22_X1 U8077 ( .A1(n7170), .A2(keyinput112), .B1(keyinput44), .B2(n7169), 
        .ZN(n7168) );
  OAI221_X1 U8078 ( .B1(n7170), .B2(keyinput112), .C1(n7169), .C2(keyinput44), 
        .A(n7168), .ZN(n7175) );
  INV_X1 U8079 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n7172) );
  AOI22_X1 U8080 ( .A1(n7173), .A2(keyinput26), .B1(n7172), .B2(keyinput122), 
        .ZN(n7171) );
  OAI221_X1 U8081 ( .B1(n7173), .B2(keyinput26), .C1(n7172), .C2(keyinput122), 
        .A(n7171), .ZN(n7174) );
  NOR4_X1 U8082 ( .A1(n7177), .A2(n7176), .A3(n7175), .A4(n7174), .ZN(n7178)
         );
  NAND4_X1 U8083 ( .A1(n7181), .A2(n7180), .A3(n7179), .A4(n7178), .ZN(n7182)
         );
  NOR3_X1 U8084 ( .A1(n7184), .A2(n7183), .A3(n7182), .ZN(n7185) );
  NAND3_X1 U8085 ( .A1(n7187), .A2(n7186), .A3(n7185), .ZN(n7188) );
  XNOR2_X1 U8086 ( .A(n7189), .B(n7188), .ZN(U2943) );
  AND2_X2 U3850 ( .A1(n3338), .A2(n3224), .ZN(n3427) );
  CLKBUF_X1 U3629 ( .A(n3434), .Z(n3214) );
  CLKBUF_X1 U3630 ( .A(n3786), .Z(n3221) );
  OAI21_X1 U3658 ( .B1(n5707), .B2(n6943), .A(n5782), .ZN(n5695) );
  AOI211_X2 U3659 ( .C1(n5017), .C2(n6571), .A(n6570), .B(n5015), .ZN(n5054)
         );
  AOI211_X2 U3671 ( .C1(n5859), .C2(n6571), .A(n6570), .B(n5857), .ZN(n5902)
         );
  NOR2_X2 U3689 ( .A1(n5714), .A2(n4731), .ZN(n6621) );
  NOR2_X2 U3811 ( .A1(n5714), .A2(n7166), .ZN(n6582) );
  NOR2_X2 U3834 ( .A1(n5714), .A2(n4721), .ZN(n6594) );
  OR2_X2 U4289 ( .A1(n6676), .A2(n6571), .ZN(n5714) );
endmodule

