

module b14_C_AntiSAT_k_128_10 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2055, n2056, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716;

  INV_X1 U2297 ( .A(n3538), .ZN(n3546) );
  CLKBUF_X3 U2298 ( .A(n2741), .Z(n2056) );
  CLKBUF_X2 U2299 ( .A(n2235), .Z(n2621) );
  INV_X1 U2300 ( .A(n3698), .ZN(n2899) );
  CLKBUF_X2 U2301 ( .A(n3702), .Z(n2058) );
  AND3_X1 U2302 ( .A1(n2341), .A2(n2141), .A3(n3960), .ZN(n2293) );
  NAND3_X1 U2303 ( .A1(n3598), .A2(n3522), .A3(n3523), .ZN(n3641) );
  NAND2_X1 U2304 ( .A1(n2780), .A2(n2779), .ZN(n2241) );
  OAI22_X1 U2305 ( .A1(n2970), .A2(n3525), .B1(n2797), .B2(n2991), .ZN(n2769)
         );
  CLKBUF_X3 U2306 ( .A(n2797), .Z(n3540) );
  NAND2_X1 U2307 ( .A1(n3834), .A2(n3771), .ZN(n2717) );
  CLKBUF_X2 U2308 ( .A(n3702), .Z(n2059) );
  CLKBUF_X2 U2309 ( .A(n2338), .Z(n3696) );
  OR2_X1 U2310 ( .A1(n3042), .A2(n2820), .ZN(n4698) );
  INV_X1 U2311 ( .A(IR_REG_31__SCAN_IN), .ZN(n2617) );
  XNOR2_X1 U2312 ( .A(n2608), .B(n2607), .ZN(n4132) );
  INV_X2 U2313 ( .A(n4479), .ZN(n3575) );
  XNOR2_X1 U2314 ( .A(n2768), .B(n2769), .ZN(n2985) );
  NAND2_X2 U2315 ( .A1(n3544), .A2(n4698), .ZN(n2746) );
  NAND2_X2 U2316 ( .A1(n2671), .A2(IR_REG_31__SCAN_IN), .ZN(n2672) );
  CLKBUF_X1 U2317 ( .A(n2741), .Z(n2055) );
  AND2_X2 U2318 ( .A1(n2327), .A2(n2328), .ZN(n2338) );
  OAI21_X1 U2319 ( .B1(n3489), .B2(n2244), .A(n2242), .ZN(n2252) );
  OAI22_X4 U2320 ( .A1(n3468), .A2(n3467), .B1(n3466), .B2(n3465), .ZN(n3489)
         );
  OAI21_X1 U2321 ( .B1(n3633), .B2(n3629), .A(n3630), .ZN(n3673) );
  NAND2_X1 U2322 ( .A1(n3448), .A2(n3447), .ZN(n3468) );
  NAND2_X1 U2323 ( .A1(n2241), .A2(n2070), .ZN(n3054) );
  AOI21_X1 U2324 ( .B1(n2229), .B2(n2766), .A(n2228), .ZN(n2227) );
  NAND2_X1 U2325 ( .A1(n3318), .A2(n4459), .ZN(n3366) );
  AND2_X1 U2326 ( .A1(n2958), .A2(n2959), .ZN(n2762) );
  AND2_X2 U2327 ( .A1(n3005), .A2(n4155), .ZN(n4479) );
  AOI21_X1 U2328 ( .B1(n3858), .B2(n3473), .A(n2723), .ZN(n2725) );
  CLKBUF_X3 U2329 ( .A(n2746), .Z(n3525) );
  BUF_X2 U2330 ( .A(n2772), .Z(n3534) );
  NAND2_X2 U2331 ( .A1(n2680), .A2(n2679), .ZN(n2718) );
  AND2_X2 U2332 ( .A1(n2798), .A2(n2717), .ZN(n3538) );
  NAND2_X1 U2333 ( .A1(n3773), .A2(n3769), .ZN(n2628) );
  XNOR2_X1 U2334 ( .A(n2606), .B(n2668), .ZN(n2719) );
  AND4_X1 U2335 ( .A1(n2367), .A2(n2366), .A3(n2365), .A4(n2364), .ZN(n3138)
         );
  NAND2_X1 U2336 ( .A1(n2670), .A2(IR_REG_31__SCAN_IN), .ZN(n2681) );
  NAND2_X1 U2338 ( .A1(n2605), .A2(IR_REG_31__SCAN_IN), .ZN(n2606) );
  INV_X1 U2339 ( .A(n3859), .ZN(n2744) );
  NAND3_X1 U2340 ( .A1(n2330), .A2(n2233), .A3(n2232), .ZN(n3859) );
  XNOR2_X1 U2341 ( .A(n2611), .B(n2610), .ZN(n3834) );
  NAND4_X1 U2342 ( .A1(n2353), .A2(n2352), .A3(n2351), .A4(n2350), .ZN(n3857)
         );
  NAND2_X1 U2343 ( .A1(n2609), .A2(IR_REG_31__SCAN_IN), .ZN(n2611) );
  INV_X1 U2344 ( .A(n2597), .ZN(n2579) );
  NOR2_X4 U2345 ( .A1(n2328), .A2(n2322), .ZN(n2235) );
  XNOR2_X1 U2346 ( .A(n2140), .B(n2316), .ZN(n2328) );
  AND2_X1 U2347 ( .A1(n2616), .A2(n2313), .ZN(n2843) );
  XNOR2_X1 U2348 ( .A(n2318), .B(n2317), .ZN(n2327) );
  NOR2_X1 U2349 ( .A1(n2433), .A2(n3162), .ZN(n2459) );
  AND2_X2 U2350 ( .A1(n2301), .A2(n2300), .ZN(n2506) );
  AND4_X1 U2351 ( .A1(n2299), .A2(n2298), .A3(n2297), .A4(n2296), .ZN(n2300)
         );
  AND4_X1 U2352 ( .A1(n2305), .A2(n2304), .A3(n2303), .A4(n2302), .ZN(n2662)
         );
  INV_X1 U2353 ( .A(IR_REG_15__SCAN_IN), .ZN(n2297) );
  NOR2_X1 U2354 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2302)
         );
  NOR2_X1 U2355 ( .A1(IR_REG_23__SCAN_IN), .A2(IR_REG_22__SCAN_IN), .ZN(n2303)
         );
  NOR2_X1 U2356 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_21__SCAN_IN), .ZN(n2304)
         );
  NOR2_X1 U2357 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2305)
         );
  INV_X1 U2358 ( .A(IR_REG_13__SCAN_IN), .ZN(n2296) );
  INV_X1 U2359 ( .A(IR_REG_25__SCAN_IN), .ZN(n2309) );
  OAI211_X1 U2360 ( .C1(n2851), .C2(n4448), .A(n2210), .B(1'b1), .ZN(n2207) );
  NAND2_X2 U2362 ( .A1(n3117), .A2(n2257), .ZN(n2255) );
  NAND2_X2 U2363 ( .A1(n3054), .A2(n3053), .ZN(n3117) );
  NAND2_X2 U2364 ( .A1(n3159), .A2(n3158), .ZN(n3206) );
  NAND2_X2 U2365 ( .A1(n2255), .A2(n2253), .ZN(n3159) );
  AND2_X1 U2366 ( .A1(n2506), .A2(n2309), .ZN(n2665) );
  NOR2_X2 U2367 ( .A1(n3283), .A2(n3151), .ZN(n3572) );
  AND2_X2 U2368 ( .A1(n2506), .A2(n2661), .ZN(n2509) );
  XNOR2_X1 U2369 ( .A(n2763), .B(n2764), .ZN(n2958) );
  NOR2_X2 U2370 ( .A1(n3366), .A2(n2109), .ZN(n4331) );
  NAND2_X2 U2371 ( .A1(n2718), .A2(n2716), .ZN(n2742) );
  NAND2_X2 U2372 ( .A1(n2718), .A2(n2717), .ZN(n2741) );
  OAI22_X1 U2373 ( .A1(n3138), .A2(n2742), .B1(n2055), .B2(n3013), .ZN(n2758)
         );
  AOI21_X2 U2374 ( .B1(n3619), .B2(n3509), .A(n2084), .ZN(n3663) );
  AOI21_X2 U2375 ( .B1(n3598), .B2(n3523), .A(n3522), .ZN(n3640) );
  NOR2_X2 U2376 ( .A1(n4375), .A2(n3604), .ZN(n2108) );
  AOI21_X2 U2377 ( .B1(n2918), .B2(n2919), .A(n2750), .ZN(n2906) );
  NOR2_X2 U2378 ( .A1(n3072), .A2(n3025), .ZN(n2107) );
  NAND2_X1 U2379 ( .A1(n3430), .A2(n3429), .ZN(n4464) );
  NAND2_X1 U2380 ( .A1(n2105), .A2(n2104), .ZN(n3702) );
  OAI22_X1 U2381 ( .A1(n3423), .A2(n2278), .B1(n3424), .B2(n2277), .ZN(n3430)
         );
  INV_X1 U2382 ( .A(n3422), .ZN(n2277) );
  NOR2_X1 U2383 ( .A1(n3425), .A2(n3422), .ZN(n2278) );
  INV_X1 U2384 ( .A(n2344), .ZN(n2200) );
  NOR2_X1 U2385 ( .A1(n2134), .A2(n3761), .ZN(n2133) );
  INV_X1 U2386 ( .A(n2135), .ZN(n2134) );
  NAND2_X1 U2387 ( .A1(n2117), .A2(n2542), .ZN(n2116) );
  INV_X1 U2388 ( .A(n2120), .ZN(n2117) );
  NAND2_X1 U2389 ( .A1(n3658), .A2(n4330), .ZN(n2124) );
  NAND2_X1 U2390 ( .A1(n2676), .A2(n2308), .ZN(n2842) );
  AND2_X1 U2391 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2308)
         );
  INV_X1 U2392 ( .A(IR_REG_17__SCAN_IN), .ZN(n2508) );
  AND2_X1 U2393 ( .A1(n3600), .A2(n3601), .ZN(n3516) );
  INV_X1 U2394 ( .A(DATAI_1_), .ZN(n2106) );
  INV_X1 U2395 ( .A(n2246), .ZN(n2244) );
  AOI21_X1 U2396 ( .B1(n2246), .B2(n2243), .A(n3656), .ZN(n2242) );
  NAND2_X1 U2397 ( .A1(n2259), .A2(n2258), .ZN(n2257) );
  INV_X1 U2398 ( .A(n3116), .ZN(n2258) );
  INV_X1 U2399 ( .A(n3115), .ZN(n2259) );
  AND2_X1 U2400 ( .A1(n2249), .A2(n2247), .ZN(n2246) );
  INV_X1 U2401 ( .A(n3654), .ZN(n2247) );
  OR2_X1 U2403 ( .A1(n2066), .A2(n4527), .ZN(n2214) );
  OR2_X1 U2404 ( .A1(n4518), .A2(n2215), .ZN(n2213) );
  OR2_X1 U2405 ( .A1(n4527), .A2(n4519), .ZN(n2215) );
  NOR2_X1 U2406 ( .A1(n4545), .A2(n2282), .ZN(n4080) );
  AOI21_X1 U2407 ( .B1(n2515), .B2(n2514), .A(n2513), .ZN(n3403) );
  NAND2_X1 U2408 ( .A1(n3435), .A2(n3458), .ZN(n2514) );
  INV_X1 U2409 ( .A(n2172), .ZN(n2170) );
  AND2_X1 U2410 ( .A1(n2077), .A2(n3487), .ZN(n2245) );
  INV_X1 U2411 ( .A(n2717), .ZN(n2716) );
  INV_X1 U2412 ( .A(n3861), .ZN(n2195) );
  AND2_X1 U2413 ( .A1(n4169), .A2(n3552), .ZN(n4151) );
  NOR2_X1 U2414 ( .A1(n2169), .A2(n3703), .ZN(n2168) );
  NOR2_X1 U2415 ( .A1(n2170), .A2(n2175), .ZN(n2169) );
  NAND2_X1 U2416 ( .A1(n2168), .A2(n2170), .ZN(n2167) );
  NOR2_X1 U2417 ( .A1(n2137), .A2(n3761), .ZN(n2131) );
  AND2_X1 U2418 ( .A1(n4204), .A2(n2653), .ZN(n3761) );
  AND2_X1 U2419 ( .A1(n2146), .A2(n3690), .ZN(n2145) );
  NAND2_X1 U2420 ( .A1(n2542), .A2(n2119), .ZN(n2118) );
  INV_X1 U2421 ( .A(n2121), .ZN(n2119) );
  AND2_X1 U2422 ( .A1(n4233), .A2(n4232), .ZN(n4294) );
  NOR2_X1 U2423 ( .A1(n2638), .A2(n2187), .ZN(n2186) );
  INV_X1 U2424 ( .A(n3803), .ZN(n2187) );
  NAND2_X1 U2425 ( .A1(n2162), .A2(n2087), .ZN(n2161) );
  INV_X1 U2426 ( .A(n2163), .ZN(n2162) );
  INV_X1 U2427 ( .A(n3790), .ZN(n2164) );
  INV_X1 U2428 ( .A(n3782), .ZN(n2177) );
  NAND2_X1 U2429 ( .A1(n3856), .A2(n3013), .ZN(n3783) );
  OR2_X1 U2430 ( .A1(n3337), .A2(n3219), .ZN(n2465) );
  NAND2_X1 U2431 ( .A1(n2627), .A2(n2719), .ZN(n3042) );
  INV_X1 U2432 ( .A(IR_REG_2__SCAN_IN), .ZN(n2341) );
  NOR2_X1 U2433 ( .A1(n2378), .A2(n2239), .ZN(n2238) );
  INV_X1 U2434 ( .A(n2310), .ZN(n2239) );
  NOR2_X1 U2435 ( .A1(n2307), .A2(n2378), .ZN(n2311) );
  INV_X1 U2436 ( .A(n2378), .ZN(n2661) );
  INV_X1 U2437 ( .A(IR_REG_11__SCAN_IN), .ZN(n2451) );
  INV_X1 U2438 ( .A(IR_REG_6__SCAN_IN), .ZN(n2400) );
  NOR2_X1 U2439 ( .A1(n2276), .A2(n3671), .ZN(n2275) );
  INV_X1 U2440 ( .A(n3630), .ZN(n2276) );
  AOI21_X1 U2441 ( .B1(n2275), .B2(n3629), .A(n2088), .ZN(n2274) );
  NAND2_X1 U2442 ( .A1(n2274), .A2(n2273), .ZN(n2272) );
  INV_X1 U2443 ( .A(n3589), .ZN(n2273) );
  INV_X1 U2444 ( .A(n3643), .ZN(n2266) );
  INV_X1 U2445 ( .A(n2272), .ZN(n2267) );
  INV_X1 U2446 ( .A(n2269), .ZN(n2264) );
  AOI21_X1 U2447 ( .B1(n2271), .B2(n2274), .A(n2270), .ZN(n2269) );
  NOR2_X1 U2448 ( .A1(n3542), .A2(n3543), .ZN(n2270) );
  NOR2_X1 U2449 ( .A1(n3589), .A2(n2275), .ZN(n2271) );
  OR2_X1 U2450 ( .A1(n2741), .A2(n3044), .ZN(n2734) );
  INV_X1 U2451 ( .A(n3443), .ZN(n3446) );
  XNOR2_X1 U2452 ( .A(n2757), .B(n3538), .ZN(n2761) );
  OR2_X1 U2453 ( .A1(n2741), .A2(n2754), .ZN(n2755) );
  NAND2_X1 U2454 ( .A1(n3115), .A2(n3116), .ZN(n2256) );
  OR2_X1 U2455 ( .A1(n2527), .A2(n2526), .ZN(n2536) );
  NAND2_X1 U2456 ( .A1(n3489), .A2(n2245), .ZN(n2248) );
  NAND2_X1 U2457 ( .A1(n2250), .A2(n2077), .ZN(n2249) );
  NAND2_X1 U2458 ( .A1(n3611), .A2(n2251), .ZN(n2250) );
  AND2_X1 U2459 ( .A1(n2543), .A2(REG3_REG_21__SCAN_IN), .ZN(n2548) );
  INV_X1 U2460 ( .A(n3838), .ZN(n2807) );
  INV_X1 U2461 ( .A(n3430), .ZN(n3427) );
  AND4_X1 U2462 ( .A1(n2376), .A2(n2375), .A3(n2374), .A4(n2373), .ZN(n2970)
         );
  NAND2_X1 U2463 ( .A1(n4439), .A2(n2322), .ZN(n2339) );
  AND2_X1 U2464 ( .A1(n2235), .A2(REG2_REG_0__SCAN_IN), .ZN(n2283) );
  OAI21_X1 U2465 ( .B1(n2344), .B2(n2101), .A(n2100), .ZN(n3885) );
  OR2_X1 U2466 ( .A1(n2343), .A2(REG2_REG_2__SCAN_IN), .ZN(n2101) );
  OAI21_X1 U2467 ( .B1(n2344), .B2(n2343), .A(REG2_REG_2__SCAN_IN), .ZN(n2100)
         );
  NAND2_X1 U2468 ( .A1(n2197), .A2(n2196), .ZN(n3879) );
  OAI21_X1 U2469 ( .B1(n2344), .B2(n2343), .A(REG1_REG_2__SCAN_IN), .ZN(n2196)
         );
  NAND2_X1 U2470 ( .A1(n2200), .A2(n2069), .ZN(n2197) );
  AOI21_X1 U2471 ( .B1(REG2_REG_5__SCAN_IN), .B2(n4447), .A(n2882), .ZN(n2864)
         );
  OAI211_X1 U2472 ( .C1(n2851), .C2(n2202), .A(n2201), .B(n2068), .ZN(n2852)
         );
  AOI21_X1 U2473 ( .B1(n2204), .B2(n2212), .A(n2203), .ZN(n2202) );
  NAND2_X1 U2474 ( .A1(n2219), .A2(n2221), .ZN(n2220) );
  AND2_X1 U2475 ( .A1(n4073), .A2(REG1_REG_8__SCAN_IN), .ZN(n2219) );
  AND3_X1 U2476 ( .A1(n2213), .A2(n2214), .A3(n2090), .ZN(n4076) );
  OAI21_X1 U2477 ( .B1(n4558), .B2(n2223), .A(n2222), .ZN(n4571) );
  NAND2_X1 U2478 ( .A1(n2226), .A2(REG1_REG_14__SCAN_IN), .ZN(n2223) );
  INV_X1 U2479 ( .A(n4572), .ZN(n2226) );
  OR2_X1 U2480 ( .A1(n4558), .A2(n4559), .ZN(n2225) );
  NAND2_X1 U2481 ( .A1(n4584), .A2(n2096), .ZN(n4605) );
  OR2_X1 U2482 ( .A1(n4639), .A2(REG2_REG_17__SCAN_IN), .ZN(n2096) );
  NAND2_X1 U2483 ( .A1(n4581), .A2(n4119), .ZN(n4596) );
  NOR2_X1 U2484 ( .A1(n4605), .A2(n4606), .ZN(n4604) );
  OR2_X1 U2485 ( .A1(n2595), .A2(n3553), .ZN(n4156) );
  OAI21_X1 U2486 ( .B1(n4161), .B2(n2594), .A(n2593), .ZN(n4139) );
  AOI21_X1 U2487 ( .B1(n2061), .B2(n2137), .A(n2083), .ZN(n2135) );
  INV_X1 U2488 ( .A(n2559), .ZN(n2136) );
  AOI22_X1 U2489 ( .A1(n4273), .A2(n2547), .B1(n4256), .B2(n4283), .ZN(n4255)
         );
  NAND2_X1 U2490 ( .A1(n2523), .A2(n2124), .ZN(n2121) );
  NAND2_X1 U2491 ( .A1(n2122), .A2(n2124), .ZN(n2120) );
  NAND2_X1 U2492 ( .A1(n3403), .A2(n3729), .ZN(n3402) );
  OR2_X1 U2493 ( .A1(n3358), .A2(n2085), .ZN(n2515) );
  NAND2_X1 U2494 ( .A1(n2497), .A2(n2281), .ZN(n3359) );
  NAND2_X1 U2495 ( .A1(n3848), .A2(n2495), .ZN(n2496) );
  NOR2_X1 U2496 ( .A1(n3359), .A2(n3755), .ZN(n3358) );
  OR2_X1 U2497 ( .A1(n2413), .A2(n2319), .ZN(n2433) );
  NAND2_X1 U2498 ( .A1(n2139), .A2(n2393), .ZN(n3079) );
  OR2_X1 U2499 ( .A1(n2969), .A2(n2968), .ZN(n2632) );
  AOI21_X1 U2500 ( .B1(n3180), .B2(n2358), .A(n2357), .ZN(n2995) );
  OR2_X1 U2501 ( .A1(n2824), .A2(D_REG_1__SCAN_IN), .ZN(n3001) );
  AND2_X1 U2502 ( .A1(n2785), .A2(n2827), .ZN(n3003) );
  NAND2_X1 U2503 ( .A1(n4345), .A2(n2112), .ZN(n4352) );
  OR2_X1 U2504 ( .A1(n4142), .A2(n4147), .ZN(n2112) );
  AOI21_X1 U2505 ( .B1(n2156), .B2(n3409), .A(n2154), .ZN(n4353) );
  INV_X1 U2506 ( .A(n2155), .ZN(n2154) );
  XNOR2_X1 U2507 ( .A(n2157), .B(n4153), .ZN(n2156) );
  AOI21_X1 U2508 ( .B1(n4169), .B2(n4325), .A(n4154), .ZN(n2155) );
  INV_X1 U2509 ( .A(IR_REG_30__SCAN_IN), .ZN(n2316) );
  OAI21_X1 U2510 ( .B1(n2816), .B2(IR_REG_29__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2140) );
  OR3_X1 U2512 ( .A1(n2409), .A2(IR_REG_7__SCAN_IN), .A3(IR_REG_8__SCAN_IN), 
        .ZN(n2439) );
  NAND2_X1 U2513 ( .A1(n2190), .A2(n2188), .ZN(n2333) );
  NAND2_X1 U2514 ( .A1(n2191), .A2(IR_REG_31__SCAN_IN), .ZN(n2190) );
  INV_X1 U2515 ( .A(n4204), .ZN(n4162) );
  AND2_X1 U2516 ( .A1(n3160), .A2(n3161), .ZN(n3158) );
  INV_X1 U2517 ( .A(n4300), .ZN(n3658) );
  INV_X1 U2518 ( .A(n4220), .ZN(n4182) );
  INV_X1 U2519 ( .A(n4472), .ZN(n3680) );
  NAND2_X1 U2520 ( .A1(n4503), .A2(n4095), .ZN(n4512) );
  NAND2_X1 U2521 ( .A1(n4102), .A2(n4540), .ZN(n4552) );
  XNOR2_X1 U2522 ( .A(n4080), .B(n4079), .ZN(n4558) );
  OR2_X1 U2523 ( .A1(n4484), .A2(n4440), .ZN(n4611) );
  INV_X1 U2524 ( .A(n4593), .ZN(n4603) );
  AOI21_X1 U2525 ( .B1(n4596), .B2(n4595), .A(n4594), .ZN(n4602) );
  INV_X1 U2526 ( .A(n4560), .ZN(n4608) );
  NOR2_X1 U2527 ( .A1(n3816), .A2(n2148), .ZN(n2147) );
  INV_X1 U2528 ( .A(n2150), .ZN(n2148) );
  NAND2_X1 U2529 ( .A1(n2147), .A2(n2153), .ZN(n2146) );
  NAND2_X1 U2530 ( .A1(n3858), .A2(n2722), .ZN(n3777) );
  INV_X1 U2531 ( .A(n2245), .ZN(n2243) );
  NOR2_X1 U2532 ( .A1(n2500), .A2(n2499), .ZN(n2516) );
  INV_X2 U2533 ( .A(n2772), .ZN(n2797) );
  NAND2_X1 U2534 ( .A1(n3883), .A2(n2858), .ZN(n2859) );
  NAND2_X1 U2535 ( .A1(n2210), .A2(n4448), .ZN(n2204) );
  NAND2_X1 U2536 ( .A1(n4447), .A2(REG1_REG_5__SCAN_IN), .ZN(n2212) );
  INV_X1 U2537 ( .A(n2206), .ZN(n2203) );
  NAND2_X1 U2538 ( .A1(n2212), .A2(n2363), .ZN(n2206) );
  AOI22_X1 U2539 ( .A1(REG2_REG_13__SCAN_IN), .A2(n4643), .B1(n4552), .B2(
        n4103), .ZN(n4104) );
  INV_X1 U2540 ( .A(IR_REG_18__SCAN_IN), .ZN(n2532) );
  NOR2_X1 U2541 ( .A1(n2174), .A2(n3726), .ZN(n2172) );
  OAI21_X1 U2542 ( .B1(n3818), .B2(n3695), .A(n3693), .ZN(n2174) );
  NAND2_X1 U2543 ( .A1(n2651), .A2(n2175), .ZN(n2173) );
  NOR2_X1 U2544 ( .A1(n3406), .A2(n3405), .ZN(n4233) );
  AOI21_X1 U2545 ( .B1(n3755), .B2(n2152), .A(n2151), .ZN(n2150) );
  INV_X1 U2546 ( .A(n3685), .ZN(n2152) );
  INV_X1 U2547 ( .A(n3813), .ZN(n2151) );
  INV_X1 U2548 ( .A(n3755), .ZN(n2153) );
  OAI21_X1 U2549 ( .B1(n3100), .B2(n2628), .A(n3773), .ZN(n2929) );
  NAND2_X1 U2550 ( .A1(n3777), .A2(n3774), .ZN(n2629) );
  NAND2_X1 U2551 ( .A1(n2744), .A2(n2334), .ZN(n3773) );
  OAI21_X1 U2552 ( .B1(n4152), .B2(n4151), .A(n4150), .ZN(n2157) );
  NOR2_X1 U2553 ( .A1(n4304), .A2(n2704), .ZN(n4266) );
  INV_X1 U2554 ( .A(IR_REG_26__SCAN_IN), .ZN(n2306) );
  INV_X1 U2555 ( .A(IR_REG_22__SCAN_IN), .ZN(n2668) );
  INV_X1 U2556 ( .A(IR_REG_20__SCAN_IN), .ZN(n2610) );
  INV_X1 U2557 ( .A(IR_REG_1__SCAN_IN), .ZN(n2191) );
  NAND2_X1 U2558 ( .A1(n2189), .A2(IR_REG_1__SCAN_IN), .ZN(n2188) );
  NAND2_X1 U2559 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2189)
         );
  INV_X1 U2560 ( .A(n2792), .ZN(n2790) );
  OAI22_X1 U2561 ( .A1(n3385), .A2(n3525), .B1(n3540), .B2(n3388), .ZN(n3422)
         );
  NAND2_X1 U2562 ( .A1(n2516), .A2(REG3_REG_18__SCAN_IN), .ZN(n2527) );
  AND2_X1 U2563 ( .A1(REG3_REG_12__SCAN_IN), .A2(REG3_REG_11__SCAN_IN), .ZN(
        n2320) );
  NOR2_X1 U2564 ( .A1(n2536), .A2(n4047), .ZN(n2543) );
  NAND2_X1 U2565 ( .A1(n2548), .A2(REG3_REG_22__SCAN_IN), .ZN(n2552) );
  INV_X1 U2566 ( .A(n2766), .ZN(n2230) );
  NAND2_X1 U2567 ( .A1(n2843), .A2(n2314), .ZN(n2104) );
  NAND2_X1 U2568 ( .A1(n2842), .A2(IR_REG_28__SCAN_IN), .ZN(n2105) );
  OR2_X1 U2569 ( .A1(n2719), .A2(n4443), .ZN(n2798) );
  INV_X1 U2570 ( .A(n3862), .ZN(n2193) );
  NAND2_X1 U2571 ( .A1(n3860), .A2(n2846), .ZN(n3878) );
  XNOR2_X1 U2572 ( .A(n2859), .B(n2897), .ZN(n2892) );
  XNOR2_X1 U2573 ( .A(n2851), .B(n4491), .ZN(n4486) );
  AOI22_X1 U2574 ( .A1(n2874), .A2(REG2_REG_6__SCAN_IN), .B1(n4446), .B2(n2865), .ZN(n2867) );
  OAI21_X1 U2575 ( .B1(n4092), .B2(n4091), .A(n4090), .ZN(n4094) );
  INV_X1 U2576 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3162) );
  NAND2_X1 U2577 ( .A1(n4511), .A2(n2081), .ZN(n4097) );
  OR2_X1 U2578 ( .A1(n4518), .A2(n4519), .ZN(n2216) );
  NOR2_X1 U2579 ( .A1(n4535), .A2(n4077), .ZN(n4547) );
  XNOR2_X1 U2580 ( .A(n4104), .B(n4079), .ZN(n4562) );
  NOR2_X1 U2581 ( .A1(n4562), .A2(n3238), .ZN(n4561) );
  NOR2_X1 U2582 ( .A1(n4571), .A2(n4083), .ZN(n4115) );
  NOR2_X1 U2583 ( .A1(n4345), .A2(n4348), .ZN(n4344) );
  AND2_X1 U2584 ( .A1(n3738), .A2(n3737), .ZN(n4153) );
  AOI21_X1 U2585 ( .B1(n2651), .B2(n2168), .A(n2166), .ZN(n2165) );
  NAND2_X1 U2586 ( .A1(n2167), .A2(n2655), .ZN(n2166) );
  INV_X1 U2587 ( .A(n3741), .ZN(n4165) );
  NAND2_X1 U2588 ( .A1(n2132), .A2(n2129), .ZN(n4161) );
  AOI21_X1 U2589 ( .B1(n2135), .B2(n2131), .A(n2130), .ZN(n2129) );
  INV_X1 U2590 ( .A(n3762), .ZN(n2130) );
  NAND2_X1 U2591 ( .A1(n2173), .A2(n2171), .ZN(n4200) );
  INV_X1 U2592 ( .A(n2174), .ZN(n2171) );
  AND2_X1 U2593 ( .A1(n2113), .A2(n2115), .ZN(n4273) );
  AND2_X1 U2594 ( .A1(n2086), .A2(n2116), .ZN(n2115) );
  OR2_X1 U2595 ( .A1(n3403), .A2(n2118), .ZN(n2113) );
  NAND2_X1 U2596 ( .A1(n2149), .A2(n2150), .ZN(n3406) );
  OR2_X1 U2597 ( .A1(n2643), .A2(n2153), .ZN(n2149) );
  NAND2_X1 U2598 ( .A1(n2643), .A2(n3685), .ZN(n3361) );
  AND2_X1 U2599 ( .A1(n3811), .A2(n3813), .ZN(n3755) );
  OR2_X1 U2600 ( .A1(n2487), .A2(n4452), .ZN(n2500) );
  NAND2_X1 U2601 ( .A1(n2126), .A2(n2125), .ZN(n3312) );
  AOI21_X1 U2602 ( .B1(n2060), .B2(n2076), .A(n2063), .ZN(n2125) );
  NAND2_X1 U2603 ( .A1(n2467), .A2(REG3_REG_13__SCAN_IN), .ZN(n2477) );
  OR2_X1 U2604 ( .A1(n2477), .A2(n2476), .ZN(n2487) );
  AOI21_X1 U2605 ( .B1(n2184), .B2(n3805), .A(n3231), .ZN(n2183) );
  INV_X1 U2606 ( .A(n2186), .ZN(n2184) );
  NAND2_X1 U2607 ( .A1(n2182), .A2(n3805), .ZN(n3687) );
  NAND2_X1 U2608 ( .A1(n3563), .A2(n2186), .ZN(n2182) );
  NAND2_X1 U2609 ( .A1(n3563), .A2(n3803), .ZN(n3217) );
  AND2_X1 U2610 ( .A1(n3216), .A2(n3803), .ZN(n3562) );
  OR2_X1 U2611 ( .A1(n3561), .A2(n3562), .ZN(n3559) );
  INV_X1 U2612 ( .A(n2454), .ZN(n3571) );
  NOR2_X1 U2613 ( .A1(n2161), .A2(n2160), .ZN(n2159) );
  NAND2_X1 U2614 ( .A1(n2158), .A2(n2161), .ZN(n3272) );
  NAND2_X1 U2615 ( .A1(n3065), .A2(n2089), .ZN(n2158) );
  AND2_X1 U2616 ( .A1(n3786), .A2(n3788), .ZN(n3727) );
  AOI21_X1 U2617 ( .B1(n2180), .B2(n2178), .A(n2177), .ZN(n2176) );
  INV_X1 U2618 ( .A(n2180), .ZN(n2179) );
  INV_X1 U2619 ( .A(n3783), .ZN(n2178) );
  INV_X1 U2620 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2384) );
  NOR2_X1 U2621 ( .A1(n2385), .A2(n2384), .ZN(n2394) );
  NAND2_X1 U2622 ( .A1(n3135), .A2(n2382), .ZN(n2138) );
  INV_X1 U2623 ( .A(n2991), .ZN(n3141) );
  AND2_X1 U2624 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2372) );
  OR2_X1 U2625 ( .A1(n3190), .A2(n3007), .ZN(n3142) );
  INV_X1 U2626 ( .A(n3858), .ZN(n3184) );
  NAND2_X1 U2627 ( .A1(n3098), .A2(n2628), .ZN(n3097) );
  NAND2_X1 U2628 ( .A1(n2729), .A2(n3096), .ZN(n3100) );
  NOR2_X1 U2629 ( .A1(n4170), .A2(n4137), .ZN(n4142) );
  NAND2_X1 U2630 ( .A1(n4187), .A2(n4171), .ZN(n4170) );
  NOR2_X1 U2631 ( .A1(n4223), .A2(n4208), .ZN(n4207) );
  AND2_X1 U2632 ( .A1(n4207), .A2(n4189), .ZN(n4187) );
  NAND2_X1 U2633 ( .A1(n2108), .A2(n4224), .ZN(n4223) );
  NAND2_X1 U2634 ( .A1(n4266), .A2(n4267), .ZN(n4375) );
  NAND2_X1 U2635 ( .A1(n2059), .A2(DATAI_20_), .ZN(n4305) );
  OR2_X1 U2636 ( .A1(n4329), .A2(n3722), .ZN(n4304) );
  NAND2_X1 U2637 ( .A1(n3458), .A2(n2110), .ZN(n2109) );
  NOR2_X1 U2638 ( .A1(n3469), .A2(n3365), .ZN(n2110) );
  NAND2_X1 U2639 ( .A1(n4331), .A2(n4330), .ZN(n4329) );
  AND2_X1 U2640 ( .A1(n3257), .A2(n3388), .ZN(n3318) );
  NAND2_X1 U2641 ( .A1(n2127), .A2(n2060), .ZN(n3230) );
  OR2_X1 U2642 ( .A1(n3244), .A2(n2076), .ZN(n2127) );
  NOR2_X1 U2643 ( .A1(n3256), .A2(n3250), .ZN(n3257) );
  NAND2_X1 U2644 ( .A1(n3572), .A2(n3571), .ZN(n3570) );
  INV_X1 U2645 ( .A(n3304), .ZN(n3219) );
  OR2_X1 U2646 ( .A1(n3570), .A2(n3219), .ZN(n3256) );
  NAND2_X1 U2647 ( .A1(n2107), .A2(n3284), .ZN(n3283) );
  NAND2_X1 U2648 ( .A1(n3074), .A2(n3073), .ZN(n3072) );
  INV_X1 U2649 ( .A(n3059), .ZN(n3025) );
  NOR2_X1 U2650 ( .A1(n3142), .A2(n3141), .ZN(n3144) );
  AND2_X1 U2651 ( .A1(n3144), .A2(n2978), .ZN(n3074) );
  NAND2_X1 U2652 ( .A1(n2745), .A2(n3044), .ZN(n3094) );
  INV_X1 U2653 ( .A(n2786), .ZN(n3004) );
  AND3_X1 U2654 ( .A1(n2697), .A2(n2696), .A3(n2785), .ZN(n2709) );
  INV_X1 U2655 ( .A(n2307), .ZN(n2240) );
  INV_X1 U2656 ( .A(IR_REG_4__SCAN_IN), .ZN(n2141) );
  INV_X1 U2657 ( .A(IR_REG_16__SCAN_IN), .ZN(n2299) );
  INV_X1 U2658 ( .A(IR_REG_14__SCAN_IN), .ZN(n2298) );
  INV_X1 U2659 ( .A(IR_REG_21__SCAN_IN), .ZN(n2613) );
  AND2_X1 U2660 ( .A1(n2456), .A2(n2453), .ZN(n4089) );
  NOR2_X1 U2661 ( .A1(n2378), .A2(IR_REG_5__SCAN_IN), .ZN(n2401) );
  MUX2_X1 U2662 ( .A(n2617), .B(n2340), .S(IR_REG_2__SCAN_IN), .Z(n2344) );
  INV_X1 U2663 ( .A(n3066), .ZN(n3073) );
  AND4_X1 U2664 ( .A1(n2417), .A2(n2416), .A3(n2415), .A4(n2414), .ZN(n3275)
         );
  NAND2_X1 U2665 ( .A1(n2268), .A2(n2274), .ZN(n3590) );
  NOR2_X1 U2666 ( .A1(n2254), .A2(n3120), .ZN(n2253) );
  INV_X1 U2667 ( .A(n2256), .ZN(n2254) );
  AOI21_X1 U2668 ( .B1(n3641), .B2(n2265), .A(n2264), .ZN(n2260) );
  NAND2_X1 U2669 ( .A1(n3640), .A2(n2267), .ZN(n2261) );
  NOR2_X1 U2670 ( .A1(n2272), .A2(n2266), .ZN(n2265) );
  AND2_X1 U2671 ( .A1(n4156), .A2(n2596), .ZN(n3582) );
  AND4_X1 U2672 ( .A1(n2399), .A2(n2398), .A3(n2397), .A4(n2396), .ZN(n3058)
         );
  INV_X1 U2673 ( .A(n3846), .ZN(n4322) );
  AND4_X1 U2674 ( .A1(n2447), .A2(n2446), .A3(n2445), .A4(n2444), .ZN(n3306)
         );
  NAND2_X1 U2675 ( .A1(n3446), .A2(n3445), .ZN(n3447) );
  INV_X1 U2676 ( .A(n3444), .ZN(n3445) );
  CLKBUF_X1 U2677 ( .A(n2956), .Z(n2957) );
  NAND2_X1 U2678 ( .A1(n2255), .A2(n2256), .ZN(n3119) );
  INV_X1 U2679 ( .A(n3677), .ZN(n4454) );
  NAND2_X1 U2680 ( .A1(n2248), .A2(n2249), .ZN(n3653) );
  INV_X1 U2681 ( .A(n4465), .ZN(n3665) );
  OR2_X1 U2682 ( .A1(n2809), .A2(n2800), .ZN(n3675) );
  NAND2_X1 U2683 ( .A1(n2592), .A2(n2591), .ZN(n4184) );
  OR2_X1 U2684 ( .A1(n3591), .A2(n2579), .ZN(n2592) );
  NAND2_X1 U2685 ( .A1(n2584), .A2(n2583), .ZN(n4204) );
  NAND2_X1 U2686 ( .A1(n2574), .A2(n2573), .ZN(n4220) );
  OR2_X1 U2687 ( .A1(n3634), .A2(n2579), .ZN(n2574) );
  OAI211_X1 U2688 ( .C1(n4285), .C2(n2339), .A(n2546), .B(n2545), .ZN(n4299)
         );
  OR2_X1 U2689 ( .A1(n2530), .A2(n2529), .ZN(n4300) );
  INV_X1 U2690 ( .A(n3564), .ZN(n3337) );
  INV_X1 U2691 ( .A(n3306), .ZN(n3850) );
  NAND4_X1 U2692 ( .A1(n2438), .A2(n2437), .A3(n2436), .A4(n2435), .ZN(n3851)
         );
  OR2_X1 U2693 ( .A1(n2408), .A2(n2407), .ZN(n3852) );
  INV_X1 U2694 ( .A(n3058), .ZN(n3853) );
  INV_X1 U2695 ( .A(n3138), .ZN(n3856) );
  OR2_X1 U2696 ( .A1(n2579), .A2(REG3_REG_3__SCAN_IN), .ZN(n2353) );
  NAND2_X1 U2697 ( .A1(n2345), .A2(n2067), .ZN(n3858) );
  AND2_X1 U2698 ( .A1(n2331), .A2(n2234), .ZN(n2233) );
  NAND2_X1 U2699 ( .A1(n2338), .A2(REG0_REG_1__SCAN_IN), .ZN(n2330) );
  NAND2_X1 U2700 ( .A1(n2235), .A2(REG2_REG_1__SCAN_IN), .ZN(n2232) );
  NOR2_X1 U2701 ( .A1(n2283), .A2(n2143), .ZN(n2335) );
  OAI21_X1 U2702 ( .B1(n2339), .B2(n2917), .A(n2142), .ZN(n2143) );
  NAND2_X1 U2703 ( .A1(n2199), .A2(n2198), .ZN(n3861) );
  NOR2_X1 U2704 ( .A1(n2211), .A2(REG1_REG_4__SCAN_IN), .ZN(n2205) );
  AND2_X1 U2705 ( .A1(n2209), .A2(n2208), .ZN(n2885) );
  INV_X1 U2706 ( .A(n2211), .ZN(n2209) );
  NAND2_X1 U2707 ( .A1(n4486), .A2(REG1_REG_4__SCAN_IN), .ZN(n2208) );
  XNOR2_X1 U2708 ( .A(n2864), .B(n4446), .ZN(n2874) );
  OR2_X1 U2709 ( .A1(n2867), .A2(n2866), .ZN(n4090) );
  AOI22_X1 U2710 ( .A1(n2875), .A2(REG1_REG_6__SCAN_IN), .B1(n4446), .B2(n2853), .ZN(n4069) );
  INV_X1 U2711 ( .A(n2220), .ZN(n4498) );
  NAND2_X1 U2712 ( .A1(n4512), .A2(n4513), .ZN(n4511) );
  NAND2_X1 U2713 ( .A1(n4073), .A2(n2218), .ZN(n2217) );
  NOR2_X1 U2714 ( .A1(n4508), .A2(n2411), .ZN(n2218) );
  XNOR2_X1 U2715 ( .A(n4097), .B(n4650), .ZN(n4523) );
  NAND2_X1 U2716 ( .A1(n2214), .A2(n2213), .ZN(n4526) );
  NOR2_X1 U2717 ( .A1(n4536), .A2(n4537), .ZN(n4535) );
  INV_X1 U2718 ( .A(n4643), .ZN(n4556) );
  INV_X1 U2719 ( .A(n2225), .ZN(n4557) );
  OAI21_X1 U2720 ( .B1(n4562), .B2(n2098), .A(n2097), .ZN(n4575) );
  NAND2_X1 U2721 ( .A1(n2099), .A2(REG2_REG_14__SCAN_IN), .ZN(n2098) );
  NAND2_X1 U2722 ( .A1(n4105), .A2(n2099), .ZN(n2097) );
  INV_X1 U2723 ( .A(n4576), .ZN(n2099) );
  INV_X1 U2724 ( .A(n4081), .ZN(n2224) );
  XNOR2_X1 U2725 ( .A(n2095), .B(n4129), .ZN(n4134) );
  NOR2_X1 U2726 ( .A1(n4604), .A2(n2094), .ZN(n2095) );
  OR2_X1 U2727 ( .A1(n4484), .A2(n4481), .ZN(n4594) );
  NAND2_X1 U2728 ( .A1(n2128), .A2(n2135), .ZN(n4178) );
  OR2_X1 U2729 ( .A1(n2560), .A2(n2286), .ZN(n2128) );
  NAND2_X1 U2730 ( .A1(n2114), .A2(n2120), .ZN(n4291) );
  OR2_X1 U2731 ( .A1(n3403), .A2(n2121), .ZN(n2114) );
  NAND2_X1 U2732 ( .A1(n3402), .A2(n2523), .ZN(n4313) );
  INV_X1 U2733 ( .A(n2515), .ZN(n3372) );
  OR2_X1 U2734 ( .A1(n4479), .A2(n3081), .ZN(n4338) );
  OAI21_X1 U2735 ( .B1(n4352), .B2(n4698), .A(n2072), .ZN(n4408) );
  NAND3_X1 U2736 ( .A1(n2240), .A2(n2236), .A3(n2506), .ZN(n2816) );
  NOR2_X1 U2737 ( .A1(n2378), .A2(n2237), .ZN(n2236) );
  NAND2_X1 U2738 ( .A1(n2310), .A2(n2314), .ZN(n2237) );
  INV_X1 U2739 ( .A(n2627), .ZN(n3771) );
  INV_X1 U2740 ( .A(n4132), .ZN(n4443) );
  XNOR2_X1 U2741 ( .A(n2457), .B(IR_REG_12__SCAN_IN), .ZN(n4645) );
  XNOR2_X1 U2742 ( .A(n2410), .B(IR_REG_9__SCAN_IN), .ZN(n4651) );
  INV_X1 U2743 ( .A(IR_REG_8__SCAN_IN), .ZN(n2421) );
  AND2_X1 U2744 ( .A1(n2368), .A2(n2356), .ZN(n4449) );
  NOR2_X1 U2745 ( .A1(n2344), .A2(n2343), .ZN(n4450) );
  NAND2_X1 U2746 ( .A1(n2955), .A2(n2766), .ZN(n2986) );
  AOI21_X1 U2747 ( .B1(n4603), .B2(n4602), .A(n4601), .ZN(n4610) );
  NAND2_X1 U2748 ( .A1(n4714), .A2(REG1_REG_28__SCAN_IN), .ZN(n2711) );
  AND2_X1 U2749 ( .A1(n2280), .A2(n3231), .ZN(n2060) );
  INV_X1 U2750 ( .A(n2745), .ZN(n2334) );
  AND3_X1 U2751 ( .A1(n2240), .A2(n2506), .A3(n2238), .ZN(n2315) );
  OR2_X1 U2752 ( .A1(n4197), .A2(n2136), .ZN(n2061) );
  OR3_X1 U2753 ( .A1(n3366), .A2(n3452), .A3(n3365), .ZN(n2062) );
  AND2_X1 U2754 ( .A1(n3385), .A2(n3388), .ZN(n2063) );
  AND2_X1 U2755 ( .A1(n3788), .A2(n3794), .ZN(n2064) );
  AND2_X1 U2756 ( .A1(n2087), .A2(n2064), .ZN(n2065) );
  INV_X1 U2757 ( .A(n4074), .ZN(n2221) );
  NAND2_X1 U2758 ( .A1(n2241), .A2(n2945), .ZN(n2789) );
  XNOR2_X1 U2759 ( .A(n2614), .B(n2613), .ZN(n2627) );
  OR2_X1 U2760 ( .A1(n4075), .A2(n4650), .ZN(n2066) );
  NAND2_X1 U2761 ( .A1(n2560), .A2(n2559), .ZN(n4195) );
  NAND2_X1 U2762 ( .A1(n3663), .A2(n3664), .ZN(n3599) );
  AND3_X1 U2763 ( .A1(n2347), .A2(n2346), .A3(n2348), .ZN(n2067) );
  INV_X1 U2764 ( .A(n2252), .ZN(n3619) );
  OR2_X1 U2765 ( .A1(n2206), .A2(n4448), .ZN(n2068) );
  INV_X1 U2766 ( .A(n2327), .ZN(n2322) );
  INV_X1 U2767 ( .A(n3044), .ZN(n3096) );
  NOR2_X1 U2768 ( .A1(n2343), .A2(REG1_REG_2__SCAN_IN), .ZN(n2069) );
  AND2_X1 U2769 ( .A1(n2790), .A2(n2945), .ZN(n2070) );
  NAND2_X1 U2770 ( .A1(n2248), .A2(n2246), .ZN(n2071) );
  INV_X1 U2771 ( .A(IR_REG_28__SCAN_IN), .ZN(n2314) );
  INV_X1 U2772 ( .A(n2075), .ZN(n2210) );
  AND2_X1 U2773 ( .A1(n4354), .A2(n4353), .ZN(n2072) );
  NAND2_X1 U2774 ( .A1(n3854), .A2(n2776), .ZN(n2073) );
  NOR2_X1 U2775 ( .A1(n4072), .A2(n4654), .ZN(n4074) );
  AND2_X1 U2776 ( .A1(n2073), .A2(n2383), .ZN(n2074) );
  INV_X1 U2777 ( .A(IR_REG_27__SCAN_IN), .ZN(n2312) );
  AND2_X1 U2778 ( .A1(n3389), .A2(n3340), .ZN(n2076) );
  NAND2_X1 U2779 ( .A1(n3497), .A2(n3496), .ZN(n2077) );
  AND2_X1 U2780 ( .A1(n2127), .A2(n2280), .ZN(n2078) );
  AND2_X1 U2781 ( .A1(n2173), .A2(n2172), .ZN(n2079) );
  NOR2_X1 U2782 ( .A1(n4561), .A2(n4105), .ZN(n2080) );
  INV_X1 U2783 ( .A(n2108), .ZN(n4245) );
  INV_X1 U2784 ( .A(n2111), .ZN(n4398) );
  NOR2_X1 U2785 ( .A1(n3366), .A2(n3365), .ZN(n2111) );
  OR2_X1 U2786 ( .A1(n4516), .A2(n4096), .ZN(n2081) );
  AND2_X1 U2787 ( .A1(n2225), .A2(n2224), .ZN(n2082) );
  AND4_X1 U2788 ( .A1(n2492), .A2(n2491), .A3(n2490), .A4(n2489), .ZN(n3433)
         );
  INV_X1 U2789 ( .A(n3433), .ZN(n3848) );
  AND2_X1 U2790 ( .A1(n4220), .A2(n4208), .ZN(n2083) );
  INV_X1 U2791 ( .A(n2286), .ZN(n2137) );
  AND2_X1 U2792 ( .A1(n3508), .A2(n3507), .ZN(n2084) );
  INV_X1 U2793 ( .A(n2523), .ZN(n2123) );
  AND2_X1 U2794 ( .A1(n3502), .A2(n3501), .ZN(n3656) );
  OAI21_X1 U2795 ( .B1(n3729), .B2(n2123), .A(n2535), .ZN(n2122) );
  AND2_X1 U2796 ( .A1(n4453), .A2(n3365), .ZN(n2085) );
  OR2_X1 U2797 ( .A1(n4322), .A2(n4305), .ZN(n2086) );
  INV_X1 U2798 ( .A(n3385), .ZN(n4455) );
  AND4_X1 U2799 ( .A1(n2482), .A2(n2481), .A3(n2480), .A4(n2479), .ZN(n3385)
         );
  AND4_X1 U2800 ( .A1(n2472), .A2(n2471), .A3(n2470), .A4(n2469), .ZN(n3389)
         );
  INV_X1 U2801 ( .A(n3805), .ZN(n2185) );
  NAND2_X1 U2802 ( .A1(n2336), .A2(n2335), .ZN(n2733) );
  NAND2_X1 U2803 ( .A1(n3067), .A2(n3059), .ZN(n2087) );
  NAND2_X1 U2804 ( .A1(n2138), .A2(n2383), .ZN(n2967) );
  INV_X1 U2805 ( .A(n3794), .ZN(n2160) );
  NAND2_X1 U2806 ( .A1(n3559), .A2(n2455), .ZN(n3215) );
  AND2_X1 U2807 ( .A1(n3533), .A2(n3532), .ZN(n2088) );
  INV_X1 U2808 ( .A(n3793), .ZN(n2181) );
  AND2_X1 U2809 ( .A1(n2087), .A2(n3788), .ZN(n2089) );
  INV_X1 U2810 ( .A(n3458), .ZN(n3452) );
  INV_X1 U2811 ( .A(n2107), .ZN(n3282) );
  NAND2_X1 U2812 ( .A1(n4089), .A2(REG1_REG_11__SCAN_IN), .ZN(n2090) );
  AND2_X1 U2813 ( .A1(n2220), .A2(n2221), .ZN(n2091) );
  AND2_X1 U2814 ( .A1(n2216), .A2(n2066), .ZN(n2092) );
  AND2_X1 U2815 ( .A1(n2851), .A2(n4448), .ZN(n2211) );
  NAND2_X1 U2816 ( .A1(n2956), .A2(n2762), .ZN(n2955) );
  NAND2_X1 U2817 ( .A1(n3097), .A2(n2337), .ZN(n2925) );
  NOR2_X1 U2818 ( .A1(n2207), .A2(n2205), .ZN(n2093) );
  INV_X1 U2819 ( .A(IR_REG_0__SCAN_IN), .ZN(n2103) );
  INV_X1 U2820 ( .A(IR_REG_3__SCAN_IN), .ZN(n3960) );
  INV_X1 U2821 ( .A(DATAI_0_), .ZN(n2102) );
  AND2_X1 U2822 ( .A1(n4128), .A2(REG2_REG_18__SCAN_IN), .ZN(n2094) );
  NAND2_X1 U2823 ( .A1(n3884), .A2(n3885), .ZN(n3883) );
  MUX2_X1 U2824 ( .A(n2103), .B(n2102), .S(n2059), .Z(n3044) );
  MUX2_X1 U2825 ( .A(n2855), .B(n2106), .S(n3702), .Z(n2745) );
  NAND3_X1 U2826 ( .A1(n3097), .A2(n2337), .A3(n2629), .ZN(n2927) );
  NAND3_X1 U2827 ( .A1(n2345), .A2(n2067), .A3(n2936), .ZN(n3774) );
  NAND2_X1 U2828 ( .A1(n3244), .A2(n2060), .ZN(n2126) );
  NAND2_X1 U2829 ( .A1(n3215), .A2(n2288), .ZN(n2466) );
  OAI21_X1 U2830 ( .B1(n3084), .B2(n2442), .A(n2441), .ZN(n3561) );
  NAND2_X1 U2831 ( .A1(n2560), .A2(n2133), .ZN(n2132) );
  NAND2_X1 U2832 ( .A1(n2138), .A2(n2074), .ZN(n2139) );
  NOR2_X1 U2833 ( .A1(n2432), .A2(n2431), .ZN(n3084) );
  NOR2_X1 U2834 ( .A1(n4575), .A2(n4107), .ZN(n4125) );
  NOR2_X1 U2835 ( .A1(n2884), .A2(n2883), .ZN(n2882) );
  NAND2_X1 U2836 ( .A1(n2995), .A2(n3728), .ZN(n2997) );
  AOI22_X1 U2837 ( .A1(n4139), .A2(n4138), .B1(n4137), .B2(n4169), .ZN(n4141)
         );
  NAND2_X1 U2838 ( .A1(n2927), .A2(n2349), .ZN(n3180) );
  NOR2_X1 U2839 ( .A1(n3079), .A2(n2425), .ZN(n2432) );
  NAND2_X1 U2840 ( .A1(n2997), .A2(n2370), .ZN(n3135) );
  NAND2_X1 U2841 ( .A1(n2816), .A2(IR_REG_31__SCAN_IN), .ZN(n2318) );
  NAND2_X2 U2842 ( .A1(n2322), .A2(n2328), .ZN(n3698) );
  NAND3_X1 U2843 ( .A1(n2322), .A2(n2328), .A3(REG1_REG_0__SCAN_IN), .ZN(n2142) );
  NAND2_X1 U2844 ( .A1(n3732), .A2(n2929), .ZN(n2928) );
  NAND2_X1 U2845 ( .A1(n2144), .A2(n2145), .ZN(n2647) );
  NAND2_X1 U2846 ( .A1(n2643), .A2(n2147), .ZN(n2144) );
  AOI21_X1 U2847 ( .B1(n3065), .B2(n2065), .A(n2159), .ZN(n2634) );
  OAI21_X1 U2848 ( .B1(n3065), .B2(n2633), .A(n3788), .ZN(n3021) );
  AOI21_X1 U2849 ( .B1(n2633), .B2(n3788), .A(n2164), .ZN(n2163) );
  INV_X1 U2850 ( .A(n2165), .ZN(n4164) );
  NOR2_X1 U2851 ( .A1(n2651), .A2(n2650), .ZN(n4215) );
  INV_X1 U2852 ( .A(n3818), .ZN(n2175) );
  OAI21_X1 U2853 ( .B1(n3006), .B2(n2179), .A(n2176), .ZN(n2969) );
  OAI21_X1 U2854 ( .B1(n3006), .B2(n2631), .A(n3783), .ZN(n3136) );
  AOI21_X1 U2855 ( .B1(n2631), .B2(n3783), .A(n2181), .ZN(n2180) );
  OAI21_X1 U2856 ( .B1(n3563), .B2(n2185), .A(n2183), .ZN(n3313) );
  NAND3_X1 U2857 ( .A1(n3879), .A2(n2194), .A3(n2192), .ZN(n3877) );
  NAND2_X1 U2858 ( .A1(n2846), .A2(n2193), .ZN(n2192) );
  NAND2_X1 U2859 ( .A1(n2195), .A2(n2846), .ZN(n2194) );
  NAND2_X1 U2860 ( .A1(n2855), .A2(REG1_REG_1__SCAN_IN), .ZN(n2198) );
  OR2_X1 U2861 ( .A1(n2855), .A2(REG1_REG_1__SCAN_IN), .ZN(n2199) );
  NAND2_X1 U2862 ( .A1(n3861), .A2(n3862), .ZN(n3860) );
  NAND3_X1 U2863 ( .A1(n2851), .A2(n2075), .A3(n2212), .ZN(n2201) );
  INV_X1 U2864 ( .A(n2216), .ZN(n4517) );
  OAI22_X1 U2865 ( .A1(n2217), .A2(n4074), .B1(n2221), .B2(n4508), .ZN(n4507)
         );
  NAND2_X1 U2866 ( .A1(n2221), .A2(n4073), .ZN(n4499) );
  NAND2_X1 U2867 ( .A1(n4081), .A2(n2226), .ZN(n2222) );
  OAI21_X1 U2868 ( .B1(n2956), .B2(n2230), .A(n2227), .ZN(n2231) );
  INV_X1 U2869 ( .A(n2985), .ZN(n2228) );
  INV_X1 U2870 ( .A(n2762), .ZN(n2229) );
  NAND2_X1 U2871 ( .A1(n2231), .A2(n2771), .ZN(n2944) );
  NAND3_X1 U2872 ( .A1(n2322), .A2(n2328), .A3(REG1_REG_1__SCAN_IN), .ZN(n2234) );
  INV_X1 U2873 ( .A(n2328), .ZN(n4439) );
  OAI21_X1 U2874 ( .B1(n3489), .B2(n3488), .A(n3487), .ZN(n3612) );
  NAND2_X1 U2875 ( .A1(n3488), .A2(n3487), .ZN(n2251) );
  INV_X1 U2876 ( .A(n3640), .ZN(n2262) );
  NAND2_X1 U2877 ( .A1(n3641), .A2(n3643), .ZN(n2263) );
  NAND2_X1 U2878 ( .A1(n2261), .A2(n2260), .ZN(n3551) );
  AND2_X2 U2879 ( .A1(n2263), .A2(n2262), .ZN(n3633) );
  NAND3_X1 U2880 ( .A1(n2263), .A2(n2262), .A3(n2275), .ZN(n2268) );
  NAND2_X1 U2881 ( .A1(n2710), .A2(n4716), .ZN(n2712) );
  OAI21_X1 U2882 ( .B1(n2710), .B2(n4703), .A(n2703), .ZN(n2708) );
  INV_X1 U2883 ( .A(IR_REG_19__SCAN_IN), .ZN(n2607) );
  NAND2_X2 U2884 ( .A1(n3206), .A2(n3205), .ZN(n3298) );
  NAND2_X1 U2885 ( .A1(n2665), .A2(n2311), .ZN(n2676) );
  XNOR2_X1 U2886 ( .A(n2743), .B(n3538), .ZN(n2749) );
  OAI22_X1 U2887 ( .A1(n2744), .A2(n2742), .B1(n2741), .B2(n2745), .ZN(n2743)
         );
  NAND2_X1 U2888 ( .A1(n4351), .A2(n4694), .ZN(n4354) );
  AND2_X1 U2889 ( .A1(n2607), .A2(n2610), .ZN(n2279) );
  OR2_X1 U2890 ( .A1(n3389), .A2(n3340), .ZN(n2280) );
  OR2_X1 U2891 ( .A1(n3848), .A2(n2495), .ZN(n2281) );
  INV_X1 U2892 ( .A(n4459), .ZN(n2495) );
  INV_X1 U2893 ( .A(n3340), .ZN(n3250) );
  AND2_X1 U2894 ( .A1(n4643), .A2(REG1_REG_13__SCAN_IN), .ZN(n2282) );
  INV_X1 U2895 ( .A(n4698), .ZN(n2707) );
  OR2_X1 U2896 ( .A1(n4240), .A2(n4267), .ZN(n2284) );
  INV_X1 U2897 ( .A(n2715), .ZN(U4043) );
  OR2_X1 U2898 ( .A1(n3584), .A2(n4435), .ZN(n2285) );
  OR2_X1 U2899 ( .A1(n2576), .A2(n2575), .ZN(n2286) );
  INV_X1 U2900 ( .A(n3232), .ZN(n3388) );
  OR2_X1 U2901 ( .A1(n4263), .A2(n3604), .ZN(n2287) );
  OR2_X1 U2902 ( .A1(n3304), .A2(n3564), .ZN(n2288) );
  AND2_X1 U2903 ( .A1(n2558), .A2(n2557), .ZN(n4218) );
  INV_X1 U2904 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2844) );
  AND2_X1 U2905 ( .A1(n2654), .A2(n3725), .ZN(n3826) );
  NAND2_X1 U2906 ( .A1(n3859), .A2(n2745), .ZN(n3769) );
  AND2_X1 U2907 ( .A1(n2309), .A2(n2312), .ZN(n2310) );
  OR2_X1 U2908 ( .A1(n2729), .A2(n2746), .ZN(n2732) );
  NAND2_X1 U2909 ( .A1(n4263), .A2(n3604), .ZN(n2559) );
  NOR2_X1 U2910 ( .A1(n2749), .A2(n2748), .ZN(n2750) );
  INV_X1 U2911 ( .A(n3675), .ZN(n4456) );
  NAND2_X1 U2912 ( .A1(n2577), .A2(REG3_REG_26__SCAN_IN), .ZN(n2585) );
  AND2_X1 U2913 ( .A1(n2567), .A2(REG3_REG_25__SCAN_IN), .ZN(n2577) );
  NAND2_X1 U2914 ( .A1(n4072), .A2(n4654), .ZN(n4073) );
  INV_X1 U2915 ( .A(n4565), .ZN(n4079) );
  OR2_X1 U2916 ( .A1(n4639), .A2(REG1_REG_17__SCAN_IN), .ZN(n4119) );
  OR2_X1 U2917 ( .A1(n4324), .A2(n3469), .ZN(n2523) );
  AND2_X1 U2918 ( .A1(n3847), .A2(n3452), .ZN(n2513) );
  NAND2_X1 U2919 ( .A1(n2372), .A2(REG3_REG_5__SCAN_IN), .ZN(n2385) );
  INV_X1 U2920 ( .A(n2629), .ZN(n3732) );
  AND2_X1 U2921 ( .A1(n4440), .A2(n2836), .ZN(n4325) );
  INV_X1 U2922 ( .A(IR_REG_29__SCAN_IN), .ZN(n2317) );
  NOR2_X1 U2923 ( .A1(n2439), .A2(IR_REG_9__SCAN_IN), .ZN(n2449) );
  OR2_X1 U2924 ( .A1(n2552), .A2(n3605), .ZN(n2561) );
  NAND2_X1 U2925 ( .A1(n3328), .A2(n3327), .ZN(n3383) );
  INV_X1 U2926 ( .A(n2776), .ZN(n2978) );
  OR2_X1 U2927 ( .A1(n2585), .A2(n3592), .ZN(n2595) );
  NOR2_X1 U2928 ( .A1(n2561), .A2(n3646), .ZN(n2567) );
  AND4_X1 U2929 ( .A1(n2326), .A2(n2325), .A3(n2324), .A4(n2323), .ZN(n3420)
         );
  AND4_X1 U2930 ( .A1(n2464), .A2(n2463), .A3(n2462), .A4(n2461), .ZN(n3564)
         );
  XNOR2_X1 U2931 ( .A(n2848), .B(n2897), .ZN(n2891) );
  NOR2_X1 U2932 ( .A1(n4547), .A2(n4546), .ZN(n4545) );
  NAND2_X1 U2933 ( .A1(n4582), .A2(n4583), .ZN(n4581) );
  INV_X1 U2934 ( .A(n4598), .ZN(n4599) );
  OR2_X1 U2935 ( .A1(n3042), .A2(n3834), .ZN(n4320) );
  INV_X1 U2936 ( .A(n4624), .ZN(n4335) );
  INV_X1 U2937 ( .A(n4325), .ZN(n4277) );
  OR2_X1 U2938 ( .A1(n4479), .A2(n4443), .ZN(n3415) );
  OR2_X1 U2939 ( .A1(n2824), .A2(D_REG_0__SCAN_IN), .ZN(n2701) );
  INV_X1 U2940 ( .A(n4321), .ZN(n4298) );
  AND2_X1 U2941 ( .A1(n2657), .A2(n2656), .ZN(n4327) );
  OR2_X1 U2942 ( .A1(n2824), .A2(n2695), .ZN(n2785) );
  OR2_X1 U2943 ( .A1(n2483), .A2(IR_REG_14__SCAN_IN), .ZN(n2485) );
  OR2_X1 U2944 ( .A1(n2809), .A2(n2808), .ZN(n3677) );
  NAND2_X1 U2945 ( .A1(n2394), .A2(REG3_REG_7__SCAN_IN), .ZN(n2413) );
  AND2_X1 U2946 ( .A1(n2459), .A2(n2320), .ZN(n2467) );
  OR2_X1 U2947 ( .A1(n3674), .A2(n2579), .ZN(n2584) );
  INV_X1 U2948 ( .A(n3420), .ZN(n4453) );
  NAND2_X1 U2949 ( .A1(n4600), .A2(n4599), .ZN(n4601) );
  OR2_X1 U2950 ( .A1(n4151), .A2(n4149), .ZN(n4138) );
  OR2_X1 U2951 ( .A1(n3000), .A2(n2805), .ZN(n4155) );
  INV_X1 U2952 ( .A(n4327), .ZN(n3409) );
  AND2_X1 U2953 ( .A1(n2701), .A2(n2700), .ZN(n2786) );
  NAND2_X1 U2954 ( .A1(n4703), .A2(n2702), .ZN(n2703) );
  AND2_X1 U2955 ( .A1(n3046), .A2(n2719), .ZN(n4675) );
  NAND2_X1 U2956 ( .A1(n2678), .A2(n4441), .ZN(n2824) );
  AND2_X1 U2957 ( .A1(n2486), .A2(n2485), .ZN(n4565) );
  NAND2_X1 U2958 ( .A1(n2380), .A2(n2379), .ZN(n2887) );
  AND2_X1 U2959 ( .A1(n2841), .A2(n2838), .ZN(n4597) );
  NAND2_X1 U2960 ( .A1(n2804), .A2(n2788), .ZN(n4465) );
  AND2_X1 U2961 ( .A1(n2799), .A2(n2901), .ZN(n4472) );
  NAND2_X1 U2962 ( .A1(n2602), .A2(n2601), .ZN(n4169) );
  OAI211_X1 U2963 ( .C1(n4307), .C2(n2579), .A(n2541), .B(n2540), .ZN(n3846)
         );
  INV_X1 U2964 ( .A(n3389), .ZN(n3849) );
  INV_X1 U2965 ( .A(n2970), .ZN(n3855) );
  INV_X1 U2966 ( .A(n4449), .ZN(n2897) );
  INV_X1 U2967 ( .A(n4645), .ZN(n4544) );
  NAND2_X1 U2968 ( .A1(n2712), .A2(n2711), .ZN(n2714) );
  INV_X1 U2969 ( .A(n4716), .ZN(n4714) );
  NAND2_X1 U2970 ( .A1(n4705), .A2(n2707), .ZN(n4435) );
  INV_X1 U2971 ( .A(n4705), .ZN(n4703) );
  INV_X1 U2972 ( .A(n4106), .ZN(n4641) );
  OR2_X1 U2973 ( .A1(n2714), .A2(n2713), .ZN(U3546) );
  NOR2_X1 U2974 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2292)
         );
  NOR2_X2 U2975 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2291)
         );
  NOR2_X2 U2976 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2290)
         );
  NOR2_X2 U2977 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2289)
         );
  AND4_X2 U2978 ( .A1(n2292), .A2(n2291), .A3(n2290), .A4(n2289), .ZN(n2301)
         );
  NOR2_X4 U2979 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2342)
         );
  NAND2_X2 U2980 ( .A1(n2293), .A2(n2342), .ZN(n2378) );
  AND2_X1 U2981 ( .A1(n2301), .A2(n2661), .ZN(n2473) );
  NAND2_X1 U2982 ( .A1(n2473), .A2(n2296), .ZN(n2483) );
  NAND2_X1 U2983 ( .A1(n2485), .A2(IR_REG_31__SCAN_IN), .ZN(n2493) );
  NAND2_X1 U2984 ( .A1(n2493), .A2(n2297), .ZN(n2294) );
  NAND2_X1 U2985 ( .A1(n2294), .A2(IR_REG_31__SCAN_IN), .ZN(n2295) );
  XNOR2_X1 U2986 ( .A(n2295), .B(IR_REG_16__SCAN_IN), .ZN(n4444) );
  NAND2_X1 U2987 ( .A1(n2662), .A2(n2306), .ZN(n2307) );
  INV_X1 U2988 ( .A(n2315), .ZN(n2616) );
  NAND2_X1 U2989 ( .A1(n2312), .A2(n2617), .ZN(n2313) );
  MUX2_X1 U2990 ( .A(n4444), .B(DATAI_16_), .S(n2058), .Z(n3365) );
  NAND2_X1 U2991 ( .A1(n3696), .A2(REG0_REG_16__SCAN_IN), .ZN(n2326) );
  NAND2_X1 U2992 ( .A1(n2235), .A2(REG2_REG_16__SCAN_IN), .ZN(n2325) );
  NAND2_X1 U2993 ( .A1(REG3_REG_8__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .ZN(
        n2319) );
  INV_X1 U2994 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2476) );
  INV_X1 U2995 ( .A(REG3_REG_15__SCAN_IN), .ZN(n4452) );
  INV_X1 U2996 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2321) );
  XNOR2_X1 U2997 ( .A(n2500), .B(n2321), .ZN(n3440) );
  OR2_X1 U2998 ( .A1(n2339), .A2(n3440), .ZN(n2324) );
  INV_X1 U2999 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4084) );
  OR2_X1 U3000 ( .A1(n3698), .A2(n4084), .ZN(n2323) );
  INV_X1 U3001 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3099) );
  OR2_X1 U3002 ( .A1(n3099), .A2(n2327), .ZN(n2329) );
  OR2_X1 U3003 ( .A1(n2329), .A2(n2328), .ZN(n2331) );
  INV_X1 U3004 ( .A(n2342), .ZN(n2332) );
  NAND2_X1 U3005 ( .A1(n2333), .A2(n2332), .ZN(n2855) );
  INV_X1 U3006 ( .A(n2855), .ZN(n4451) );
  NAND2_X1 U3007 ( .A1(n2338), .A2(REG0_REG_0__SCAN_IN), .ZN(n2336) );
  INV_X1 U3008 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2917) );
  INV_X1 U3009 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2736) );
  AND2_X1 U3010 ( .A1(n2733), .A2(n3096), .ZN(n3098) );
  NAND2_X1 U3011 ( .A1(n3859), .A2(n2334), .ZN(n2337) );
  NAND2_X1 U3012 ( .A1(n2338), .A2(REG0_REG_2__SCAN_IN), .ZN(n2348) );
  NAND2_X1 U3013 ( .A1(n2235), .A2(REG2_REG_2__SCAN_IN), .ZN(n2347) );
  INV_X1 U3014 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2911) );
  OR2_X1 U3015 ( .A1(n2339), .A2(n2911), .ZN(n2346) );
  OR2_X1 U3016 ( .A1(n3698), .A2(n2844), .ZN(n2345) );
  NOR2_X1 U3017 ( .A1(n2342), .A2(n2617), .ZN(n2340) );
  NAND2_X1 U3018 ( .A1(n2342), .A2(n2341), .ZN(n2354) );
  INV_X1 U3019 ( .A(n2354), .ZN(n2343) );
  MUX2_X1 U3020 ( .A(n4450), .B(DATAI_2_), .S(n2058), .Z(n2936) );
  INV_X1 U3021 ( .A(n2936), .ZN(n2722) );
  NAND2_X1 U3022 ( .A1(n3184), .A2(n2722), .ZN(n2349) );
  AND2_X1 U3023 ( .A1(n4439), .A2(n2322), .ZN(n2597) );
  NAND2_X1 U3024 ( .A1(n2899), .A2(REG1_REG_3__SCAN_IN), .ZN(n2352) );
  NAND2_X1 U3025 ( .A1(n3696), .A2(REG0_REG_3__SCAN_IN), .ZN(n2351) );
  NAND2_X1 U3026 ( .A1(n2235), .A2(REG2_REG_3__SCAN_IN), .ZN(n2350) );
  NAND2_X1 U3027 ( .A1(n2354), .A2(IR_REG_31__SCAN_IN), .ZN(n2355) );
  NAND2_X1 U3028 ( .A1(n2355), .A2(n3960), .ZN(n2368) );
  OR2_X1 U3029 ( .A1(n2355), .A2(n3960), .ZN(n2356) );
  MUX2_X1 U3030 ( .A(n4449), .B(DATAI_3_), .S(n2059), .Z(n3182) );
  NAND2_X1 U3031 ( .A1(n3857), .A2(n3182), .ZN(n2358) );
  NOR2_X1 U3032 ( .A1(n3857), .A2(n3182), .ZN(n2357) );
  NAND2_X1 U3033 ( .A1(n2621), .A2(REG2_REG_4__SCAN_IN), .ZN(n2367) );
  NAND2_X1 U3034 ( .A1(n2338), .A2(REG0_REG_4__SCAN_IN), .ZN(n2366) );
  INV_X1 U3035 ( .A(n2372), .ZN(n2362) );
  INV_X1 U3036 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2360) );
  INV_X1 U3037 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2359) );
  NAND2_X1 U3038 ( .A1(n2360), .A2(n2359), .ZN(n2361) );
  NAND2_X1 U3039 ( .A1(n2362), .A2(n2361), .ZN(n3015) );
  OR2_X1 U3040 ( .A1(n2339), .A2(n3015), .ZN(n2365) );
  INV_X1 U3041 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2363) );
  OR2_X1 U3042 ( .A1(n3698), .A2(n2363), .ZN(n2364) );
  NAND2_X1 U3043 ( .A1(n2368), .A2(IR_REG_31__SCAN_IN), .ZN(n2369) );
  XNOR2_X1 U3044 ( .A(n2369), .B(IR_REG_4__SCAN_IN), .ZN(n4448) );
  MUX2_X1 U3045 ( .A(n4448), .B(DATAI_4_), .S(n2058), .Z(n3007) );
  NAND2_X1 U3046 ( .A1(n3138), .A2(n3007), .ZN(n3780) );
  INV_X1 U3047 ( .A(n3007), .ZN(n3013) );
  NAND2_X1 U3048 ( .A1(n3780), .A2(n3783), .ZN(n3728) );
  NAND2_X1 U3049 ( .A1(n3856), .A2(n3007), .ZN(n2370) );
  NAND2_X1 U3050 ( .A1(n3696), .A2(REG0_REG_5__SCAN_IN), .ZN(n2376) );
  NAND2_X1 U3051 ( .A1(n2235), .A2(REG2_REG_5__SCAN_IN), .ZN(n2375) );
  INV_X1 U3052 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2371) );
  OR2_X1 U3053 ( .A1(n3698), .A2(n2371), .ZN(n2374) );
  OAI21_X1 U3054 ( .B1(n2372), .B2(REG3_REG_5__SCAN_IN), .A(n2385), .ZN(n2987)
         );
  OR2_X1 U3055 ( .A1(n2579), .A2(n2987), .ZN(n2373) );
  NAND2_X1 U3056 ( .A1(n2378), .A2(IR_REG_31__SCAN_IN), .ZN(n2377) );
  MUX2_X1 U3057 ( .A(IR_REG_31__SCAN_IN), .B(n2377), .S(IR_REG_5__SCAN_IN), 
        .Z(n2380) );
  INV_X1 U3058 ( .A(n2401), .ZN(n2379) );
  INV_X1 U3059 ( .A(DATAI_5_), .ZN(n2381) );
  MUX2_X1 U3060 ( .A(n2887), .B(n2381), .S(n2059), .Z(n2991) );
  NAND2_X1 U3061 ( .A1(n2970), .A2(n2991), .ZN(n2382) );
  NAND2_X1 U3062 ( .A1(n3855), .A2(n3141), .ZN(n2383) );
  AND2_X1 U3063 ( .A1(n2385), .A2(n2384), .ZN(n2386) );
  NOR2_X1 U3064 ( .A1(n2394), .A2(n2386), .ZN(n4612) );
  INV_X1 U3065 ( .A(n4612), .ZN(n2387) );
  OR2_X1 U3066 ( .A1(n2339), .A2(n2387), .ZN(n2391) );
  NAND2_X1 U3067 ( .A1(n2899), .A2(REG1_REG_6__SCAN_IN), .ZN(n2390) );
  NAND2_X1 U3068 ( .A1(n2621), .A2(REG2_REG_6__SCAN_IN), .ZN(n2389) );
  NAND2_X1 U3069 ( .A1(n3696), .A2(REG0_REG_6__SCAN_IN), .ZN(n2388) );
  NAND4_X1 U3070 ( .A1(n2391), .A2(n2390), .A3(n2389), .A4(n2388), .ZN(n3854)
         );
  OR2_X1 U3071 ( .A1(n2401), .A2(n2617), .ZN(n2392) );
  XNOR2_X1 U3072 ( .A(n2392), .B(IR_REG_6__SCAN_IN), .ZN(n4446) );
  MUX2_X1 U3073 ( .A(n4446), .B(DATAI_6_), .S(n2058), .Z(n2776) );
  INV_X1 U3074 ( .A(n3854), .ZN(n3069) );
  NAND2_X1 U3075 ( .A1(n3069), .A2(n2978), .ZN(n2393) );
  NAND2_X1 U3076 ( .A1(n2621), .A2(REG2_REG_7__SCAN_IN), .ZN(n2399) );
  NAND2_X1 U3077 ( .A1(n3696), .A2(REG0_REG_7__SCAN_IN), .ZN(n2398) );
  OR2_X1 U3078 ( .A1(n2394), .A2(REG3_REG_7__SCAN_IN), .ZN(n2395) );
  NAND2_X1 U3079 ( .A1(n2413), .A2(n2395), .ZN(n3075) );
  OR2_X1 U3080 ( .A1(n2579), .A2(n3075), .ZN(n2397) );
  INV_X1 U3081 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4070) );
  OR2_X1 U3082 ( .A1(n3698), .A2(n4070), .ZN(n2396) );
  NAND2_X1 U3083 ( .A1(n2401), .A2(n2400), .ZN(n2409) );
  NAND2_X1 U3084 ( .A1(n2409), .A2(IR_REG_31__SCAN_IN), .ZN(n2419) );
  XNOR2_X1 U3085 ( .A(n2419), .B(IR_REG_7__SCAN_IN), .ZN(n4445) );
  MUX2_X1 U3086 ( .A(n4445), .B(DATAI_7_), .S(n2059), .Z(n3066) );
  NAND2_X1 U3087 ( .A1(n3058), .A2(n3066), .ZN(n3786) );
  NAND2_X1 U3088 ( .A1(n3853), .A2(n3073), .ZN(n3788) );
  NAND2_X1 U3089 ( .A1(n2621), .A2(REG2_REG_9__SCAN_IN), .ZN(n2403) );
  NAND2_X1 U3090 ( .A1(n3696), .A2(REG0_REG_9__SCAN_IN), .ZN(n2402) );
  NAND2_X1 U3091 ( .A1(n2403), .A2(n2402), .ZN(n2408) );
  INV_X1 U3092 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2412) );
  INV_X1 U3093 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2404) );
  OAI21_X1 U3094 ( .B1(n2413), .B2(n2412), .A(n2404), .ZN(n2405) );
  NAND2_X1 U3095 ( .A1(n2405), .A2(n2433), .ZN(n3285) );
  INV_X1 U3096 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2406) );
  OAI22_X1 U3097 ( .A1(n2579), .A2(n3285), .B1(n3698), .B2(n2406), .ZN(n2407)
         );
  NAND2_X1 U3098 ( .A1(n2439), .A2(IR_REG_31__SCAN_IN), .ZN(n2410) );
  MUX2_X1 U3099 ( .A(n4651), .B(DATAI_9_), .S(n2059), .Z(n3273) );
  AND2_X1 U3100 ( .A1(n3852), .A2(n3273), .ZN(n2427) );
  NAND2_X1 U3101 ( .A1(n3696), .A2(REG0_REG_8__SCAN_IN), .ZN(n2417) );
  NAND2_X1 U3102 ( .A1(n2621), .A2(REG2_REG_8__SCAN_IN), .ZN(n2416) );
  INV_X1 U3103 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2411) );
  OR2_X1 U3104 ( .A1(n3698), .A2(n2411), .ZN(n2415) );
  XNOR2_X1 U3105 ( .A(n2413), .B(n2412), .ZN(n3127) );
  OR2_X1 U3106 ( .A1(n2339), .A2(n3127), .ZN(n2414) );
  INV_X1 U3107 ( .A(IR_REG_7__SCAN_IN), .ZN(n2418) );
  NAND2_X1 U3108 ( .A1(n2419), .A2(n2418), .ZN(n2420) );
  NAND2_X1 U3109 ( .A1(n2420), .A2(IR_REG_31__SCAN_IN), .ZN(n2422) );
  XNOR2_X1 U3110 ( .A(n2422), .B(n2421), .ZN(n4654) );
  INV_X1 U3111 ( .A(DATAI_8_), .ZN(n4653) );
  MUX2_X1 U3112 ( .A(n4654), .B(n4653), .S(n2058), .Z(n3059) );
  NAND2_X1 U3113 ( .A1(n3275), .A2(n3059), .ZN(n3279) );
  INV_X1 U3114 ( .A(n3852), .ZN(n3060) );
  INV_X1 U3115 ( .A(n3273), .ZN(n3284) );
  NAND2_X1 U3116 ( .A1(n3060), .A2(n3284), .ZN(n2423) );
  AND2_X1 U3117 ( .A1(n3279), .A2(n2423), .ZN(n2424) );
  NOR2_X1 U3118 ( .A1(n2427), .A2(n2424), .ZN(n2430) );
  OR2_X1 U3119 ( .A1(n3727), .A2(n2430), .ZN(n2425) );
  NAND2_X1 U3120 ( .A1(n3853), .A2(n3066), .ZN(n3019) );
  INV_X1 U3121 ( .A(n3275), .ZN(n3067) );
  NAND2_X1 U3122 ( .A1(n3067), .A2(n3025), .ZN(n2426) );
  AND2_X1 U3123 ( .A1(n3019), .A2(n2426), .ZN(n3278) );
  INV_X1 U3124 ( .A(n2427), .ZN(n2428) );
  AND2_X1 U3125 ( .A1(n3278), .A2(n2428), .ZN(n2429) );
  NOR2_X1 U3126 ( .A1(n2430), .A2(n2429), .ZN(n2431) );
  AND2_X1 U3127 ( .A1(n2433), .A2(n3162), .ZN(n2434) );
  OR2_X1 U3128 ( .A1(n2434), .A2(n2459), .ZN(n3173) );
  OR2_X1 U3129 ( .A1(n2579), .A2(n3173), .ZN(n2438) );
  NAND2_X1 U3130 ( .A1(n2899), .A2(REG1_REG_10__SCAN_IN), .ZN(n2437) );
  NAND2_X1 U3131 ( .A1(n3696), .A2(REG0_REG_10__SCAN_IN), .ZN(n2436) );
  NAND2_X1 U3132 ( .A1(n2621), .A2(REG2_REG_10__SCAN_IN), .ZN(n2435) );
  OR2_X1 U3133 ( .A1(n2449), .A2(n2617), .ZN(n2440) );
  XNOR2_X1 U3134 ( .A(n2440), .B(IR_REG_10__SCAN_IN), .ZN(n4098) );
  MUX2_X1 U3135 ( .A(n4098), .B(DATAI_10_), .S(n2059), .Z(n3151) );
  NOR2_X1 U3136 ( .A1(n3851), .A2(n3151), .ZN(n2442) );
  NAND2_X1 U3137 ( .A1(n3851), .A2(n3151), .ZN(n2441) );
  NAND2_X1 U3138 ( .A1(n3696), .A2(REG0_REG_11__SCAN_IN), .ZN(n2447) );
  NAND2_X1 U3139 ( .A1(n2621), .A2(REG2_REG_11__SCAN_IN), .ZN(n2446) );
  INV_X1 U3140 ( .A(REG1_REG_11__SCAN_IN), .ZN(n2443) );
  OR2_X1 U3141 ( .A1(n3698), .A2(n2443), .ZN(n2445) );
  XNOR2_X1 U3142 ( .A(n2459), .B(REG3_REG_11__SCAN_IN), .ZN(n3573) );
  OR2_X1 U3143 ( .A1(n2339), .A2(n3573), .ZN(n2444) );
  INV_X1 U3144 ( .A(IR_REG_10__SCAN_IN), .ZN(n2448) );
  NAND2_X1 U3145 ( .A1(n2449), .A2(n2448), .ZN(n2450) );
  NAND2_X1 U3146 ( .A1(n2450), .A2(IR_REG_31__SCAN_IN), .ZN(n2452) );
  NAND2_X1 U3147 ( .A1(n2452), .A2(n2451), .ZN(n2456) );
  OR2_X1 U31480 ( .A1(n2452), .A2(n2451), .ZN(n2453) );
  MUX2_X1 U31490 ( .A(n4089), .B(DATAI_11_), .S(n2059), .Z(n2454) );
  NAND2_X1 U3150 ( .A1(n3306), .A2(n2454), .ZN(n3216) );
  NAND2_X1 U3151 ( .A1(n3850), .A2(n3571), .ZN(n3803) );
  NAND2_X1 U3152 ( .A1(n3306), .A2(n3571), .ZN(n2455) );
  NAND2_X1 U3153 ( .A1(n2456), .A2(IR_REG_31__SCAN_IN), .ZN(n2457) );
  INV_X1 U3154 ( .A(DATAI_12_), .ZN(n2458) );
  MUX2_X1 U3155 ( .A(n4544), .B(n2458), .S(n2059), .Z(n3304) );
  NAND2_X1 U3156 ( .A1(n2621), .A2(REG2_REG_12__SCAN_IN), .ZN(n2464) );
  NAND2_X1 U3157 ( .A1(n3696), .A2(REG0_REG_12__SCAN_IN), .ZN(n2463) );
  AOI21_X1 U3158 ( .B1(n2459), .B2(REG3_REG_11__SCAN_IN), .A(
        REG3_REG_12__SCAN_IN), .ZN(n2460) );
  OR2_X1 U3159 ( .A1(n2467), .A2(n2460), .ZN(n3311) );
  OR2_X1 U3160 ( .A1(n2579), .A2(n3311), .ZN(n2462) );
  INV_X1 U3161 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4537) );
  OR2_X1 U3162 ( .A1(n3698), .A2(n4537), .ZN(n2461) );
  NAND2_X1 U3163 ( .A1(n2466), .A2(n2465), .ZN(n3244) );
  NAND2_X1 U3164 ( .A1(n2621), .A2(REG2_REG_13__SCAN_IN), .ZN(n2472) );
  NAND2_X1 U3165 ( .A1(n2338), .A2(REG0_REG_13__SCAN_IN), .ZN(n2471) );
  OR2_X1 U3166 ( .A1(n2467), .A2(REG3_REG_13__SCAN_IN), .ZN(n2468) );
  NAND2_X1 U3167 ( .A1(n2477), .A2(n2468), .ZN(n3260) );
  OR2_X1 U3168 ( .A1(n2339), .A2(n3260), .ZN(n2470) );
  INV_X1 U3169 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4078) );
  OR2_X1 U3170 ( .A1(n3698), .A2(n4078), .ZN(n2469) );
  OR2_X1 U3171 ( .A1(n2473), .A2(n2617), .ZN(n2474) );
  XNOR2_X1 U3172 ( .A(n2474), .B(IR_REG_13__SCAN_IN), .ZN(n4643) );
  INV_X1 U3173 ( .A(DATAI_13_), .ZN(n2475) );
  MUX2_X1 U3174 ( .A(n4556), .B(n2475), .S(n2058), .Z(n3340) );
  NAND2_X1 U3175 ( .A1(n3696), .A2(REG0_REG_14__SCAN_IN), .ZN(n2482) );
  NAND2_X1 U3176 ( .A1(n2621), .A2(REG2_REG_14__SCAN_IN), .ZN(n2481) );
  INV_X1 U3177 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4559) );
  OR2_X1 U3178 ( .A1(n3698), .A2(n4559), .ZN(n2480) );
  NAND2_X1 U3179 ( .A1(n2477), .A2(n2476), .ZN(n2478) );
  NAND2_X1 U3180 ( .A1(n2487), .A2(n2478), .ZN(n3394) );
  OR2_X1 U3181 ( .A1(n2339), .A2(n3394), .ZN(n2479) );
  NAND2_X1 U3182 ( .A1(n2483), .A2(IR_REG_31__SCAN_IN), .ZN(n2484) );
  MUX2_X1 U3183 ( .A(IR_REG_31__SCAN_IN), .B(n2484), .S(IR_REG_14__SCAN_IN), 
        .Z(n2486) );
  MUX2_X1 U3184 ( .A(n4565), .B(DATAI_14_), .S(n2058), .Z(n3232) );
  NAND2_X1 U3185 ( .A1(n3385), .A2(n3232), .ZN(n3683) );
  NAND2_X1 U3186 ( .A1(n4455), .A2(n3388), .ZN(n3684) );
  NAND2_X1 U3187 ( .A1(n3683), .A2(n3684), .ZN(n3231) );
  NAND2_X1 U3188 ( .A1(n2338), .A2(REG0_REG_15__SCAN_IN), .ZN(n2492) );
  NAND2_X1 U3189 ( .A1(n2621), .A2(REG2_REG_15__SCAN_IN), .ZN(n2491) );
  NAND2_X1 U3190 ( .A1(n2487), .A2(n4452), .ZN(n2488) );
  NAND2_X1 U3191 ( .A1(n2500), .A2(n2488), .ZN(n4471) );
  OR2_X1 U3192 ( .A1(n2579), .A2(n4471), .ZN(n2490) );
  INV_X1 U3193 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4082) );
  OR2_X1 U3194 ( .A1(n3698), .A2(n4082), .ZN(n2489) );
  XNOR2_X1 U3195 ( .A(n2493), .B(IR_REG_15__SCAN_IN), .ZN(n4106) );
  INV_X1 U3196 ( .A(DATAI_15_), .ZN(n2494) );
  MUX2_X1 U3197 ( .A(n4641), .B(n2494), .S(n2059), .Z(n4459) );
  NAND2_X1 U3198 ( .A1(n3312), .A2(n2496), .ZN(n2497) );
  NAND2_X1 U3199 ( .A1(n3420), .A2(n3365), .ZN(n3811) );
  INV_X1 U3200 ( .A(n3365), .ZN(n3434) );
  NAND2_X1 U3201 ( .A1(n4453), .A2(n3434), .ZN(n3813) );
  INV_X1 U3202 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4118) );
  OR2_X1 U3203 ( .A1(n3698), .A2(n4118), .ZN(n2505) );
  INV_X1 U3204 ( .A(n2500), .ZN(n2498) );
  AOI21_X1 U3205 ( .B1(n2498), .B2(REG3_REG_16__SCAN_IN), .A(
        REG3_REG_17__SCAN_IN), .ZN(n2501) );
  NAND2_X1 U3206 ( .A1(REG3_REG_16__SCAN_IN), .A2(REG3_REG_17__SCAN_IN), .ZN(
        n2499) );
  OR2_X1 U3207 ( .A1(n2501), .A2(n2516), .ZN(n3376) );
  OR2_X1 U3208 ( .A1(n2339), .A2(n3376), .ZN(n2504) );
  NAND2_X1 U3209 ( .A1(n3696), .A2(REG0_REG_17__SCAN_IN), .ZN(n2503) );
  NAND2_X1 U32100 ( .A1(n2235), .A2(REG2_REG_17__SCAN_IN), .ZN(n2502) );
  NAND4_X1 U32110 ( .A1(n2505), .A2(n2504), .A3(n2503), .A4(n2502), .ZN(n3847)
         );
  INV_X1 U32120 ( .A(n3847), .ZN(n3435) );
  NOR2_X1 U32130 ( .A1(n2509), .A2(n2617), .ZN(n2507) );
  MUX2_X1 U32140 ( .A(n2617), .B(n2507), .S(IR_REG_17__SCAN_IN), .Z(n2511) );
  NAND2_X1 U32150 ( .A1(n2509), .A2(n2508), .ZN(n2531) );
  OR2_X1 U32160 ( .A1(n2511), .A2(n2533), .ZN(n4592) );
  INV_X1 U32170 ( .A(DATAI_17_), .ZN(n2512) );
  MUX2_X1 U32180 ( .A(n4592), .B(n2512), .S(n2058), .Z(n3458) );
  INV_X1 U32190 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4114) );
  OR2_X1 U32200 ( .A1(n3698), .A2(n4114), .ZN(n2521) );
  OR2_X1 U32210 ( .A1(n2516), .A2(REG3_REG_18__SCAN_IN), .ZN(n2517) );
  NAND2_X1 U32220 ( .A1(n2527), .A2(n2517), .ZN(n3413) );
  OR2_X1 U32230 ( .A1(n2339), .A2(n3413), .ZN(n2520) );
  NAND2_X1 U32240 ( .A1(n3696), .A2(REG0_REG_18__SCAN_IN), .ZN(n2519) );
  NAND2_X1 U32250 ( .A1(n2235), .A2(REG2_REG_18__SCAN_IN), .ZN(n2518) );
  NAND4_X1 U32260 ( .A1(n2521), .A2(n2520), .A3(n2519), .A4(n2518), .ZN(n4324)
         );
  INV_X1 U32270 ( .A(n4324), .ZN(n3614) );
  NAND2_X1 U32280 ( .A1(n2531), .A2(IR_REG_31__SCAN_IN), .ZN(n2522) );
  XNOR2_X1 U32290 ( .A(n2522), .B(IR_REG_18__SCAN_IN), .ZN(n4128) );
  INV_X1 U32300 ( .A(n4128), .ZN(n4638) );
  INV_X1 U32310 ( .A(DATAI_18_), .ZN(n4637) );
  MUX2_X1 U32320 ( .A(n4638), .B(n4637), .S(n2059), .Z(n3482) );
  INV_X1 U32330 ( .A(n3482), .ZN(n3469) );
  NAND2_X1 U32340 ( .A1(n3614), .A2(n3469), .ZN(n4316) );
  NAND2_X1 U32350 ( .A1(n4324), .A2(n3482), .ZN(n4314) );
  NAND2_X1 U32360 ( .A1(n4316), .A2(n4314), .ZN(n3729) );
  NAND2_X1 U32370 ( .A1(n2235), .A2(REG2_REG_19__SCAN_IN), .ZN(n2525) );
  NAND2_X1 U32380 ( .A1(n3696), .A2(REG0_REG_19__SCAN_IN), .ZN(n2524) );
  NAND2_X1 U32390 ( .A1(n2525), .A2(n2524), .ZN(n2530) );
  INV_X1 U32400 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2526) );
  NAND2_X1 U32410 ( .A1(n2527), .A2(n2526), .ZN(n2528) );
  NAND2_X1 U32420 ( .A1(n2536), .A2(n2528), .ZN(n4332) );
  INV_X1 U32430 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4390) );
  OAI22_X1 U32440 ( .A1(n2339), .A2(n4332), .B1(n3698), .B2(n4390), .ZN(n2529)
         );
  INV_X1 U32450 ( .A(n2531), .ZN(n2533) );
  NAND2_X1 U32460 ( .A1(n2533), .A2(n2532), .ZN(n2603) );
  NAND2_X1 U32470 ( .A1(n2603), .A2(IR_REG_31__SCAN_IN), .ZN(n2608) );
  INV_X1 U32480 ( .A(DATAI_19_), .ZN(n2534) );
  MUX2_X1 U32490 ( .A(n4132), .B(n2534), .S(n2058), .Z(n4330) );
  INV_X1 U32500 ( .A(n4330), .ZN(n3490) );
  NAND2_X1 U32510 ( .A1(n4300), .A2(n3490), .ZN(n2535) );
  INV_X1 U32520 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4047) );
  AND2_X1 U32530 ( .A1(n2536), .A2(n4047), .ZN(n2537) );
  OR2_X1 U32540 ( .A1(n2537), .A2(n2543), .ZN(n4307) );
  NAND2_X1 U32550 ( .A1(n2621), .A2(REG2_REG_20__SCAN_IN), .ZN(n2539) );
  NAND2_X1 U32560 ( .A1(n3696), .A2(REG0_REG_20__SCAN_IN), .ZN(n2538) );
  AND2_X1 U32570 ( .A1(n2539), .A2(n2538), .ZN(n2541) );
  NAND2_X1 U32580 ( .A1(n2899), .A2(REG1_REG_20__SCAN_IN), .ZN(n2540) );
  NAND2_X1 U32590 ( .A1(n4322), .A2(n4305), .ZN(n2542) );
  NOR2_X1 U32600 ( .A1(n2543), .A2(REG3_REG_21__SCAN_IN), .ZN(n2544) );
  OR2_X1 U32610 ( .A1(n2548), .A2(n2544), .ZN(n4285) );
  AOI22_X1 U32620 ( .A1(n2235), .A2(REG2_REG_21__SCAN_IN), .B1(n3696), .B2(
        REG0_REG_21__SCAN_IN), .ZN(n2546) );
  INV_X1 U32630 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4382) );
  OR2_X1 U32640 ( .A1(n3698), .A2(n4382), .ZN(n2545) );
  NAND2_X1 U32650 ( .A1(n2058), .A2(DATAI_21_), .ZN(n4283) );
  INV_X1 U32660 ( .A(n4283), .ZN(n2704) );
  NAND2_X1 U32670 ( .A1(n4299), .A2(n2704), .ZN(n2547) );
  INV_X1 U32680 ( .A(n4299), .ZN(n4256) );
  OR2_X1 U32690 ( .A1(n2548), .A2(REG3_REG_22__SCAN_IN), .ZN(n2549) );
  NAND2_X1 U32700 ( .A1(n2552), .A2(n2549), .ZN(n4264) );
  AOI22_X1 U32710 ( .A1(n2899), .A2(REG1_REG_22__SCAN_IN), .B1(n3696), .B2(
        REG0_REG_22__SCAN_IN), .ZN(n2551) );
  NAND2_X1 U32720 ( .A1(n2621), .A2(REG2_REG_22__SCAN_IN), .ZN(n2550) );
  OAI211_X1 U32730 ( .C1(n4264), .C2(n2579), .A(n2551), .B(n2550), .ZN(n4279)
         );
  NAND2_X1 U32740 ( .A1(n2058), .A2(DATAI_22_), .ZN(n4267) );
  OR2_X1 U32750 ( .A1(n4279), .A2(n4267), .ZN(n2646) );
  NAND2_X1 U32760 ( .A1(n4279), .A2(n4267), .ZN(n2648) );
  NAND2_X1 U32770 ( .A1(n2646), .A2(n2648), .ZN(n4258) );
  NAND2_X1 U32780 ( .A1(n4255), .A2(n4258), .ZN(n4254) );
  INV_X1 U32790 ( .A(n4279), .ZN(n4240) );
  NAND2_X1 U32800 ( .A1(n4254), .A2(n2284), .ZN(n4231) );
  INV_X1 U32810 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3605) );
  NAND2_X1 U32820 ( .A1(n2552), .A2(n3605), .ZN(n2553) );
  NAND2_X1 U32830 ( .A1(n2561), .A2(n2553), .ZN(n4248) );
  OR2_X1 U32840 ( .A1(n4248), .A2(n2579), .ZN(n2558) );
  INV_X1 U32850 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4373) );
  NAND2_X1 U32860 ( .A1(n3696), .A2(REG0_REG_23__SCAN_IN), .ZN(n2555) );
  NAND2_X1 U32870 ( .A1(n2621), .A2(REG2_REG_23__SCAN_IN), .ZN(n2554) );
  OAI211_X1 U32880 ( .C1(n3698), .C2(n4373), .A(n2555), .B(n2554), .ZN(n2556)
         );
  INV_X1 U32890 ( .A(n2556), .ZN(n2557) );
  INV_X1 U32900 ( .A(n4218), .ZN(n4263) );
  AND2_X1 U32910 ( .A1(n2058), .A2(DATAI_23_), .ZN(n3604) );
  NAND2_X1 U32920 ( .A1(n4231), .A2(n2287), .ZN(n2560) );
  INV_X1 U32930 ( .A(n3604), .ZN(n4246) );
  INV_X1 U32940 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3646) );
  AND2_X1 U32950 ( .A1(n2561), .A2(n3646), .ZN(n2562) );
  OR2_X1 U32960 ( .A1(n2562), .A2(n2567), .ZN(n4225) );
  INV_X1 U32970 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4369) );
  NAND2_X1 U32980 ( .A1(n2235), .A2(REG2_REG_24__SCAN_IN), .ZN(n2564) );
  NAND2_X1 U32990 ( .A1(n3696), .A2(REG0_REG_24__SCAN_IN), .ZN(n2563) );
  OAI211_X1 U33000 ( .C1(n4369), .C2(n3698), .A(n2564), .B(n2563), .ZN(n2565)
         );
  INV_X1 U33010 ( .A(n2565), .ZN(n2566) );
  OAI21_X1 U33020 ( .B1(n4225), .B2(n2579), .A(n2566), .ZN(n4242) );
  INV_X1 U33030 ( .A(n4242), .ZN(n4202) );
  NAND2_X1 U33040 ( .A1(n2059), .A2(DATAI_24_), .ZN(n4224) );
  NOR2_X1 U33050 ( .A1(n4202), .A2(n4224), .ZN(n4197) );
  NOR2_X1 U33060 ( .A1(n2567), .A2(REG3_REG_25__SCAN_IN), .ZN(n2568) );
  OR2_X1 U33070 ( .A1(n2577), .A2(n2568), .ZN(n3634) );
  INV_X1 U33080 ( .A(REG1_REG_25__SCAN_IN), .ZN(n2571) );
  NAND2_X1 U33090 ( .A1(n2338), .A2(REG0_REG_25__SCAN_IN), .ZN(n2570) );
  NAND2_X1 U33100 ( .A1(n2621), .A2(REG2_REG_25__SCAN_IN), .ZN(n2569) );
  OAI211_X1 U33110 ( .C1(n3698), .C2(n2571), .A(n2570), .B(n2569), .ZN(n2572)
         );
  INV_X1 U33120 ( .A(n2572), .ZN(n2573) );
  AND2_X1 U33130 ( .A1(n2059), .A2(DATAI_25_), .ZN(n4208) );
  NOR2_X1 U33140 ( .A1(n4220), .A2(n4208), .ZN(n2576) );
  INV_X1 U33150 ( .A(n4224), .ZN(n4196) );
  NOR2_X1 U33160 ( .A1(n4242), .A2(n4196), .ZN(n2575) );
  OR2_X1 U33170 ( .A1(n2577), .A2(REG3_REG_26__SCAN_IN), .ZN(n2578) );
  NAND2_X1 U33180 ( .A1(n2585), .A2(n2578), .ZN(n3674) );
  INV_X1 U33190 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4361) );
  NAND2_X1 U33200 ( .A1(n3696), .A2(REG0_REG_26__SCAN_IN), .ZN(n2581) );
  NAND2_X1 U33210 ( .A1(n2621), .A2(REG2_REG_26__SCAN_IN), .ZN(n2580) );
  OAI211_X1 U33220 ( .C1(n3698), .C2(n4361), .A(n2581), .B(n2580), .ZN(n2582)
         );
  INV_X1 U33230 ( .A(n2582), .ZN(n2583) );
  NAND2_X1 U33240 ( .A1(n2058), .A2(DATAI_26_), .ZN(n4189) );
  INV_X1 U33250 ( .A(n4189), .ZN(n2653) );
  NAND2_X1 U33260 ( .A1(n4162), .A2(n4189), .ZN(n3762) );
  INV_X1 U33270 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3592) );
  NAND2_X1 U33280 ( .A1(n2585), .A2(n3592), .ZN(n2586) );
  NAND2_X1 U33290 ( .A1(n2595), .A2(n2586), .ZN(n3591) );
  INV_X1 U33300 ( .A(REG1_REG_27__SCAN_IN), .ZN(n2589) );
  NAND2_X1 U33310 ( .A1(n2235), .A2(REG2_REG_27__SCAN_IN), .ZN(n2588) );
  NAND2_X1 U33320 ( .A1(n3696), .A2(REG0_REG_27__SCAN_IN), .ZN(n2587) );
  OAI211_X1 U33330 ( .C1(n3698), .C2(n2589), .A(n2588), .B(n2587), .ZN(n2590)
         );
  INV_X1 U33340 ( .A(n2590), .ZN(n2591) );
  AND2_X1 U33350 ( .A1(n2058), .A2(DATAI_27_), .ZN(n3822) );
  NOR2_X1 U33360 ( .A1(n4184), .A2(n3822), .ZN(n2594) );
  NAND2_X1 U33370 ( .A1(n4184), .A2(n3822), .ZN(n2593) );
  INV_X1 U33380 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3553) );
  NAND2_X1 U33390 ( .A1(n2595), .A2(n3553), .ZN(n2596) );
  NAND2_X1 U33400 ( .A1(n3582), .A2(n2597), .ZN(n2602) );
  INV_X1 U33410 ( .A(REG1_REG_28__SCAN_IN), .ZN(n3906) );
  NAND2_X1 U33420 ( .A1(n3696), .A2(REG0_REG_28__SCAN_IN), .ZN(n2599) );
  NAND2_X1 U33430 ( .A1(n2621), .A2(REG2_REG_28__SCAN_IN), .ZN(n2598) );
  OAI211_X1 U33440 ( .C1(n3698), .C2(n3906), .A(n2599), .B(n2598), .ZN(n2600)
         );
  INV_X1 U33450 ( .A(n2600), .ZN(n2601) );
  NAND2_X1 U33460 ( .A1(n2059), .A2(DATAI_28_), .ZN(n3552) );
  NOR2_X1 U33470 ( .A1(n4169), .A2(n3552), .ZN(n4149) );
  XNOR2_X1 U33480 ( .A(n4139), .B(n4138), .ZN(n3588) );
  INV_X1 U33490 ( .A(n2603), .ZN(n2604) );
  NAND2_X1 U33500 ( .A1(n2604), .A2(n2279), .ZN(n2612) );
  NOR2_X2 U33510 ( .A1(n2612), .A2(IR_REG_21__SCAN_IN), .ZN(n2669) );
  INV_X1 U33520 ( .A(n2669), .ZN(n2605) );
  INV_X1 U3353 ( .A(n2719), .ZN(n4442) );
  NAND2_X1 U33540 ( .A1(n2608), .A2(n2607), .ZN(n2609) );
  NAND2_X1 U3355 ( .A1(n2612), .A2(IR_REG_31__SCAN_IN), .ZN(n2614) );
  XNOR2_X1 U3356 ( .A(n4442), .B(n2717), .ZN(n2615) );
  NAND2_X1 U3357 ( .A1(n2615), .A2(n4132), .ZN(n3565) );
  AND2_X1 U3358 ( .A1(n3834), .A2(n4443), .ZN(n3046) );
  INV_X1 U3359 ( .A(n4675), .ZN(n4699) );
  NAND2_X1 U3360 ( .A1(n3565), .A2(n4699), .ZN(n4694) );
  INV_X1 U3361 ( .A(n4694), .ZN(n4678) );
  NOR2_X1 U3362 ( .A1(n2315), .A2(n2617), .ZN(n2618) );
  MUX2_X1 U3363 ( .A(n2617), .B(n2618), .S(IR_REG_28__SCAN_IN), .Z(n2619) );
  INV_X1 U3364 ( .A(n2619), .ZN(n2620) );
  NAND2_X1 U3365 ( .A1(n2620), .A2(n2816), .ZN(n3871) );
  INV_X1 U3366 ( .A(n3871), .ZN(n4440) );
  NAND2_X1 U3367 ( .A1(n4442), .A2(n3771), .ZN(n2787) );
  INV_X1 U3368 ( .A(n2787), .ZN(n2836) );
  INV_X1 U3369 ( .A(REG1_REG_29__SCAN_IN), .ZN(n3905) );
  NAND2_X1 U3370 ( .A1(n2621), .A2(REG2_REG_29__SCAN_IN), .ZN(n2623) );
  NAND2_X1 U3371 ( .A1(n3696), .A2(REG0_REG_29__SCAN_IN), .ZN(n2622) );
  OAI211_X1 U3372 ( .C1(n3905), .C2(n3698), .A(n2623), .B(n2622), .ZN(n2624)
         );
  INV_X1 U3373 ( .A(n2624), .ZN(n2625) );
  OAI21_X1 U3374 ( .B1(n4156), .B2(n2579), .A(n2625), .ZN(n3844) );
  INV_X1 U3375 ( .A(n3844), .ZN(n3554) );
  NAND2_X1 U3376 ( .A1(n3871), .A2(n2836), .ZN(n4321) );
  OAI22_X1 U3377 ( .A1(n3554), .A2(n4321), .B1(n3552), .B2(n4320), .ZN(n2660)
         );
  NAND2_X1 U3378 ( .A1(n2928), .A2(n3774), .ZN(n3181) );
  INV_X1 U3379 ( .A(n3857), .ZN(n2933) );
  NAND2_X1 U3380 ( .A1(n2933), .A2(n3182), .ZN(n3779) );
  NAND2_X1 U3381 ( .A1(n3857), .A2(n2754), .ZN(n3776) );
  AND2_X1 U3382 ( .A1(n3779), .A2(n3776), .ZN(n3733) );
  NAND2_X1 U3383 ( .A1(n3181), .A2(n3733), .ZN(n2630) );
  NAND2_X1 U3384 ( .A1(n2630), .A2(n3779), .ZN(n3006) );
  INV_X1 U3385 ( .A(n3780), .ZN(n2631) );
  NAND2_X1 U3386 ( .A1(n2970), .A2(n3141), .ZN(n3793) );
  NAND2_X1 U3387 ( .A1(n3855), .A2(n2991), .ZN(n3782) );
  AND2_X1 U3388 ( .A1(n3854), .A2(n2978), .ZN(n2968) );
  NAND2_X1 U3389 ( .A1(n3069), .A2(n2776), .ZN(n3785) );
  NAND2_X1 U3390 ( .A1(n2632), .A2(n3785), .ZN(n3065) );
  INV_X1 U3391 ( .A(n3786), .ZN(n2633) );
  NAND2_X1 U3392 ( .A1(n3275), .A2(n3025), .ZN(n3790) );
  NAND2_X1 U3393 ( .A1(n3852), .A2(n3284), .ZN(n3794) );
  NAND2_X1 U3394 ( .A1(n3060), .A2(n3273), .ZN(n3789) );
  NAND2_X1 U3395 ( .A1(n2634), .A2(n3789), .ZN(n3085) );
  INV_X1 U3396 ( .A(n3151), .ZN(n3165) );
  NAND2_X1 U3397 ( .A1(n3851), .A2(n3165), .ZN(n3802) );
  NAND2_X1 U3398 ( .A1(n3085), .A2(n3802), .ZN(n2636) );
  INV_X1 U3399 ( .A(n3851), .ZN(n2635) );
  NAND2_X1 U3400 ( .A1(n2635), .A2(n3151), .ZN(n3796) );
  NAND2_X1 U3401 ( .A1(n2636), .A2(n3796), .ZN(n3563) );
  NAND2_X1 U3402 ( .A1(n3337), .A2(n3304), .ZN(n3246) );
  NAND2_X1 U3403 ( .A1(n3849), .A2(n3340), .ZN(n2637) );
  NAND2_X1 U3404 ( .A1(n3246), .A2(n2637), .ZN(n2638) );
  INV_X1 U3405 ( .A(n2638), .ZN(n3804) );
  NAND2_X1 U3406 ( .A1(n3564), .A2(n3219), .ZN(n3245) );
  NAND2_X1 U3407 ( .A1(n3216), .A2(n3245), .ZN(n2640) );
  NOR2_X1 U3408 ( .A1(n3849), .A2(n3340), .ZN(n2639) );
  AOI21_X1 U3409 ( .B1(n3804), .B2(n2640), .A(n2639), .ZN(n3805) );
  INV_X1 U3410 ( .A(n3231), .ZN(n3754) );
  NAND2_X1 U3411 ( .A1(n3433), .A2(n2495), .ZN(n3686) );
  NAND2_X1 U3412 ( .A1(n3848), .A2(n4459), .ZN(n3685) );
  NAND2_X1 U3413 ( .A1(n3686), .A2(n3685), .ZN(n3752) );
  INV_X1 U3414 ( .A(n3683), .ZN(n2641) );
  NOR2_X1 U3415 ( .A1(n3752), .A2(n2641), .ZN(n2642) );
  NAND2_X1 U3416 ( .A1(n3313), .A2(n2642), .ZN(n2643) );
  NAND2_X1 U3417 ( .A1(n4300), .A2(n4330), .ZN(n3719) );
  AND2_X1 U3418 ( .A1(n3719), .A2(n4314), .ZN(n4232) );
  NAND2_X1 U3419 ( .A1(n3847), .A2(n3458), .ZN(n3404) );
  NAND2_X1 U3420 ( .A1(n3846), .A2(n4305), .ZN(n4235) );
  NAND3_X1 U3421 ( .A1(n4232), .A2(n3404), .A3(n4235), .ZN(n3816) );
  NAND2_X1 U3422 ( .A1(n3435), .A2(n3452), .ZN(n3407) );
  NAND2_X1 U3423 ( .A1(n3407), .A2(n4316), .ZN(n2644) );
  NOR2_X1 U3424 ( .A1(n4300), .A2(n4330), .ZN(n3720) );
  AOI21_X1 U3425 ( .B1(n4232), .B2(n2644), .A(n3720), .ZN(n4292) );
  OAI21_X1 U3426 ( .B1(n4305), .B2(n3846), .A(n4292), .ZN(n2645) );
  NAND2_X1 U3427 ( .A1(n2645), .A2(n4235), .ZN(n3815) );
  INV_X1 U3428 ( .A(n3815), .ZN(n4234) );
  OR2_X1 U3429 ( .A1(n4299), .A2(n4283), .ZN(n3716) );
  INV_X1 U3430 ( .A(n3716), .ZN(n4236) );
  NOR2_X1 U3431 ( .A1(n4234), .A2(n4236), .ZN(n3690) );
  NAND2_X1 U3432 ( .A1(n4299), .A2(n4283), .ZN(n3821) );
  INV_X1 U3433 ( .A(n2646), .ZN(n4237) );
  AOI21_X1 U3434 ( .B1(n2647), .B2(n3821), .A(n4237), .ZN(n2651) );
  NOR2_X1 U3435 ( .A1(n4218), .A2(n3604), .ZN(n3718) );
  INV_X1 U3436 ( .A(n2648), .ZN(n2649) );
  NOR2_X1 U3437 ( .A1(n3718), .A2(n2649), .ZN(n3695) );
  INV_X1 U3438 ( .A(n3695), .ZN(n2650) );
  OR2_X1 U3439 ( .A1(n4242), .A2(n4224), .ZN(n2652) );
  NAND2_X1 U3440 ( .A1(n4218), .A2(n3604), .ZN(n3717) );
  NAND2_X1 U3441 ( .A1(n2652), .A2(n3717), .ZN(n3818) );
  NAND2_X1 U3442 ( .A1(n4242), .A2(n4224), .ZN(n3693) );
  INV_X1 U3443 ( .A(n4208), .ZN(n4201) );
  NAND2_X1 U3444 ( .A1(n4220), .A2(n4201), .ZN(n3694) );
  INV_X1 U3445 ( .A(n3694), .ZN(n3726) );
  NAND2_X1 U3446 ( .A1(n4162), .A2(n2653), .ZN(n2654) );
  NAND2_X1 U3447 ( .A1(n4182), .A2(n4208), .ZN(n3725) );
  INV_X1 U3448 ( .A(n3826), .ZN(n3703) );
  AND2_X1 U3449 ( .A1(n4204), .A2(n4189), .ZN(n3707) );
  INV_X1 U3450 ( .A(n3707), .ZN(n2655) );
  XNOR2_X1 U3451 ( .A(n4184), .B(n3822), .ZN(n3741) );
  NOR2_X1 U3452 ( .A1(n4164), .A2(n4165), .ZN(n4163) );
  INV_X1 U3453 ( .A(n3822), .ZN(n4171) );
  NOR2_X1 U3454 ( .A1(n4184), .A2(n4171), .ZN(n3708) );
  NOR2_X1 U3455 ( .A1(n4163), .A2(n3708), .ZN(n4152) );
  XOR2_X1 U3456 ( .A(n4138), .B(n4152), .Z(n2658) );
  NAND2_X1 U3457 ( .A1(n4442), .A2(n4443), .ZN(n2657) );
  INV_X1 U34580 ( .A(n3834), .ZN(n2820) );
  NAND2_X1 U34590 ( .A1(n2820), .A2(n3771), .ZN(n2656) );
  NOR2_X1 U3460 ( .A1(n2658), .A2(n4327), .ZN(n2659) );
  AOI211_X1 U3461 ( .C1(n4325), .C2(n4184), .A(n2660), .B(n2659), .ZN(n3581)
         );
  OAI21_X1 U3462 ( .B1(n3588), .B2(n4678), .A(n3581), .ZN(n2710) );
  AND2_X1 U3463 ( .A1(n2662), .A2(n2661), .ZN(n2666) );
  NAND2_X1 U3464 ( .A1(n2506), .A2(n2666), .ZN(n2663) );
  NAND2_X1 U3465 ( .A1(n2663), .A2(IR_REG_31__SCAN_IN), .ZN(n2664) );
  MUX2_X1 U3466 ( .A(IR_REG_31__SCAN_IN), .B(n2664), .S(IR_REG_25__SCAN_IN), 
        .Z(n2667) );
  NAND2_X1 U34670 ( .A1(n2666), .A2(n2665), .ZN(n2674) );
  NAND2_X1 U3468 ( .A1(n2667), .A2(n2674), .ZN(n2815) );
  NAND2_X1 U34690 ( .A1(n2815), .A2(B_REG_SCAN_IN), .ZN(n2673) );
  NAND2_X1 U3470 ( .A1(n2669), .A2(n2668), .ZN(n2670) );
  INV_X1 U34710 ( .A(IR_REG_23__SCAN_IN), .ZN(n2682) );
  NAND2_X1 U3472 ( .A1(n2681), .A2(n2682), .ZN(n2671) );
  XNOR2_X2 U34730 ( .A(n2672), .B(IR_REG_24__SCAN_IN), .ZN(n2680) );
  MUX2_X1 U3474 ( .A(n2673), .B(B_REG_SCAN_IN), .S(n2680), .Z(n2678) );
  NAND2_X1 U34750 ( .A1(n2674), .A2(IR_REG_31__SCAN_IN), .ZN(n2675) );
  MUX2_X1 U3476 ( .A(IR_REG_31__SCAN_IN), .B(n2675), .S(IR_REG_26__SCAN_IN), 
        .Z(n2677) );
  NAND2_X1 U34770 ( .A1(n2677), .A2(n2676), .ZN(n2698) );
  INV_X1 U3478 ( .A(n2698), .ZN(n4441) );
  NAND2_X1 U34790 ( .A1(n2698), .A2(n2815), .ZN(n2827) );
  NAND2_X1 U3480 ( .A1(n3001), .A2(n2827), .ZN(n2697) );
  NOR2_X1 U34810 ( .A1(n2698), .A2(n2815), .ZN(n2679) );
  XNOR2_X1 U3482 ( .A(n2681), .B(n2682), .ZN(n2835) );
  NAND2_X1 U34830 ( .A1(n2835), .A2(STATE_REG_SCAN_IN), .ZN(n4635) );
  INV_X1 U3484 ( .A(n4635), .ZN(n2828) );
  NAND2_X1 U34850 ( .A1(n2718), .A2(n2828), .ZN(n3000) );
  NAND2_X1 U3486 ( .A1(n4675), .A2(n2627), .ZN(n2805) );
  AND2_X1 U34870 ( .A1(n3834), .A2(n4132), .ZN(n2683) );
  OR2_X1 U3488 ( .A1(n2787), .A2(n2683), .ZN(n2998) );
  NAND2_X1 U34890 ( .A1(n2805), .A2(n2998), .ZN(n2684) );
  NOR2_X1 U3490 ( .A1(n3000), .A2(n2684), .ZN(n2696) );
  NOR4_X1 U34910 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_15__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2688) );
  NOR4_X1 U3492 ( .A1(D_REG_9__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2687) );
  NOR4_X1 U34930 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2686) );
  NOR4_X1 U3494 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2685) );
  NAND4_X1 U34950 ( .A1(n2688), .A2(n2687), .A3(n2686), .A4(n2685), .ZN(n2694)
         );
  NOR2_X1 U3496 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_20__SCAN_IN), .ZN(n2692)
         );
  NOR4_X1 U34970 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2691) );
  NOR4_X1 U3498 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_5__SCAN_IN), .A3(
        D_REG_7__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2690) );
  NOR4_X1 U34990 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_2__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2689) );
  NAND4_X1 U3500 ( .A1(n2692), .A2(n2691), .A3(n2690), .A4(n2689), .ZN(n2693)
         );
  NOR2_X1 U35010 ( .A1(n2694), .A2(n2693), .ZN(n2695) );
  INV_X1 U3502 ( .A(n2680), .ZN(n2699) );
  NAND2_X1 U35030 ( .A1(n2699), .A2(n2698), .ZN(n2700) );
  AND2_X2 U3504 ( .A1(n2709), .A2(n3004), .ZN(n4705) );
  INV_X1 U35050 ( .A(REG0_REG_28__SCAN_IN), .ZN(n2702) );
  NAND2_X1 U35060 ( .A1(n3188), .A2(n2754), .ZN(n3190) );
  INV_X1 U35070 ( .A(n4305), .ZN(n3722) );
  INV_X1 U35080 ( .A(n4170), .ZN(n2706) );
  INV_X1 U35090 ( .A(n3552), .ZN(n4137) );
  INV_X1 U35100 ( .A(n4142), .ZN(n2705) );
  OAI21_X1 U35110 ( .B1(n2706), .B2(n3552), .A(n2705), .ZN(n3584) );
  NAND2_X1 U35120 ( .A1(n2708), .A2(n2285), .ZN(U3514) );
  AND2_X2 U35130 ( .A1(n2709), .A2(n2786), .ZN(n4716) );
  NAND2_X1 U35140 ( .A1(n4716), .A2(n2707), .ZN(n4392) );
  NOR2_X1 U35150 ( .A1(n3584), .A2(n4392), .ZN(n2713) );
  OR2_X1 U35160 ( .A1(n2718), .A2(n4635), .ZN(n2715) );
  INV_X2 U35170 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X2 U35180 ( .A(n2742), .ZN(n2772) );
  OAI22_X1 U35190 ( .A1(n3058), .A2(n3540), .B1(n2056), .B2(n3073), .ZN(n2720)
         );
  XNOR2_X1 U35200 ( .A(n2720), .B(n3546), .ZN(n3052) );
  OAI22_X1 U35210 ( .A1(n3058), .A2(n3525), .B1(n3540), .B2(n3073), .ZN(n3051)
         );
  XNOR2_X1 U35220 ( .A(n3052), .B(n3051), .ZN(n2792) );
  OAI22_X1 U35230 ( .A1(n3184), .A2(n2742), .B1(n2741), .B2(n2722), .ZN(n2721)
         );
  XNOR2_X1 U35240 ( .A(n2721), .B(n3538), .ZN(n2724) );
  INV_X1 U35250 ( .A(n2746), .ZN(n3473) );
  NOR2_X1 U35260 ( .A1(n2722), .A2(n2742), .ZN(n2723) );
  NAND2_X1 U35270 ( .A1(n2724), .A2(n2725), .ZN(n2751) );
  INV_X1 U35280 ( .A(n2724), .ZN(n2727) );
  INV_X1 U35290 ( .A(n2725), .ZN(n2726) );
  NAND2_X1 U35300 ( .A1(n2727), .A2(n2726), .ZN(n2728) );
  AND2_X1 U35310 ( .A1(n2751), .A2(n2728), .ZN(n2905) );
  INV_X1 U35320 ( .A(n2733), .ZN(n2729) );
  INV_X1 U35330 ( .A(n2718), .ZN(n2730) );
  AOI22_X1 U35340 ( .A1(n2772), .A2(n3096), .B1(n2730), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2731) );
  NAND2_X1 U35350 ( .A1(n2732), .A2(n2731), .ZN(n2912) );
  NAND2_X1 U35360 ( .A1(n2733), .A2(n2772), .ZN(n2735) );
  AND2_X1 U35370 ( .A1(n2735), .A2(n2734), .ZN(n2738) );
  OR2_X1 U35380 ( .A1(n2718), .A2(n2736), .ZN(n2737) );
  NAND2_X1 U35390 ( .A1(n2738), .A2(n2737), .ZN(n2914) );
  NAND2_X1 U35400 ( .A1(n2912), .A2(n2914), .ZN(n2740) );
  NAND2_X1 U35410 ( .A1(n2738), .A2(n3538), .ZN(n2739) );
  NAND2_X1 U35420 ( .A1(n2740), .A2(n2739), .ZN(n2918) );
  OAI22_X1 U35430 ( .A1(n2746), .A2(n2744), .B1(n2742), .B2(n2745), .ZN(n2747)
         );
  XNOR2_X1 U35440 ( .A(n2749), .B(n2747), .ZN(n2919) );
  INV_X1 U35450 ( .A(n2747), .ZN(n2748) );
  NAND2_X1 U35460 ( .A1(n2905), .A2(n2906), .ZN(n2904) );
  NAND2_X1 U35470 ( .A1(n2904), .A2(n2751), .ZN(n3033) );
  INV_X2 U35480 ( .A(n2746), .ZN(n3545) );
  NAND2_X1 U35490 ( .A1(n3857), .A2(n3545), .ZN(n2753) );
  NAND2_X1 U35500 ( .A1(n3534), .A2(n3182), .ZN(n2752) );
  NAND2_X1 U35510 ( .A1(n2753), .A2(n2752), .ZN(n2759) );
  NAND2_X1 U35520 ( .A1(n3857), .A2(n3534), .ZN(n2756) );
  INV_X1 U35530 ( .A(n3182), .ZN(n2754) );
  NAND2_X1 U35540 ( .A1(n2756), .A2(n2755), .ZN(n2757) );
  XNOR2_X1 U35550 ( .A(n2759), .B(n2761), .ZN(n3034) );
  NAND2_X1 U35560 ( .A1(n3033), .A2(n3034), .ZN(n2956) );
  XNOR2_X1 U35570 ( .A(n2758), .B(n3538), .ZN(n2763) );
  OAI22_X1 U35580 ( .A1(n3138), .A2(n2746), .B1(n2742), .B2(n3013), .ZN(n2764)
         );
  INV_X1 U35590 ( .A(n2759), .ZN(n2760) );
  NAND2_X1 U35600 ( .A1(n2761), .A2(n2760), .ZN(n2959) );
  INV_X1 U35610 ( .A(n2763), .ZN(n2765) );
  NAND2_X1 U35620 ( .A1(n2765), .A2(n2764), .ZN(n2766) );
  OAI22_X1 U35630 ( .A1(n2970), .A2(n2742), .B1(n2056), .B2(n2991), .ZN(n2767)
         );
  XNOR2_X1 U35640 ( .A(n2767), .B(n3538), .ZN(n2768) );
  INV_X1 U35650 ( .A(n2768), .ZN(n2770) );
  NAND2_X1 U35660 ( .A1(n2770), .A2(n2769), .ZN(n2771) );
  INV_X1 U35670 ( .A(n2944), .ZN(n2780) );
  NAND2_X1 U35680 ( .A1(n3854), .A2(n3534), .ZN(n2774) );
  INV_X2 U35690 ( .A(n2741), .ZN(n3544) );
  NAND2_X1 U35700 ( .A1(n3544), .A2(n2776), .ZN(n2773) );
  NAND2_X1 U35710 ( .A1(n2774), .A2(n2773), .ZN(n2775) );
  XNOR2_X1 U35720 ( .A(n2775), .B(n3546), .ZN(n2781) );
  NAND2_X1 U35730 ( .A1(n3854), .A2(n3545), .ZN(n2778) );
  NAND2_X1 U35740 ( .A1(n3534), .A2(n2776), .ZN(n2777) );
  NAND2_X1 U35750 ( .A1(n2778), .A2(n2777), .ZN(n2782) );
  AND2_X1 U35760 ( .A1(n2781), .A2(n2782), .ZN(n2946) );
  INV_X1 U35770 ( .A(n2946), .ZN(n2779) );
  INV_X1 U35780 ( .A(n2781), .ZN(n2784) );
  INV_X1 U35790 ( .A(n2782), .ZN(n2783) );
  NAND2_X1 U35800 ( .A1(n2784), .A2(n2783), .ZN(n2945) );
  NAND3_X1 U35810 ( .A1(n3003), .A2(n2786), .A3(n3001), .ZN(n2809) );
  INV_X1 U3582 ( .A(n2809), .ZN(n2804) );
  OAI211_X1 U3583 ( .C1(n3042), .C2(n4132), .A(n4320), .B(n2787), .ZN(n2793)
         );
  NOR2_X1 U3584 ( .A1(n3000), .A2(n2793), .ZN(n2788) );
  INV_X1 U3585 ( .A(n3054), .ZN(n2791) );
  AOI211_X1 U3586 ( .C1(n2792), .C2(n2789), .A(n4465), .B(n2791), .ZN(n2813)
         );
  NAND2_X1 U3587 ( .A1(n2793), .A2(n4320), .ZN(n2794) );
  NAND2_X1 U3588 ( .A1(n2809), .A2(n2794), .ZN(n2795) );
  NAND2_X1 U3589 ( .A1(n2795), .A2(n2998), .ZN(n2902) );
  NAND2_X1 U3590 ( .A1(n2718), .A2(n2835), .ZN(n2796) );
  OAI21_X1 U3591 ( .B1(n2902), .B2(n2796), .A(STATE_REG_SCAN_IN), .ZN(n2799)
         );
  OR3_X1 U3592 ( .A1(n3540), .A2(n2798), .A3(n4635), .ZN(n3838) );
  NAND2_X1 U3593 ( .A1(n2809), .A2(n2807), .ZN(n2901) );
  NOR2_X1 U3594 ( .A1(n4472), .A2(n3075), .ZN(n2812) );
  NAND2_X1 U3595 ( .A1(n2807), .A2(n4440), .ZN(n2800) );
  INV_X1 U3596 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2801) );
  NOR2_X1 U3597 ( .A1(STATE_REG_SCAN_IN), .A2(n2801), .ZN(n2868) );
  INV_X1 U3598 ( .A(n2868), .ZN(n2802) );
  OAI21_X1 U3599 ( .B1(n3675), .B2(n3069), .A(n2802), .ZN(n2811) );
  NOR2_X1 U3600 ( .A1(n3000), .A2(n4320), .ZN(n2803) );
  NAND2_X1 U3601 ( .A1(n2804), .A2(n2803), .ZN(n2806) );
  AND2_X2 U3602 ( .A1(n2806), .A2(n4155), .ZN(n4460) );
  NAND2_X1 U3603 ( .A1(n2807), .A2(n3871), .ZN(n2808) );
  OAI22_X1 U3604 ( .A1(n4460), .A2(n3073), .B1(n3275), .B2(n3677), .ZN(n2810)
         );
  OR4_X1 U3605 ( .A1(n2813), .A2(n2812), .A3(n2811), .A4(n2810), .ZN(U3210) );
  NAND2_X1 U3606 ( .A1(U3149), .A2(DATAI_25_), .ZN(n2814) );
  OAI21_X1 U3607 ( .B1(n2815), .B2(U3149), .A(n2814), .ZN(U3327) );
  INV_X1 U3608 ( .A(DATAI_31_), .ZN(n2819) );
  OR2_X1 U3609 ( .A1(n2816), .A2(IR_REG_29__SCAN_IN), .ZN(n2817) );
  OR4_X1 U3610 ( .A1(n2817), .A2(IR_REG_30__SCAN_IN), .A3(n2617), .A4(U3149), 
        .ZN(n2818) );
  OAI21_X1 U3611 ( .B1(STATE_REG_SCAN_IN), .B2(n2819), .A(n2818), .ZN(U3321)
         );
  INV_X1 U3612 ( .A(DATAI_20_), .ZN(n4048) );
  NAND2_X1 U3613 ( .A1(n2820), .A2(STATE_REG_SCAN_IN), .ZN(n2821) );
  OAI21_X1 U3614 ( .B1(STATE_REG_SCAN_IN), .B2(n4048), .A(n2821), .ZN(U3332)
         );
  INV_X1 U3615 ( .A(DATAI_21_), .ZN(n4054) );
  NAND2_X1 U3616 ( .A1(n3771), .A2(STATE_REG_SCAN_IN), .ZN(n2822) );
  OAI21_X1 U3617 ( .B1(STATE_REG_SCAN_IN), .B2(n4054), .A(n2822), .ZN(U3331)
         );
  INV_X1 U3618 ( .A(n3000), .ZN(n2823) );
  NAND2_X1 U3619 ( .A1(n2824), .A2(n2823), .ZN(n4632) );
  INV_X1 U3620 ( .A(D_REG_0__SCAN_IN), .ZN(n2826) );
  NOR3_X1 U3621 ( .A1(n2680), .A2(n4635), .A3(n4441), .ZN(n2825) );
  AOI21_X1 U3622 ( .B1(n4632), .B2(n2826), .A(n2825), .ZN(U3458) );
  INV_X1 U3623 ( .A(D_REG_1__SCAN_IN), .ZN(n2830) );
  INV_X1 U3624 ( .A(n2827), .ZN(n2829) );
  AOI22_X1 U3625 ( .A1(n4632), .A2(n2830), .B1(n2829), .B2(n2828), .ZN(U3459)
         );
  INV_X1 U3626 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n3894) );
  NAND2_X1 U3627 ( .A1(n3337), .A2(U4043), .ZN(n2831) );
  OAI21_X1 U3628 ( .B1(U4043), .B2(n3894), .A(n2831), .ZN(U3562) );
  INV_X1 U3629 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n4037) );
  NAND2_X1 U3630 ( .A1(n2733), .A2(U4043), .ZN(n2832) );
  OAI21_X1 U3631 ( .B1(U4043), .B2(n4037), .A(n2832), .ZN(U3550) );
  INV_X1 U3632 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n3890) );
  NAND2_X1 U3633 ( .A1(n4324), .A2(U4043), .ZN(n2833) );
  OAI21_X1 U3634 ( .B1(U4043), .B2(n3890), .A(n2833), .ZN(U3568) );
  INV_X1 U3635 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n3895) );
  NAND2_X1 U3636 ( .A1(n3067), .A2(U4043), .ZN(n2834) );
  OAI21_X1 U3637 ( .B1(U4043), .B2(n3895), .A(n2834), .ZN(U3558) );
  OR2_X1 U3638 ( .A1(n2835), .A2(U3149), .ZN(n3841) );
  NAND2_X1 U3639 ( .A1(n3000), .A2(n3841), .ZN(n2841) );
  NAND2_X1 U3640 ( .A1(n2836), .A2(n2835), .ZN(n2837) );
  AND2_X1 U3641 ( .A1(n2837), .A2(n2058), .ZN(n2840) );
  INV_X1 U3642 ( .A(n2840), .ZN(n2838) );
  NOR2_X1 U3643 ( .A1(n4597), .A2(U4043), .ZN(U3148) );
  INV_X1 U3644 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n4053) );
  NAND2_X1 U3645 ( .A1(n4453), .A2(U4043), .ZN(n2839) );
  OAI21_X1 U3646 ( .B1(U4043), .B2(n4053), .A(n2839), .ZN(U3566) );
  NAND2_X1 U3647 ( .A1(n2841), .A2(n2840), .ZN(n4484) );
  NAND2_X1 U3648 ( .A1(n2843), .A2(n2842), .ZN(n4145) );
  INV_X1 U3649 ( .A(n4145), .ZN(n4481) );
  INV_X1 U3650 ( .A(n2887), .ZN(n4447) );
  INV_X1 U3651 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2845) );
  AND2_X1 U3652 ( .A1(REG1_REG_0__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n3862)
         );
  NAND2_X1 U3653 ( .A1(n4451), .A2(REG1_REG_1__SCAN_IN), .ZN(n2846) );
  NAND2_X1 U3654 ( .A1(n4450), .A2(REG1_REG_2__SCAN_IN), .ZN(n2847) );
  NAND2_X1 U3655 ( .A1(n3877), .A2(n2847), .ZN(n2848) );
  NAND2_X1 U3656 ( .A1(n2891), .A2(REG1_REG_3__SCAN_IN), .ZN(n2850) );
  NAND2_X1 U3657 ( .A1(n2848), .A2(n4449), .ZN(n2849) );
  NAND2_X1 U3658 ( .A1(n2850), .A2(n2849), .ZN(n2851) );
  INV_X1 U3659 ( .A(n4448), .ZN(n4491) );
  MUX2_X1 U3660 ( .A(REG1_REG_5__SCAN_IN), .B(n2371), .S(n2887), .Z(n2075) );
  XNOR2_X1 U3661 ( .A(n2852), .B(n4446), .ZN(n2875) );
  INV_X1 U3662 ( .A(n2852), .ZN(n2853) );
  MUX2_X1 U3663 ( .A(n4070), .B(REG1_REG_7__SCAN_IN), .S(n4445), .Z(n2854) );
  XNOR2_X1 U3664 ( .A(n4069), .B(n2854), .ZN(n2873) );
  INV_X1 U3665 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2856) );
  MUX2_X1 U3666 ( .A(REG2_REG_1__SCAN_IN), .B(n2856), .S(n2855), .Z(n3863) );
  NAND2_X1 U3667 ( .A1(REG2_REG_0__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n3872) );
  NAND2_X1 U3668 ( .A1(n4451), .A2(REG2_REG_1__SCAN_IN), .ZN(n2857) );
  OAI21_X1 U3669 ( .B1(n3863), .B2(n3872), .A(n2857), .ZN(n3884) );
  NAND2_X1 U3670 ( .A1(n4450), .A2(REG2_REG_2__SCAN_IN), .ZN(n2858) );
  NAND2_X1 U3671 ( .A1(n2892), .A2(REG2_REG_3__SCAN_IN), .ZN(n2861) );
  NAND2_X1 U3672 ( .A1(n2859), .A2(n4449), .ZN(n2860) );
  NAND2_X1 U3673 ( .A1(n2861), .A2(n2860), .ZN(n2862) );
  XNOR2_X1 U3674 ( .A(n2862), .B(n4491), .ZN(n4492) );
  AOI22_X1 U3675 ( .A1(n4492), .A2(REG2_REG_4__SCAN_IN), .B1(n4448), .B2(n2862), .ZN(n2884) );
  INV_X1 U3676 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2863) );
  MUX2_X1 U3677 ( .A(REG2_REG_5__SCAN_IN), .B(n2863), .S(n2887), .Z(n2883) );
  INV_X1 U3678 ( .A(n2864), .ZN(n2865) );
  INV_X1 U3679 ( .A(REG2_REG_7__SCAN_IN), .ZN(n4092) );
  MUX2_X1 U3680 ( .A(n4092), .B(REG2_REG_7__SCAN_IN), .S(n4445), .Z(n2866) );
  OR2_X1 U3681 ( .A1(n3871), .A2(n4145), .ZN(n3873) );
  OR2_X1 U3682 ( .A1(n4484), .A2(n3873), .ZN(n4560) );
  AOI21_X1 U3683 ( .B1(n2867), .B2(n2866), .A(n4560), .ZN(n2871) );
  INV_X1 U3684 ( .A(n4445), .ZN(n4091) );
  AOI21_X1 U3685 ( .B1(n4597), .B2(ADDR_REG_7__SCAN_IN), .A(n2868), .ZN(n2869)
         );
  OAI21_X1 U3686 ( .B1(n4611), .B2(n4091), .A(n2869), .ZN(n2870) );
  AOI21_X1 U3687 ( .B1(n2871), .B2(n4090), .A(n2870), .ZN(n2872) );
  OAI21_X1 U3688 ( .B1(n4594), .B2(n2873), .A(n2872), .ZN(U3247) );
  XNOR2_X1 U3689 ( .A(n2874), .B(REG2_REG_6__SCAN_IN), .ZN(n2881) );
  XOR2_X1 U3690 ( .A(REG1_REG_6__SCAN_IN), .B(n2875), .Z(n2879) );
  INV_X1 U3691 ( .A(n4594), .ZN(n4589) );
  INV_X1 U3692 ( .A(n4446), .ZN(n2877) );
  AND2_X1 U3693 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n2949) );
  AOI21_X1 U3694 ( .B1(n4597), .B2(ADDR_REG_6__SCAN_IN), .A(n2949), .ZN(n2876)
         );
  OAI21_X1 U3695 ( .B1(n4611), .B2(n2877), .A(n2876), .ZN(n2878) );
  AOI21_X1 U3696 ( .B1(n2879), .B2(n4589), .A(n2878), .ZN(n2880) );
  OAI21_X1 U3697 ( .B1(n2881), .B2(n4560), .A(n2880), .ZN(U3246) );
  AOI211_X1 U3698 ( .C1(n2884), .C2(n2883), .A(n2882), .B(n4560), .ZN(n2890)
         );
  AOI211_X1 U3699 ( .C1(n2885), .C2(n2075), .A(n2093), .B(n4594), .ZN(n2889)
         );
  AND2_X1 U3700 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n2988) );
  AOI21_X1 U3701 ( .B1(n4597), .B2(ADDR_REG_5__SCAN_IN), .A(n2988), .ZN(n2886)
         );
  OAI21_X1 U3702 ( .B1(n4611), .B2(n2887), .A(n2886), .ZN(n2888) );
  OR3_X1 U3703 ( .A1(n2890), .A2(n2889), .A3(n2888), .ZN(U3245) );
  XOR2_X1 U3704 ( .A(n2891), .B(REG1_REG_3__SCAN_IN), .Z(n2894) );
  XOR2_X1 U3705 ( .A(REG2_REG_3__SCAN_IN), .B(n2892), .Z(n2893) );
  AOI22_X1 U3706 ( .A1(n4589), .A2(n2894), .B1(n4608), .B2(n2893), .ZN(n2896)
         );
  NOR2_X1 U3707 ( .A1(STATE_REG_SCAN_IN), .A2(n2360), .ZN(n3036) );
  AOI21_X1 U3708 ( .B1(n4597), .B2(ADDR_REG_3__SCAN_IN), .A(n3036), .ZN(n2895)
         );
  OAI211_X1 U3709 ( .C1(n2897), .C2(n4611), .A(n2896), .B(n2895), .ZN(U3243)
         );
  INV_X1 U3710 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n3897) );
  NAND2_X1 U3711 ( .A1(n4299), .A2(U4043), .ZN(n2898) );
  OAI21_X1 U3712 ( .B1(U4043), .B2(n3897), .A(n2898), .ZN(U3571) );
  AOI222_X1 U3713 ( .A1(n2235), .A2(REG2_REG_30__SCAN_IN), .B1(n2899), .B2(
        REG1_REG_30__SCAN_IN), .C1(n3696), .C2(REG0_REG_30__SCAN_IN), .ZN(
        n4148) );
  INV_X2 U3714 ( .A(U4043), .ZN(n3875) );
  NAND2_X1 U3715 ( .A1(n3875), .A2(DATAO_REG_30__SCAN_IN), .ZN(n2900) );
  OAI21_X1 U3716 ( .B1(n4148), .B2(n3875), .A(n2900), .ZN(U3580) );
  INV_X1 U3717 ( .A(n2901), .ZN(n2903) );
  NOR3_X1 U3718 ( .A1(n2903), .A2(n2902), .A3(n3000), .ZN(n2920) );
  OAI21_X1 U3719 ( .B1(n2906), .B2(n2905), .A(n2904), .ZN(n2907) );
  NAND2_X1 U3720 ( .A1(n2907), .A2(n3665), .ZN(n2910) );
  INV_X1 U3721 ( .A(n4460), .ZN(n3645) );
  OAI22_X1 U3722 ( .A1(n2933), .A2(n3677), .B1(n3675), .B2(n2744), .ZN(n2908)
         );
  AOI21_X1 U3723 ( .B1(n3645), .B2(n2936), .A(n2908), .ZN(n2909) );
  OAI211_X1 U3724 ( .C1(n2920), .C2(n2911), .A(n2910), .B(n2909), .ZN(U3234)
         );
  INV_X1 U3725 ( .A(n2912), .ZN(n2913) );
  XNOR2_X1 U3726 ( .A(n2914), .B(n2913), .ZN(n3869) );
  AOI22_X1 U3727 ( .A1(n3665), .A2(n3869), .B1(n4454), .B2(n3859), .ZN(n2916)
         );
  NAND2_X1 U3728 ( .A1(n3645), .A2(n3096), .ZN(n2915) );
  OAI211_X1 U3729 ( .C1(n2920), .C2(n2917), .A(n2916), .B(n2915), .ZN(U3229)
         );
  XNOR2_X1 U3730 ( .A(n2919), .B(n2918), .ZN(n2924) );
  OAI22_X1 U3731 ( .A1(n2729), .A2(n3675), .B1(n3677), .B2(n3184), .ZN(n2922)
         );
  NOR2_X1 U3732 ( .A1(n2920), .A2(n3099), .ZN(n2921) );
  AOI211_X1 U3733 ( .C1(n2334), .C2(n3645), .A(n2922), .B(n2921), .ZN(n2923)
         );
  OAI21_X1 U3734 ( .B1(n2924), .B2(n4465), .A(n2923), .ZN(U3219) );
  NAND2_X1 U3735 ( .A1(n2925), .A2(n3732), .ZN(n2926) );
  NAND2_X1 U3736 ( .A1(n2927), .A2(n2926), .ZN(n4621) );
  INV_X1 U3737 ( .A(n4621), .ZN(n2935) );
  INV_X1 U3738 ( .A(n3565), .ZN(n2975) );
  OAI21_X1 U3739 ( .B1(n3732), .B2(n2929), .A(n2928), .ZN(n2930) );
  NAND2_X1 U3740 ( .A1(n2930), .A2(n3409), .ZN(n2932) );
  INV_X1 U3741 ( .A(n4320), .ZN(n4347) );
  AOI22_X1 U3742 ( .A1(n3859), .A2(n4325), .B1(n2936), .B2(n4347), .ZN(n2931)
         );
  OAI211_X1 U3743 ( .C1(n2933), .C2(n4321), .A(n2932), .B(n2931), .ZN(n2934)
         );
  AOI21_X1 U3744 ( .B1(n2975), .B2(n4621), .A(n2934), .ZN(n4627) );
  OAI21_X1 U3745 ( .B1(n2935), .B2(n4699), .A(n4627), .ZN(n2942) );
  AND2_X1 U3746 ( .A1(n3094), .A2(n2936), .ZN(n2937) );
  OR2_X1 U3747 ( .A1(n2937), .A2(n3188), .ZN(n4620) );
  OAI22_X1 U3748 ( .A1(n4392), .A2(n4620), .B1(n4716), .B2(n2844), .ZN(n2938)
         );
  AOI21_X1 U3749 ( .B1(n2942), .B2(n4716), .A(n2938), .ZN(n2939) );
  INV_X1 U3750 ( .A(n2939), .ZN(U3520) );
  INV_X1 U3751 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2940) );
  OAI22_X1 U3752 ( .A1(n4435), .A2(n4620), .B1(n4705), .B2(n2940), .ZN(n2941)
         );
  AOI21_X1 U3753 ( .B1(n2942), .B2(n4705), .A(n2941), .ZN(n2943) );
  INV_X1 U3754 ( .A(n2943), .ZN(U3471) );
  INV_X1 U3755 ( .A(n2945), .ZN(n2947) );
  NOR2_X1 U3756 ( .A1(n2947), .A2(n2946), .ZN(n2948) );
  XNOR2_X1 U3757 ( .A(n2944), .B(n2948), .ZN(n2954) );
  AOI21_X1 U3758 ( .B1(n4454), .B2(n3853), .A(n2949), .ZN(n2951) );
  NAND2_X1 U3759 ( .A1(n4456), .A2(n3855), .ZN(n2950) );
  OAI211_X1 U3760 ( .C1(n4460), .C2(n2978), .A(n2951), .B(n2950), .ZN(n2952)
         );
  AOI21_X1 U3761 ( .B1(n3680), .B2(n4612), .A(n2952), .ZN(n2953) );
  OAI21_X1 U3762 ( .B1(n2954), .B2(n4465), .A(n2953), .ZN(U3236) );
  NAND2_X1 U3763 ( .A1(n2955), .A2(n3665), .ZN(n2966) );
  AOI21_X1 U3764 ( .B1(n2957), .B2(n2959), .A(n2958), .ZN(n2965) );
  INV_X1 U3765 ( .A(n3015), .ZN(n2963) );
  AND2_X1 U3766 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n4488) );
  AOI21_X1 U3767 ( .B1(n4454), .B2(n3855), .A(n4488), .ZN(n2961) );
  NAND2_X1 U3768 ( .A1(n4456), .A2(n3857), .ZN(n2960) );
  OAI211_X1 U3769 ( .C1(n4460), .C2(n3013), .A(n2961), .B(n2960), .ZN(n2962)
         );
  AOI21_X1 U3770 ( .B1(n3680), .B2(n2963), .A(n2962), .ZN(n2964) );
  OAI21_X1 U3771 ( .B1(n2966), .B2(n2965), .A(n2964), .ZN(U3227) );
  INV_X1 U3772 ( .A(n2968), .ZN(n3795) );
  AND2_X1 U3773 ( .A1(n3795), .A2(n3785), .ZN(n3756) );
  XNOR2_X1 U3774 ( .A(n2967), .B(n3756), .ZN(n4615) );
  INV_X1 U3775 ( .A(n4615), .ZN(n2976) );
  XNOR2_X1 U3776 ( .A(n2969), .B(n3756), .ZN(n2973) );
  OAI22_X1 U3777 ( .A1(n2970), .A2(n4277), .B1(n2978), .B2(n4320), .ZN(n2971)
         );
  AOI21_X1 U3778 ( .B1(n4298), .B2(n3853), .A(n2971), .ZN(n2972) );
  OAI21_X1 U3779 ( .B1(n2973), .B2(n4327), .A(n2972), .ZN(n2974) );
  AOI21_X1 U3780 ( .B1(n2975), .B2(n4615), .A(n2974), .ZN(n4618) );
  OAI21_X1 U3781 ( .B1(n4699), .B2(n2976), .A(n4618), .ZN(n2983) );
  INV_X1 U3782 ( .A(n3074), .ZN(n2977) );
  OAI21_X1 U3783 ( .B1(n3144), .B2(n2978), .A(n2977), .ZN(n4613) );
  INV_X1 U3784 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2979) );
  OAI22_X1 U3785 ( .A1(n4613), .A2(n4392), .B1(n4716), .B2(n2979), .ZN(n2980)
         );
  AOI21_X1 U3786 ( .B1(n2983), .B2(n4716), .A(n2980), .ZN(n2981) );
  INV_X1 U3787 ( .A(n2981), .ZN(U3524) );
  INV_X1 U3788 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3915) );
  OAI22_X1 U3789 ( .A1(n4613), .A2(n4435), .B1(n4705), .B2(n3915), .ZN(n2982)
         );
  AOI21_X1 U3790 ( .B1(n2983), .B2(n4705), .A(n2982), .ZN(n2984) );
  INV_X1 U3791 ( .A(n2984), .ZN(U3479) );
  XNOR2_X1 U3792 ( .A(n2986), .B(n2985), .ZN(n2994) );
  INV_X1 U3793 ( .A(n2987), .ZN(n3145) );
  AOI21_X1 U3794 ( .B1(n4454), .B2(n3854), .A(n2988), .ZN(n2990) );
  NAND2_X1 U3795 ( .A1(n4456), .A2(n3856), .ZN(n2989) );
  OAI211_X1 U3796 ( .C1(n4460), .C2(n2991), .A(n2990), .B(n2989), .ZN(n2992)
         );
  AOI21_X1 U3797 ( .B1(n3680), .B2(n3145), .A(n2992), .ZN(n2993) );
  OAI21_X1 U3798 ( .B1(n2994), .B2(n4465), .A(n2993), .ZN(U3224) );
  OR2_X1 U3799 ( .A1(n2995), .A2(n3728), .ZN(n2996) );
  NAND2_X1 U3800 ( .A1(n2997), .A2(n2996), .ZN(n4671) );
  INV_X1 U3801 ( .A(n2998), .ZN(n2999) );
  NOR2_X1 U3802 ( .A1(n3000), .A2(n2999), .ZN(n3002) );
  NAND4_X1 U3803 ( .A1(n3004), .A2(n3003), .A3(n3002), .A4(n3001), .ZN(n3005)
         );
  OR2_X1 U3804 ( .A1(n2717), .A2(n4132), .ZN(n3080) );
  OR2_X1 U3805 ( .A1(n4479), .A2(n3080), .ZN(n3580) );
  XOR2_X1 U3806 ( .A(n3728), .B(n3006), .Z(n3011) );
  AOI22_X1 U3807 ( .A1(n3857), .A2(n4325), .B1(n3007), .B2(n4347), .ZN(n3009)
         );
  NAND2_X1 U3808 ( .A1(n3855), .A2(n4298), .ZN(n3008) );
  OAI211_X1 U3809 ( .C1(n4671), .C2(n3565), .A(n3009), .B(n3008), .ZN(n3010)
         );
  AOI21_X1 U3810 ( .B1(n3011), .B2(n3409), .A(n3010), .ZN(n3012) );
  INV_X1 U3811 ( .A(n3012), .ZN(n4673) );
  INV_X1 U3812 ( .A(n3190), .ZN(n3014) );
  OAI211_X1 U3813 ( .C1(n3014), .C2(n3013), .A(n2707), .B(n3142), .ZN(n4672)
         );
  OAI22_X1 U3814 ( .A1(n4672), .A2(n4443), .B1(n4155), .B2(n3015), .ZN(n3016)
         );
  OAI21_X1 U3815 ( .B1(n4673), .B2(n3016), .A(n3575), .ZN(n3018) );
  NAND2_X1 U3816 ( .A1(n4479), .A2(REG2_REG_4__SCAN_IN), .ZN(n3017) );
  OAI211_X1 U3817 ( .C1(n4671), .C2(n3580), .A(n3018), .B(n3017), .ZN(U3286)
         );
  OR2_X1 U3818 ( .A1(n3079), .A2(n3727), .ZN(n4686) );
  NAND2_X1 U3819 ( .A1(n4686), .A2(n3019), .ZN(n3020) );
  NAND2_X1 U3820 ( .A1(n2087), .A2(n3790), .ZN(n3746) );
  XNOR2_X1 U3821 ( .A(n3020), .B(n3746), .ZN(n3129) );
  XNOR2_X1 U3822 ( .A(n3021), .B(n3746), .ZN(n3024) );
  AOI22_X1 U3823 ( .A1(n3852), .A2(n4298), .B1(n4347), .B2(n3025), .ZN(n3022)
         );
  OAI21_X1 U3824 ( .B1(n3058), .B2(n4277), .A(n3022), .ZN(n3023) );
  AOI21_X1 U3825 ( .B1(n3024), .B2(n3409), .A(n3023), .ZN(n3134) );
  OAI21_X1 U3826 ( .B1(n3129), .B2(n4678), .A(n3134), .ZN(n3031) );
  NAND2_X1 U3827 ( .A1(n3072), .A2(n3025), .ZN(n3026) );
  NAND2_X1 U3828 ( .A1(n3282), .A2(n3026), .ZN(n3126) );
  INV_X1 U3829 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3027) );
  OAI22_X1 U3830 ( .A1(n3126), .A2(n4435), .B1(n4705), .B2(n3027), .ZN(n3028)
         );
  AOI21_X1 U3831 ( .B1(n3031), .B2(n4705), .A(n3028), .ZN(n3029) );
  INV_X1 U3832 ( .A(n3029), .ZN(U3483) );
  OAI22_X1 U3833 ( .A1(n3126), .A2(n4392), .B1(n4716), .B2(n2411), .ZN(n3030)
         );
  AOI21_X1 U3834 ( .B1(n3031), .B2(n4716), .A(n3030), .ZN(n3032) );
  INV_X1 U3835 ( .A(n3032), .ZN(U3526) );
  OAI21_X1 U3836 ( .B1(n3034), .B2(n3033), .A(n2957), .ZN(n3040) );
  OAI22_X1 U3837 ( .A1(n4460), .A2(n2754), .B1(n3184), .B2(n3675), .ZN(n3035)
         );
  INV_X1 U3838 ( .A(n3035), .ZN(n3038) );
  AOI21_X1 U3839 ( .B1(n4454), .B2(n3856), .A(n3036), .ZN(n3037) );
  OAI211_X1 U3840 ( .C1(n4472), .C2(REG3_REG_3__SCAN_IN), .A(n3038), .B(n3037), 
        .ZN(n3039) );
  AOI21_X1 U3841 ( .B1(n3040), .B2(n3665), .A(n3039), .ZN(n3041) );
  INV_X1 U3842 ( .A(n3041), .ZN(U3215) );
  INV_X1 U3843 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3050) );
  INV_X1 U3844 ( .A(n3042), .ZN(n3043) );
  NAND2_X1 U3845 ( .A1(n3096), .A2(n3043), .ZN(n4655) );
  NAND2_X1 U3846 ( .A1(n2733), .A2(n3044), .ZN(n3770) );
  NAND2_X1 U3847 ( .A1(n3100), .A2(n3770), .ZN(n4659) );
  NAND2_X1 U3848 ( .A1(n3565), .A2(n4327), .ZN(n3045) );
  AOI22_X1 U3849 ( .A1(n4659), .A2(n3045), .B1(n4298), .B2(n3859), .ZN(n4656)
         );
  OAI21_X1 U3850 ( .B1(n3046), .B2(n4655), .A(n4656), .ZN(n3047) );
  INV_X1 U3851 ( .A(n4155), .ZN(n4619) );
  AOI22_X1 U3852 ( .A1(n3575), .A2(n3047), .B1(REG3_REG_0__SCAN_IN), .B2(n4619), .ZN(n3049) );
  INV_X1 U3853 ( .A(n3580), .ZN(n4622) );
  NAND2_X1 U3854 ( .A1(n4622), .A2(n4659), .ZN(n3048) );
  OAI211_X1 U3855 ( .C1(n3575), .C2(n3050), .A(n3049), .B(n3048), .ZN(U3290)
         );
  NAND2_X1 U3856 ( .A1(n3052), .A2(n3051), .ZN(n3053) );
  OAI22_X1 U3857 ( .A1(n3275), .A2(n3540), .B1(n2056), .B2(n3059), .ZN(n3055)
         );
  XNOR2_X1 U3858 ( .A(n3055), .B(n3546), .ZN(n3115) );
  OAI22_X1 U3859 ( .A1(n3275), .A2(n3525), .B1(n3540), .B2(n3059), .ZN(n3116)
         );
  XNOR2_X1 U3860 ( .A(n3115), .B(n3116), .ZN(n3056) );
  XNOR2_X1 U3861 ( .A(n3117), .B(n3056), .ZN(n3057) );
  NAND2_X1 U3862 ( .A1(n3057), .A2(n3665), .ZN(n3064) );
  OAI22_X1 U3863 ( .A1(n4460), .A2(n3059), .B1(n3058), .B2(n3675), .ZN(n3062)
         );
  NAND2_X1 U3864 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n4500) );
  OAI21_X1 U3865 ( .B1(n3677), .B2(n3060), .A(n4500), .ZN(n3061) );
  NOR2_X1 U3866 ( .A1(n3062), .A2(n3061), .ZN(n3063) );
  OAI211_X1 U3867 ( .C1(n4472), .C2(n3127), .A(n3064), .B(n3063), .ZN(U3218)
         );
  XNOR2_X1 U3868 ( .A(n3065), .B(n3727), .ZN(n3071) );
  AOI22_X1 U3869 ( .A1(n3067), .A2(n4298), .B1(n4347), .B2(n3066), .ZN(n3068)
         );
  OAI21_X1 U3870 ( .B1(n3069), .B2(n4277), .A(n3068), .ZN(n3070) );
  AOI21_X1 U3871 ( .B1(n3071), .B2(n3409), .A(n3070), .ZN(n4689) );
  OAI211_X1 U3872 ( .C1(n3074), .C2(n3073), .A(n2707), .B(n3072), .ZN(n4688)
         );
  INV_X1 U3873 ( .A(n4688), .ZN(n3078) );
  INV_X1 U3874 ( .A(n3415), .ZN(n3077) );
  OAI22_X1 U3875 ( .A1(n3575), .A2(n4092), .B1(n3075), .B2(n4155), .ZN(n3076)
         );
  AOI21_X1 U3876 ( .B1(n3078), .B2(n3077), .A(n3076), .ZN(n3083) );
  NAND2_X1 U3877 ( .A1(n3079), .A2(n3727), .ZN(n4685) );
  AND2_X1 U3878 ( .A1(n3565), .A2(n3080), .ZN(n3081) );
  INV_X1 U3879 ( .A(n4338), .ZN(n3288) );
  NAND3_X1 U3880 ( .A1(n4686), .A2(n4685), .A3(n3288), .ZN(n3082) );
  OAI211_X1 U3881 ( .C1(n4689), .C2(n4479), .A(n3083), .B(n3082), .ZN(U3283)
         );
  NAND2_X1 U3882 ( .A1(n3796), .A2(n3802), .ZN(n3745) );
  XNOR2_X1 U3883 ( .A(n3084), .B(n3745), .ZN(n3171) );
  XNOR2_X1 U3884 ( .A(n3085), .B(n3745), .ZN(n3088) );
  OAI22_X1 U3885 ( .A1(n3306), .A2(n4321), .B1(n4320), .B2(n3165), .ZN(n3086)
         );
  AOI21_X1 U3886 ( .B1(n4325), .B2(n3852), .A(n3086), .ZN(n3087) );
  OAI21_X1 U3887 ( .B1(n3088), .B2(n4327), .A(n3087), .ZN(n3172) );
  AOI21_X1 U3888 ( .B1(n4694), .B2(n3171), .A(n3172), .ZN(n3093) );
  AOI21_X1 U3889 ( .B1(n3151), .B2(n3283), .A(n3572), .ZN(n3176) );
  INV_X1 U3890 ( .A(n4392), .ZN(n3089) );
  AOI22_X1 U3891 ( .A1(n3176), .A2(n3089), .B1(n4714), .B2(
        REG1_REG_10__SCAN_IN), .ZN(n3090) );
  OAI21_X1 U3892 ( .B1(n3093), .B2(n4714), .A(n3090), .ZN(U3528) );
  INV_X1 U3893 ( .A(n4435), .ZN(n3091) );
  AOI22_X1 U3894 ( .A1(n3176), .A2(n3091), .B1(n4703), .B2(
        REG0_REG_10__SCAN_IN), .ZN(n3092) );
  OAI21_X1 U3895 ( .B1(n3093), .B2(n4703), .A(n3092), .ZN(U3487) );
  NOR2_X2 U3896 ( .A1(n3415), .A2(n4698), .ZN(n4624) );
  INV_X1 U3897 ( .A(n3094), .ZN(n3095) );
  AOI21_X1 U3898 ( .B1(n2334), .B2(n3096), .A(n3095), .ZN(n4664) );
  OAI21_X1 U3899 ( .B1(n2628), .B2(n3098), .A(n3097), .ZN(n4661) );
  OAI22_X1 U3900 ( .A1(n3580), .A2(n4661), .B1(n3099), .B2(n4155), .ZN(n3108)
         );
  INV_X1 U3901 ( .A(n3100), .ZN(n3772) );
  XNOR2_X1 U3902 ( .A(n2628), .B(n3772), .ZN(n3106) );
  OR2_X1 U3903 ( .A1(n4661), .A2(n3565), .ZN(n3105) );
  NAND2_X1 U3904 ( .A1(n2334), .A2(n4347), .ZN(n3102) );
  NAND2_X1 U3905 ( .A1(n2733), .A2(n4325), .ZN(n3101) );
  OAI211_X1 U3906 ( .C1(n3184), .C2(n4321), .A(n3102), .B(n3101), .ZN(n3103)
         );
  INV_X1 U3907 ( .A(n3103), .ZN(n3104) );
  OAI211_X1 U3908 ( .C1(n3106), .C2(n4327), .A(n3105), .B(n3104), .ZN(n4662)
         );
  MUX2_X1 U3909 ( .A(n4662), .B(REG2_REG_1__SCAN_IN), .S(n4479), .Z(n3107) );
  AOI211_X1 U3910 ( .C1(n4624), .C2(n4664), .A(n3108), .B(n3107), .ZN(n3109)
         );
  INV_X1 U3911 ( .A(n3109), .ZN(U3289) );
  NAND2_X1 U3912 ( .A1(n3852), .A2(n3534), .ZN(n3111) );
  NAND2_X1 U3913 ( .A1(n3544), .A2(n3273), .ZN(n3110) );
  NAND2_X1 U3914 ( .A1(n3111), .A2(n3110), .ZN(n3112) );
  XNOR2_X1 U3915 ( .A(n3112), .B(n3546), .ZN(n3154) );
  NAND2_X1 U3916 ( .A1(n3852), .A2(n3545), .ZN(n3114) );
  NAND2_X1 U3917 ( .A1(n3534), .A2(n3273), .ZN(n3113) );
  NAND2_X1 U3918 ( .A1(n3114), .A2(n3113), .ZN(n3155) );
  XNOR2_X1 U3919 ( .A(n3154), .B(n3155), .ZN(n3120) );
  INV_X1 U3920 ( .A(n3159), .ZN(n3118) );
  AOI21_X1 U3921 ( .B1(n3120), .B2(n3119), .A(n3118), .ZN(n3125) );
  AND2_X1 U3922 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4509) );
  OAI22_X1 U3923 ( .A1(n4460), .A2(n3284), .B1(n3275), .B2(n3675), .ZN(n3121)
         );
  AOI211_X1 U3924 ( .C1(n4454), .C2(n3851), .A(n4509), .B(n3121), .ZN(n3124)
         );
  INV_X1 U3925 ( .A(n3285), .ZN(n3122) );
  NAND2_X1 U3926 ( .A1(n3680), .A2(n3122), .ZN(n3123) );
  OAI211_X1 U3927 ( .C1(n3125), .C2(n4465), .A(n3124), .B(n3123), .ZN(U3228)
         );
  INV_X1 U3928 ( .A(n3126), .ZN(n3132) );
  INV_X1 U3929 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3128) );
  OAI22_X1 U3930 ( .A1(n3575), .A2(n3128), .B1(n3127), .B2(n4155), .ZN(n3131)
         );
  NOR2_X1 U3931 ( .A1(n3129), .A2(n4338), .ZN(n3130) );
  AOI211_X1 U3932 ( .C1(n3132), .C2(n4624), .A(n3131), .B(n3130), .ZN(n3133)
         );
  OAI21_X1 U3933 ( .B1(n4479), .B2(n3134), .A(n3133), .ZN(U3282) );
  NAND2_X1 U3934 ( .A1(n3793), .A2(n3782), .ZN(n3744) );
  XNOR2_X1 U3935 ( .A(n3135), .B(n3744), .ZN(n4679) );
  XNOR2_X1 U3936 ( .A(n3136), .B(n3744), .ZN(n3140) );
  AOI22_X1 U3937 ( .A1(n3854), .A2(n4298), .B1(n4347), .B2(n3141), .ZN(n3137)
         );
  OAI21_X1 U3938 ( .B1(n3138), .B2(n4277), .A(n3137), .ZN(n3139) );
  AOI21_X1 U3939 ( .B1(n3140), .B2(n3409), .A(n3139), .ZN(n4680) );
  MUX2_X1 U3940 ( .A(n2863), .B(n4680), .S(n3575), .Z(n3147) );
  AND2_X1 U3941 ( .A1(n3142), .A2(n3141), .ZN(n3143) );
  NOR2_X1 U3942 ( .A1(n3144), .A2(n3143), .ZN(n4683) );
  AOI22_X1 U3943 ( .A1(n4624), .A2(n4683), .B1(n3145), .B2(n4619), .ZN(n3146)
         );
  OAI211_X1 U3944 ( .C1(n4338), .C2(n4679), .A(n3147), .B(n3146), .ZN(U3285)
         );
  NAND2_X1 U3945 ( .A1(n3851), .A2(n3534), .ZN(n3149) );
  NAND2_X1 U3946 ( .A1(n3544), .A2(n3151), .ZN(n3148) );
  NAND2_X1 U3947 ( .A1(n3149), .A2(n3148), .ZN(n3150) );
  XNOR2_X1 U3948 ( .A(n3150), .B(n3538), .ZN(n3202) );
  NAND2_X1 U3949 ( .A1(n3851), .A2(n3545), .ZN(n3153) );
  NAND2_X1 U3950 ( .A1(n3534), .A2(n3151), .ZN(n3152) );
  NAND2_X1 U3951 ( .A1(n3153), .A2(n3152), .ZN(n3203) );
  XNOR2_X1 U3952 ( .A(n3202), .B(n3203), .ZN(n3160) );
  INV_X1 U3953 ( .A(n3154), .ZN(n3157) );
  INV_X1 U3954 ( .A(n3155), .ZN(n3156) );
  NAND2_X1 U3955 ( .A1(n3157), .A2(n3156), .ZN(n3161) );
  NAND2_X1 U3956 ( .A1(n3206), .A2(n3665), .ZN(n3170) );
  AOI21_X1 U3957 ( .B1(n3159), .B2(n3161), .A(n3160), .ZN(n3169) );
  INV_X1 U3958 ( .A(n3173), .ZN(n3167) );
  NOR2_X1 U3959 ( .A1(STATE_REG_SCAN_IN), .A2(n3162), .ZN(n4521) );
  AOI21_X1 U3960 ( .B1(n4456), .B2(n3852), .A(n4521), .ZN(n3164) );
  NAND2_X1 U3961 ( .A1(n4454), .A2(n3850), .ZN(n3163) );
  OAI211_X1 U3962 ( .C1(n4460), .C2(n3165), .A(n3164), .B(n3163), .ZN(n3166)
         );
  AOI21_X1 U3963 ( .B1(n3680), .B2(n3167), .A(n3166), .ZN(n3168) );
  OAI21_X1 U3964 ( .B1(n3170), .B2(n3169), .A(n3168), .ZN(U3214) );
  INV_X1 U3965 ( .A(n3171), .ZN(n3179) );
  NAND2_X1 U3966 ( .A1(n3172), .A2(n3575), .ZN(n3178) );
  INV_X1 U3967 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3174) );
  OAI22_X1 U3968 ( .A1(n3575), .A2(n3174), .B1(n3173), .B2(n4155), .ZN(n3175)
         );
  AOI21_X1 U3969 ( .B1(n3176), .B2(n4624), .A(n3175), .ZN(n3177) );
  OAI211_X1 U3970 ( .C1(n4338), .C2(n3179), .A(n3178), .B(n3177), .ZN(U3280)
         );
  XNOR2_X1 U3971 ( .A(n3180), .B(n3733), .ZN(n4667) );
  XNOR2_X1 U3972 ( .A(n3181), .B(n3733), .ZN(n3186) );
  AOI22_X1 U3973 ( .A1(n3856), .A2(n4298), .B1(n4347), .B2(n3182), .ZN(n3183)
         );
  OAI21_X1 U3974 ( .B1(n3184), .B2(n4277), .A(n3183), .ZN(n3185) );
  AOI21_X1 U3975 ( .B1(n3186), .B2(n3409), .A(n3185), .ZN(n3187) );
  OAI21_X1 U3976 ( .B1(n4667), .B2(n3565), .A(n3187), .ZN(n4669) );
  AOI22_X1 U3977 ( .A1(n4479), .A2(REG2_REG_3__SCAN_IN), .B1(n4619), .B2(n2360), .ZN(n3193) );
  OR2_X1 U3978 ( .A1(n3188), .A2(n2754), .ZN(n3189) );
  NAND2_X1 U3979 ( .A1(n3190), .A2(n3189), .ZN(n4666) );
  INV_X1 U3980 ( .A(n4666), .ZN(n3191) );
  NAND2_X1 U3981 ( .A1(n4624), .A2(n3191), .ZN(n3192) );
  OAI211_X1 U3982 ( .C1(n4667), .C2(n3580), .A(n3193), .B(n3192), .ZN(n3194)
         );
  AOI21_X1 U3983 ( .B1(n4669), .B2(n3575), .A(n3194), .ZN(n3195) );
  INV_X1 U3984 ( .A(n3195), .ZN(U3287) );
  OAI22_X1 U3985 ( .A1(n3306), .A2(n3540), .B1(n2056), .B2(n3571), .ZN(n3196)
         );
  XNOR2_X1 U3986 ( .A(n3196), .B(n3538), .ZN(n3201) );
  INV_X1 U3987 ( .A(n3201), .ZN(n3199) );
  NOR2_X1 U3988 ( .A1(n3571), .A2(n3540), .ZN(n3197) );
  AOI21_X1 U3989 ( .B1(n3850), .B2(n3545), .A(n3197), .ZN(n3200) );
  INV_X1 U3990 ( .A(n3200), .ZN(n3198) );
  NAND2_X1 U3991 ( .A1(n3199), .A2(n3198), .ZN(n3299) );
  NAND2_X1 U3992 ( .A1(n3201), .A2(n3200), .ZN(n3297) );
  NAND2_X1 U3993 ( .A1(n3299), .A2(n3297), .ZN(n3207) );
  INV_X1 U3994 ( .A(n3202), .ZN(n3204) );
  NAND2_X1 U3995 ( .A1(n3204), .A2(n3203), .ZN(n3205) );
  XOR2_X1 U3996 ( .A(n3207), .B(n3298), .Z(n3213) );
  INV_X1 U3997 ( .A(n3573), .ZN(n3211) );
  AND2_X1 U3998 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4528) );
  AOI21_X1 U3999 ( .B1(n4456), .B2(n3851), .A(n4528), .ZN(n3209) );
  NAND2_X1 U4000 ( .A1(n4454), .A2(n3337), .ZN(n3208) );
  OAI211_X1 U4001 ( .C1(n4460), .C2(n3571), .A(n3209), .B(n3208), .ZN(n3210)
         );
  AOI21_X1 U4002 ( .B1(n3680), .B2(n3211), .A(n3210), .ZN(n3212) );
  OAI21_X1 U4003 ( .B1(n3213), .B2(n4465), .A(n3212), .ZN(U3233) );
  NAND2_X1 U4004 ( .A1(n3570), .A2(n3219), .ZN(n3214) );
  NAND2_X1 U4005 ( .A1(n3256), .A2(n3214), .ZN(n3267) );
  NAND2_X1 U4006 ( .A1(n3245), .A2(n3246), .ZN(n3747) );
  XNOR2_X1 U4007 ( .A(n3215), .B(n3747), .ZN(n3269) );
  NAND2_X1 U4008 ( .A1(n3269), .A2(n4694), .ZN(n3224) );
  NAND2_X1 U4009 ( .A1(n3217), .A2(n3216), .ZN(n3248) );
  INV_X1 U4010 ( .A(n3747), .ZN(n3218) );
  XNOR2_X1 U4011 ( .A(n3248), .B(n3218), .ZN(n3223) );
  NAND2_X1 U4012 ( .A1(n3850), .A2(n4325), .ZN(n3221) );
  NAND2_X1 U4013 ( .A1(n3219), .A2(n4347), .ZN(n3220) );
  OAI211_X1 U4014 ( .C1(n3389), .C2(n4321), .A(n3221), .B(n3220), .ZN(n3222)
         );
  AOI21_X1 U4015 ( .B1(n3223), .B2(n3409), .A(n3222), .ZN(n3271) );
  NAND2_X1 U4016 ( .A1(n3224), .A2(n3271), .ZN(n3227) );
  MUX2_X1 U4017 ( .A(n3227), .B(REG1_REG_12__SCAN_IN), .S(n4714), .Z(n3225) );
  INV_X1 U4018 ( .A(n3225), .ZN(n3226) );
  OAI21_X1 U4019 ( .B1(n4392), .B2(n3267), .A(n3226), .ZN(U3530) );
  MUX2_X1 U4020 ( .A(REG0_REG_12__SCAN_IN), .B(n3227), .S(n4705), .Z(n3228) );
  INV_X1 U4021 ( .A(n3228), .ZN(n3229) );
  OAI21_X1 U4022 ( .B1(n3267), .B2(n4435), .A(n3229), .ZN(U3491) );
  OAI21_X1 U4023 ( .B1(n2078), .B2(n3231), .A(n3230), .ZN(n3353) );
  INV_X1 U4024 ( .A(n3353), .ZN(n3243) );
  OAI21_X1 U4025 ( .B1(n3754), .B2(n3687), .A(n3313), .ZN(n3235) );
  AOI22_X1 U4026 ( .A1(n3848), .A2(n4298), .B1(n4347), .B2(n3232), .ZN(n3233)
         );
  OAI21_X1 U4027 ( .B1(n3389), .B2(n4277), .A(n3233), .ZN(n3234) );
  AOI21_X1 U4028 ( .B1(n3235), .B2(n3409), .A(n3234), .ZN(n3236) );
  OAI21_X1 U4029 ( .B1(n3243), .B2(n3565), .A(n3236), .ZN(n3352) );
  NAND2_X1 U4030 ( .A1(n3352), .A2(n3575), .ZN(n3242) );
  INV_X1 U4031 ( .A(n3318), .ZN(n3237) );
  OAI21_X1 U4032 ( .B1(n3257), .B2(n3388), .A(n3237), .ZN(n3357) );
  INV_X1 U4033 ( .A(n3357), .ZN(n3240) );
  INV_X1 U4034 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3238) );
  OAI22_X1 U4035 ( .A1(n3575), .A2(n3238), .B1(n3394), .B2(n4155), .ZN(n3239)
         );
  AOI21_X1 U4036 ( .B1(n3240), .B2(n4624), .A(n3239), .ZN(n3241) );
  OAI211_X1 U4037 ( .C1(n3243), .C2(n3580), .A(n3242), .B(n3241), .ZN(U3276)
         );
  XNOR2_X1 U4038 ( .A(n3389), .B(n3250), .ZN(n3758) );
  XOR2_X1 U4039 ( .A(n3758), .B(n3244), .Z(n3255) );
  INV_X1 U4040 ( .A(n3245), .ZN(n3247) );
  OAI21_X1 U4041 ( .B1(n3248), .B2(n3247), .A(n3246), .ZN(n3249) );
  XNOR2_X1 U4042 ( .A(n3249), .B(n3758), .ZN(n3253) );
  AOI22_X1 U40430 ( .A1(n4455), .A2(n4298), .B1(n4347), .B2(n3250), .ZN(n3251)
         );
  OAI21_X1 U4044 ( .B1(n3564), .B2(n4277), .A(n3251), .ZN(n3252) );
  AOI21_X1 U4045 ( .B1(n3253), .B2(n3409), .A(n3252), .ZN(n3254) );
  OAI21_X1 U4046 ( .B1(n3255), .B2(n3565), .A(n3254), .ZN(n3290) );
  INV_X1 U4047 ( .A(n3290), .ZN(n3264) );
  INV_X1 U4048 ( .A(n3255), .ZN(n3291) );
  INV_X1 U4049 ( .A(n3256), .ZN(n3259) );
  INV_X1 U4050 ( .A(n3257), .ZN(n3258) );
  OAI21_X1 U4051 ( .B1(n3259), .B2(n3340), .A(n3258), .ZN(n3296) );
  INV_X1 U4052 ( .A(n3260), .ZN(n3342) );
  AOI22_X1 U4053 ( .A1(n4479), .A2(REG2_REG_13__SCAN_IN), .B1(n3342), .B2(
        n4619), .ZN(n3261) );
  OAI21_X1 U4054 ( .B1(n3296), .B2(n4335), .A(n3261), .ZN(n3262) );
  AOI21_X1 U4055 ( .B1(n3291), .B2(n4622), .A(n3262), .ZN(n3263) );
  OAI21_X1 U4056 ( .B1(n3264), .B2(n4479), .A(n3263), .ZN(U3277) );
  NOR2_X1 U4057 ( .A1(n4155), .A2(n3311), .ZN(n3265) );
  AOI21_X1 U4058 ( .B1(n4479), .B2(REG2_REG_12__SCAN_IN), .A(n3265), .ZN(n3266) );
  OAI21_X1 U4059 ( .B1(n3267), .B2(n4335), .A(n3266), .ZN(n3268) );
  AOI21_X1 U4060 ( .B1(n3269), .B2(n3288), .A(n3268), .ZN(n3270) );
  OAI21_X1 U4061 ( .B1(n4479), .B2(n3271), .A(n3270), .ZN(U3278) );
  NAND2_X1 U4062 ( .A1(n3789), .A2(n3794), .ZN(n3734) );
  XOR2_X1 U4063 ( .A(n3734), .B(n3272), .Z(n3277) );
  AOI22_X1 U4064 ( .A1(n3851), .A2(n4298), .B1(n4347), .B2(n3273), .ZN(n3274)
         );
  OAI21_X1 U4065 ( .B1(n3275), .B2(n4277), .A(n3274), .ZN(n3276) );
  AOI21_X1 U4066 ( .B1(n3277), .B2(n3409), .A(n3276), .ZN(n4691) );
  NAND2_X1 U4067 ( .A1(n4686), .A2(n3278), .ZN(n3280) );
  AND2_X1 U4068 ( .A1(n3280), .A2(n3279), .ZN(n3281) );
  XOR2_X1 U4069 ( .A(n3734), .B(n3281), .Z(n4695) );
  OAI21_X1 U4070 ( .B1(n2107), .B2(n3284), .A(n3283), .ZN(n4692) );
  NOR2_X1 U4071 ( .A1(n4692), .A2(n4335), .ZN(n3287) );
  INV_X1 U4072 ( .A(REG2_REG_9__SCAN_IN), .ZN(n4096) );
  OAI22_X1 U4073 ( .A1(n3575), .A2(n4096), .B1(n3285), .B2(n4155), .ZN(n3286)
         );
  AOI211_X1 U4074 ( .C1(n4695), .C2(n3288), .A(n3287), .B(n3286), .ZN(n3289)
         );
  OAI21_X1 U4075 ( .B1(n4479), .B2(n4691), .A(n3289), .ZN(U3281) );
  AOI21_X1 U4076 ( .B1(n4675), .B2(n3291), .A(n3290), .ZN(n3293) );
  MUX2_X1 U4077 ( .A(n4078), .B(n3293), .S(n4716), .Z(n3292) );
  OAI21_X1 U4078 ( .B1(n4392), .B2(n3296), .A(n3292), .ZN(U3531) );
  INV_X1 U4079 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3294) );
  MUX2_X1 U4080 ( .A(n3294), .B(n3293), .S(n4705), .Z(n3295) );
  OAI21_X1 U4081 ( .B1(n3296), .B2(n4435), .A(n3295), .ZN(U3493) );
  NAND2_X1 U4082 ( .A1(n3298), .A2(n3297), .ZN(n3300) );
  NAND2_X1 U4083 ( .A1(n3300), .A2(n3299), .ZN(n3326) );
  OAI22_X1 U4084 ( .A1(n3564), .A2(n3540), .B1(n2056), .B2(n3304), .ZN(n3301)
         );
  XNOR2_X1 U4085 ( .A(n3301), .B(n3546), .ZN(n3325) );
  OAI22_X1 U4086 ( .A1(n3564), .A2(n3525), .B1(n3540), .B2(n3304), .ZN(n3324)
         );
  XNOR2_X1 U4087 ( .A(n3325), .B(n3324), .ZN(n3302) );
  XNOR2_X1 U4088 ( .A(n3326), .B(n3302), .ZN(n3303) );
  NAND2_X1 U4089 ( .A1(n3303), .A2(n3665), .ZN(n3310) );
  OAI22_X1 U4090 ( .A1(n4460), .A2(n3304), .B1(n3389), .B2(n3677), .ZN(n3308)
         );
  INV_X1 U4091 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4010) );
  NOR2_X1 U4092 ( .A1(n4010), .A2(STATE_REG_SCAN_IN), .ZN(n4538) );
  INV_X1 U4093 ( .A(n4538), .ZN(n3305) );
  OAI21_X1 U4094 ( .B1(n3675), .B2(n3306), .A(n3305), .ZN(n3307) );
  NOR2_X1 U4095 ( .A1(n3308), .A2(n3307), .ZN(n3309) );
  OAI211_X1 U4096 ( .C1(n4472), .C2(n3311), .A(n3310), .B(n3309), .ZN(U3221)
         );
  XNOR2_X1 U4097 ( .A(n3312), .B(n3752), .ZN(n3346) );
  INV_X1 U4098 ( .A(n3346), .ZN(n3323) );
  NAND2_X1 U4099 ( .A1(n3313), .A2(n3683), .ZN(n3314) );
  XNOR2_X1 U4100 ( .A(n3314), .B(n3752), .ZN(n3317) );
  OAI22_X1 U4101 ( .A1(n3420), .A2(n4321), .B1(n4459), .B2(n4320), .ZN(n3315)
         );
  AOI21_X1 U4102 ( .B1(n4325), .B2(n4455), .A(n3315), .ZN(n3316) );
  OAI21_X1 U4103 ( .B1(n3317), .B2(n4327), .A(n3316), .ZN(n3345) );
  OAI21_X1 U4104 ( .B1(n3318), .B2(n4459), .A(n3366), .ZN(n3351) );
  NOR2_X1 U4105 ( .A1(n3351), .A2(n4335), .ZN(n3321) );
  INV_X1 U4106 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3319) );
  OAI22_X1 U4107 ( .A1(n3575), .A2(n3319), .B1(n4471), .B2(n4155), .ZN(n3320)
         );
  AOI211_X1 U4108 ( .C1(n3345), .C2(n3575), .A(n3321), .B(n3320), .ZN(n3322)
         );
  OAI21_X1 U4109 ( .B1(n3323), .B2(n4338), .A(n3322), .ZN(U3275) );
  OAI21_X1 U4110 ( .B1(n3326), .B2(n3325), .A(n3324), .ZN(n3328) );
  NAND2_X1 U4111 ( .A1(n3326), .A2(n3325), .ZN(n3327) );
  OAI22_X1 U4112 ( .A1(n3389), .A2(n3540), .B1(n2056), .B2(n3340), .ZN(n3329)
         );
  XNOR2_X1 U4113 ( .A(n3329), .B(n3546), .ZN(n3333) );
  INV_X1 U4114 ( .A(n3333), .ZN(n3331) );
  OAI22_X1 U4115 ( .A1(n3389), .A2(n3525), .B1(n3540), .B2(n3340), .ZN(n3332)
         );
  INV_X1 U4116 ( .A(n3332), .ZN(n3330) );
  NAND2_X1 U4117 ( .A1(n3331), .A2(n3330), .ZN(n3381) );
  INV_X1 U4118 ( .A(n3381), .ZN(n3334) );
  AND2_X1 U4119 ( .A1(n3333), .A2(n3332), .ZN(n3382) );
  NOR2_X1 U4120 ( .A1(n3334), .A2(n3382), .ZN(n3335) );
  XNOR2_X1 U4121 ( .A(n3383), .B(n3335), .ZN(n3344) );
  INV_X1 U4122 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3336) );
  NOR2_X1 U4123 ( .A1(STATE_REG_SCAN_IN), .A2(n3336), .ZN(n4548) );
  AOI21_X1 U4124 ( .B1(n4456), .B2(n3337), .A(n4548), .ZN(n3339) );
  NAND2_X1 U4125 ( .A1(n4454), .A2(n4455), .ZN(n3338) );
  OAI211_X1 U4126 ( .C1(n4460), .C2(n3340), .A(n3339), .B(n3338), .ZN(n3341)
         );
  AOI21_X1 U4127 ( .B1(n3680), .B2(n3342), .A(n3341), .ZN(n3343) );
  OAI21_X1 U4128 ( .B1(n3344), .B2(n4465), .A(n3343), .ZN(U3231) );
  INV_X1 U4129 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3347) );
  AOI21_X1 U4130 ( .B1(n3346), .B2(n4694), .A(n3345), .ZN(n3349) );
  MUX2_X1 U4131 ( .A(n3347), .B(n3349), .S(n4705), .Z(n3348) );
  OAI21_X1 U4132 ( .B1(n3351), .B2(n4435), .A(n3348), .ZN(U3497) );
  MUX2_X1 U4133 ( .A(n4082), .B(n3349), .S(n4716), .Z(n3350) );
  OAI21_X1 U4134 ( .B1(n4392), .B2(n3351), .A(n3350), .ZN(U3533) );
  INV_X1 U4135 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4039) );
  AOI21_X1 U4136 ( .B1(n4675), .B2(n3353), .A(n3352), .ZN(n3355) );
  MUX2_X1 U4137 ( .A(n4039), .B(n3355), .S(n4705), .Z(n3354) );
  OAI21_X1 U4138 ( .B1(n3357), .B2(n4435), .A(n3354), .ZN(U3495) );
  MUX2_X1 U4139 ( .A(n4559), .B(n3355), .S(n4716), .Z(n3356) );
  OAI21_X1 U4140 ( .B1(n4392), .B2(n3357), .A(n3356), .ZN(U3532) );
  AOI21_X1 U4141 ( .B1(n3755), .B2(n3359), .A(n3358), .ZN(n3360) );
  INV_X1 U4142 ( .A(n3360), .ZN(n4401) );
  XOR2_X1 U4143 ( .A(n3755), .B(n3361), .Z(n3364) );
  AOI22_X1 U4144 ( .A1(n3847), .A2(n4298), .B1(n4347), .B2(n3365), .ZN(n3362)
         );
  OAI21_X1 U4145 ( .B1(n3433), .B2(n4277), .A(n3362), .ZN(n3363) );
  AOI21_X1 U4146 ( .B1(n3364), .B2(n3409), .A(n3363), .ZN(n4400) );
  INV_X1 U4147 ( .A(n4400), .ZN(n3370) );
  NAND2_X1 U4148 ( .A1(n3366), .A2(n3365), .ZN(n4397) );
  AND3_X1 U4149 ( .A1(n4398), .A2(n4624), .A3(n4397), .ZN(n3369) );
  INV_X1 U4150 ( .A(REG2_REG_16__SCAN_IN), .ZN(n3367) );
  OAI22_X1 U4151 ( .A1(n3575), .A2(n3367), .B1(n3440), .B2(n4155), .ZN(n3368)
         );
  AOI211_X1 U4152 ( .C1(n3370), .C2(n3575), .A(n3369), .B(n3368), .ZN(n3371)
         );
  OAI21_X1 U4153 ( .B1(n4401), .B2(n4338), .A(n3371), .ZN(U3274) );
  NAND2_X1 U4154 ( .A1(n3407), .A2(n3404), .ZN(n3743) );
  XNOR2_X1 U4155 ( .A(n3372), .B(n3743), .ZN(n3396) );
  INV_X1 U4156 ( .A(n3396), .ZN(n3380) );
  XOR2_X1 U4157 ( .A(n3743), .B(n3406), .Z(n3375) );
  OAI22_X1 U4158 ( .A1(n3614), .A2(n4321), .B1(n4320), .B2(n3458), .ZN(n3373)
         );
  AOI21_X1 U4159 ( .B1(n4325), .B2(n4453), .A(n3373), .ZN(n3374) );
  OAI21_X1 U4160 ( .B1(n3375), .B2(n4327), .A(n3374), .ZN(n3395) );
  OAI21_X1 U4161 ( .B1(n2111), .B2(n3458), .A(n2062), .ZN(n3401) );
  INV_X1 U4162 ( .A(n3376), .ZN(n3460) );
  AOI22_X1 U4163 ( .A1(n4479), .A2(REG2_REG_17__SCAN_IN), .B1(n3460), .B2(
        n4619), .ZN(n3377) );
  OAI21_X1 U4164 ( .B1(n3401), .B2(n4335), .A(n3377), .ZN(n3378) );
  AOI21_X1 U4165 ( .B1(n3395), .B2(n3575), .A(n3378), .ZN(n3379) );
  OAI21_X1 U4166 ( .B1(n3380), .B2(n4338), .A(n3379), .ZN(U3273) );
  OAI21_X2 U4167 ( .B1(n3383), .B2(n3382), .A(n3381), .ZN(n3423) );
  OAI22_X1 U4168 ( .A1(n3385), .A2(n3540), .B1(n2056), .B2(n3388), .ZN(n3384)
         );
  XNOR2_X1 U4169 ( .A(n3384), .B(n3538), .ZN(n3424) );
  XNOR2_X1 U4170 ( .A(n3424), .B(n3422), .ZN(n3386) );
  XNOR2_X1 U4171 ( .A(n3423), .B(n3386), .ZN(n3387) );
  NAND2_X1 U4172 ( .A1(n3387), .A2(n3665), .ZN(n3393) );
  OAI22_X1 U4173 ( .A1(n4460), .A2(n3388), .B1(n3433), .B2(n3677), .ZN(n3391)
         );
  NAND2_X1 U4174 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4567) );
  OAI21_X1 U4175 ( .B1(n3675), .B2(n3389), .A(n4567), .ZN(n3390) );
  NOR2_X1 U4176 ( .A1(n3391), .A2(n3390), .ZN(n3392) );
  OAI211_X1 U4177 ( .C1(n4472), .C2(n3394), .A(n3393), .B(n3392), .ZN(U3212)
         );
  INV_X1 U4178 ( .A(REG0_REG_17__SCAN_IN), .ZN(n3397) );
  AOI21_X1 U4179 ( .B1(n3396), .B2(n4694), .A(n3395), .ZN(n3399) );
  MUX2_X1 U4180 ( .A(n3397), .B(n3399), .S(n4705), .Z(n3398) );
  OAI21_X1 U4181 ( .B1(n3401), .B2(n4435), .A(n3398), .ZN(U3501) );
  MUX2_X1 U4182 ( .A(n4118), .B(n3399), .S(n4716), .Z(n3400) );
  OAI21_X1 U4183 ( .B1(n4392), .B2(n3401), .A(n3400), .ZN(U3535) );
  OAI21_X1 U4184 ( .B1(n3403), .B2(n3729), .A(n3402), .ZN(n4395) );
  INV_X1 U4185 ( .A(n4395), .ZN(n3419) );
  INV_X1 U4186 ( .A(n3404), .ZN(n3405) );
  INV_X1 U4187 ( .A(n3407), .ZN(n3408) );
  NOR2_X1 U4188 ( .A1(n4233), .A2(n3408), .ZN(n4317) );
  XNOR2_X1 U4189 ( .A(n4317), .B(n3729), .ZN(n3410) );
  NAND2_X1 U4190 ( .A1(n3410), .A2(n3409), .ZN(n3412) );
  AOI22_X1 U4191 ( .A1(n4300), .A2(n4298), .B1(n3469), .B2(n4347), .ZN(n3411)
         );
  OAI211_X1 U4192 ( .C1(n3435), .C2(n4277), .A(n3412), .B(n3411), .ZN(n4393)
         );
  AOI211_X1 U4193 ( .C1(n3469), .C2(n2062), .A(n4698), .B(n4331), .ZN(n4394)
         );
  INV_X1 U4194 ( .A(n4394), .ZN(n3416) );
  INV_X1 U4195 ( .A(n3413), .ZN(n3484) );
  AOI22_X1 U4196 ( .A1(n4479), .A2(REG2_REG_18__SCAN_IN), .B1(n3484), .B2(
        n4619), .ZN(n3414) );
  OAI21_X1 U4197 ( .B1(n3416), .B2(n3415), .A(n3414), .ZN(n3417) );
  AOI21_X1 U4198 ( .B1(n4393), .B2(n3575), .A(n3417), .ZN(n3418) );
  OAI21_X1 U4199 ( .B1(n3419), .B2(n4338), .A(n3418), .ZN(U3272) );
  OAI22_X1 U4200 ( .A1(n3420), .A2(n3525), .B1(n3540), .B2(n3434), .ZN(n3444)
         );
  OAI22_X1 U4201 ( .A1(n3420), .A2(n3540), .B1(n2056), .B2(n3434), .ZN(n3421)
         );
  XNOR2_X1 U4202 ( .A(n3421), .B(n3546), .ZN(n3443) );
  XOR2_X1 U4203 ( .A(n3444), .B(n3443), .Z(n3441) );
  INV_X1 U4204 ( .A(n3424), .ZN(n3425) );
  OAI22_X1 U4205 ( .A1(n3433), .A2(n3540), .B1(n2056), .B2(n4459), .ZN(n3426)
         );
  XNOR2_X1 U4206 ( .A(n3426), .B(n3538), .ZN(n3428) );
  NAND2_X1 U4207 ( .A1(n3427), .A2(n3428), .ZN(n4462) );
  OAI22_X1 U4208 ( .A1(n3433), .A2(n3525), .B1(n3540), .B2(n4459), .ZN(n4463)
         );
  NAND2_X1 U4209 ( .A1(n4462), .A2(n4463), .ZN(n3442) );
  INV_X1 U4210 ( .A(n3428), .ZN(n3429) );
  NAND2_X1 U4211 ( .A1(n3442), .A2(n4464), .ZN(n3431) );
  XOR2_X1 U4212 ( .A(n3441), .B(n3431), .Z(n3432) );
  NAND2_X1 U4213 ( .A1(n3432), .A2(n3665), .ZN(n3439) );
  OAI22_X1 U4214 ( .A1(n4460), .A2(n3434), .B1(n3433), .B2(n3675), .ZN(n3437)
         );
  NAND2_X1 U4215 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4087) );
  OAI21_X1 U4216 ( .B1(n3677), .B2(n3435), .A(n4087), .ZN(n3436) );
  NOR2_X1 U4217 ( .A1(n3437), .A2(n3436), .ZN(n3438) );
  OAI211_X1 U4218 ( .C1(n4472), .C2(n3440), .A(n3439), .B(n3438), .ZN(U3223)
         );
  NAND3_X1 U4219 ( .A1(n3442), .A2(n4464), .A3(n3441), .ZN(n3448) );
  NAND2_X1 U4220 ( .A1(n3847), .A2(n2772), .ZN(n3450) );
  NAND2_X1 U4221 ( .A1(n3544), .A2(n3452), .ZN(n3449) );
  NAND2_X1 U4222 ( .A1(n3450), .A2(n3449), .ZN(n3451) );
  XNOR2_X1 U4223 ( .A(n3451), .B(n3546), .ZN(n3463) );
  NAND2_X1 U4224 ( .A1(n3545), .A2(n3847), .ZN(n3454) );
  NAND2_X1 U4225 ( .A1(n2772), .A2(n3452), .ZN(n3453) );
  NAND2_X1 U4226 ( .A1(n3454), .A2(n3453), .ZN(n3464) );
  XNOR2_X1 U4227 ( .A(n3463), .B(n3464), .ZN(n3455) );
  XNOR2_X1 U4228 ( .A(n3468), .B(n3455), .ZN(n3462) );
  AND2_X1 U4229 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4580) );
  AOI21_X1 U4230 ( .B1(n4454), .B2(n4324), .A(n4580), .ZN(n3457) );
  NAND2_X1 U4231 ( .A1(n4456), .A2(n4453), .ZN(n3456) );
  OAI211_X1 U4232 ( .C1(n4460), .C2(n3458), .A(n3457), .B(n3456), .ZN(n3459)
         );
  AOI21_X1 U4233 ( .B1(n3680), .B2(n3460), .A(n3459), .ZN(n3461) );
  OAI21_X1 U4234 ( .B1(n3462), .B2(n4465), .A(n3461), .ZN(U3225) );
  NOR2_X1 U4235 ( .A1(n3463), .A2(n3464), .ZN(n3467) );
  INV_X1 U4236 ( .A(n3463), .ZN(n3466) );
  INV_X1 U4237 ( .A(n3464), .ZN(n3465) );
  NAND2_X1 U4238 ( .A1(n4324), .A2(n2772), .ZN(n3471) );
  NAND2_X1 U4239 ( .A1(n3544), .A2(n3469), .ZN(n3470) );
  NAND2_X1 U4240 ( .A1(n3471), .A2(n3470), .ZN(n3472) );
  XNOR2_X1 U4241 ( .A(n3472), .B(n3538), .ZN(n3476) );
  NOR2_X1 U4242 ( .A1(n3540), .A2(n3482), .ZN(n3474) );
  AOI21_X1 U4243 ( .B1(n3545), .B2(n4324), .A(n3474), .ZN(n3475) );
  NOR2_X1 U4244 ( .A1(n3476), .A2(n3475), .ZN(n3488) );
  NAND2_X1 U4245 ( .A1(n3476), .A2(n3475), .ZN(n3487) );
  INV_X1 U4246 ( .A(n3487), .ZN(n3477) );
  NOR2_X1 U4247 ( .A1(n3488), .A2(n3477), .ZN(n3478) );
  XNOR2_X1 U4248 ( .A(n3489), .B(n3478), .ZN(n3486) );
  INV_X1 U4249 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3479) );
  NOR2_X1 U4250 ( .A1(STATE_REG_SCAN_IN), .A2(n3479), .ZN(n4598) );
  AOI21_X1 U4251 ( .B1(n4454), .B2(n4300), .A(n4598), .ZN(n3481) );
  NAND2_X1 U4252 ( .A1(n4456), .A2(n3847), .ZN(n3480) );
  OAI211_X1 U4253 ( .C1(n4460), .C2(n3482), .A(n3481), .B(n3480), .ZN(n3483)
         );
  AOI21_X1 U4254 ( .B1(n3680), .B2(n3484), .A(n3483), .ZN(n3485) );
  OAI21_X1 U4255 ( .B1(n3486), .B2(n4465), .A(n3485), .ZN(U3235) );
  OAI22_X1 U4256 ( .A1(n3658), .A2(n3525), .B1(n3540), .B2(n4330), .ZN(n3495)
         );
  NAND2_X1 U4257 ( .A1(n4300), .A2(n2772), .ZN(n3492) );
  NAND2_X1 U4258 ( .A1(n3544), .A2(n3490), .ZN(n3491) );
  NAND2_X1 U4259 ( .A1(n3492), .A2(n3491), .ZN(n3493) );
  XNOR2_X1 U4260 ( .A(n3493), .B(n3546), .ZN(n3494) );
  XOR2_X1 U4261 ( .A(n3495), .B(n3494), .Z(n3611) );
  INV_X1 U4262 ( .A(n3494), .ZN(n3497) );
  INV_X1 U4263 ( .A(n3495), .ZN(n3496) );
  NOR2_X1 U4264 ( .A1(n2056), .A2(n4305), .ZN(n3498) );
  AOI21_X1 U4265 ( .B1(n3846), .B2(n2772), .A(n3498), .ZN(n3499) );
  XNOR2_X1 U4266 ( .A(n3499), .B(n3546), .ZN(n3502) );
  NOR2_X1 U4267 ( .A1(n3540), .A2(n4305), .ZN(n3500) );
  AOI21_X1 U4268 ( .B1(n3846), .B2(n3545), .A(n3500), .ZN(n3501) );
  NOR2_X1 U4269 ( .A1(n3502), .A2(n3501), .ZN(n3654) );
  NAND2_X1 U4270 ( .A1(n4299), .A2(n2772), .ZN(n3504) );
  OR2_X1 U4271 ( .A1(n2056), .A2(n4283), .ZN(n3503) );
  NAND2_X1 U4272 ( .A1(n3504), .A2(n3503), .ZN(n3505) );
  XNOR2_X1 U4273 ( .A(n3505), .B(n3538), .ZN(n3621) );
  NOR2_X1 U4274 ( .A1(n3540), .A2(n4283), .ZN(n3506) );
  AOI21_X1 U4275 ( .B1(n4299), .B2(n3545), .A(n3506), .ZN(n3620) );
  NAND2_X1 U4276 ( .A1(n3621), .A2(n3620), .ZN(n3509) );
  INV_X1 U4277 ( .A(n3621), .ZN(n3508) );
  INV_X1 U4278 ( .A(n3620), .ZN(n3507) );
  OAI22_X1 U4279 ( .A1(n4240), .A2(n3525), .B1(n3540), .B2(n4267), .ZN(n3513)
         );
  OAI22_X1 U4280 ( .A1(n4240), .A2(n3540), .B1(n2056), .B2(n4267), .ZN(n3510)
         );
  XNOR2_X1 U4281 ( .A(n3510), .B(n3546), .ZN(n3512) );
  XOR2_X1 U4282 ( .A(n3513), .B(n3512), .Z(n3664) );
  OAI22_X1 U4283 ( .A1(n4218), .A2(n3540), .B1(n2056), .B2(n4246), .ZN(n3511)
         );
  XNOR2_X1 U4284 ( .A(n3511), .B(n3538), .ZN(n3518) );
  OAI22_X1 U4285 ( .A1(n4218), .A2(n3525), .B1(n3540), .B2(n4246), .ZN(n3519)
         );
  XNOR2_X1 U4286 ( .A(n3518), .B(n3519), .ZN(n3600) );
  INV_X1 U4287 ( .A(n3512), .ZN(n3515) );
  INV_X1 U4288 ( .A(n3513), .ZN(n3514) );
  NAND2_X1 U4289 ( .A1(n3515), .A2(n3514), .ZN(n3601) );
  NAND2_X2 U4290 ( .A1(n3599), .A2(n3516), .ZN(n3598) );
  NOR2_X1 U4291 ( .A1(n2797), .A2(n4224), .ZN(n3517) );
  AOI21_X1 U4292 ( .B1(n4242), .B2(n3545), .A(n3517), .ZN(n3522) );
  INV_X1 U4293 ( .A(n3518), .ZN(n3520) );
  NAND2_X1 U4294 ( .A1(n3520), .A2(n3519), .ZN(n3523) );
  OAI22_X1 U4295 ( .A1(n4202), .A2(n2797), .B1(n2056), .B2(n4224), .ZN(n3521)
         );
  XNOR2_X1 U4296 ( .A(n3521), .B(n3546), .ZN(n3643) );
  OAI22_X1 U4297 ( .A1(n4182), .A2(n3540), .B1(n2056), .B2(n4201), .ZN(n3524)
         );
  XNOR2_X1 U4298 ( .A(n3524), .B(n3546), .ZN(n3527) );
  OAI22_X1 U4299 ( .A1(n4182), .A2(n3525), .B1(n3540), .B2(n4201), .ZN(n3526)
         );
  NOR2_X1 U4300 ( .A1(n3527), .A2(n3526), .ZN(n3629) );
  NAND2_X1 U4301 ( .A1(n3527), .A2(n3526), .ZN(n3630) );
  NAND2_X1 U4302 ( .A1(n4204), .A2(n2772), .ZN(n3529) );
  OR2_X1 U4303 ( .A1(n2056), .A2(n4189), .ZN(n3528) );
  NAND2_X1 U4304 ( .A1(n3529), .A2(n3528), .ZN(n3530) );
  XNOR2_X1 U4305 ( .A(n3530), .B(n3538), .ZN(n3533) );
  NOR2_X1 U4306 ( .A1(n3540), .A2(n4189), .ZN(n3531) );
  AOI21_X1 U4307 ( .B1(n4204), .B2(n3545), .A(n3531), .ZN(n3532) );
  NOR2_X1 U4308 ( .A1(n3533), .A2(n3532), .ZN(n3671) );
  NAND2_X1 U4309 ( .A1(n4184), .A2(n2772), .ZN(n3537) );
  OR2_X1 U4310 ( .A1(n2056), .A2(n4171), .ZN(n3536) );
  NAND2_X1 U4311 ( .A1(n3537), .A2(n3536), .ZN(n3539) );
  XNOR2_X1 U4312 ( .A(n3539), .B(n3538), .ZN(n3542) );
  NOR2_X1 U4313 ( .A1(n2797), .A2(n4171), .ZN(n3541) );
  AOI21_X1 U4314 ( .B1(n4184), .B2(n3545), .A(n3541), .ZN(n3543) );
  XNOR2_X1 U4315 ( .A(n3542), .B(n3543), .ZN(n3589) );
  AOI22_X1 U4316 ( .A1(n4169), .A2(n2772), .B1(n3544), .B2(n4137), .ZN(n3549)
         );
  AOI22_X1 U4317 ( .A1(n4169), .A2(n3545), .B1(n2772), .B2(n4137), .ZN(n3547)
         );
  XNOR2_X1 U4318 ( .A(n3547), .B(n3546), .ZN(n3548) );
  XOR2_X1 U4319 ( .A(n3549), .B(n3548), .Z(n3550) );
  XNOR2_X1 U4320 ( .A(n3551), .B(n3550), .ZN(n3558) );
  INV_X1 U4321 ( .A(n4184), .ZN(n3823) );
  OAI22_X1 U4322 ( .A1(n3823), .A2(n3675), .B1(n4460), .B2(n3552), .ZN(n3556)
         );
  OAI22_X1 U4323 ( .A1(n3554), .A2(n3677), .B1(STATE_REG_SCAN_IN), .B2(n3553), 
        .ZN(n3555) );
  AOI211_X1 U4324 ( .C1(n3582), .C2(n3680), .A(n3556), .B(n3555), .ZN(n3557)
         );
  OAI21_X1 U4325 ( .B1(n3558), .B2(n4465), .A(n3557), .ZN(U3217) );
  INV_X1 U4326 ( .A(n3559), .ZN(n3560) );
  AOI21_X1 U4327 ( .B1(n3562), .B2(n3561), .A(n3560), .ZN(n4700) );
  INV_X1 U4328 ( .A(n3562), .ZN(n3731) );
  XNOR2_X1 U4329 ( .A(n3563), .B(n3731), .ZN(n3569) );
  OAI22_X1 U4330 ( .A1(n3564), .A2(n4321), .B1(n4320), .B2(n3571), .ZN(n3567)
         );
  NOR2_X1 U4331 ( .A1(n4700), .A2(n3565), .ZN(n3566) );
  AOI211_X1 U4332 ( .C1(n4325), .C2(n3851), .A(n3567), .B(n3566), .ZN(n3568)
         );
  OAI21_X1 U4333 ( .B1(n4327), .B2(n3569), .A(n3568), .ZN(n4702) );
  NAND2_X1 U4334 ( .A1(n4702), .A2(n3575), .ZN(n3579) );
  OAI21_X1 U4335 ( .B1(n3572), .B2(n3571), .A(n3570), .ZN(n4697) );
  INV_X1 U4336 ( .A(n4697), .ZN(n3577) );
  INV_X1 U4337 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3574) );
  OAI22_X1 U4338 ( .A1(n3575), .A2(n3574), .B1(n3573), .B2(n4155), .ZN(n3576)
         );
  AOI21_X1 U4339 ( .B1(n3577), .B2(n4624), .A(n3576), .ZN(n3578) );
  OAI211_X1 U4340 ( .C1(n4700), .C2(n3580), .A(n3579), .B(n3578), .ZN(U3279)
         );
  INV_X1 U4341 ( .A(n3581), .ZN(n3586) );
  AOI22_X1 U4342 ( .A1(n3582), .A2(n4619), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4479), .ZN(n3583) );
  OAI21_X1 U4343 ( .B1(n3584), .B2(n4335), .A(n3583), .ZN(n3585) );
  AOI21_X1 U4344 ( .B1(n3586), .B2(n3575), .A(n3585), .ZN(n3587) );
  OAI21_X1 U4345 ( .B1(n3588), .B2(n4338), .A(n3587), .ZN(U3262) );
  XNOR2_X1 U4346 ( .A(n3590), .B(n3589), .ZN(n3597) );
  INV_X1 U4347 ( .A(n3591), .ZN(n4172) );
  OAI22_X1 U4348 ( .A1(n4162), .A2(n3675), .B1(STATE_REG_SCAN_IN), .B2(n3592), 
        .ZN(n3595) );
  INV_X1 U4349 ( .A(n4169), .ZN(n3593) );
  OAI22_X1 U4350 ( .A1(n3593), .A2(n3677), .B1(n4460), .B2(n4171), .ZN(n3594)
         );
  AOI211_X1 U4351 ( .C1(n4172), .C2(n3680), .A(n3595), .B(n3594), .ZN(n3596)
         );
  OAI21_X1 U4352 ( .B1(n3597), .B2(n4465), .A(n3596), .ZN(U3211) );
  INV_X1 U4353 ( .A(n3598), .ZN(n3603) );
  AOI21_X1 U4354 ( .B1(n3599), .B2(n3601), .A(n3600), .ZN(n3602) );
  NOR3_X1 U4355 ( .A1(n3603), .A2(n3602), .A3(n4465), .ZN(n3610) );
  AOI22_X1 U4356 ( .A1(n3645), .A2(n3604), .B1(n4454), .B2(n4242), .ZN(n3608)
         );
  OAI22_X1 U4357 ( .A1(n3675), .A2(n4240), .B1(STATE_REG_SCAN_IN), .B2(n3605), 
        .ZN(n3606) );
  INV_X1 U4358 ( .A(n3606), .ZN(n3607) );
  OAI211_X1 U4359 ( .C1(n4472), .C2(n4248), .A(n3608), .B(n3607), .ZN(n3609)
         );
  OR2_X1 U4360 ( .A1(n3610), .A2(n3609), .ZN(U3213) );
  XNOR2_X1 U4361 ( .A(n3612), .B(n3611), .ZN(n3613) );
  NAND2_X1 U4362 ( .A1(n3613), .A2(n3665), .ZN(n3618) );
  OAI22_X1 U4363 ( .A1(n4460), .A2(n4330), .B1(n4322), .B2(n3677), .ZN(n3616)
         );
  NAND2_X1 U4364 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4131) );
  OAI21_X1 U4365 ( .B1(n3675), .B2(n3614), .A(n4131), .ZN(n3615) );
  NOR2_X1 U4366 ( .A1(n3616), .A2(n3615), .ZN(n3617) );
  OAI211_X1 U4367 ( .C1(n4472), .C2(n4332), .A(n3618), .B(n3617), .ZN(U3216)
         );
  XNOR2_X1 U4368 ( .A(n3621), .B(n3620), .ZN(n3622) );
  XNOR2_X1 U4369 ( .A(n3619), .B(n3622), .ZN(n3623) );
  NAND2_X1 U4370 ( .A1(n3623), .A2(n3665), .ZN(n3628) );
  OAI22_X1 U4371 ( .A1(n4460), .A2(n4283), .B1(n4240), .B2(n3677), .ZN(n3626)
         );
  INV_X1 U4372 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3624) );
  OAI22_X1 U4373 ( .A1(n3675), .A2(n4322), .B1(STATE_REG_SCAN_IN), .B2(n3624), 
        .ZN(n3625) );
  NOR2_X1 U4374 ( .A1(n3626), .A2(n3625), .ZN(n3627) );
  OAI211_X1 U4375 ( .C1(n4472), .C2(n4285), .A(n3628), .B(n3627), .ZN(U3220)
         );
  INV_X1 U4376 ( .A(n3629), .ZN(n3631) );
  NAND2_X1 U4377 ( .A1(n3631), .A2(n3630), .ZN(n3632) );
  XNOR2_X1 U4378 ( .A(n3633), .B(n3632), .ZN(n3639) );
  INV_X1 U4379 ( .A(n3634), .ZN(n4209) );
  INV_X1 U4380 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3635) );
  OAI22_X1 U4381 ( .A1(n4202), .A2(n3675), .B1(STATE_REG_SCAN_IN), .B2(n3635), 
        .ZN(n3637) );
  OAI22_X1 U4382 ( .A1(n4162), .A2(n3677), .B1(n4460), .B2(n4201), .ZN(n3636)
         );
  AOI211_X1 U4383 ( .C1(n4209), .C2(n3680), .A(n3637), .B(n3636), .ZN(n3638)
         );
  OAI21_X1 U4384 ( .B1(n3639), .B2(n4465), .A(n3638), .ZN(U3222) );
  INV_X1 U4385 ( .A(n3641), .ZN(n3642) );
  NOR2_X1 U4386 ( .A1(n3640), .A2(n3642), .ZN(n3644) );
  XNOR2_X1 U4387 ( .A(n3644), .B(n3643), .ZN(n3652) );
  AOI22_X1 U4388 ( .A1(n3645), .A2(n4196), .B1(n4220), .B2(n4454), .ZN(n3649)
         );
  OAI22_X1 U4389 ( .A1(n3675), .A2(n4218), .B1(STATE_REG_SCAN_IN), .B2(n3646), 
        .ZN(n3647) );
  INV_X1 U4390 ( .A(n3647), .ZN(n3648) );
  OAI211_X1 U4391 ( .C1(n4472), .C2(n4225), .A(n3649), .B(n3648), .ZN(n3650)
         );
  INV_X1 U4392 ( .A(n3650), .ZN(n3651) );
  OAI21_X1 U4393 ( .B1(n3652), .B2(n4465), .A(n3651), .ZN(U3226) );
  OAI21_X1 U4394 ( .B1(n3656), .B2(n3654), .A(n3653), .ZN(n3655) );
  OAI21_X1 U4395 ( .B1(n2071), .B2(n3656), .A(n3655), .ZN(n3657) );
  NAND2_X1 U4396 ( .A1(n3657), .A2(n3665), .ZN(n3662) );
  OAI22_X1 U4397 ( .A1(n4460), .A2(n4305), .B1(n4256), .B2(n3677), .ZN(n3660)
         );
  OAI22_X1 U4398 ( .A1(n3675), .A2(n3658), .B1(STATE_REG_SCAN_IN), .B2(n4047), 
        .ZN(n3659) );
  NOR2_X1 U4399 ( .A1(n3660), .A2(n3659), .ZN(n3661) );
  OAI211_X1 U4400 ( .C1(n4472), .C2(n4307), .A(n3662), .B(n3661), .ZN(U3230)
         );
  OAI21_X1 U4401 ( .B1(n3664), .B2(n3663), .A(n3599), .ZN(n3666) );
  NAND2_X1 U4402 ( .A1(n3666), .A2(n3665), .ZN(n3670) );
  OAI22_X1 U4403 ( .A1(n4460), .A2(n4267), .B1(n4218), .B2(n3677), .ZN(n3668)
         );
  INV_X1 U4404 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4026) );
  OAI22_X1 U4405 ( .A1(n3675), .A2(n4256), .B1(STATE_REG_SCAN_IN), .B2(n4026), 
        .ZN(n3667) );
  NOR2_X1 U4406 ( .A1(n3668), .A2(n3667), .ZN(n3669) );
  OAI211_X1 U4407 ( .C1(n4472), .C2(n4264), .A(n3670), .B(n3669), .ZN(U3232)
         );
  NOR2_X1 U4408 ( .A1(n3671), .A2(n2088), .ZN(n3672) );
  XNOR2_X1 U4409 ( .A(n3673), .B(n3672), .ZN(n3682) );
  INV_X1 U4410 ( .A(n3674), .ZN(n4190) );
  OAI22_X1 U4411 ( .A1(n4182), .A2(n3675), .B1(n4460), .B2(n4189), .ZN(n3679)
         );
  INV_X1 U4412 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3676) );
  OAI22_X1 U4413 ( .A1(n3823), .A2(n3677), .B1(STATE_REG_SCAN_IN), .B2(n3676), 
        .ZN(n3678) );
  AOI211_X1 U4414 ( .C1(n4190), .C2(n3680), .A(n3679), .B(n3678), .ZN(n3681)
         );
  OAI21_X1 U4415 ( .B1(n3682), .B2(n4465), .A(n3681), .ZN(U3237) );
  NAND2_X1 U4416 ( .A1(n3683), .A2(n3686), .ZN(n3807) );
  NAND2_X1 U4417 ( .A1(n3685), .A2(n3684), .ZN(n3792) );
  NAND2_X1 U4418 ( .A1(n3792), .A2(n3686), .ZN(n3806) );
  OAI21_X1 U4419 ( .B1(n3687), .B2(n3807), .A(n3806), .ZN(n3688) );
  NAND2_X1 U4420 ( .A1(n3688), .A2(n3811), .ZN(n3689) );
  NAND2_X1 U4421 ( .A1(n3689), .A2(n3813), .ZN(n3691) );
  OAI21_X1 U4422 ( .B1(n3816), .B2(n3691), .A(n3690), .ZN(n3692) );
  AOI211_X1 U4423 ( .C1(n3821), .C2(n3692), .A(n4237), .B(n3818), .ZN(n3706)
         );
  OAI211_X1 U4424 ( .C1(n3695), .C2(n3818), .A(n3694), .B(n3693), .ZN(n3825)
         );
  AND2_X1 U4425 ( .A1(n2058), .A2(DATAI_30_), .ZN(n4348) );
  NAND2_X1 U4426 ( .A1(n2235), .A2(REG2_REG_31__SCAN_IN), .ZN(n3701) );
  NAND2_X1 U4427 ( .A1(n3696), .A2(REG0_REG_31__SCAN_IN), .ZN(n3700) );
  INV_X1 U4428 ( .A(REG1_REG_31__SCAN_IN), .ZN(n3697) );
  OR2_X1 U4429 ( .A1(n3698), .A2(n3697), .ZN(n3699) );
  AND3_X1 U4430 ( .A1(n3701), .A2(n3700), .A3(n3699), .ZN(n4341) );
  INV_X1 U4431 ( .A(n4341), .ZN(n3843) );
  AND2_X1 U4432 ( .A1(n2059), .A2(DATAI_31_), .ZN(n4342) );
  INV_X1 U4433 ( .A(n4342), .ZN(n3713) );
  AND2_X1 U4434 ( .A1(n3843), .A2(n3713), .ZN(n3831) );
  AOI21_X1 U4435 ( .B1(n4148), .B2(n4348), .A(n3831), .ZN(n3740) );
  NAND2_X1 U4436 ( .A1(n2059), .A2(DATAI_29_), .ZN(n4147) );
  OR2_X1 U4437 ( .A1(n3844), .A2(n4147), .ZN(n3737) );
  INV_X1 U4438 ( .A(n3737), .ZN(n3704) );
  NOR4_X1 U4439 ( .A1(n3704), .A2(n4149), .A3(n3708), .A4(n3703), .ZN(n3705)
         );
  OAI211_X1 U4440 ( .C1(n3706), .C2(n3825), .A(n3740), .B(n3705), .ZN(n3715)
         );
  NOR2_X1 U4441 ( .A1(n4148), .A2(n4348), .ZN(n3739) );
  OR2_X1 U4442 ( .A1(n3739), .A2(n4341), .ZN(n3712) );
  AND2_X1 U4443 ( .A1(n3844), .A2(n4147), .ZN(n3736) );
  NOR3_X1 U4444 ( .A1(n3736), .A2(n4151), .A3(n3707), .ZN(n3829) );
  NOR2_X1 U4445 ( .A1(n4149), .A2(n3708), .ZN(n3710) );
  OR2_X1 U4446 ( .A1(n3736), .A2(n4151), .ZN(n3709) );
  OAI211_X1 U4447 ( .C1(n3710), .C2(n3709), .A(n3740), .B(n3737), .ZN(n3832)
         );
  AOI21_X1 U4448 ( .B1(n3741), .B2(n3829), .A(n3832), .ZN(n3711) );
  AOI21_X1 U4449 ( .B1(n4342), .B2(n3712), .A(n3711), .ZN(n3714) );
  AOI22_X1 U4450 ( .A1(n3715), .A2(n3714), .B1(n4348), .B2(n3713), .ZN(n3768)
         );
  INV_X1 U4451 ( .A(n4138), .ZN(n3766) );
  NAND2_X1 U4452 ( .A1(n3716), .A2(n3821), .ZN(n4275) );
  INV_X1 U4453 ( .A(n3717), .ZN(n4214) );
  NOR2_X1 U4454 ( .A1(n3718), .A2(n4214), .ZN(n4238) );
  XNOR2_X1 U4455 ( .A(n4242), .B(n4196), .ZN(n4216) );
  INV_X1 U4456 ( .A(n3719), .ZN(n3721) );
  OR2_X1 U4457 ( .A1(n3721), .A2(n3720), .ZN(n4318) );
  INV_X1 U4458 ( .A(n4318), .ZN(n3723) );
  XNOR2_X1 U4459 ( .A(n3846), .B(n3722), .ZN(n4295) );
  NAND4_X1 U4460 ( .A1(n4238), .A2(n4216), .A3(n3723), .A4(n4295), .ZN(n3724)
         );
  NOR3_X1 U4461 ( .A1(n4258), .A2(n4275), .A3(n3724), .ZN(n3765) );
  INV_X1 U4462 ( .A(n3725), .ZN(n4179) );
  NOR2_X1 U4463 ( .A1(n4179), .A2(n3726), .ZN(n4199) );
  INV_X1 U4464 ( .A(n4199), .ZN(n3760) );
  INV_X1 U4465 ( .A(n3727), .ZN(n3730) );
  NOR4_X1 U4466 ( .A1(n3731), .A2(n3730), .A3(n3729), .A4(n3728), .ZN(n3751)
         );
  INV_X1 U4467 ( .A(n3733), .ZN(n3735) );
  NOR4_X1 U4468 ( .A1(n2629), .A2(n3735), .A3(n2628), .A4(n3734), .ZN(n3750)
         );
  INV_X1 U4469 ( .A(n3736), .ZN(n3738) );
  AOI21_X1 U4470 ( .B1(n4342), .B2(n4341), .A(n3739), .ZN(n3830) );
  NAND4_X1 U4471 ( .A1(n4153), .A2(n3741), .A3(n3740), .A4(n3830), .ZN(n3742)
         );
  NOR3_X1 U4472 ( .A1(n3743), .A2(n4659), .A3(n3742), .ZN(n3749) );
  NOR4_X1 U4473 ( .A1(n3747), .A2(n3746), .A3(n3745), .A4(n3744), .ZN(n3748)
         );
  NAND4_X1 U4474 ( .A1(n3751), .A2(n3750), .A3(n3749), .A4(n3748), .ZN(n3759)
         );
  INV_X1 U4475 ( .A(n3752), .ZN(n3753) );
  NAND4_X1 U4476 ( .A1(n3756), .A2(n3755), .A3(n3754), .A4(n3753), .ZN(n3757)
         );
  NOR4_X1 U4477 ( .A1(n3760), .A2(n3759), .A3(n3758), .A4(n3757), .ZN(n3764)
         );
  INV_X1 U4478 ( .A(n3761), .ZN(n3763) );
  NAND2_X1 U4479 ( .A1(n3763), .A2(n3762), .ZN(n4180) );
  NAND4_X1 U4480 ( .A1(n3766), .A2(n3765), .A3(n3764), .A4(n4180), .ZN(n3767)
         );
  MUX2_X1 U4481 ( .A(n3768), .B(n3767), .S(n2627), .Z(n3836) );
  OAI211_X1 U4482 ( .C1(n3772), .C2(n3771), .A(n3770), .B(n3769), .ZN(n3775)
         );
  NAND3_X1 U4483 ( .A1(n3775), .A2(n3774), .A3(n3773), .ZN(n3778) );
  NAND3_X1 U4484 ( .A1(n3778), .A2(n3777), .A3(n3776), .ZN(n3781) );
  NAND3_X1 U4485 ( .A1(n3781), .A2(n3780), .A3(n3779), .ZN(n3784) );
  NAND4_X1 U4486 ( .A1(n3784), .A2(n3783), .A3(n3795), .A4(n3782), .ZN(n3787)
         );
  AND3_X1 U4487 ( .A1(n3787), .A2(n3786), .A3(n3785), .ZN(n3791) );
  NAND2_X1 U4488 ( .A1(n2087), .A2(n3788), .ZN(n3797) );
  OAI211_X1 U4489 ( .C1(n3791), .C2(n3797), .A(n3790), .B(n3789), .ZN(n3801)
         );
  NOR2_X1 U4490 ( .A1(n2160), .A2(n3792), .ZN(n3800) );
  NAND3_X1 U4491 ( .A1(n3795), .A2(n2181), .A3(n3794), .ZN(n3798) );
  OAI21_X1 U4492 ( .B1(n3798), .B2(n3797), .A(n3796), .ZN(n3799) );
  AOI22_X1 U4493 ( .A1(n3801), .A2(n3800), .B1(n3806), .B2(n3799), .ZN(n3810)
         );
  NAND3_X1 U4494 ( .A1(n3804), .A2(n3803), .A3(n3802), .ZN(n3809) );
  OAI21_X1 U4495 ( .B1(n2185), .B2(n3807), .A(n3806), .ZN(n3808) );
  OAI21_X1 U4496 ( .B1(n3810), .B2(n3809), .A(n3808), .ZN(n3814) );
  INV_X1 U4497 ( .A(n3811), .ZN(n3812) );
  AOI21_X1 U4498 ( .B1(n3814), .B2(n3813), .A(n3812), .ZN(n3817) );
  OAI21_X1 U4499 ( .B1(n3817), .B2(n3816), .A(n3815), .ZN(n3820) );
  OR2_X1 U4500 ( .A1(n3818), .A2(n4237), .ZN(n3819) );
  AOI211_X1 U4501 ( .C1(n3821), .C2(n3820), .A(n4236), .B(n3819), .ZN(n3827)
         );
  NOR2_X1 U4502 ( .A1(n3823), .A2(n3822), .ZN(n3824) );
  AOI221_X1 U4503 ( .B1(n3827), .B2(n3826), .C1(n3825), .C2(n3826), .A(n3824), 
        .ZN(n3828) );
  AND2_X1 U4504 ( .A1(n3829), .A2(n3828), .ZN(n3833) );
  OAI22_X1 U4505 ( .A1(n3833), .A2(n3832), .B1(n3831), .B2(n3830), .ZN(n3835)
         );
  MUX2_X1 U4506 ( .A(n3836), .B(n3835), .S(n3834), .Z(n3837) );
  XNOR2_X1 U4507 ( .A(n3837), .B(n4132), .ZN(n3842) );
  NOR2_X1 U4508 ( .A1(n3838), .A2(n3873), .ZN(n3840) );
  OAI21_X1 U4509 ( .B1(n3841), .B2(n4442), .A(B_REG_SCAN_IN), .ZN(n3839) );
  OAI22_X1 U4510 ( .A1(n3842), .A2(n3841), .B1(n3840), .B2(n3839), .ZN(U3239)
         );
  MUX2_X1 U4511 ( .A(n3843), .B(DATAO_REG_31__SCAN_IN), .S(n3875), .Z(U3581)
         );
  MUX2_X1 U4512 ( .A(n3844), .B(DATAO_REG_29__SCAN_IN), .S(n3875), .Z(U3579)
         );
  MUX2_X1 U4513 ( .A(n4169), .B(DATAO_REG_28__SCAN_IN), .S(n3875), .Z(U3578)
         );
  MUX2_X1 U4514 ( .A(n4184), .B(DATAO_REG_27__SCAN_IN), .S(n3875), .Z(U3577)
         );
  MUX2_X1 U4515 ( .A(n4204), .B(DATAO_REG_26__SCAN_IN), .S(n3875), .Z(U3576)
         );
  MUX2_X1 U4516 ( .A(n4220), .B(DATAO_REG_25__SCAN_IN), .S(n3875), .Z(U3575)
         );
  MUX2_X1 U4517 ( .A(n4242), .B(DATAO_REG_24__SCAN_IN), .S(n3875), .Z(U3574)
         );
  MUX2_X1 U4518 ( .A(n4263), .B(DATAO_REG_23__SCAN_IN), .S(n3875), .Z(U3573)
         );
  MUX2_X1 U4519 ( .A(DATAO_REG_22__SCAN_IN), .B(n4279), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4520 ( .A(n3846), .B(DATAO_REG_20__SCAN_IN), .S(n3875), .Z(U3570)
         );
  MUX2_X1 U4521 ( .A(n4300), .B(DATAO_REG_19__SCAN_IN), .S(n3875), .Z(U3569)
         );
  MUX2_X1 U4522 ( .A(n3847), .B(DATAO_REG_17__SCAN_IN), .S(n3875), .Z(U3567)
         );
  MUX2_X1 U4523 ( .A(n3848), .B(DATAO_REG_15__SCAN_IN), .S(n3875), .Z(U3565)
         );
  MUX2_X1 U4524 ( .A(n4455), .B(DATAO_REG_14__SCAN_IN), .S(n3875), .Z(U3564)
         );
  MUX2_X1 U4525 ( .A(n3849), .B(DATAO_REG_13__SCAN_IN), .S(n3875), .Z(U3563)
         );
  MUX2_X1 U4526 ( .A(n3850), .B(DATAO_REG_11__SCAN_IN), .S(n3875), .Z(U3561)
         );
  MUX2_X1 U4527 ( .A(n3851), .B(DATAO_REG_10__SCAN_IN), .S(n3875), .Z(U3560)
         );
  MUX2_X1 U4528 ( .A(n3852), .B(DATAO_REG_9__SCAN_IN), .S(n3875), .Z(U3559) );
  MUX2_X1 U4529 ( .A(n3853), .B(DATAO_REG_7__SCAN_IN), .S(n3875), .Z(U3557) );
  MUX2_X1 U4530 ( .A(n3854), .B(DATAO_REG_6__SCAN_IN), .S(n3875), .Z(U3556) );
  MUX2_X1 U4531 ( .A(n3855), .B(DATAO_REG_5__SCAN_IN), .S(n3875), .Z(U3555) );
  MUX2_X1 U4532 ( .A(n3856), .B(DATAO_REG_4__SCAN_IN), .S(n3875), .Z(U3554) );
  MUX2_X1 U4533 ( .A(n3857), .B(DATAO_REG_3__SCAN_IN), .S(n3875), .Z(U3553) );
  MUX2_X1 U4534 ( .A(n3858), .B(DATAO_REG_2__SCAN_IN), .S(n3875), .Z(U3552) );
  MUX2_X1 U4535 ( .A(n3859), .B(DATAO_REG_1__SCAN_IN), .S(n3875), .Z(U3551) );
  OAI211_X1 U4536 ( .C1(n3862), .C2(n3861), .A(n4589), .B(n3860), .ZN(n3868)
         );
  INV_X1 U4537 ( .A(n4611), .ZN(n4566) );
  NAND2_X1 U4538 ( .A1(n4566), .A2(n4451), .ZN(n3867) );
  XOR2_X1 U4539 ( .A(n3863), .B(n3872), .Z(n3864) );
  NAND2_X1 U4540 ( .A1(n4608), .A2(n3864), .ZN(n3866) );
  AOI22_X1 U4541 ( .A1(n4597), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3865) );
  NAND4_X1 U4542 ( .A1(n3868), .A2(n3867), .A3(n3866), .A4(n3865), .ZN(U3241)
         );
  NOR3_X1 U4543 ( .A1(n3869), .A2(n4481), .A3(n3871), .ZN(n3876) );
  NOR2_X1 U4544 ( .A1(n4145), .A2(REG2_REG_0__SCAN_IN), .ZN(n3870) );
  NOR2_X1 U4545 ( .A1(n3871), .A2(n3870), .ZN(n4480) );
  OAI22_X1 U4546 ( .A1(n4480), .A2(IR_REG_0__SCAN_IN), .B1(n3873), .B2(n3872), 
        .ZN(n3874) );
  OR3_X1 U4547 ( .A1(n3876), .A2(n3875), .A3(n3874), .ZN(n4496) );
  AOI22_X1 U4548 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4597), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3888) );
  INV_X1 U4549 ( .A(n4450), .ZN(n3881) );
  OAI21_X1 U4550 ( .B1(n3879), .B2(n3878), .A(n3877), .ZN(n3880) );
  OAI22_X1 U4551 ( .A1(n3881), .A2(n4611), .B1(n4594), .B2(n3880), .ZN(n3882)
         );
  INV_X1 U4552 ( .A(n3882), .ZN(n3887) );
  OAI211_X1 U4553 ( .C1(n3885), .C2(n3884), .A(n4608), .B(n3883), .ZN(n3886)
         );
  NAND4_X1 U4554 ( .A1(n4496), .A2(n3888), .A3(n3887), .A4(n3886), .ZN(n4068)
         );
  AOI22_X1 U4555 ( .A1(n3890), .A2(keyinput66), .B1(keyinput71), .B2(n4053), 
        .ZN(n3889) );
  OAI221_X1 U4556 ( .B1(n3890), .B2(keyinput66), .C1(n4053), .C2(keyinput71), 
        .A(n3889), .ZN(n3901) );
  INV_X1 U4557 ( .A(REG1_REG_22__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4558 ( .A1(n4382), .A2(keyinput119), .B1(n3892), .B2(keyinput90), 
        .ZN(n3891) );
  OAI221_X1 U4559 ( .B1(n4382), .B2(keyinput119), .C1(n3892), .C2(keyinput90), 
        .A(n3891), .ZN(n3900) );
  AOI22_X1 U4560 ( .A1(n3895), .A2(keyinput102), .B1(keyinput81), .B2(n3894), 
        .ZN(n3893) );
  OAI221_X1 U4561 ( .B1(n3895), .B2(keyinput102), .C1(n3894), .C2(keyinput81), 
        .A(n3893), .ZN(n3899) );
  INV_X1 U4562 ( .A(ADDR_REG_14__SCAN_IN), .ZN(n4569) );
  AOI22_X1 U4563 ( .A1(n3897), .A2(keyinput96), .B1(n4569), .B2(keyinput92), 
        .ZN(n3896) );
  OAI221_X1 U4564 ( .B1(n3897), .B2(keyinput96), .C1(n4569), .C2(keyinput92), 
        .A(n3896), .ZN(n3898) );
  NOR4_X1 U4565 ( .A1(n3901), .A2(n3900), .A3(n3899), .A4(n3898), .ZN(n3935)
         );
  AOI22_X1 U4566 ( .A1(n4070), .A2(keyinput89), .B1(keyinput84), .B2(n2371), 
        .ZN(n3902) );
  OAI221_X1 U4567 ( .B1(n4070), .B2(keyinput89), .C1(n2371), .C2(keyinput84), 
        .A(n3902), .ZN(n3912) );
  INV_X1 U4568 ( .A(REG2_REG_6__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U4569 ( .A1(n3174), .A2(keyinput117), .B1(keyinput88), .B2(n4024), 
        .ZN(n3903) );
  OAI221_X1 U4570 ( .B1(n3174), .B2(keyinput117), .C1(n4024), .C2(keyinput88), 
        .A(n3903), .ZN(n3911) );
  AOI22_X1 U4571 ( .A1(n3906), .A2(keyinput104), .B1(n3905), .B2(keyinput113), 
        .ZN(n3904) );
  OAI221_X1 U4572 ( .B1(n3906), .B2(keyinput104), .C1(n3905), .C2(keyinput113), 
        .A(n3904), .ZN(n3910) );
  INV_X1 U4573 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4012) );
  XOR2_X1 U4574 ( .A(n4012), .B(keyinput111), .Z(n3908) );
  XNOR2_X1 U4575 ( .A(REG2_REG_0__SCAN_IN), .B(keyinput107), .ZN(n3907) );
  NAND2_X1 U4576 ( .A1(n3908), .A2(n3907), .ZN(n3909) );
  NOR4_X1 U4577 ( .A1(n3912), .A2(n3911), .A3(n3910), .A4(n3909), .ZN(n3934)
         );
  INV_X1 U4578 ( .A(D_REG_11__SCAN_IN), .ZN(n4631) );
  AOI22_X1 U4579 ( .A1(n4039), .A2(keyinput65), .B1(n4631), .B2(keyinput69), 
        .ZN(n3913) );
  OAI221_X1 U4580 ( .B1(n4039), .B2(keyinput65), .C1(n4631), .C2(keyinput69), 
        .A(n3913), .ZN(n3921) );
  INV_X1 U4581 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U4582 ( .A1(n3915), .A2(keyinput74), .B1(n4028), .B2(keyinput116), 
        .ZN(n3914) );
  OAI221_X1 U4583 ( .B1(n3915), .B2(keyinput74), .C1(n4028), .C2(keyinput116), 
        .A(n3914), .ZN(n3920) );
  INV_X1 U4584 ( .A(D_REG_23__SCAN_IN), .ZN(n4629) );
  INV_X1 U4585 ( .A(D_REG_20__SCAN_IN), .ZN(n4630) );
  AOI22_X1 U4586 ( .A1(n4629), .A2(keyinput124), .B1(n4630), .B2(keyinput68), 
        .ZN(n3916) );
  OAI221_X1 U4587 ( .B1(n4629), .B2(keyinput124), .C1(n4630), .C2(keyinput68), 
        .A(n3916), .ZN(n3919) );
  INV_X1 U4588 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4677) );
  INV_X1 U4589 ( .A(D_REG_31__SCAN_IN), .ZN(n4628) );
  AOI22_X1 U4590 ( .A1(n4677), .A2(keyinput67), .B1(n4628), .B2(keyinput80), 
        .ZN(n3917) );
  OAI221_X1 U4591 ( .B1(n4677), .B2(keyinput67), .C1(n4628), .C2(keyinput80), 
        .A(n3917), .ZN(n3918) );
  NOR4_X1 U4592 ( .A1(n3921), .A2(n3920), .A3(n3919), .A4(n3918), .ZN(n3933)
         );
  AOI22_X1 U4593 ( .A1(n4054), .A2(keyinput78), .B1(keyinput91), .B2(n4048), 
        .ZN(n3922) );
  OAI221_X1 U4594 ( .B1(n4054), .B2(keyinput78), .C1(n4048), .C2(keyinput91), 
        .A(n3922), .ZN(n3931) );
  INV_X1 U4595 ( .A(DATAI_26_), .ZN(n3924) );
  AOI22_X1 U4596 ( .A1(n3924), .A2(keyinput127), .B1(keyinput94), .B2(n2102), 
        .ZN(n3923) );
  OAI221_X1 U4597 ( .B1(n3924), .B2(keyinput127), .C1(n2102), .C2(keyinput94), 
        .A(n3923), .ZN(n3930) );
  AOI22_X1 U4598 ( .A1(n4037), .A2(keyinput76), .B1(n4047), .B2(keyinput86), 
        .ZN(n3925) );
  OAI221_X1 U4599 ( .B1(n4037), .B2(keyinput76), .C1(n4047), .C2(keyinput86), 
        .A(n3925), .ZN(n3929) );
  XOR2_X1 U4600 ( .A(n4010), .B(keyinput95), .Z(n3927) );
  XNOR2_X1 U4601 ( .A(IR_REG_4__SCAN_IN), .B(keyinput87), .ZN(n3926) );
  NAND2_X1 U4602 ( .A1(n3927), .A2(n3926), .ZN(n3928) );
  NOR4_X1 U4603 ( .A1(n3931), .A2(n3930), .A3(n3929), .A4(n3928), .ZN(n3932)
         );
  AND4_X1 U4604 ( .A1(n3935), .A2(n3934), .A3(n3933), .A4(n3932), .ZN(n4066)
         );
  OAI22_X1 U4605 ( .A1(B_REG_SCAN_IN), .A2(keyinput121), .B1(
        ADDR_REG_3__SCAN_IN), .B2(keyinput109), .ZN(n3936) );
  AOI221_X1 U4606 ( .B1(B_REG_SCAN_IN), .B2(keyinput121), .C1(keyinput109), 
        .C2(ADDR_REG_3__SCAN_IN), .A(n3936), .ZN(n3943) );
  OAI22_X1 U4607 ( .A1(REG3_REG_22__SCAN_IN), .A2(keyinput64), .B1(
        REG3_REG_9__SCAN_IN), .B2(keyinput112), .ZN(n3937) );
  AOI221_X1 U4608 ( .B1(REG3_REG_22__SCAN_IN), .B2(keyinput64), .C1(
        keyinput112), .C2(REG3_REG_9__SCAN_IN), .A(n3937), .ZN(n3942) );
  OAI22_X1 U4609 ( .A1(IR_REG_0__SCAN_IN), .A2(keyinput82), .B1(keyinput75), 
        .B2(DATAO_REG_6__SCAN_IN), .ZN(n3938) );
  AOI221_X1 U4610 ( .B1(IR_REG_0__SCAN_IN), .B2(keyinput82), .C1(
        DATAO_REG_6__SCAN_IN), .C2(keyinput75), .A(n3938), .ZN(n3941) );
  OAI22_X1 U4611 ( .A1(ADDR_REG_13__SCAN_IN), .A2(keyinput110), .B1(keyinput70), .B2(ADDR_REG_10__SCAN_IN), .ZN(n3939) );
  AOI221_X1 U4612 ( .B1(ADDR_REG_13__SCAN_IN), .B2(keyinput110), .C1(
        ADDR_REG_10__SCAN_IN), .C2(keyinput70), .A(n3939), .ZN(n3940) );
  NAND4_X1 U4613 ( .A1(n3943), .A2(n3942), .A3(n3941), .A4(n3940), .ZN(n3972)
         );
  OAI22_X1 U4614 ( .A1(REG2_REG_17__SCAN_IN), .A2(keyinput79), .B1(
        REG2_REG_14__SCAN_IN), .B2(keyinput73), .ZN(n3944) );
  AOI221_X1 U4615 ( .B1(REG2_REG_17__SCAN_IN), .B2(keyinput79), .C1(keyinput73), .C2(REG2_REG_14__SCAN_IN), .A(n3944), .ZN(n3951) );
  OAI22_X1 U4616 ( .A1(REG2_REG_28__SCAN_IN), .A2(keyinput101), .B1(keyinput99), .B2(REG2_REG_12__SCAN_IN), .ZN(n3945) );
  AOI221_X1 U4617 ( .B1(REG2_REG_28__SCAN_IN), .B2(keyinput101), .C1(
        REG2_REG_12__SCAN_IN), .C2(keyinput99), .A(n3945), .ZN(n3950) );
  OAI22_X1 U4618 ( .A1(DATAO_REG_20__SCAN_IN), .A2(keyinput118), .B1(
        DATAO_REG_17__SCAN_IN), .B2(keyinput77), .ZN(n3946) );
  AOI221_X1 U4619 ( .B1(DATAO_REG_20__SCAN_IN), .B2(keyinput118), .C1(
        keyinput77), .C2(DATAO_REG_17__SCAN_IN), .A(n3946), .ZN(n3949) );
  OAI22_X1 U4620 ( .A1(REG1_REG_16__SCAN_IN), .A2(keyinput100), .B1(
        REG1_REG_6__SCAN_IN), .B2(keyinput122), .ZN(n3947) );
  AOI221_X1 U4621 ( .B1(REG1_REG_16__SCAN_IN), .B2(keyinput100), .C1(
        keyinput122), .C2(REG1_REG_6__SCAN_IN), .A(n3947), .ZN(n3948) );
  NAND4_X1 U4622 ( .A1(n3951), .A2(n3950), .A3(n3949), .A4(n3948), .ZN(n3971)
         );
  OAI22_X1 U4623 ( .A1(REG0_REG_27__SCAN_IN), .A2(keyinput108), .B1(keyinput97), .B2(REG1_REG_1__SCAN_IN), .ZN(n3952) );
  AOI221_X1 U4624 ( .B1(REG0_REG_27__SCAN_IN), .B2(keyinput108), .C1(
        REG1_REG_1__SCAN_IN), .C2(keyinput97), .A(n3952), .ZN(n3959) );
  OAI22_X1 U4625 ( .A1(REG0_REG_12__SCAN_IN), .A2(keyinput93), .B1(keyinput106), .B2(REG0_REG_11__SCAN_IN), .ZN(n3953) );
  AOI221_X1 U4626 ( .B1(REG0_REG_12__SCAN_IN), .B2(keyinput93), .C1(
        REG0_REG_11__SCAN_IN), .C2(keyinput106), .A(n3953), .ZN(n3958) );
  OAI22_X1 U4627 ( .A1(D_REG_6__SCAN_IN), .A2(keyinput114), .B1(
        D_REG_2__SCAN_IN), .B2(keyinput126), .ZN(n3954) );
  AOI221_X1 U4628 ( .B1(D_REG_6__SCAN_IN), .B2(keyinput114), .C1(keyinput126), 
        .C2(D_REG_2__SCAN_IN), .A(n3954), .ZN(n3957) );
  OAI22_X1 U4629 ( .A1(D_REG_19__SCAN_IN), .A2(keyinput125), .B1(keyinput115), 
        .B2(REG0_REG_26__SCAN_IN), .ZN(n3955) );
  AOI221_X1 U4630 ( .B1(D_REG_19__SCAN_IN), .B2(keyinput125), .C1(
        REG0_REG_26__SCAN_IN), .C2(keyinput115), .A(n3955), .ZN(n3956) );
  NAND4_X1 U4631 ( .A1(n3959), .A2(n3958), .A3(n3957), .A4(n3956), .ZN(n3970)
         );
  OAI22_X1 U4632 ( .A1(IR_REG_14__SCAN_IN), .A2(keyinput105), .B1(
        IR_REG_3__SCAN_IN), .B2(keyinput103), .ZN(n3961) );
  AOI221_X1 U4633 ( .B1(IR_REG_14__SCAN_IN), .B2(keyinput105), .C1(keyinput103), .C2(IR_REG_3__SCAN_IN), .A(n3961), .ZN(n3968) );
  OAI22_X1 U4634 ( .A1(IR_REG_16__SCAN_IN), .A2(keyinput123), .B1(keyinput72), 
        .B2(REG3_REG_1__SCAN_IN), .ZN(n3962) );
  AOI221_X1 U4635 ( .B1(IR_REG_16__SCAN_IN), .B2(keyinput123), .C1(
        REG3_REG_1__SCAN_IN), .C2(keyinput72), .A(n3962), .ZN(n3967) );
  OAI22_X1 U4636 ( .A1(DATAI_11_), .A2(keyinput98), .B1(keyinput120), .B2(
        DATAI_4_), .ZN(n3963) );
  AOI221_X1 U4637 ( .B1(DATAI_11_), .B2(keyinput98), .C1(DATAI_4_), .C2(
        keyinput120), .A(n3963), .ZN(n3966) );
  OAI22_X1 U4638 ( .A1(DATAI_25_), .A2(keyinput85), .B1(DATAI_1_), .B2(
        keyinput83), .ZN(n3964) );
  AOI221_X1 U4639 ( .B1(DATAI_25_), .B2(keyinput85), .C1(keyinput83), .C2(
        DATAI_1_), .A(n3964), .ZN(n3965) );
  NAND4_X1 U4640 ( .A1(n3968), .A2(n3967), .A3(n3966), .A4(n3965), .ZN(n3969)
         );
  NOR4_X1 U4641 ( .A1(n3972), .A2(n3971), .A3(n3970), .A4(n3969), .ZN(n4065)
         );
  AOI22_X1 U4642 ( .A1(REG2_REG_10__SCAN_IN), .A2(keyinput53), .B1(
        D_REG_19__SCAN_IN), .B2(keyinput61), .ZN(n3973) );
  OAI221_X1 U4643 ( .B1(REG2_REG_10__SCAN_IN), .B2(keyinput53), .C1(
        D_REG_19__SCAN_IN), .C2(keyinput61), .A(n3973), .ZN(n3980) );
  AOI22_X1 U4644 ( .A1(ADDR_REG_3__SCAN_IN), .A2(keyinput45), .B1(
        B_REG_SCAN_IN), .B2(keyinput57), .ZN(n3974) );
  OAI221_X1 U4645 ( .B1(ADDR_REG_3__SCAN_IN), .B2(keyinput45), .C1(
        B_REG_SCAN_IN), .C2(keyinput57), .A(n3974), .ZN(n3979) );
  AOI22_X1 U4646 ( .A1(DATAO_REG_17__SCAN_IN), .A2(keyinput13), .B1(
        IR_REG_14__SCAN_IN), .B2(keyinput41), .ZN(n3975) );
  OAI221_X1 U4647 ( .B1(DATAO_REG_17__SCAN_IN), .B2(keyinput13), .C1(
        IR_REG_14__SCAN_IN), .C2(keyinput41), .A(n3975), .ZN(n3978) );
  AOI22_X1 U4648 ( .A1(DATAO_REG_12__SCAN_IN), .A2(keyinput17), .B1(
        REG1_REG_29__SCAN_IN), .B2(keyinput49), .ZN(n3976) );
  OAI221_X1 U4649 ( .B1(DATAO_REG_12__SCAN_IN), .B2(keyinput17), .C1(
        REG1_REG_29__SCAN_IN), .C2(keyinput49), .A(n3976), .ZN(n3977) );
  NOR4_X1 U4650 ( .A1(n3980), .A2(n3979), .A3(n3978), .A4(n3977), .ZN(n4008)
         );
  AOI22_X1 U4651 ( .A1(DATAI_4_), .A2(keyinput56), .B1(DATAI_26_), .B2(
        keyinput63), .ZN(n3981) );
  OAI221_X1 U4652 ( .B1(DATAI_4_), .B2(keyinput56), .C1(DATAI_26_), .C2(
        keyinput63), .A(n3981), .ZN(n3988) );
  AOI22_X1 U4653 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput8), .B1(
        REG3_REG_9__SCAN_IN), .B2(keyinput48), .ZN(n3982) );
  OAI221_X1 U4654 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput8), .C1(
        REG3_REG_9__SCAN_IN), .C2(keyinput48), .A(n3982), .ZN(n3987) );
  AOI22_X1 U4655 ( .A1(REG1_REG_28__SCAN_IN), .A2(keyinput40), .B1(
        D_REG_20__SCAN_IN), .B2(keyinput4), .ZN(n3983) );
  OAI221_X1 U4656 ( .B1(REG1_REG_28__SCAN_IN), .B2(keyinput40), .C1(
        D_REG_20__SCAN_IN), .C2(keyinput4), .A(n3983), .ZN(n3986) );
  AOI22_X1 U4657 ( .A1(DATAO_REG_21__SCAN_IN), .A2(keyinput32), .B1(
        ADDR_REG_14__SCAN_IN), .B2(keyinput28), .ZN(n3984) );
  OAI221_X1 U4658 ( .B1(DATAO_REG_21__SCAN_IN), .B2(keyinput32), .C1(
        ADDR_REG_14__SCAN_IN), .C2(keyinput28), .A(n3984), .ZN(n3985) );
  NOR4_X1 U4659 ( .A1(n3988), .A2(n3987), .A3(n3986), .A4(n3985), .ZN(n4007)
         );
  AOI22_X1 U4660 ( .A1(REG1_REG_6__SCAN_IN), .A2(keyinput58), .B1(
        D_REG_6__SCAN_IN), .B2(keyinput50), .ZN(n3989) );
  OAI221_X1 U4661 ( .B1(REG1_REG_6__SCAN_IN), .B2(keyinput58), .C1(
        D_REG_6__SCAN_IN), .C2(keyinput50), .A(n3989), .ZN(n3996) );
  AOI22_X1 U4662 ( .A1(DATAO_REG_20__SCAN_IN), .A2(keyinput54), .B1(
        REG0_REG_11__SCAN_IN), .B2(keyinput42), .ZN(n3990) );
  OAI221_X1 U4663 ( .B1(DATAO_REG_20__SCAN_IN), .B2(keyinput54), .C1(
        REG0_REG_11__SCAN_IN), .C2(keyinput42), .A(n3990), .ZN(n3995) );
  AOI22_X1 U4664 ( .A1(DATAO_REG_8__SCAN_IN), .A2(keyinput38), .B1(DATAI_0_), 
        .B2(keyinput30), .ZN(n3991) );
  OAI221_X1 U4665 ( .B1(DATAO_REG_8__SCAN_IN), .B2(keyinput38), .C1(DATAI_0_), 
        .C2(keyinput30), .A(n3991), .ZN(n3994) );
  AOI22_X1 U4666 ( .A1(ADDR_REG_10__SCAN_IN), .A2(keyinput6), .B1(
        REG1_REG_22__SCAN_IN), .B2(keyinput26), .ZN(n3992) );
  OAI221_X1 U4667 ( .B1(ADDR_REG_10__SCAN_IN), .B2(keyinput6), .C1(
        REG1_REG_22__SCAN_IN), .C2(keyinput26), .A(n3992), .ZN(n3993) );
  NOR4_X1 U4668 ( .A1(n3996), .A2(n3995), .A3(n3994), .A4(n3993), .ZN(n4006)
         );
  AOI22_X1 U4669 ( .A1(DATAO_REG_18__SCAN_IN), .A2(keyinput2), .B1(
        REG0_REG_6__SCAN_IN), .B2(keyinput10), .ZN(n3997) );
  OAI221_X1 U4670 ( .B1(DATAO_REG_18__SCAN_IN), .B2(keyinput2), .C1(
        REG0_REG_6__SCAN_IN), .C2(keyinput10), .A(n3997), .ZN(n4004) );
  AOI22_X1 U4671 ( .A1(DATAO_REG_6__SCAN_IN), .A2(keyinput11), .B1(DATAI_1_), 
        .B2(keyinput19), .ZN(n3998) );
  OAI221_X1 U4672 ( .B1(DATAO_REG_6__SCAN_IN), .B2(keyinput11), .C1(DATAI_1_), 
        .C2(keyinput19), .A(n3998), .ZN(n4003) );
  AOI22_X1 U4673 ( .A1(REG0_REG_4__SCAN_IN), .A2(keyinput3), .B1(
        REG2_REG_12__SCAN_IN), .B2(keyinput35), .ZN(n3999) );
  OAI221_X1 U4674 ( .B1(REG0_REG_4__SCAN_IN), .B2(keyinput3), .C1(
        REG2_REG_12__SCAN_IN), .C2(keyinput35), .A(n3999), .ZN(n4002) );
  AOI22_X1 U4675 ( .A1(REG1_REG_21__SCAN_IN), .A2(keyinput55), .B1(
        IR_REG_4__SCAN_IN), .B2(keyinput23), .ZN(n4000) );
  OAI221_X1 U4676 ( .B1(REG1_REG_21__SCAN_IN), .B2(keyinput55), .C1(
        IR_REG_4__SCAN_IN), .C2(keyinput23), .A(n4000), .ZN(n4001) );
  NOR4_X1 U4677 ( .A1(n4004), .A2(n4003), .A3(n4002), .A4(n4001), .ZN(n4005)
         );
  NAND4_X1 U4678 ( .A1(n4008), .A2(n4007), .A3(n4006), .A4(n4005), .ZN(n4064)
         );
  INV_X1 U4679 ( .A(DATAI_11_), .ZN(n4647) );
  AOI22_X1 U4680 ( .A1(n4647), .A2(keyinput34), .B1(n4010), .B2(keyinput31), 
        .ZN(n4009) );
  OAI221_X1 U4681 ( .B1(n4647), .B2(keyinput34), .C1(n4010), .C2(keyinput31), 
        .A(n4009), .ZN(n4020) );
  INV_X1 U4682 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4683 ( .A1(n4013), .A2(keyinput46), .B1(n4012), .B2(keyinput47), 
        .ZN(n4011) );
  OAI221_X1 U4684 ( .B1(n4013), .B2(keyinput46), .C1(n4012), .C2(keyinput47), 
        .A(n4011), .ZN(n4019) );
  XNOR2_X1 U4685 ( .A(IR_REG_16__SCAN_IN), .B(keyinput59), .ZN(n4017) );
  XNOR2_X1 U4686 ( .A(REG0_REG_26__SCAN_IN), .B(keyinput51), .ZN(n4016) );
  XNOR2_X1 U4687 ( .A(REG2_REG_0__SCAN_IN), .B(keyinput43), .ZN(n4015) );
  XNOR2_X1 U4688 ( .A(IR_REG_3__SCAN_IN), .B(keyinput39), .ZN(n4014) );
  NAND4_X1 U4689 ( .A1(n4017), .A2(n4016), .A3(n4015), .A4(n4014), .ZN(n4018)
         );
  NOR3_X1 U4690 ( .A1(n4020), .A2(n4019), .A3(n4018), .ZN(n4062) );
  INV_X1 U4691 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U4692 ( .A1(n4084), .A2(keyinput36), .B1(n4022), .B2(keyinput44), 
        .ZN(n4021) );
  OAI221_X1 U4693 ( .B1(n4084), .B2(keyinput36), .C1(n4022), .C2(keyinput44), 
        .A(n4021), .ZN(n4032) );
  AOI22_X1 U4694 ( .A1(n4024), .A2(keyinput24), .B1(n4628), .B2(keyinput16), 
        .ZN(n4023) );
  OAI221_X1 U4695 ( .B1(n4024), .B2(keyinput24), .C1(n4628), .C2(keyinput16), 
        .A(n4023), .ZN(n4031) );
  INV_X1 U4696 ( .A(D_REG_2__SCAN_IN), .ZN(n4633) );
  AOI22_X1 U4697 ( .A1(n4026), .A2(keyinput0), .B1(n4633), .B2(keyinput62), 
        .ZN(n4025) );
  OAI221_X1 U4698 ( .B1(n4026), .B2(keyinput0), .C1(n4633), .C2(keyinput62), 
        .A(n4025), .ZN(n4030) );
  AOI22_X1 U4699 ( .A1(n4028), .A2(keyinput52), .B1(n4629), .B2(keyinput60), 
        .ZN(n4027) );
  OAI221_X1 U4700 ( .B1(n4028), .B2(keyinput52), .C1(n4629), .C2(keyinput60), 
        .A(n4027), .ZN(n4029) );
  NOR4_X1 U4701 ( .A1(n4032), .A2(n4031), .A3(n4030), .A4(n4029), .ZN(n4061)
         );
  INV_X1 U4702 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4034) );
  AOI22_X1 U4703 ( .A1(n3238), .A2(keyinput9), .B1(keyinput29), .B2(n4034), 
        .ZN(n4033) );
  OAI221_X1 U4704 ( .B1(n3238), .B2(keyinput9), .C1(n4034), .C2(keyinput29), 
        .A(n4033), .ZN(n4043) );
  AOI22_X1 U4705 ( .A1(n4070), .A2(keyinput25), .B1(keyinput20), .B2(n2371), 
        .ZN(n4035) );
  OAI221_X1 U4706 ( .B1(n4070), .B2(keyinput25), .C1(n2371), .C2(keyinput20), 
        .A(n4035), .ZN(n4042) );
  AOI22_X1 U4707 ( .A1(n4631), .A2(keyinput5), .B1(keyinput12), .B2(n4037), 
        .ZN(n4036) );
  OAI221_X1 U4708 ( .B1(n4631), .B2(keyinput5), .C1(n4037), .C2(keyinput12), 
        .A(n4036), .ZN(n4041) );
  AOI22_X1 U4709 ( .A1(n2845), .A2(keyinput33), .B1(n4039), .B2(keyinput1), 
        .ZN(n4038) );
  OAI221_X1 U4710 ( .B1(n2845), .B2(keyinput33), .C1(n4039), .C2(keyinput1), 
        .A(n4038), .ZN(n4040) );
  NOR4_X1 U4711 ( .A1(n4043), .A2(n4042), .A3(n4041), .A4(n4040), .ZN(n4060)
         );
  INV_X1 U4712 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U4713 ( .A1(n2103), .A2(keyinput18), .B1(keyinput15), .B2(n4045), 
        .ZN(n4044) );
  OAI221_X1 U4714 ( .B1(n2103), .B2(keyinput18), .C1(n4045), .C2(keyinput15), 
        .A(n4044), .ZN(n4058) );
  AOI22_X1 U4715 ( .A1(n4048), .A2(keyinput27), .B1(n4047), .B2(keyinput22), 
        .ZN(n4046) );
  OAI221_X1 U4716 ( .B1(n4048), .B2(keyinput27), .C1(n4047), .C2(keyinput22), 
        .A(n4046), .ZN(n4057) );
  INV_X1 U4717 ( .A(REG2_REG_28__SCAN_IN), .ZN(n4051) );
  INV_X1 U4718 ( .A(DATAI_25_), .ZN(n4050) );
  AOI22_X1 U4719 ( .A1(n4051), .A2(keyinput37), .B1(keyinput21), .B2(n4050), 
        .ZN(n4049) );
  OAI221_X1 U4720 ( .B1(n4051), .B2(keyinput37), .C1(n4050), .C2(keyinput21), 
        .A(n4049), .ZN(n4056) );
  AOI22_X1 U4721 ( .A1(n4054), .A2(keyinput14), .B1(keyinput7), .B2(n4053), 
        .ZN(n4052) );
  OAI221_X1 U4722 ( .B1(n4054), .B2(keyinput14), .C1(n4053), .C2(keyinput7), 
        .A(n4052), .ZN(n4055) );
  NOR4_X1 U4723 ( .A1(n4058), .A2(n4057), .A3(n4056), .A4(n4055), .ZN(n4059)
         );
  NAND4_X1 U4724 ( .A1(n4062), .A2(n4061), .A3(n4060), .A4(n4059), .ZN(n4063)
         );
  AOI211_X1 U4725 ( .C1(n4066), .C2(n4065), .A(n4064), .B(n4063), .ZN(n4067)
         );
  XOR2_X1 U4726 ( .A(n4068), .B(n4067), .Z(U3242) );
  OAI21_X1 U4727 ( .B1(n4070), .B2(n4091), .A(n4069), .ZN(n4071) );
  OAI21_X1 U4728 ( .B1(REG1_REG_7__SCAN_IN), .B2(n4445), .A(n4071), .ZN(n4072)
         );
  INV_X1 U4729 ( .A(n4651), .ZN(n4516) );
  AOI22_X1 U4730 ( .A1(n4651), .A2(n2406), .B1(REG1_REG_9__SCAN_IN), .B2(n4516), .ZN(n4508) );
  AOI21_X1 U4731 ( .B1(REG1_REG_9__SCAN_IN), .B2(n4651), .A(n4507), .ZN(n4075)
         );
  INV_X1 U4732 ( .A(n4098), .ZN(n4650) );
  INV_X1 U4733 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4519) );
  XNOR2_X1 U4734 ( .A(n4650), .B(n4075), .ZN(n4518) );
  INV_X1 U4735 ( .A(n4089), .ZN(n4648) );
  AOI22_X1 U4736 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4648), .B1(n4089), .B2(
        n2443), .ZN(n4527) );
  XOR2_X1 U4737 ( .A(n4076), .B(n4645), .Z(n4536) );
  NOR2_X1 U4738 ( .A1(n4076), .A2(n4544), .ZN(n4077) );
  AOI22_X1 U4739 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4556), .B1(n4643), .B2(
        n4078), .ZN(n4546) );
  NOR2_X1 U4740 ( .A1(n4080), .A2(n4079), .ZN(n4081) );
  AOI22_X1 U4741 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4641), .B1(n4106), .B2(
        n4082), .ZN(n4572) );
  AND2_X1 U4742 ( .A1(n4106), .A2(REG1_REG_15__SCAN_IN), .ZN(n4083) );
  XNOR2_X1 U4743 ( .A(n4115), .B(n4444), .ZN(n4085) );
  NAND2_X1 U4744 ( .A1(n4085), .A2(n4084), .ZN(n4116) );
  OAI21_X1 U4745 ( .B1(n4085), .B2(n4084), .A(n4116), .ZN(n4086) );
  NAND2_X1 U4746 ( .A1(n4086), .A2(n4589), .ZN(n4113) );
  INV_X1 U4747 ( .A(n4087), .ZN(n4088) );
  AOI21_X1 U4748 ( .B1(n4597), .B2(ADDR_REG_16__SCAN_IN), .A(n4088), .ZN(n4112) );
  NAND2_X1 U4749 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4089), .ZN(n4100) );
  AOI22_X1 U4750 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4089), .B1(n4648), .B2(
        n3574), .ZN(n4532) );
  AOI22_X1 U4751 ( .A1(n4651), .A2(REG2_REG_9__SCAN_IN), .B1(n4096), .B2(n4516), .ZN(n4513) );
  INV_X1 U4752 ( .A(n4654), .ZN(n4093) );
  NAND2_X1 U4753 ( .A1(n4094), .A2(n4093), .ZN(n4095) );
  XNOR2_X1 U4754 ( .A(n4094), .B(n4654), .ZN(n4504) );
  NAND2_X1 U4755 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4504), .ZN(n4503) );
  NAND2_X1 U4756 ( .A1(n4098), .A2(n4097), .ZN(n4099) );
  NAND2_X1 U4757 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4523), .ZN(n4522) );
  NAND2_X1 U4758 ( .A1(n4099), .A2(n4522), .ZN(n4531) );
  NAND2_X1 U4759 ( .A1(n4532), .A2(n4531), .ZN(n4530) );
  NAND2_X1 U4760 ( .A1(n4100), .A2(n4530), .ZN(n4101) );
  NAND2_X1 U4761 ( .A1(n4645), .A2(n4101), .ZN(n4102) );
  XNOR2_X1 U4762 ( .A(n4101), .B(n4544), .ZN(n4541) );
  NAND2_X1 U4763 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4541), .ZN(n4540) );
  INV_X1 U4764 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4550) );
  NAND2_X1 U4765 ( .A1(n4550), .A2(n4556), .ZN(n4103) );
  NOR2_X1 U4766 ( .A1(n4104), .A2(n4079), .ZN(n4105) );
  AOI22_X1 U4767 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4641), .B1(n4106), .B2(
        n3319), .ZN(n4576) );
  AND2_X1 U4768 ( .A1(n4106), .A2(REG2_REG_15__SCAN_IN), .ZN(n4107) );
  XNOR2_X1 U4769 ( .A(n4125), .B(n4444), .ZN(n4108) );
  NAND2_X1 U4770 ( .A1(n4108), .A2(n3367), .ZN(n4126) );
  OAI21_X1 U4771 ( .B1(n4108), .B2(n3367), .A(n4126), .ZN(n4109) );
  NAND2_X1 U4772 ( .A1(n4109), .A2(n4608), .ZN(n4111) );
  NAND2_X1 U4773 ( .A1(n4566), .A2(n4444), .ZN(n4110) );
  NAND4_X1 U4774 ( .A1(n4113), .A2(n4112), .A3(n4111), .A4(n4110), .ZN(U3256)
         );
  AOI22_X1 U4775 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4638), .B1(n4128), .B2(
        n4114), .ZN(n4595) );
  INV_X1 U4776 ( .A(n4444), .ZN(n4124) );
  NAND2_X1 U4777 ( .A1(n4115), .A2(n4124), .ZN(n4117) );
  NAND2_X1 U4778 ( .A1(n4117), .A2(n4116), .ZN(n4582) );
  INV_X1 U4779 ( .A(n4592), .ZN(n4639) );
  AOI22_X1 U4780 ( .A1(n4639), .A2(REG1_REG_17__SCAN_IN), .B1(n4118), .B2(
        n4592), .ZN(n4583) );
  NOR2_X1 U4781 ( .A1(n4595), .A2(n4596), .ZN(n4593) );
  AOI21_X1 U4782 ( .B1(REG1_REG_18__SCAN_IN), .B2(n4128), .A(n4593), .ZN(n4121) );
  XNOR2_X1 U4783 ( .A(n4132), .B(n4390), .ZN(n4120) );
  XNOR2_X1 U4784 ( .A(n4121), .B(n4120), .ZN(n4136) );
  NAND2_X1 U4785 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4128), .ZN(n4122) );
  OAI21_X1 U4786 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4128), .A(n4122), .ZN(n4606) );
  NOR2_X1 U4787 ( .A1(n4639), .A2(REG2_REG_17__SCAN_IN), .ZN(n4123) );
  AOI21_X1 U4788 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4639), .A(n4123), .ZN(n4586) );
  NAND2_X1 U4789 ( .A1(n4125), .A2(n4124), .ZN(n4127) );
  NAND2_X1 U4790 ( .A1(n4127), .A2(n4126), .ZN(n4585) );
  NAND2_X1 U4791 ( .A1(n4586), .A2(n4585), .ZN(n4584) );
  XNOR2_X1 U4792 ( .A(n4132), .B(REG2_REG_19__SCAN_IN), .ZN(n4129) );
  NAND2_X1 U4793 ( .A1(n4597), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4130) );
  OAI211_X1 U4794 ( .C1(n4611), .C2(n4132), .A(n4131), .B(n4130), .ZN(n4133)
         );
  AOI21_X1 U4795 ( .B1(n4134), .B2(n4608), .A(n4133), .ZN(n4135) );
  OAI21_X1 U4796 ( .B1(n4136), .B2(n4594), .A(n4135), .ZN(U3259) );
  INV_X1 U4797 ( .A(n4153), .ZN(n4140) );
  XNOR2_X1 U4798 ( .A(n4141), .B(n4140), .ZN(n4351) );
  INV_X1 U4799 ( .A(n4351), .ZN(n4160) );
  NAND2_X1 U4800 ( .A1(n4142), .A2(n4147), .ZN(n4345) );
  INV_X1 U4801 ( .A(n4352), .ZN(n4143) );
  AOI22_X1 U4802 ( .A1(n4143), .A2(n4624), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4479), .ZN(n4159) );
  INV_X1 U4803 ( .A(B_REG_SCAN_IN), .ZN(n4144) );
  NOR2_X1 U4804 ( .A1(n4145), .A2(n4144), .ZN(n4146) );
  OR2_X1 U4805 ( .A1(n4321), .A2(n4146), .ZN(n4340) );
  OAI22_X1 U4806 ( .A1(n4148), .A2(n4340), .B1(n4320), .B2(n4147), .ZN(n4154)
         );
  INV_X1 U4807 ( .A(n4149), .ZN(n4150) );
  OAI21_X1 U4808 ( .B1(n4156), .B2(n4155), .A(n4353), .ZN(n4157) );
  NAND2_X1 U4809 ( .A1(n4157), .A2(n3575), .ZN(n4158) );
  OAI211_X1 U4810 ( .C1(n4160), .C2(n4338), .A(n4159), .B(n4158), .ZN(U3354)
         );
  XNOR2_X1 U4811 ( .A(n4161), .B(n4165), .ZN(n4355) );
  INV_X1 U4812 ( .A(n4355), .ZN(n4177) );
  OAI22_X1 U4813 ( .A1(n4162), .A2(n4277), .B1(n4171), .B2(n4320), .ZN(n4168)
         );
  AOI21_X1 U4814 ( .B1(n4165), .B2(n4164), .A(n4163), .ZN(n4166) );
  NOR2_X1 U4815 ( .A1(n4166), .A2(n4327), .ZN(n4167) );
  AOI211_X1 U4816 ( .C1(n4298), .C2(n4169), .A(n4168), .B(n4167), .ZN(n4356)
         );
  INV_X1 U4817 ( .A(n4356), .ZN(n4175) );
  OAI21_X1 U4818 ( .B1(n4187), .B2(n4171), .A(n4170), .ZN(n4358) );
  AOI22_X1 U4819 ( .A1(n4172), .A2(n4619), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4479), .ZN(n4173) );
  OAI21_X1 U4820 ( .B1(n4358), .B2(n4335), .A(n4173), .ZN(n4174) );
  AOI21_X1 U4821 ( .B1(n4175), .B2(n3575), .A(n4174), .ZN(n4176) );
  OAI21_X1 U4822 ( .B1(n4177), .B2(n4338), .A(n4176), .ZN(U3263) );
  XNOR2_X1 U4823 ( .A(n4178), .B(n4180), .ZN(n4360) );
  INV_X1 U4824 ( .A(n4360), .ZN(n4194) );
  NOR2_X1 U4825 ( .A1(n2079), .A2(n4179), .ZN(n4181) );
  XNOR2_X1 U4826 ( .A(n4181), .B(n4180), .ZN(n4186) );
  OAI22_X1 U4827 ( .A1(n4182), .A2(n4277), .B1(n4189), .B2(n4320), .ZN(n4183)
         );
  AOI21_X1 U4828 ( .B1(n4298), .B2(n4184), .A(n4183), .ZN(n4185) );
  OAI21_X1 U4829 ( .B1(n4186), .B2(n4327), .A(n4185), .ZN(n4359) );
  INV_X1 U4830 ( .A(n4187), .ZN(n4188) );
  OAI21_X1 U4831 ( .B1(n4207), .B2(n4189), .A(n4188), .ZN(n4413) );
  AOI22_X1 U4832 ( .A1(n4190), .A2(n4619), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4479), .ZN(n4191) );
  OAI21_X1 U4833 ( .B1(n4413), .B2(n4335), .A(n4191), .ZN(n4192) );
  AOI21_X1 U4834 ( .B1(n4359), .B2(n3575), .A(n4192), .ZN(n4193) );
  OAI21_X1 U4835 ( .B1(n4194), .B2(n4338), .A(n4193), .ZN(U3264) );
  OAI22_X1 U4836 ( .A1(n4195), .A2(n4197), .B1(n4196), .B2(n4242), .ZN(n4198)
         );
  XNOR2_X1 U4837 ( .A(n4198), .B(n4199), .ZN(n4366) );
  XNOR2_X1 U4838 ( .A(n4200), .B(n4199), .ZN(n4206) );
  OAI22_X1 U4839 ( .A1(n4202), .A2(n4277), .B1(n4201), .B2(n4320), .ZN(n4203)
         );
  AOI21_X1 U4840 ( .B1(n4298), .B2(n4204), .A(n4203), .ZN(n4205) );
  OAI21_X1 U4841 ( .B1(n4206), .B2(n4327), .A(n4205), .ZN(n4363) );
  AOI21_X1 U4842 ( .B1(n4208), .B2(n4223), .A(n4207), .ZN(n4364) );
  INV_X1 U4843 ( .A(n4364), .ZN(n4211) );
  AOI22_X1 U4844 ( .A1(n4209), .A2(n4619), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4479), .ZN(n4210) );
  OAI21_X1 U4845 ( .B1(n4211), .B2(n4335), .A(n4210), .ZN(n4212) );
  AOI21_X1 U4846 ( .B1(n4363), .B2(n3575), .A(n4212), .ZN(n4213) );
  OAI21_X1 U4847 ( .B1(n4366), .B2(n4338), .A(n4213), .ZN(U3265) );
  XNOR2_X1 U4848 ( .A(n4195), .B(n4216), .ZN(n4368) );
  INV_X1 U4849 ( .A(n4368), .ZN(n4230) );
  NOR2_X1 U4850 ( .A1(n4215), .A2(n4214), .ZN(n4217) );
  XNOR2_X1 U4851 ( .A(n4217), .B(n4216), .ZN(n4222) );
  OAI22_X1 U4852 ( .A1(n4218), .A2(n4277), .B1(n4320), .B2(n4224), .ZN(n4219)
         );
  AOI21_X1 U4853 ( .B1(n4220), .B2(n4298), .A(n4219), .ZN(n4221) );
  OAI21_X1 U4854 ( .B1(n4222), .B2(n4327), .A(n4221), .ZN(n4367) );
  OAI21_X1 U4855 ( .B1(n2108), .B2(n4224), .A(n4223), .ZN(n4418) );
  INV_X1 U4856 ( .A(n4225), .ZN(n4226) );
  AOI22_X1 U4857 ( .A1(n4479), .A2(REG2_REG_24__SCAN_IN), .B1(n4226), .B2(
        n4619), .ZN(n4227) );
  OAI21_X1 U4858 ( .B1(n4418), .B2(n4335), .A(n4227), .ZN(n4228) );
  AOI21_X1 U4859 ( .B1(n4367), .B2(n3575), .A(n4228), .ZN(n4229) );
  OAI21_X1 U4860 ( .B1(n4230), .B2(n4338), .A(n4229), .ZN(U3266) );
  XNOR2_X1 U4861 ( .A(n4231), .B(n4238), .ZN(n4372) );
  INV_X1 U4862 ( .A(n4372), .ZN(n4253) );
  AOI21_X1 U4863 ( .B1(n4294), .B2(n4235), .A(n4234), .ZN(n4276) );
  NOR2_X1 U4864 ( .A1(n4276), .A2(n4275), .ZN(n4274) );
  NOR2_X1 U4865 ( .A1(n4274), .A2(n4236), .ZN(n4259) );
  NOR2_X1 U4866 ( .A1(n4259), .A2(n4258), .ZN(n4257) );
  NOR2_X1 U4867 ( .A1(n4257), .A2(n4237), .ZN(n4239) );
  XNOR2_X1 U4868 ( .A(n4239), .B(n4238), .ZN(n4244) );
  OAI22_X1 U4869 ( .A1(n4240), .A2(n4277), .B1(n4320), .B2(n4246), .ZN(n4241)
         );
  AOI21_X1 U4870 ( .B1(n4242), .B2(n4298), .A(n4241), .ZN(n4243) );
  OAI21_X1 U4871 ( .B1(n4244), .B2(n4327), .A(n4243), .ZN(n4371) );
  INV_X1 U4872 ( .A(n4375), .ZN(n4247) );
  OAI21_X1 U4873 ( .B1(n4247), .B2(n4246), .A(n4245), .ZN(n4422) );
  INV_X1 U4874 ( .A(n4248), .ZN(n4249) );
  AOI22_X1 U4875 ( .A1(n4479), .A2(REG2_REG_23__SCAN_IN), .B1(n4249), .B2(
        n4619), .ZN(n4250) );
  OAI21_X1 U4876 ( .B1(n4422), .B2(n4335), .A(n4250), .ZN(n4251) );
  AOI21_X1 U4877 ( .B1(n4371), .B2(n3575), .A(n4251), .ZN(n4252) );
  OAI21_X1 U4878 ( .B1(n4253), .B2(n4338), .A(n4252), .ZN(U3267) );
  OAI21_X1 U4879 ( .B1(n4255), .B2(n4258), .A(n4254), .ZN(n4379) );
  OAI22_X1 U4880 ( .A1(n4256), .A2(n4277), .B1(n4267), .B2(n4320), .ZN(n4262)
         );
  AOI21_X1 U4881 ( .B1(n4259), .B2(n4258), .A(n4257), .ZN(n4260) );
  NOR2_X1 U4882 ( .A1(n4260), .A2(n4327), .ZN(n4261) );
  AOI211_X1 U4883 ( .C1(n4298), .C2(n4263), .A(n4262), .B(n4261), .ZN(n4378)
         );
  INV_X1 U4884 ( .A(n4264), .ZN(n4265) );
  AOI22_X1 U4885 ( .A1(n4479), .A2(REG2_REG_22__SCAN_IN), .B1(n4265), .B2(
        n4619), .ZN(n4270) );
  INV_X1 U4886 ( .A(n4266), .ZN(n4282) );
  INV_X1 U4887 ( .A(n4267), .ZN(n4268) );
  NAND2_X1 U4888 ( .A1(n4282), .A2(n4268), .ZN(n4376) );
  NAND3_X1 U4889 ( .A1(n4376), .A2(n4624), .A3(n4375), .ZN(n4269) );
  OAI211_X1 U4890 ( .C1(n4378), .C2(n4479), .A(n4270), .B(n4269), .ZN(n4271)
         );
  INV_X1 U4891 ( .A(n4271), .ZN(n4272) );
  OAI21_X1 U4892 ( .B1(n4379), .B2(n4338), .A(n4272), .ZN(U3268) );
  XNOR2_X1 U4893 ( .A(n4273), .B(n4275), .ZN(n4381) );
  INV_X1 U4894 ( .A(n4381), .ZN(n4290) );
  AOI21_X1 U4895 ( .B1(n4276), .B2(n4275), .A(n4274), .ZN(n4281) );
  OAI22_X1 U4896 ( .A1(n4322), .A2(n4277), .B1(n4283), .B2(n4320), .ZN(n4278)
         );
  AOI21_X1 U4897 ( .B1(n4298), .B2(n4279), .A(n4278), .ZN(n4280) );
  OAI21_X1 U4898 ( .B1(n4281), .B2(n4327), .A(n4280), .ZN(n4380) );
  INV_X1 U4899 ( .A(n4304), .ZN(n4284) );
  OAI21_X1 U4900 ( .B1(n4284), .B2(n4283), .A(n4282), .ZN(n4427) );
  INV_X1 U4901 ( .A(n4285), .ZN(n4286) );
  AOI22_X1 U4902 ( .A1(n4479), .A2(REG2_REG_21__SCAN_IN), .B1(n4286), .B2(
        n4619), .ZN(n4287) );
  OAI21_X1 U4903 ( .B1(n4427), .B2(n4335), .A(n4287), .ZN(n4288) );
  AOI21_X1 U4904 ( .B1(n4380), .B2(n3575), .A(n4288), .ZN(n4289) );
  OAI21_X1 U4905 ( .B1(n4290), .B2(n4338), .A(n4289), .ZN(U3269) );
  XNOR2_X1 U4906 ( .A(n4291), .B(n4295), .ZN(n4385) );
  INV_X1 U4907 ( .A(n4385), .ZN(n4312) );
  INV_X1 U4908 ( .A(n4292), .ZN(n4293) );
  NOR2_X1 U4909 ( .A1(n4294), .A2(n4293), .ZN(n4296) );
  XNOR2_X1 U4910 ( .A(n4296), .B(n4295), .ZN(n4303) );
  NOR2_X1 U4911 ( .A1(n4320), .A2(n4305), .ZN(n4297) );
  AOI21_X1 U4912 ( .B1(n4299), .B2(n4298), .A(n4297), .ZN(n4302) );
  NAND2_X1 U4913 ( .A1(n4300), .A2(n4325), .ZN(n4301) );
  OAI211_X1 U4914 ( .C1(n4303), .C2(n4327), .A(n4302), .B(n4301), .ZN(n4384)
         );
  INV_X1 U4915 ( .A(n4329), .ZN(n4306) );
  OAI21_X1 U4916 ( .B1(n4306), .B2(n4305), .A(n4304), .ZN(n4431) );
  INV_X1 U4917 ( .A(n4307), .ZN(n4308) );
  AOI22_X1 U4918 ( .A1(n4479), .A2(REG2_REG_20__SCAN_IN), .B1(n4308), .B2(
        n4619), .ZN(n4309) );
  OAI21_X1 U4919 ( .B1(n4431), .B2(n4335), .A(n4309), .ZN(n4310) );
  AOI21_X1 U4920 ( .B1(n4384), .B2(n3575), .A(n4310), .ZN(n4311) );
  OAI21_X1 U4921 ( .B1(n4312), .B2(n4338), .A(n4311), .ZN(U3270) );
  XNOR2_X1 U4922 ( .A(n4313), .B(n4318), .ZN(n4389) );
  INV_X1 U4923 ( .A(n4389), .ZN(n4339) );
  INV_X1 U4924 ( .A(n4314), .ZN(n4315) );
  AOI21_X1 U4925 ( .B1(n4317), .B2(n4316), .A(n4315), .ZN(n4319) );
  XNOR2_X1 U4926 ( .A(n4319), .B(n4318), .ZN(n4328) );
  OAI22_X1 U4927 ( .A1(n4322), .A2(n4321), .B1(n4320), .B2(n4330), .ZN(n4323)
         );
  AOI21_X1 U4928 ( .B1(n4325), .B2(n4324), .A(n4323), .ZN(n4326) );
  OAI21_X1 U4929 ( .B1(n4328), .B2(n4327), .A(n4326), .ZN(n4388) );
  OAI21_X1 U4930 ( .B1(n4331), .B2(n4330), .A(n4329), .ZN(n4436) );
  INV_X1 U4931 ( .A(n4332), .ZN(n4333) );
  AOI22_X1 U4932 ( .A1(n4479), .A2(REG2_REG_19__SCAN_IN), .B1(n4333), .B2(
        n4619), .ZN(n4334) );
  OAI21_X1 U4933 ( .B1(n4436), .B2(n4335), .A(n4334), .ZN(n4336) );
  AOI21_X1 U4934 ( .B1(n4388), .B2(n3575), .A(n4336), .ZN(n4337) );
  OAI21_X1 U4935 ( .B1(n4339), .B2(n4338), .A(n4337), .ZN(U3271) );
  XNOR2_X1 U4936 ( .A(n4344), .B(n4342), .ZN(n4473) );
  INV_X1 U4937 ( .A(n4473), .ZN(n4404) );
  NOR2_X1 U4938 ( .A1(n4341), .A2(n4340), .ZN(n4346) );
  AOI21_X1 U4939 ( .B1(n4342), .B2(n4347), .A(n4346), .ZN(n4475) );
  MUX2_X1 U4940 ( .A(n3697), .B(n4475), .S(n4716), .Z(n4343) );
  OAI21_X1 U4941 ( .B1(n4404), .B2(n4392), .A(n4343), .ZN(U3549) );
  AOI21_X1 U4942 ( .B1(n4348), .B2(n4345), .A(n4344), .ZN(n4476) );
  INV_X1 U4943 ( .A(n4476), .ZN(n4407) );
  INV_X1 U4944 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4349) );
  AOI21_X1 U4945 ( .B1(n4348), .B2(n4347), .A(n4346), .ZN(n4478) );
  MUX2_X1 U4946 ( .A(n4349), .B(n4478), .S(n4716), .Z(n4350) );
  OAI21_X1 U4947 ( .B1(n4407), .B2(n4392), .A(n4350), .ZN(U3548) );
  MUX2_X1 U4948 ( .A(REG1_REG_29__SCAN_IN), .B(n4408), .S(n4716), .Z(U3547) );
  NAND2_X1 U4949 ( .A1(n4355), .A2(n4694), .ZN(n4357) );
  OAI211_X1 U4950 ( .C1(n4698), .C2(n4358), .A(n4357), .B(n4356), .ZN(n4409)
         );
  MUX2_X1 U4951 ( .A(REG1_REG_27__SCAN_IN), .B(n4409), .S(n4716), .Z(U3545) );
  AOI21_X1 U4952 ( .B1(n4360), .B2(n4694), .A(n4359), .ZN(n4410) );
  MUX2_X1 U4953 ( .A(n4361), .B(n4410), .S(n4716), .Z(n4362) );
  OAI21_X1 U4954 ( .B1(n4392), .B2(n4413), .A(n4362), .ZN(U3544) );
  AOI21_X1 U4955 ( .B1(n2707), .B2(n4364), .A(n4363), .ZN(n4365) );
  OAI21_X1 U4956 ( .B1(n4366), .B2(n4678), .A(n4365), .ZN(n4414) );
  MUX2_X1 U4957 ( .A(REG1_REG_25__SCAN_IN), .B(n4414), .S(n4716), .Z(U3543) );
  AOI21_X1 U4958 ( .B1(n4368), .B2(n4694), .A(n4367), .ZN(n4415) );
  MUX2_X1 U4959 ( .A(n4369), .B(n4415), .S(n4716), .Z(n4370) );
  OAI21_X1 U4960 ( .B1(n4392), .B2(n4418), .A(n4370), .ZN(U3542) );
  AOI21_X1 U4961 ( .B1(n4372), .B2(n4694), .A(n4371), .ZN(n4419) );
  MUX2_X1 U4962 ( .A(n4373), .B(n4419), .S(n4716), .Z(n4374) );
  OAI21_X1 U4963 ( .B1(n4392), .B2(n4422), .A(n4374), .ZN(U3541) );
  NAND3_X1 U4964 ( .A1(n4376), .A2(n2707), .A3(n4375), .ZN(n4377) );
  OAI211_X1 U4965 ( .C1(n4379), .C2(n4678), .A(n4378), .B(n4377), .ZN(n4423)
         );
  MUX2_X1 U4966 ( .A(REG1_REG_22__SCAN_IN), .B(n4423), .S(n4716), .Z(U3540) );
  AOI21_X1 U4967 ( .B1(n4381), .B2(n4694), .A(n4380), .ZN(n4424) );
  MUX2_X1 U4968 ( .A(n4382), .B(n4424), .S(n4716), .Z(n4383) );
  OAI21_X1 U4969 ( .B1(n4392), .B2(n4427), .A(n4383), .ZN(U3539) );
  INV_X1 U4970 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4386) );
  AOI21_X1 U4971 ( .B1(n4385), .B2(n4694), .A(n4384), .ZN(n4428) );
  MUX2_X1 U4972 ( .A(n4386), .B(n4428), .S(n4716), .Z(n4387) );
  OAI21_X1 U4973 ( .B1(n4392), .B2(n4431), .A(n4387), .ZN(U3538) );
  AOI21_X1 U4974 ( .B1(n4389), .B2(n4694), .A(n4388), .ZN(n4432) );
  MUX2_X1 U4975 ( .A(n4390), .B(n4432), .S(n4716), .Z(n4391) );
  OAI21_X1 U4976 ( .B1(n4392), .B2(n4436), .A(n4391), .ZN(U3537) );
  AOI211_X1 U4977 ( .C1(n4395), .C2(n4694), .A(n4394), .B(n4393), .ZN(n4396)
         );
  INV_X1 U4978 ( .A(n4396), .ZN(n4437) );
  MUX2_X1 U4979 ( .A(REG1_REG_18__SCAN_IN), .B(n4437), .S(n4716), .Z(U3536) );
  NAND3_X1 U4980 ( .A1(n4398), .A2(n2707), .A3(n4397), .ZN(n4399) );
  OAI211_X1 U4981 ( .C1(n4401), .C2(n4678), .A(n4400), .B(n4399), .ZN(n4438)
         );
  MUX2_X1 U4982 ( .A(REG1_REG_16__SCAN_IN), .B(n4438), .S(n4716), .Z(U3534) );
  INV_X1 U4983 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4402) );
  MUX2_X1 U4984 ( .A(n4402), .B(n4475), .S(n4705), .Z(n4403) );
  OAI21_X1 U4985 ( .B1(n4404), .B2(n4435), .A(n4403), .ZN(U3517) );
  INV_X1 U4986 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4405) );
  MUX2_X1 U4987 ( .A(n4405), .B(n4478), .S(n4705), .Z(n4406) );
  OAI21_X1 U4988 ( .B1(n4407), .B2(n4435), .A(n4406), .ZN(U3516) );
  MUX2_X1 U4989 ( .A(REG0_REG_29__SCAN_IN), .B(n4408), .S(n4705), .Z(U3515) );
  MUX2_X1 U4990 ( .A(REG0_REG_27__SCAN_IN), .B(n4409), .S(n4705), .Z(U3513) );
  INV_X1 U4991 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4411) );
  MUX2_X1 U4992 ( .A(n4411), .B(n4410), .S(n4705), .Z(n4412) );
  OAI21_X1 U4993 ( .B1(n4413), .B2(n4435), .A(n4412), .ZN(U3512) );
  MUX2_X1 U4994 ( .A(REG0_REG_25__SCAN_IN), .B(n4414), .S(n4705), .Z(U3511) );
  INV_X1 U4995 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4416) );
  MUX2_X1 U4996 ( .A(n4416), .B(n4415), .S(n4705), .Z(n4417) );
  OAI21_X1 U4997 ( .B1(n4418), .B2(n4435), .A(n4417), .ZN(U3510) );
  INV_X1 U4998 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4420) );
  MUX2_X1 U4999 ( .A(n4420), .B(n4419), .S(n4705), .Z(n4421) );
  OAI21_X1 U5000 ( .B1(n4422), .B2(n4435), .A(n4421), .ZN(U3509) );
  MUX2_X1 U5001 ( .A(REG0_REG_22__SCAN_IN), .B(n4423), .S(n4705), .Z(U3508) );
  INV_X1 U5002 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4425) );
  MUX2_X1 U5003 ( .A(n4425), .B(n4424), .S(n4705), .Z(n4426) );
  OAI21_X1 U5004 ( .B1(n4427), .B2(n4435), .A(n4426), .ZN(U3507) );
  INV_X1 U5005 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4429) );
  MUX2_X1 U5006 ( .A(n4429), .B(n4428), .S(n4705), .Z(n4430) );
  OAI21_X1 U5007 ( .B1(n4431), .B2(n4435), .A(n4430), .ZN(U3506) );
  INV_X1 U5008 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4433) );
  MUX2_X1 U5009 ( .A(n4433), .B(n4432), .S(n4705), .Z(n4434) );
  OAI21_X1 U5010 ( .B1(n4436), .B2(n4435), .A(n4434), .ZN(U3505) );
  MUX2_X1 U5011 ( .A(REG0_REG_18__SCAN_IN), .B(n4437), .S(n4705), .Z(U3503) );
  MUX2_X1 U5012 ( .A(REG0_REG_16__SCAN_IN), .B(n4438), .S(n4705), .Z(U3499) );
  MUX2_X1 U5013 ( .A(n4439), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U5014 ( .A(n2322), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5015 ( .A(DATAI_28_), .B(n4440), .S(STATE_REG_SCAN_IN), .Z(U3324)
         );
  MUX2_X1 U5016 ( .A(DATAI_27_), .B(n4481), .S(STATE_REG_SCAN_IN), .Z(U3325)
         );
  MUX2_X1 U5017 ( .A(n4441), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5018 ( .A(n2680), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U5019 ( .A(DATAI_22_), .B(n4442), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U5020 ( .A(DATAI_19_), .B(n4443), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U5021 ( .A(n4444), .B(DATAI_16_), .S(U3149), .Z(U3336) );
  MUX2_X1 U5022 ( .A(DATAI_7_), .B(n4445), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U5023 ( .A(n4446), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5024 ( .A(n4447), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5025 ( .A(DATAI_4_), .B(n4448), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5026 ( .A(n4449), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5027 ( .A(DATAI_2_), .B(n4450), .S(STATE_REG_SCAN_IN), .Z(U3350) );
  MUX2_X1 U5028 ( .A(n4451), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  NOR2_X1 U5029 ( .A1(STATE_REG_SCAN_IN), .A2(n4452), .ZN(n4574) );
  AOI21_X1 U5030 ( .B1(n4454), .B2(n4453), .A(n4574), .ZN(n4458) );
  NAND2_X1 U5031 ( .A1(n4456), .A2(n4455), .ZN(n4457) );
  OAI211_X1 U5032 ( .C1(n4460), .C2(n4459), .A(n4458), .B(n4457), .ZN(n4461)
         );
  INV_X1 U5033 ( .A(n4461), .ZN(n4470) );
  INV_X1 U5034 ( .A(n4464), .ZN(n4468) );
  AOI21_X1 U5035 ( .B1(n4462), .B2(n4464), .A(n4463), .ZN(n4466) );
  NOR2_X1 U5036 ( .A1(n4466), .A2(n4465), .ZN(n4467) );
  OAI21_X1 U5037 ( .B1(n4468), .B2(n3442), .A(n4467), .ZN(n4469) );
  OAI211_X1 U5038 ( .C1(n4472), .C2(n4471), .A(n4470), .B(n4469), .ZN(U3238)
         );
  AOI22_X1 U5039 ( .A1(n4473), .A2(n4624), .B1(n4479), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n4474) );
  OAI21_X1 U5040 ( .B1(n4479), .B2(n4475), .A(n4474), .ZN(U3260) );
  AOI22_X1 U5041 ( .A1(n4476), .A2(n4624), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4479), .ZN(n4477) );
  OAI21_X1 U5042 ( .B1(n4479), .B2(n4478), .A(n4477), .ZN(U3261) );
  OAI21_X1 U5043 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4481), .A(n4480), .ZN(n4482)
         );
  XNOR2_X1 U5044 ( .A(n4482), .B(n2103), .ZN(n4485) );
  AOI22_X1 U5045 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4597), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4483) );
  OAI21_X1 U5046 ( .B1(n4485), .B2(n4484), .A(n4483), .ZN(U3240) );
  XNOR2_X1 U5047 ( .A(n4486), .B(REG1_REG_4__SCAN_IN), .ZN(n4487) );
  OR2_X1 U5048 ( .A1(n4594), .A2(n4487), .ZN(n4490) );
  AOI21_X1 U5049 ( .B1(n4597), .B2(ADDR_REG_4__SCAN_IN), .A(n4488), .ZN(n4489)
         );
  OAI211_X1 U5050 ( .C1(n4611), .C2(n4491), .A(n4490), .B(n4489), .ZN(n4495)
         );
  XNOR2_X1 U5051 ( .A(n4492), .B(REG2_REG_4__SCAN_IN), .ZN(n4493) );
  NOR2_X1 U5052 ( .A1(n4560), .A2(n4493), .ZN(n4494) );
  NOR2_X1 U5053 ( .A1(n4495), .A2(n4494), .ZN(n4497) );
  NAND2_X1 U5054 ( .A1(n4497), .A2(n4496), .ZN(U3244) );
  AOI211_X1 U5055 ( .C1(n2411), .C2(n4499), .A(n4498), .B(n4594), .ZN(n4502)
         );
  INV_X1 U5056 ( .A(n4500), .ZN(n4501) );
  AOI211_X1 U5057 ( .C1(n4597), .C2(ADDR_REG_8__SCAN_IN), .A(n4502), .B(n4501), 
        .ZN(n4506) );
  OAI211_X1 U5058 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4504), .A(n4608), .B(n4503), 
        .ZN(n4505) );
  OAI211_X1 U5059 ( .C1(n4611), .C2(n4654), .A(n4506), .B(n4505), .ZN(U3248)
         );
  AOI211_X1 U5060 ( .C1(n2091), .C2(n4508), .A(n4507), .B(n4594), .ZN(n4510)
         );
  AOI211_X1 U5061 ( .C1(n4597), .C2(ADDR_REG_9__SCAN_IN), .A(n4510), .B(n4509), 
        .ZN(n4515) );
  OAI211_X1 U5062 ( .C1(n4513), .C2(n4512), .A(n4608), .B(n4511), .ZN(n4514)
         );
  OAI211_X1 U5063 ( .C1(n4611), .C2(n4516), .A(n4515), .B(n4514), .ZN(U3249)
         );
  AOI211_X1 U5064 ( .C1(n4519), .C2(n4518), .A(n4517), .B(n4594), .ZN(n4520)
         );
  AOI211_X1 U5065 ( .C1(n4597), .C2(ADDR_REG_10__SCAN_IN), .A(n4521), .B(n4520), .ZN(n4525) );
  OAI211_X1 U5066 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4523), .A(n4608), .B(n4522), .ZN(n4524) );
  OAI211_X1 U5067 ( .C1(n4611), .C2(n4650), .A(n4525), .B(n4524), .ZN(U3250)
         );
  AOI211_X1 U5068 ( .C1(n2092), .C2(n4527), .A(n4526), .B(n4594), .ZN(n4529)
         );
  AOI211_X1 U5069 ( .C1(n4597), .C2(ADDR_REG_11__SCAN_IN), .A(n4529), .B(n4528), .ZN(n4534) );
  OAI211_X1 U5070 ( .C1(n4532), .C2(n4531), .A(n4608), .B(n4530), .ZN(n4533)
         );
  OAI211_X1 U5071 ( .C1(n4611), .C2(n4648), .A(n4534), .B(n4533), .ZN(U3251)
         );
  AOI211_X1 U5072 ( .C1(n4537), .C2(n4536), .A(n4535), .B(n4594), .ZN(n4539)
         );
  AOI211_X1 U5073 ( .C1(n4597), .C2(ADDR_REG_12__SCAN_IN), .A(n4539), .B(n4538), .ZN(n4543) );
  OAI211_X1 U5074 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4541), .A(n4608), .B(n4540), .ZN(n4542) );
  OAI211_X1 U5075 ( .C1(n4611), .C2(n4544), .A(n4543), .B(n4542), .ZN(U3252)
         );
  AOI211_X1 U5076 ( .C1(n4547), .C2(n4546), .A(n4545), .B(n4594), .ZN(n4549)
         );
  AOI211_X1 U5077 ( .C1(n4597), .C2(ADDR_REG_13__SCAN_IN), .A(n4549), .B(n4548), .ZN(n4555) );
  AOI22_X1 U5078 ( .A1(REG2_REG_13__SCAN_IN), .A2(n4643), .B1(n4556), .B2(
        n4550), .ZN(n4553) );
  AOI21_X1 U5079 ( .B1(n4553), .B2(n4552), .A(n4560), .ZN(n4551) );
  OAI21_X1 U5080 ( .B1(n4553), .B2(n4552), .A(n4551), .ZN(n4554) );
  OAI211_X1 U5081 ( .C1(n4611), .C2(n4556), .A(n4555), .B(n4554), .ZN(U3253)
         );
  INV_X1 U5082 ( .A(n4597), .ZN(n4570) );
  AOI211_X1 U5083 ( .C1(n4559), .C2(n4558), .A(n4557), .B(n4594), .ZN(n4564)
         );
  AOI211_X1 U5084 ( .C1(n3238), .C2(n4562), .A(n4561), .B(n4560), .ZN(n4563)
         );
  AOI211_X1 U5085 ( .C1(n4566), .C2(n4565), .A(n4564), .B(n4563), .ZN(n4568)
         );
  OAI211_X1 U5086 ( .C1(n4570), .C2(n4569), .A(n4568), .B(n4567), .ZN(U3254)
         );
  AOI211_X1 U5087 ( .C1(n2082), .C2(n4572), .A(n4571), .B(n4594), .ZN(n4573)
         );
  AOI211_X1 U5088 ( .C1(n4597), .C2(ADDR_REG_15__SCAN_IN), .A(n4574), .B(n4573), .ZN(n4579) );
  AOI21_X1 U5089 ( .B1(n4576), .B2(n2080), .A(n4575), .ZN(n4577) );
  NAND2_X1 U5090 ( .A1(n4608), .A2(n4577), .ZN(n4578) );
  OAI211_X1 U5091 ( .C1(n4611), .C2(n4641), .A(n4579), .B(n4578), .ZN(U3255)
         );
  AOI21_X1 U5092 ( .B1(n4597), .B2(ADDR_REG_17__SCAN_IN), .A(n4580), .ZN(n4591) );
  OAI21_X1 U5093 ( .B1(n4583), .B2(n4582), .A(n4581), .ZN(n4588) );
  OAI21_X1 U5094 ( .B1(n4586), .B2(n4585), .A(n4584), .ZN(n4587) );
  AOI22_X1 U5095 ( .A1(n4589), .A2(n4588), .B1(n4608), .B2(n4587), .ZN(n4590)
         );
  OAI211_X1 U5096 ( .C1(n4592), .C2(n4611), .A(n4591), .B(n4590), .ZN(U3257)
         );
  NAND2_X1 U5097 ( .A1(n4597), .A2(ADDR_REG_18__SCAN_IN), .ZN(n4600) );
  AOI21_X1 U5098 ( .B1(n4606), .B2(n4605), .A(n4604), .ZN(n4607) );
  NAND2_X1 U5099 ( .A1(n4608), .A2(n4607), .ZN(n4609) );
  OAI211_X1 U5100 ( .C1(n4611), .C2(n4638), .A(n4610), .B(n4609), .ZN(U3258)
         );
  AOI22_X1 U5101 ( .A1(n4612), .A2(n4619), .B1(REG2_REG_6__SCAN_IN), .B2(n4479), .ZN(n4617) );
  INV_X1 U5102 ( .A(n4613), .ZN(n4614) );
  AOI22_X1 U5103 ( .A1(n4615), .A2(n4622), .B1(n4624), .B2(n4614), .ZN(n4616)
         );
  OAI211_X1 U5104 ( .C1(n4479), .C2(n4618), .A(n4617), .B(n4616), .ZN(U3284)
         );
  AOI22_X1 U5105 ( .A1(REG3_REG_2__SCAN_IN), .A2(n4619), .B1(
        REG2_REG_2__SCAN_IN), .B2(n4479), .ZN(n4626) );
  INV_X1 U5106 ( .A(n4620), .ZN(n4623) );
  AOI22_X1 U5107 ( .A1(n4624), .A2(n4623), .B1(n4622), .B2(n4621), .ZN(n4625)
         );
  OAI211_X1 U5108 ( .C1(n4479), .C2(n4627), .A(n4626), .B(n4625), .ZN(U3288)
         );
  INV_X1 U5109 ( .A(n4632), .ZN(n4634) );
  NOR2_X1 U5110 ( .A1(n4634), .A2(n4628), .ZN(U3291) );
  AND2_X1 U5111 ( .A1(D_REG_30__SCAN_IN), .A2(n4632), .ZN(U3292) );
  AND2_X1 U5112 ( .A1(D_REG_29__SCAN_IN), .A2(n4632), .ZN(U3293) );
  AND2_X1 U5113 ( .A1(D_REG_28__SCAN_IN), .A2(n4632), .ZN(U3294) );
  AND2_X1 U5114 ( .A1(D_REG_27__SCAN_IN), .A2(n4632), .ZN(U3295) );
  AND2_X1 U5115 ( .A1(D_REG_26__SCAN_IN), .A2(n4632), .ZN(U3296) );
  AND2_X1 U5116 ( .A1(D_REG_25__SCAN_IN), .A2(n4632), .ZN(U3297) );
  AND2_X1 U5117 ( .A1(D_REG_24__SCAN_IN), .A2(n4632), .ZN(U3298) );
  NOR2_X1 U5118 ( .A1(n4634), .A2(n4629), .ZN(U3299) );
  AND2_X1 U5119 ( .A1(D_REG_22__SCAN_IN), .A2(n4632), .ZN(U3300) );
  AND2_X1 U5120 ( .A1(D_REG_21__SCAN_IN), .A2(n4632), .ZN(U3301) );
  NOR2_X1 U5121 ( .A1(n4634), .A2(n4630), .ZN(U3302) );
  AND2_X1 U5122 ( .A1(n4632), .A2(D_REG_19__SCAN_IN), .ZN(U3303) );
  AND2_X1 U5123 ( .A1(D_REG_18__SCAN_IN), .A2(n4632), .ZN(U3304) );
  AND2_X1 U5124 ( .A1(D_REG_17__SCAN_IN), .A2(n4632), .ZN(U3305) );
  AND2_X1 U5125 ( .A1(D_REG_16__SCAN_IN), .A2(n4632), .ZN(U3306) );
  AND2_X1 U5126 ( .A1(D_REG_15__SCAN_IN), .A2(n4632), .ZN(U3307) );
  AND2_X1 U5127 ( .A1(D_REG_14__SCAN_IN), .A2(n4632), .ZN(U3308) );
  AND2_X1 U5128 ( .A1(D_REG_13__SCAN_IN), .A2(n4632), .ZN(U3309) );
  AND2_X1 U5129 ( .A1(D_REG_12__SCAN_IN), .A2(n4632), .ZN(U3310) );
  NOR2_X1 U5130 ( .A1(n4634), .A2(n4631), .ZN(U3311) );
  AND2_X1 U5131 ( .A1(D_REG_10__SCAN_IN), .A2(n4632), .ZN(U3312) );
  AND2_X1 U5132 ( .A1(D_REG_9__SCAN_IN), .A2(n4632), .ZN(U3313) );
  AND2_X1 U5133 ( .A1(D_REG_8__SCAN_IN), .A2(n4632), .ZN(U3314) );
  AND2_X1 U5134 ( .A1(D_REG_7__SCAN_IN), .A2(n4632), .ZN(U3315) );
  AND2_X1 U5135 ( .A1(n4632), .A2(D_REG_6__SCAN_IN), .ZN(U3316) );
  AND2_X1 U5136 ( .A1(D_REG_5__SCAN_IN), .A2(n4632), .ZN(U3317) );
  AND2_X1 U5137 ( .A1(D_REG_4__SCAN_IN), .A2(n4632), .ZN(U3318) );
  AND2_X1 U5138 ( .A1(D_REG_3__SCAN_IN), .A2(n4632), .ZN(U3319) );
  NOR2_X1 U5139 ( .A1(n4634), .A2(n4633), .ZN(U3320) );
  OAI21_X1 U5140 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4635), .ZN(
        n4636) );
  INV_X1 U5141 ( .A(n4636), .ZN(U3329) );
  AOI22_X1 U5142 ( .A1(STATE_REG_SCAN_IN), .A2(n4638), .B1(n4637), .B2(U3149), 
        .ZN(U3334) );
  OAI22_X1 U5143 ( .A1(U3149), .A2(n4639), .B1(DATAI_17_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4640) );
  INV_X1 U5144 ( .A(n4640), .ZN(U3335) );
  AOI22_X1 U5145 ( .A1(STATE_REG_SCAN_IN), .A2(n4641), .B1(n2494), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5146 ( .A(DATAI_14_), .ZN(n4642) );
  AOI22_X1 U5147 ( .A1(STATE_REG_SCAN_IN), .A2(n4079), .B1(n4642), .B2(U3149), 
        .ZN(U3338) );
  OAI22_X1 U5148 ( .A1(U3149), .A2(n4643), .B1(DATAI_13_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4644) );
  INV_X1 U5149 ( .A(n4644), .ZN(U3339) );
  OAI22_X1 U5150 ( .A1(U3149), .A2(n4645), .B1(DATAI_12_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4646) );
  INV_X1 U5151 ( .A(n4646), .ZN(U3340) );
  AOI22_X1 U5152 ( .A1(STATE_REG_SCAN_IN), .A2(n4648), .B1(n4647), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5153 ( .A(DATAI_10_), .ZN(n4649) );
  AOI22_X1 U5154 ( .A1(STATE_REG_SCAN_IN), .A2(n4650), .B1(n4649), .B2(U3149), 
        .ZN(U3342) );
  OAI22_X1 U5155 ( .A1(U3149), .A2(n4651), .B1(DATAI_9_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4652) );
  INV_X1 U5156 ( .A(n4652), .ZN(U3343) );
  AOI22_X1 U5157 ( .A1(STATE_REG_SCAN_IN), .A2(n4654), .B1(n4653), .B2(U3149), 
        .ZN(U3344) );
  AOI22_X1 U5158 ( .A1(STATE_REG_SCAN_IN), .A2(n2103), .B1(n2102), .B2(U3149), 
        .ZN(U3352) );
  INV_X1 U5159 ( .A(n4655), .ZN(n4658) );
  INV_X1 U5160 ( .A(n4656), .ZN(n4657) );
  AOI211_X1 U5161 ( .C1(n4675), .C2(n4659), .A(n4658), .B(n4657), .ZN(n4706)
         );
  INV_X1 U5162 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4660) );
  AOI22_X1 U5163 ( .A1(n4705), .A2(n4706), .B1(n4660), .B2(n4703), .ZN(U3467)
         );
  NOR2_X1 U5164 ( .A1(n4661), .A2(n4699), .ZN(n4663) );
  AOI211_X1 U5165 ( .C1(n2707), .C2(n4664), .A(n4663), .B(n4662), .ZN(n4707)
         );
  INV_X1 U5166 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4665) );
  AOI22_X1 U5167 ( .A1(n4705), .A2(n4707), .B1(n4665), .B2(n4703), .ZN(U3469)
         );
  OAI22_X1 U5168 ( .A1(n4667), .A2(n4699), .B1(n4698), .B2(n4666), .ZN(n4668)
         );
  NOR2_X1 U5169 ( .A1(n4669), .A2(n4668), .ZN(n4709) );
  INV_X1 U5170 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4670) );
  AOI22_X1 U5171 ( .A1(n4705), .A2(n4709), .B1(n4670), .B2(n4703), .ZN(U3473)
         );
  INV_X1 U5172 ( .A(n4671), .ZN(n4676) );
  INV_X1 U5173 ( .A(n4672), .ZN(n4674) );
  AOI211_X1 U5174 ( .C1(n4676), .C2(n4675), .A(n4674), .B(n4673), .ZN(n4710)
         );
  AOI22_X1 U5175 ( .A1(n4705), .A2(n4710), .B1(n4677), .B2(n4703), .ZN(U3475)
         );
  NOR2_X1 U5176 ( .A1(n4679), .A2(n4678), .ZN(n4682) );
  INV_X1 U5177 ( .A(n4680), .ZN(n4681) );
  AOI211_X1 U5178 ( .C1(n2707), .C2(n4683), .A(n4682), .B(n4681), .ZN(n4711)
         );
  INV_X1 U5179 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4684) );
  AOI22_X1 U5180 ( .A1(n4705), .A2(n4711), .B1(n4684), .B2(n4703), .ZN(U3477)
         );
  NAND3_X1 U5181 ( .A1(n4686), .A2(n4685), .A3(n4694), .ZN(n4687) );
  AND3_X1 U5182 ( .A1(n4689), .A2(n4688), .A3(n4687), .ZN(n4712) );
  INV_X1 U5183 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4690) );
  AOI22_X1 U5184 ( .A1(n4705), .A2(n4712), .B1(n4690), .B2(n4703), .ZN(U3481)
         );
  OAI21_X1 U5185 ( .B1(n4698), .B2(n4692), .A(n4691), .ZN(n4693) );
  AOI21_X1 U5186 ( .B1(n4695), .B2(n4694), .A(n4693), .ZN(n4713) );
  INV_X1 U5187 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4696) );
  AOI22_X1 U5188 ( .A1(n4705), .A2(n4713), .B1(n4696), .B2(n4703), .ZN(U3485)
         );
  OAI22_X1 U5189 ( .A1(n4700), .A2(n4699), .B1(n4698), .B2(n4697), .ZN(n4701)
         );
  NOR2_X1 U5190 ( .A1(n4702), .A2(n4701), .ZN(n4715) );
  INV_X1 U5191 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4704) );
  AOI22_X1 U5192 ( .A1(n4705), .A2(n4715), .B1(n4704), .B2(n4703), .ZN(U3489)
         );
  AOI22_X1 U5193 ( .A1(n4716), .A2(n4706), .B1(n2736), .B2(n4714), .ZN(U3518)
         );
  AOI22_X1 U5194 ( .A1(n4716), .A2(n4707), .B1(n2845), .B2(n4714), .ZN(U3519)
         );
  INV_X1 U5195 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4708) );
  AOI22_X1 U5196 ( .A1(n4716), .A2(n4709), .B1(n4708), .B2(n4714), .ZN(U3521)
         );
  AOI22_X1 U5197 ( .A1(n4716), .A2(n4710), .B1(n2363), .B2(n4714), .ZN(U3522)
         );
  AOI22_X1 U5198 ( .A1(n4716), .A2(n4711), .B1(n2371), .B2(n4714), .ZN(U3523)
         );
  AOI22_X1 U5199 ( .A1(n4716), .A2(n4712), .B1(n4070), .B2(n4714), .ZN(U3525)
         );
  AOI22_X1 U5200 ( .A1(n4716), .A2(n4713), .B1(n2406), .B2(n4714), .ZN(U3527)
         );
  AOI22_X1 U5201 ( .A1(n4716), .A2(n4715), .B1(n2443), .B2(n4714), .ZN(U3529)
         );
  NOR2_X2 U2337 ( .A1(n3094), .A2(n2936), .ZN(n3188) );
endmodule

