

module b14_C_AntiSAT_k_128_5 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669;

  INV_X1 U2293 ( .A(n3193), .ZN(n3195) );
  XNOR2_X1 U2294 ( .A(n2337), .B(IR_REG_1__SCAN_IN), .ZN(n4277) );
  INV_X1 U2295 ( .A(n2661), .ZN(n2051) );
  AND2_X1 U2296 ( .A1(n2788), .A2(n2978), .ZN(n2734) );
  NAND2_X1 U2297 ( .A1(n2096), .A2(n3652), .ZN(n3308) );
  AND2_X1 U2298 ( .A1(n3622), .A2(n3619), .ZN(n3603) );
  INV_X1 U2299 ( .A(n2734), .ZN(n2746) );
  NAND4_X1 U2300 ( .A1(n2370), .A2(n2369), .A3(n2368), .A4(n2367), .ZN(n3050)
         );
  INV_X1 U2301 ( .A(n3418), .ZN(n2973) );
  NAND2_X1 U2302 ( .A1(n3193), .A2(n3140), .ZN(n3206) );
  NAND2_X2 U2303 ( .A1(n3359), .A2(n3669), .ZN(n3958) );
  NOR2_X1 U2304 ( .A1(n2332), .A2(n2331), .ZN(n2366) );
  CLKBUF_X3 U2305 ( .A(n2366), .Z(n2668) );
  OAI21_X1 U2306 ( .B1(n3044), .B2(n2061), .A(n2101), .ZN(n3111) );
  INV_X1 U2307 ( .A(n2052), .ZN(n2054) );
  INV_X2 U2308 ( .A(n2383), .ZN(n2052) );
  NOR2_X1 U2309 ( .A1(n4370), .A2(n2214), .ZN(n2213) );
  INV_X1 U2310 ( .A(n2193), .ZN(n4370) );
  OR2_X1 U2311 ( .A1(n4371), .A2(n4372), .ZN(n2193) );
  NAND2_X1 U2312 ( .A1(n2118), .A2(n2119), .ZN(n3825) );
  NAND2_X1 U2313 ( .A1(n3857), .A2(n2076), .ZN(n2118) );
  OAI21_X1 U2314 ( .B1(n3877), .B2(n3347), .A(n3346), .ZN(n3857) );
  NAND2_X1 U2315 ( .A1(n4356), .A2(n4058), .ZN(n4355) );
  XNOR2_X1 U2316 ( .A(n3770), .B(n2572), .ZN(n4356) );
  NAND2_X1 U2317 ( .A1(n4077), .A2(n3544), .ZN(n4062) );
  NOR2_X1 U2318 ( .A1(n4343), .A2(n2091), .ZN(n3770) );
  AOI21_X1 U2319 ( .B1(n4034), .B2(n3334), .A(n3333), .ZN(n4017) );
  AOI21_X1 U2320 ( .B1(n3786), .B2(REG1_REG_13__SCAN_IN), .A(n4314), .ZN(n3787) );
  AOI21_X1 U2321 ( .B1(n4075), .B2(n3332), .A(n2081), .ZN(n4052) );
  NAND2_X1 U2322 ( .A1(n2075), .A2(n2120), .ZN(n2119) );
  NAND2_X1 U2323 ( .A1(n3350), .A2(n2121), .ZN(n2120) );
  AOI21_X1 U2324 ( .B1(n3783), .B2(REG1_REG_11__SCAN_IN), .A(n4295), .ZN(n3784) );
  AOI21_X1 U2325 ( .B1(n2145), .B2(n2150), .A(n2144), .ZN(n2143) );
  OAI21_X1 U2326 ( .B1(n3113), .B2(n3112), .A(n3640), .ZN(n3127) );
  XNOR2_X1 U2327 ( .A(n2895), .B(n2908), .ZN(n2905) );
  AND2_X1 U2328 ( .A1(n2247), .A2(n3000), .ZN(n2246) );
  OAI22_X1 U2329 ( .A1(n3111), .A2(n2105), .B1(n2103), .B2(n3110), .ZN(n3136)
         );
  NOR2_X2 U2330 ( .A1(n2791), .A2(n4392), .ZN(n2792) );
  NOR2_X2 U2332 ( .A1(n2845), .A2(n2844), .ZN(n4351) );
  OR2_X2 U2333 ( .A1(n2745), .A2(n4443), .ZN(n2748) );
  NAND2_X2 U2334 ( .A1(n2348), .A2(n2978), .ZN(n2745) );
  INV_X1 U2335 ( .A(n3070), .ZN(n3712) );
  INV_X1 U2336 ( .A(n3115), .ZN(n3711) );
  OR2_X1 U2337 ( .A1(n2856), .A2(n2855), .ZN(n2189) );
  NAND2_X1 U2338 ( .A1(n2430), .A2(n2273), .ZN(n3708) );
  AND4_X1 U2339 ( .A1(n2396), .A2(n2395), .A3(n2394), .A4(n2393), .ZN(n3115)
         );
  AND4_X1 U2340 ( .A1(n2387), .A2(n2386), .A3(n2385), .A4(n2384), .ZN(n3070)
         );
  AND2_X1 U2341 ( .A1(n2426), .A2(n2425), .ZN(n2430) );
  NAND2_X1 U2342 ( .A1(n2185), .A2(n2851), .ZN(n2852) );
  INV_X2 U2343 ( .A(n2052), .ZN(n2053) );
  INV_X1 U2344 ( .A(n2052), .ZN(n2056) );
  INV_X1 U2345 ( .A(n2052), .ZN(n2055) );
  AND3_X1 U2346 ( .A1(n2074), .A2(n2266), .A3(n2267), .ZN(n2179) );
  AND2_X1 U2347 ( .A1(n2270), .A2(n2288), .ZN(n2269) );
  AND2_X1 U2348 ( .A1(n2286), .A2(n2287), .ZN(n2270) );
  AND2_X1 U2349 ( .A1(n2272), .A2(n2281), .ZN(n2251) );
  AND3_X1 U2350 ( .A1(n4502), .A2(n2557), .A3(n2568), .ZN(n2282) );
  AND2_X1 U2351 ( .A1(n2284), .A2(n2283), .ZN(n2266) );
  AND2_X1 U2352 ( .A1(n2285), .A2(n2268), .ZN(n2267) );
  INV_X1 U2353 ( .A(IR_REG_16__SCAN_IN), .ZN(n4502) );
  INV_X1 U2354 ( .A(IR_REG_22__SCAN_IN), .ZN(n2285) );
  NOR2_X1 U2355 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2319)
         );
  NOR2_X1 U2356 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2284)
         );
  INV_X1 U2357 ( .A(IR_REG_18__SCAN_IN), .ZN(n2283) );
  NOR2_X1 U2358 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2099)
         );
  NOR2_X1 U2359 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2098)
         );
  NOR2_X1 U2360 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2097)
         );
  NOR2_X1 U2361 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2100)
         );
  INV_X1 U2362 ( .A(IR_REG_23__SCAN_IN), .ZN(n2772) );
  NAND2_X1 U2363 ( .A1(n3264), .A2(n3649), .ZN(n2096) );
  AND2_X1 U2364 ( .A1(n2332), .A2(n2331), .ZN(n2383) );
  XNOR2_X2 U2365 ( .A(n2095), .B(n2289), .ZN(n2332) );
  INV_X1 U2366 ( .A(IR_REG_21__SCAN_IN), .ZN(n2268) );
  NAND2_X1 U2367 ( .A1(n2861), .A2(n2860), .ZN(n2863) );
  NAND2_X1 U2368 ( .A1(n2279), .A2(n2066), .ZN(n2155) );
  AND2_X1 U2369 ( .A1(n3451), .A2(n2239), .ZN(n2238) );
  OR2_X1 U2370 ( .A1(n2579), .A2(n2240), .ZN(n2239) );
  INV_X1 U2371 ( .A(n3515), .ZN(n2240) );
  AND2_X1 U2372 ( .A1(n3822), .A2(n3351), .ZN(n3809) );
  AOI21_X1 U2373 ( .B1(n2115), .B2(n2113), .A(n2057), .ZN(n2111) );
  INV_X1 U2374 ( .A(n2102), .ZN(n2101) );
  OAI21_X1 U2375 ( .B1(n2061), .B2(n3043), .A(n3045), .ZN(n2102) );
  NOR2_X1 U2376 ( .A1(n3986), .A2(n3339), .ZN(n3950) );
  INV_X1 U2377 ( .A(IR_REG_17__SCAN_IN), .ZN(n2178) );
  NAND2_X1 U2378 ( .A1(n2249), .A2(n2248), .ZN(n2247) );
  INV_X1 U2379 ( .A(n2957), .ZN(n2248) );
  INV_X1 U2380 ( .A(n2956), .ZN(n2249) );
  AND2_X1 U2381 ( .A1(n2331), .A2(REG0_REG_1__SCAN_IN), .ZN(n2094) );
  OR2_X1 U2382 ( .A1(n2948), .A2(n2407), .ZN(n2279) );
  NOR2_X1 U2383 ( .A1(n2994), .A2(n2157), .ZN(n2156) );
  INV_X1 U2384 ( .A(n2381), .ZN(n2157) );
  OR2_X1 U2385 ( .A1(n2724), .A2(n2709), .ZN(n3507) );
  AND2_X1 U2386 ( .A1(n2332), .A2(n2294), .ZN(n2682) );
  NAND2_X1 U2388 ( .A1(n2756), .A2(n2311), .ZN(n2348) );
  OAI21_X1 U2389 ( .B1(n3747), .B2(n2862), .A(n2864), .ZN(n2865) );
  XNOR2_X1 U2390 ( .A(n2852), .B(n2184), .ZN(n2853) );
  INV_X1 U2391 ( .A(n4274), .ZN(n2184) );
  OR2_X1 U2392 ( .A1(n4383), .A2(n3686), .ZN(n4059) );
  INV_X1 U2393 ( .A(IR_REG_3__SCAN_IN), .ZN(n2371) );
  OR2_X1 U2394 ( .A1(n3808), .A2(n4373), .ZN(n2208) );
  INV_X1 U2395 ( .A(n2690), .ZN(n2166) );
  INV_X1 U2396 ( .A(n2169), .ZN(n2167) );
  INV_X1 U2397 ( .A(n2089), .ZN(n2164) );
  INV_X1 U2398 ( .A(n2676), .ZN(n2168) );
  INV_X1 U2399 ( .A(n2748), .ZN(n2737) );
  NAND2_X1 U2400 ( .A1(n2148), .A2(n3381), .ZN(n2580) );
  OR2_X1 U2401 ( .A1(n3380), .A2(n3382), .ZN(n2148) );
  INV_X1 U2402 ( .A(IR_REG_28__SCAN_IN), .ZN(n2325) );
  OR2_X1 U2403 ( .A1(n2801), .A2(n2322), .ZN(n2324) );
  INV_X1 U2404 ( .A(IR_REG_27__SCAN_IN), .ZN(n2322) );
  OR2_X1 U2405 ( .A1(n2790), .A2(n4269), .ZN(n2788) );
  AND2_X1 U2406 ( .A1(n2695), .A2(REG3_REG_25__SCAN_IN), .ZN(n2708) );
  NOR2_X1 U2407 ( .A1(n2680), .A2(n3471), .ZN(n2695) );
  AOI21_X1 U2408 ( .B1(REG1_REG_9__SCAN_IN), .B2(n3778), .A(n3777), .ZN(n3780)
         );
  INV_X1 U2409 ( .A(n3826), .ZN(n2125) );
  OR2_X1 U2410 ( .A1(n3215), .A2(n3221), .ZN(n3216) );
  NAND2_X1 U2411 ( .A1(n3626), .A2(n3623), .ZN(n2106) );
  INV_X1 U2412 ( .A(n4384), .ZN(n2974) );
  AND2_X1 U2413 ( .A1(n3335), .A2(n4007), .ZN(n2175) );
  OR2_X1 U2414 ( .A1(n4054), .A2(n4055), .ZN(n4042) );
  AND2_X1 U2415 ( .A1(n2183), .A2(n3309), .ZN(n2182) );
  AND2_X1 U2416 ( .A1(n3277), .A2(n3266), .ZN(n2183) );
  INV_X1 U2417 ( .A(IR_REG_24__SCAN_IN), .ZN(n2309) );
  AND2_X1 U2418 ( .A1(n2266), .A2(n2267), .ZN(n2265) );
  AND2_X1 U2419 ( .A1(n2251), .A2(n2282), .ZN(n2139) );
  INV_X1 U2420 ( .A(n2253), .ZN(n2252) );
  NOR2_X1 U2421 ( .A1(n3489), .A2(n2170), .ZN(n2169) );
  INV_X1 U2422 ( .A(n3424), .ZN(n2170) );
  AND2_X1 U2423 ( .A1(n2771), .A2(n3037), .ZN(n2782) );
  NAND2_X1 U2424 ( .A1(n2262), .A2(n2261), .ZN(n2257) );
  INV_X1 U2425 ( .A(n3230), .ZN(n2261) );
  INV_X1 U2426 ( .A(n3229), .ZN(n2262) );
  INV_X1 U2427 ( .A(n3256), .ZN(n2259) );
  AND2_X1 U2428 ( .A1(n2492), .A2(n2264), .ZN(n2263) );
  NAND2_X1 U2429 ( .A1(n3229), .A2(n3230), .ZN(n2264) );
  OR2_X1 U2430 ( .A1(n2508), .A2(n2507), .ZN(n2523) );
  AND2_X1 U2431 ( .A1(n2146), .A2(n2235), .ZN(n2145) );
  AOI21_X1 U2432 ( .B1(n2238), .B2(n2241), .A(n2236), .ZN(n2235) );
  NAND2_X1 U2433 ( .A1(n2149), .A2(n2147), .ZN(n2146) );
  INV_X1 U2434 ( .A(n2581), .ZN(n2236) );
  NAND2_X1 U2435 ( .A1(n3382), .A2(n3381), .ZN(n2151) );
  NAND2_X1 U2436 ( .A1(n3439), .A2(n3437), .ZN(n2707) );
  AND4_X1 U2437 ( .A1(n2567), .A2(n2566), .A3(n2565), .A4(n2564), .ZN(n3517)
         );
  OR2_X1 U2438 ( .A1(n3739), .A2(n2834), .ZN(n2836) );
  NAND2_X1 U2439 ( .A1(n2849), .A2(REG2_REG_3__SCAN_IN), .ZN(n2185) );
  NAND2_X1 U2440 ( .A1(n2897), .A2(n2896), .ZN(n2202) );
  NAND2_X1 U2441 ( .A1(n3760), .A2(n2079), .ZN(n3762) );
  OR2_X1 U2442 ( .A1(n4326), .A2(n2228), .ZN(n2226) );
  OR2_X1 U2443 ( .A1(n4340), .A2(n4327), .ZN(n2228) );
  OR2_X1 U2444 ( .A1(n2060), .A2(n4340), .ZN(n2227) );
  OR2_X1 U2445 ( .A1(n4326), .A2(n4327), .ZN(n2229) );
  AND2_X1 U2446 ( .A1(n2744), .A2(n2743), .ZN(n3822) );
  OR2_X1 U2447 ( .A1(n2738), .A2(n2793), .ZN(n2794) );
  AND2_X1 U2448 ( .A1(n2125), .A2(n3823), .ZN(n2124) );
  NOR2_X1 U2449 ( .A1(n3823), .A2(n2125), .ZN(n2123) );
  NOR2_X1 U2450 ( .A1(n3827), .A2(n3828), .ZN(n4130) );
  AOI21_X1 U2451 ( .B1(n2136), .B2(n2134), .A(n2083), .ZN(n2133) );
  INV_X1 U2452 ( .A(n2136), .ZN(n2135) );
  INV_X1 U2453 ( .A(n3341), .ZN(n2134) );
  INV_X1 U2454 ( .A(n3700), .ZN(n3924) );
  OR2_X1 U2455 ( .A1(n3337), .A2(n3338), .ZN(n2113) );
  INV_X1 U2456 ( .A(n3942), .ZN(n3975) );
  AND4_X1 U2457 ( .A1(n2634), .A2(n2633), .A3(n2632), .A4(n2631), .ZN(n3999)
         );
  AOI21_X1 U2458 ( .B1(n2130), .B2(n2128), .A(n2070), .ZN(n2127) );
  INV_X1 U2459 ( .A(n2130), .ZN(n2129) );
  NAND2_X1 U2460 ( .A1(n3175), .A2(n3633), .ZN(n3176) );
  NAND2_X1 U2461 ( .A1(n3732), .A2(n2972), .ZN(n4388) );
  OR2_X1 U2462 ( .A1(n3850), .A2(n3351), .ZN(n3827) );
  AND2_X1 U2463 ( .A1(n3949), .A2(n2059), .ZN(n3868) );
  NAND2_X1 U2464 ( .A1(n3949), .A2(n2058), .ZN(n3890) );
  AND2_X1 U2465 ( .A1(n3950), .A2(n3491), .ZN(n3949) );
  INV_X1 U2466 ( .A(n3411), .ZN(n4007) );
  NAND2_X1 U2467 ( .A1(n4043), .A2(n2175), .ZN(n4006) );
  NOR2_X1 U2468 ( .A1(n4042), .A2(n3462), .ZN(n4043) );
  NOR2_X1 U2469 ( .A1(n4111), .A2(n3331), .ZN(n4085) );
  AND2_X1 U2470 ( .A1(n2330), .A2(n3686), .ZN(n4443) );
  AND3_X1 U2471 ( .A1(n3031), .A2(n3030), .A3(n3029), .ZN(n3038) );
  OR2_X1 U2472 ( .A1(n2300), .A2(n2820), .ZN(n2801) );
  INV_X1 U2473 ( .A(n2319), .ZN(n2197) );
  INV_X1 U2474 ( .A(n2250), .ZN(n2244) );
  NAND2_X1 U2475 ( .A1(n2959), .A2(n2247), .ZN(n2245) );
  NAND2_X1 U2476 ( .A1(n2682), .A2(REG1_REG_2__SCAN_IN), .ZN(n2296) );
  AOI21_X1 U2477 ( .B1(n2246), .B2(n2250), .A(n2078), .ZN(n2242) );
  AOI21_X1 U2478 ( .B1(n2382), .B2(n2063), .A(n2153), .ZN(n2243) );
  OAI21_X1 U2479 ( .B1(n2433), .B2(n2339), .A(n2338), .ZN(n3418) );
  AND4_X2 U2480 ( .A1(n2335), .A2(n2336), .A3(n2334), .A4(n2333), .ZN(n2340)
         );
  NAND2_X1 U2481 ( .A1(n2332), .A2(n2094), .ZN(n2335) );
  NAND2_X1 U2482 ( .A1(n2707), .A2(n3438), .ZN(n2162) );
  OAI21_X1 U2483 ( .B1(n3507), .B2(n2714), .A(n2713), .ZN(n3887) );
  OR2_X1 U2484 ( .A1(n3533), .A2(n2365), .ZN(n2370) );
  NOR2_X1 U2485 ( .A1(n2905), .A2(n2441), .ZN(n2904) );
  XNOR2_X1 U2486 ( .A(n3762), .B(n4416), .ZN(n4292) );
  NAND2_X1 U2487 ( .A1(n4292), .A2(REG2_REG_10__SCAN_IN), .ZN(n4291) );
  OR2_X1 U2488 ( .A1(n3808), .A2(n2212), .ZN(n2210) );
  INV_X1 U2489 ( .A(n3804), .ZN(n2212) );
  OR2_X1 U2490 ( .A1(n3808), .A2(n2221), .ZN(n2211) );
  NAND2_X1 U2491 ( .A1(n2213), .A2(n2208), .ZN(n2206) );
  NAND2_X1 U2492 ( .A1(n3804), .A2(n2222), .ZN(n2214) );
  AND2_X1 U2493 ( .A1(n4396), .A2(n3063), .ZN(n4005) );
  OR2_X1 U2494 ( .A1(n3024), .A2(n3022), .ZN(n4115) );
  XNOR2_X1 U2495 ( .A(n2389), .B(IR_REG_4__SCAN_IN), .ZN(n4274) );
  NOR2_X1 U2496 ( .A1(n2560), .A2(n3515), .ZN(n2241) );
  INV_X1 U2497 ( .A(IR_REG_13__SCAN_IN), .ZN(n2281) );
  AND3_X1 U2498 ( .A1(n2226), .A2(n2227), .A3(n2092), .ZN(n3790) );
  INV_X1 U2499 ( .A(n3348), .ZN(n2121) );
  AOI21_X1 U2500 ( .B1(n3938), .B2(n3341), .A(n2084), .ZN(n2136) );
  AOI21_X1 U2501 ( .B1(n3599), .B2(n3285), .A(n2068), .ZN(n2130) );
  INV_X1 U2502 ( .A(n3285), .ZN(n2128) );
  NOR2_X1 U2503 ( .A1(n4268), .A2(n3579), .ZN(n2984) );
  INV_X1 U2504 ( .A(n2984), .ZN(n2978) );
  AND2_X1 U2505 ( .A1(n2433), .A2(DATAI_28_), .ZN(n3351) );
  NOR2_X1 U2506 ( .A1(n3908), .A2(n3363), .ZN(n2181) );
  NAND2_X1 U2507 ( .A1(n3711), .A2(n3108), .ZN(n2104) );
  NOR2_X1 U2508 ( .A1(n2465), .A2(IR_REG_9__SCAN_IN), .ZN(n2501) );
  INV_X1 U2509 ( .A(IR_REG_6__SCAN_IN), .ZN(n2431) );
  AND2_X1 U2510 ( .A1(n2433), .A2(DATAI_27_), .ZN(n3613) );
  AOI21_X1 U2511 ( .B1(n3096), .B2(n3095), .A(n2161), .ZN(n2158) );
  INV_X1 U2512 ( .A(n3169), .ZN(n2161) );
  XNOR2_X1 U2513 ( .A(n2377), .B(n2746), .ZN(n2378) );
  NAND2_X1 U2514 ( .A1(n2376), .A2(n2375), .ZN(n2377) );
  NOR2_X1 U2515 ( .A1(n3505), .A2(n2231), .ZN(n2230) );
  INV_X1 U2516 ( .A(n3438), .ZN(n2231) );
  INV_X1 U2517 ( .A(n2246), .ZN(n2154) );
  AND2_X1 U2518 ( .A1(n2956), .A2(n2957), .ZN(n2250) );
  INV_X1 U2519 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2438) );
  AOI21_X1 U2520 ( .B1(n2975), .B2(n2051), .A(n2352), .ZN(n2354) );
  NOR2_X1 U2521 ( .A1(n2562), .A2(n2561), .ZN(n2582) );
  OAI21_X1 U2522 ( .B1(n3430), .B2(n2069), .A(n2165), .ZN(n2693) );
  AOI21_X1 U2523 ( .B1(n2676), .B2(n2167), .A(n2166), .ZN(n2165) );
  OR2_X1 U2524 ( .A1(n2347), .A2(n2748), .ZN(n2351) );
  AND2_X1 U2525 ( .A1(n2626), .A2(n3405), .ZN(n2627) );
  NAND2_X1 U2526 ( .A1(n2163), .A2(n2089), .ZN(n2171) );
  XNOR2_X1 U2527 ( .A(n2329), .B(n2746), .ZN(n2360) );
  OAI22_X1 U2528 ( .A1(n3006), .A2(n2661), .B1(n3042), .B2(n2745), .ZN(n2329)
         );
  INV_X1 U2529 ( .A(n3459), .ZN(n2144) );
  NAND2_X1 U2530 ( .A1(n2598), .A2(REG3_REG_18__SCAN_IN), .ZN(n2609) );
  INV_X1 U2531 ( .A(n3708), .ZN(n3129) );
  INV_X1 U2532 ( .A(n2782), .ZN(n2800) );
  INV_X1 U2533 ( .A(n2580), .ZN(n2237) );
  INV_X1 U2534 ( .A(n4084), .ZN(n3354) );
  NAND2_X1 U2535 ( .A1(n2324), .A2(n2323), .ZN(n2172) );
  OR3_X1 U2536 ( .A1(n2661), .A2(n2811), .A3(n2788), .ZN(n2799) );
  XNOR2_X1 U2537 ( .A(n2863), .B(n4274), .ZN(n3747) );
  NAND2_X1 U2538 ( .A1(n2189), .A2(n2188), .ZN(n2187) );
  NAND2_X1 U2539 ( .A1(n4273), .A2(REG2_REG_5__SCAN_IN), .ZN(n2188) );
  AOI21_X1 U2540 ( .B1(n2913), .B2(REG2_REG_6__SCAN_IN), .A(n2186), .ZN(n2880)
         );
  AND2_X1 U2541 ( .A1(n2187), .A2(n4272), .ZN(n2186) );
  XNOR2_X1 U2542 ( .A(n3780), .B(n4416), .ZN(n4286) );
  NOR2_X1 U2543 ( .A1(n4286), .A2(n4287), .ZN(n4285) );
  INV_X1 U2544 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3324) );
  NAND2_X1 U2545 ( .A1(n4355), .A2(n3771), .ZN(n3772) );
  AOI22_X1 U2546 ( .A1(n2217), .A2(n4363), .B1(n3800), .B2(n2090), .ZN(n2216)
         );
  INV_X1 U2547 ( .A(n3595), .ZN(n3828) );
  AND2_X1 U2548 ( .A1(n2794), .A2(n2739), .ZN(n3833) );
  INV_X1 U2549 ( .A(n3491), .ZN(n3951) );
  AND4_X1 U2550 ( .A1(n2672), .A2(n2671), .A3(n2670), .A4(n2669), .ZN(n3945)
         );
  NOR2_X1 U2551 ( .A1(n2640), .A2(n3432), .ZN(n2655) );
  NAND2_X1 U2552 ( .A1(n2138), .A2(n2137), .ZN(n3937) );
  AOI21_X1 U2553 ( .B1(n2111), .B2(n2112), .A(n2082), .ZN(n2109) );
  INV_X1 U2554 ( .A(n2113), .ZN(n2112) );
  OR2_X1 U2555 ( .A1(n2609), .A2(n3409), .ZN(n2629) );
  NAND2_X1 U2556 ( .A1(n4038), .A2(n3335), .ZN(n3336) );
  NAND2_X1 U2557 ( .A1(n4051), .A2(n2077), .ZN(n4034) );
  AND4_X1 U2558 ( .A1(n2587), .A2(n2586), .A3(n2585), .A4(n2584), .ZN(n4061)
         );
  NAND2_X1 U2559 ( .A1(n4052), .A2(n4066), .ZN(n4051) );
  NAND2_X1 U2560 ( .A1(n3330), .A2(n2107), .ZN(n4075) );
  NAND2_X1 U2561 ( .A1(n4083), .A2(n3385), .ZN(n2107) );
  AND4_X1 U2562 ( .A1(n2556), .A2(n2555), .A3(n2554), .A4(n2553), .ZN(n3452)
         );
  NAND2_X1 U2563 ( .A1(n3263), .A2(n3277), .ZN(n3285) );
  NAND2_X1 U2564 ( .A1(n2132), .A2(n2131), .ZN(n3286) );
  AND4_X1 U2565 ( .A1(n2528), .A2(n2527), .A3(n2526), .A4(n2525), .ZN(n3384)
         );
  AND2_X1 U2566 ( .A1(n3305), .A2(n3307), .ZN(n3599) );
  AND4_X1 U2567 ( .A1(n2514), .A2(n2513), .A3(n2512), .A4(n2511), .ZN(n4105)
         );
  INV_X1 U2568 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2475) );
  NOR2_X1 U2569 ( .A1(n2476), .A2(n2475), .ZN(n2493) );
  INV_X1 U2570 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2891) );
  INV_X1 U2571 ( .A(n3190), .ZN(n3183) );
  AND4_X1 U2572 ( .A1(n2445), .A2(n2444), .A3(n2443), .A4(n2442), .ZN(n3182)
         );
  NAND2_X1 U2573 ( .A1(n3128), .A2(n3628), .ZN(n3155) );
  NOR2_X1 U2574 ( .A1(n2411), .A2(n2410), .ZN(n2423) );
  NAND2_X1 U2575 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2411) );
  INV_X1 U2576 ( .A(n4388), .ZN(n4101) );
  OR2_X1 U2577 ( .A1(n3085), .A2(n3064), .ZN(n3073) );
  NAND2_X1 U2578 ( .A1(n3049), .A2(n3622), .ZN(n3068) );
  INV_X1 U2579 ( .A(n4071), .ZN(n4104) );
  NAND2_X1 U2580 ( .A1(n2093), .A2(n3604), .ZN(n3047) );
  NAND2_X1 U2581 ( .A1(n2976), .A2(n3602), .ZN(n3008) );
  AND2_X1 U2582 ( .A1(n4264), .A2(n2972), .ZN(n4071) );
  INV_X1 U2583 ( .A(n4065), .ZN(n4386) );
  INV_X1 U2584 ( .A(n4059), .ZN(n4135) );
  INV_X1 U2585 ( .A(n3903), .ZN(n3908) );
  NAND2_X1 U2586 ( .A1(n3949), .A2(n2181), .ZN(n3910) );
  NAND2_X1 U2587 ( .A1(n3949), .A2(n3928), .ZN(n3930) );
  NAND2_X1 U2588 ( .A1(n4043), .A2(n2088), .ZN(n3986) );
  NAND2_X1 U2589 ( .A1(n3224), .A2(n2080), .ZN(n4111) );
  NAND2_X1 U2590 ( .A1(n3224), .A2(n2182), .ZN(n4110) );
  NAND2_X1 U2591 ( .A1(n3224), .A2(n2183), .ZN(n3313) );
  NOR2_X1 U2592 ( .A1(n3193), .A2(n3218), .ZN(n3224) );
  AND2_X1 U2593 ( .A1(n3224), .A2(n3266), .ZN(n3278) );
  INV_X1 U2594 ( .A(n3181), .ZN(n3187) );
  OR2_X1 U2595 ( .A1(n3159), .A2(n3187), .ZN(n3193) );
  NAND2_X1 U2596 ( .A1(n4109), .A2(n4427), .ZN(n4453) );
  INV_X1 U2597 ( .A(n3134), .ZN(n3118) );
  AND2_X1 U2598 ( .A1(n3119), .A2(n3118), .ZN(n3161) );
  NOR2_X1 U2599 ( .A1(n3073), .A2(n3108), .ZN(n3119) );
  NOR2_X1 U2600 ( .A1(n3033), .A2(n3034), .ZN(n3087) );
  NAND2_X1 U2601 ( .A1(n2290), .A2(IR_REG_31__SCAN_IN), .ZN(n2292) );
  XNOR2_X1 U2602 ( .A(n2803), .B(IR_REG_28__SCAN_IN), .ZN(n3732) );
  NAND2_X1 U2603 ( .A1(n2179), .A2(n2177), .ZN(n2176) );
  NOR2_X1 U2604 ( .A1(n2180), .A2(IR_REG_17__SCAN_IN), .ZN(n2177) );
  INV_X1 U2605 ( .A(n2270), .ZN(n2180) );
  XNOR2_X1 U2606 ( .A(n2310), .B(n2309), .ZN(n2769) );
  NAND2_X1 U2607 ( .A1(n2308), .A2(IR_REG_31__SCAN_IN), .ZN(n2310) );
  XNOR2_X1 U2608 ( .A(n2327), .B(n2285), .ZN(n2790) );
  XNOR2_X1 U2609 ( .A(n2318), .B(n2317), .ZN(n3686) );
  INV_X1 U2610 ( .A(IR_REG_20__SCAN_IN), .ZN(n2317) );
  NAND2_X1 U2611 ( .A1(n2606), .A2(IR_REG_31__SCAN_IN), .ZN(n2328) );
  NAND2_X1 U2612 ( .A1(n2590), .A2(n2283), .ZN(n2606) );
  INV_X1 U2613 ( .A(IR_REG_15__SCAN_IN), .ZN(n2568) );
  AND3_X1 U2614 ( .A1(n2252), .A2(n2321), .A3(n2272), .ZN(n2529) );
  AND2_X1 U2615 ( .A1(n2515), .A2(n2505), .ZN(n3783) );
  NOR2_X1 U2616 ( .A1(n2397), .A2(IR_REG_5__SCAN_IN), .ZN(n2432) );
  INV_X1 U2617 ( .A(n3138), .ZN(n3160) );
  INV_X1 U2618 ( .A(n3613), .ZN(n3851) );
  NAND2_X1 U2619 ( .A1(n2234), .A2(n3504), .ZN(n3374) );
  AND2_X1 U2620 ( .A1(n2738), .A2(n2725), .ZN(n3852) );
  INV_X1 U2621 ( .A(n3080), .ZN(n3086) );
  INV_X1 U2622 ( .A(n2777), .ZN(n2778) );
  NAND2_X1 U2623 ( .A1(n2234), .A2(n2232), .ZN(n2777) );
  NOR2_X1 U2624 ( .A1(n3373), .A2(n2233), .ZN(n2232) );
  NAND2_X1 U2625 ( .A1(n3476), .A2(n3479), .ZN(n3430) );
  AND2_X1 U2626 ( .A1(n2782), .A2(n2774), .ZN(n3428) );
  INV_X1 U2627 ( .A(n2257), .ZN(n2254) );
  INV_X1 U2628 ( .A(n4055), .ZN(n4060) );
  INV_X1 U2629 ( .A(n3106), .ZN(n3108) );
  OR2_X1 U2630 ( .A1(n3380), .A2(n2150), .ZN(n2142) );
  NAND2_X1 U2631 ( .A1(n2433), .A2(DATAI_24_), .ZN(n3903) );
  INV_X1 U2632 ( .A(n3064), .ZN(n3055) );
  OR2_X1 U2633 ( .A1(n3094), .A2(n3096), .ZN(n2160) );
  INV_X1 U2634 ( .A(DATAI_0_), .ZN(n2173) );
  NAND2_X1 U2635 ( .A1(n2804), .A2(n3732), .ZN(n3518) );
  INV_X1 U2636 ( .A(n2256), .ZN(n2255) );
  NAND2_X1 U2637 ( .A1(n2263), .A2(n2259), .ZN(n2258) );
  OAI21_X1 U2638 ( .B1(n3256), .B2(n2257), .A(n3255), .ZN(n2256) );
  NAND2_X1 U2639 ( .A1(n2433), .A2(DATAI_22_), .ZN(n3491) );
  NAND2_X1 U2640 ( .A1(n2171), .A2(n3424), .ZN(n3488) );
  NAND2_X1 U2641 ( .A1(n3240), .A2(n2492), .ZN(n3232) );
  NAND2_X1 U2642 ( .A1(n2152), .A2(n2155), .ZN(n2959) );
  NAND2_X1 U2643 ( .A1(n2382), .A2(n2087), .ZN(n2152) );
  INV_X1 U2644 ( .A(n2792), .ZN(n3521) );
  OAI211_X1 U2645 ( .C1(n3441), .C2(n2714), .A(n2698), .B(n2697), .ZN(n3905)
         );
  OAI211_X1 U2646 ( .C1(n3470), .C2(n2714), .A(n2684), .B(n2683), .ZN(n3700)
         );
  INV_X1 U2647 ( .A(n3945), .ZN(n3701) );
  NAND4_X1 U2648 ( .A1(n2660), .A2(n2659), .A3(n2658), .A4(n2657), .ZN(n3960)
         );
  NAND4_X1 U2649 ( .A1(n2645), .A2(n2644), .A3(n2643), .A4(n2642), .ZN(n3942)
         );
  NAND4_X1 U2650 ( .A1(n2614), .A2(n2613), .A3(n2612), .A4(n2611), .ZN(n4021)
         );
  INV_X1 U2651 ( .A(n3452), .ZN(n4070) );
  INV_X1 U2652 ( .A(n3384), .ZN(n3704) );
  OR2_X1 U2653 ( .A1(n2348), .A2(n2811), .ZN(n3709) );
  AND2_X1 U2654 ( .A1(n2843), .A2(n2844), .ZN(n3716) );
  INV_X1 U2655 ( .A(n2853), .ZN(n3752) );
  XNOR2_X1 U2656 ( .A(n2187), .B(n2916), .ZN(n2913) );
  XNOR2_X1 U2657 ( .A(n2874), .B(n2916), .ZN(n2914) );
  NAND2_X1 U2658 ( .A1(n2198), .A2(n2875), .ZN(n2892) );
  NAND2_X1 U2659 ( .A1(n2200), .A2(REG1_REG_8__SCAN_IN), .ZN(n2199) );
  INV_X1 U2660 ( .A(n2202), .ZN(n2201) );
  OAI21_X1 U2661 ( .B1(n4286), .B2(n2224), .A(n2223), .ZN(n4295) );
  NAND2_X1 U2662 ( .A1(n2225), .A2(REG1_REG_10__SCAN_IN), .ZN(n2224) );
  NAND2_X1 U2663 ( .A1(n3781), .A2(n2225), .ZN(n2223) );
  INV_X1 U2664 ( .A(n4296), .ZN(n2225) );
  NAND2_X1 U2665 ( .A1(n4291), .A2(n3763), .ZN(n4300) );
  NAND2_X1 U2666 ( .A1(n2227), .A2(n2226), .ZN(n4339) );
  AND2_X1 U2667 ( .A1(n3716), .A2(n3692), .ZN(n4373) );
  AOI21_X1 U2668 ( .B1(n4369), .B2(n2062), .A(n4368), .ZN(n4374) );
  AOI21_X1 U2669 ( .B1(n4364), .B2(n4363), .A(n4362), .ZN(n4369) );
  NAND2_X1 U2670 ( .A1(n4335), .A2(n4402), .ZN(n2190) );
  NAND2_X1 U2671 ( .A1(n2216), .A2(n2219), .ZN(n2215) );
  OR2_X1 U2672 ( .A1(n4363), .A2(n2220), .ZN(n2219) );
  INV_X1 U2673 ( .A(n3800), .ZN(n2220) );
  XNOR2_X1 U2674 ( .A(n4131), .B(n4125), .ZN(n4278) );
  AOI21_X1 U2675 ( .B1(n4136), .B2(n4133), .A(n4132), .ZN(n4282) );
  NAND2_X1 U2676 ( .A1(n3820), .A2(n3826), .ZN(n2126) );
  AOI21_X1 U2677 ( .B1(n3824), .B2(n2124), .A(n2123), .ZN(n2122) );
  NAND2_X1 U2678 ( .A1(n3825), .A2(n2124), .ZN(n2117) );
  AOI21_X1 U2679 ( .B1(n3857), .B2(n3349), .A(n3348), .ZN(n3841) );
  NAND2_X1 U2680 ( .A1(n2110), .A2(n2113), .ZN(n3973) );
  NAND2_X1 U2681 ( .A1(n4015), .A2(n2114), .ZN(n2110) );
  AND2_X1 U2682 ( .A1(n4118), .A2(n3807), .ZN(n4027) );
  NAND2_X1 U2683 ( .A1(n3044), .A2(n3043), .ZN(n3078) );
  AND2_X1 U2684 ( .A1(n4027), .A2(n4443), .ZN(n4378) );
  OAI21_X1 U2685 ( .B1(n2969), .B2(n3037), .A(n4115), .ZN(n4396) );
  INV_X1 U2686 ( .A(n4115), .ZN(n4392) );
  INV_X1 U2687 ( .A(n4474), .ZN(n4472) );
  INV_X1 U2688 ( .A(n4278), .ZN(n4209) );
  OAI21_X1 U2689 ( .B1(n3871), .B2(n3870), .A(n3869), .ZN(n4218) );
  AND2_X1 U2690 ( .A1(n4043), .A2(n3335), .ZN(n4008) );
  AND2_X2 U2691 ( .A1(n3038), .A2(n3032), .ZN(n4463) );
  AND2_X1 U2692 ( .A1(n2770), .A2(n2769), .ZN(n2825) );
  NAND2_X1 U2693 ( .A1(n2926), .A2(n3026), .ZN(n4399) );
  INV_X1 U2694 ( .A(IR_REG_30__SCAN_IN), .ZN(n2289) );
  OR2_X1 U2695 ( .A1(n2819), .A2(n2820), .ZN(n2095) );
  INV_X1 U2696 ( .A(n3732), .ZN(n4264) );
  NAND2_X1 U2697 ( .A1(n2306), .A2(n2305), .ZN(n2815) );
  AOI21_X1 U2698 ( .B1(n2304), .B2(IR_REG_25__SCAN_IN), .A(n2303), .ZN(n2305)
         );
  AND2_X1 U2699 ( .A1(n2820), .A2(n2286), .ZN(n2303) );
  AND2_X1 U2700 ( .A1(n2831), .A2(STATE_REG_SCAN_IN), .ZN(n4400) );
  INV_X1 U2701 ( .A(n3686), .ZN(n4268) );
  XNOR2_X1 U2702 ( .A(n2328), .B(IR_REG_19__SCAN_IN), .ZN(n4269) );
  AND2_X1 U2703 ( .A1(n2388), .A2(n2373), .ZN(n4275) );
  NAND2_X1 U2704 ( .A1(n2196), .A2(n2195), .ZN(n2194) );
  NAND2_X1 U2705 ( .A1(n2820), .A2(n2280), .ZN(n2195) );
  XNOR2_X1 U2706 ( .A(n2162), .B(n3506), .ZN(n3513) );
  INV_X1 U2707 ( .A(n2189), .ZN(n2878) );
  INV_X1 U2708 ( .A(n2208), .ZN(n2207) );
  OAI21_X1 U2709 ( .B1(n4370), .B2(n2211), .A(n2210), .ZN(n2209) );
  NAND2_X2 U2710 ( .A1(n2984), .A2(n2348), .ZN(n2661) );
  INV_X2 U2711 ( .A(n2682), .ZN(n3533) );
  NAND2_X1 U2712 ( .A1(n2580), .A2(n2579), .ZN(n3448) );
  OAI21_X1 U2713 ( .B1(n2260), .B2(n2258), .A(n2255), .ZN(n3320) );
  INV_X1 U2714 ( .A(n3504), .ZN(n2233) );
  AND2_X1 U2715 ( .A1(n3999), .A2(n3974), .ZN(n2057) );
  INV_X1 U2716 ( .A(n4083), .ZN(n4102) );
  AND4_X1 U2717 ( .A1(n2543), .A2(n2542), .A3(n2541), .A4(n2540), .ZN(n4083)
         );
  AND2_X1 U2718 ( .A1(n3716), .A2(n3732), .ZN(n4335) );
  AND2_X1 U2719 ( .A1(n2181), .A2(n3891), .ZN(n2058) );
  AND2_X1 U2720 ( .A1(n2058), .A2(n3870), .ZN(n2059) );
  OAI211_X1 U2721 ( .C1(n3533), .C2(n4464), .A(n2271), .B(n2346), .ZN(n2975)
         );
  OR2_X1 U2722 ( .A1(n3787), .A2(n4409), .ZN(n2060) );
  INV_X1 U2723 ( .A(n2340), .ZN(n2971) );
  AND2_X1 U2724 ( .A1(n3050), .A2(n3080), .ZN(n2061) );
  XNOR2_X1 U2725 ( .A(n2292), .B(n2291), .ZN(n2331) );
  NAND2_X1 U2726 ( .A1(n3937), .A2(n3341), .ZN(n3916) );
  OR2_X1 U2727 ( .A1(n4364), .A2(n4363), .ZN(n2062) );
  AND3_X1 U2728 ( .A1(n2297), .A2(n2296), .A3(n2295), .ZN(n3006) );
  AND3_X1 U2729 ( .A1(n2156), .A2(n2246), .A3(n2279), .ZN(n2063) );
  AND3_X1 U2730 ( .A1(n2282), .A2(n2251), .A3(n2178), .ZN(n2064) );
  NAND2_X1 U2731 ( .A1(n2590), .A2(n2266), .ZN(n2312) );
  NAND2_X1 U2732 ( .A1(n2590), .A2(n2265), .ZN(n2307) );
  NAND2_X1 U2733 ( .A1(n3392), .A2(n2676), .ZN(n3391) );
  OR2_X1 U2734 ( .A1(n2312), .A2(IR_REG_21__SCAN_IN), .ZN(n2065) );
  NAND2_X1 U2735 ( .A1(n2946), .A2(n2406), .ZN(n2066) );
  NAND2_X1 U2736 ( .A1(n4271), .A2(REG1_REG_7__SCAN_IN), .ZN(n2067) );
  AND2_X1 U2737 ( .A1(n3288), .A2(n3287), .ZN(n2068) );
  INV_X1 U2738 ( .A(n3263), .ZN(n3705) );
  AND4_X1 U2739 ( .A1(n2499), .A2(n2498), .A3(n2497), .A4(n2496), .ZN(n3263)
         );
  OR2_X1 U2740 ( .A1(n2168), .A2(n2164), .ZN(n2069) );
  NOR2_X1 U2741 ( .A1(n3288), .A2(n3287), .ZN(n2070) );
  AND2_X1 U2742 ( .A1(n4374), .A2(n2190), .ZN(n2071) );
  AND2_X1 U2743 ( .A1(n2875), .A2(n2067), .ZN(n2072) );
  NAND2_X1 U2744 ( .A1(n3391), .A2(n2686), .ZN(n3467) );
  AND2_X1 U2745 ( .A1(n2229), .A2(n2060), .ZN(n2073) );
  INV_X1 U2746 ( .A(n2899), .ZN(n2200) );
  AND2_X1 U2747 ( .A1(n2772), .A2(n2309), .ZN(n2074) );
  OR2_X1 U2748 ( .A1(n3867), .A2(n3851), .ZN(n2075) );
  INV_X1 U2749 ( .A(n3284), .ZN(n3277) );
  AND3_X1 U2750 ( .A1(n2252), .A2(n2251), .A3(n2321), .ZN(n2544) );
  INV_X1 U2751 ( .A(n2150), .ZN(n2149) );
  NAND2_X1 U2752 ( .A1(n2238), .A2(n2151), .ZN(n2150) );
  NOR2_X1 U2753 ( .A1(n2588), .A2(IR_REG_17__SCAN_IN), .ZN(n2590) );
  INV_X1 U2754 ( .A(n4112), .ZN(n4100) );
  AND2_X1 U2755 ( .A1(n2075), .A2(n3349), .ZN(n2076) );
  OR2_X1 U2756 ( .A1(n3517), .A2(n4060), .ZN(n2077) );
  AND2_X1 U2757 ( .A1(n2437), .A2(n2436), .ZN(n2078) );
  OR2_X1 U2758 ( .A1(n4666), .A2(n3761), .ZN(n2079) );
  AND2_X1 U2759 ( .A1(n2182), .A2(n4112), .ZN(n2080) );
  AND2_X1 U2760 ( .A1(n3452), .A2(n3354), .ZN(n2081) );
  AND2_X1 U2761 ( .A1(n3921), .A2(n3361), .ZN(n3938) );
  AND2_X1 U2762 ( .A1(n3961), .A2(n3984), .ZN(n2082) );
  AND2_X1 U2763 ( .A1(n3701), .A2(n3363), .ZN(n2083) );
  INV_X1 U2764 ( .A(n4038), .ZN(n3702) );
  AND4_X1 U2765 ( .A1(n2603), .A2(n2602), .A3(n2601), .A4(n2600), .ZN(n4038)
         );
  INV_X1 U2766 ( .A(n2115), .ZN(n2114) );
  OR2_X1 U2767 ( .A1(n3809), .A2(n3811), .ZN(n3820) );
  NOR2_X1 U2768 ( .A1(n3701), .A2(n3363), .ZN(n2084) );
  NAND2_X1 U2769 ( .A1(n2237), .A2(n2560), .ZN(n3447) );
  NAND2_X1 U2770 ( .A1(n2142), .A2(n2145), .ZN(n3457) );
  OAI22_X1 U2771 ( .A1(n3136), .A2(n3135), .B1(n3134), .B2(n3710), .ZN(n3217)
         );
  NAND2_X1 U2772 ( .A1(n2382), .A2(n2381), .ZN(n2945) );
  NOR2_X1 U2773 ( .A1(n2301), .A2(n2300), .ZN(n2756) );
  INV_X1 U2774 ( .A(n2106), .ZN(n3105) );
  INV_X1 U2775 ( .A(n4025), .ZN(n3335) );
  NAND2_X1 U2776 ( .A1(n2243), .A2(n2242), .ZN(n3094) );
  NAND2_X1 U2777 ( .A1(n3286), .A2(n3285), .ZN(n3304) );
  NAND2_X1 U2778 ( .A1(n2245), .A2(n2244), .ZN(n2999) );
  NAND2_X1 U2779 ( .A1(n2160), .A2(n3095), .ZN(n3168) );
  NOR2_X1 U2780 ( .A1(n4285), .A2(n3781), .ZN(n2085) );
  NOR2_X1 U2781 ( .A1(n2904), .A2(n2201), .ZN(n2086) );
  NAND2_X1 U2782 ( .A1(n2487), .A2(n2486), .ZN(n3240) );
  INV_X1 U2783 ( .A(n3974), .ZN(n3984) );
  NAND2_X1 U2784 ( .A1(n2433), .A2(DATAI_20_), .ZN(n3974) );
  AND2_X1 U2785 ( .A1(n2156), .A2(n2279), .ZN(n2087) );
  INV_X1 U2786 ( .A(n3363), .ZN(n3928) );
  AND2_X1 U2787 ( .A1(n2433), .A2(DATAI_23_), .ZN(n3363) );
  AND2_X1 U2788 ( .A1(n2175), .A2(n3974), .ZN(n2088) );
  NAND2_X1 U2789 ( .A1(n2650), .A2(n2651), .ZN(n2089) );
  AND2_X1 U2790 ( .A1(n4402), .A2(REG1_REG_18__SCAN_IN), .ZN(n2090) );
  AND2_X1 U2791 ( .A1(n3789), .A2(REG2_REG_15__SCAN_IN), .ZN(n2091) );
  NAND2_X1 U2792 ( .A1(n3789), .A2(REG1_REG_15__SCAN_IN), .ZN(n2092) );
  INV_X1 U2793 ( .A(n3381), .ZN(n2147) );
  INV_X1 U2794 ( .A(n3870), .ZN(n3864) );
  INV_X1 U2795 ( .A(n3891), .ZN(n3342) );
  NAND2_X1 U2796 ( .A1(n2433), .A2(DATAI_25_), .ZN(n3891) );
  INV_X1 U2797 ( .A(n4359), .ZN(n4362) );
  INV_X1 U2798 ( .A(n2218), .ZN(n2217) );
  OR2_X1 U2799 ( .A1(n3800), .A2(n2090), .ZN(n2218) );
  INV_X1 U2800 ( .A(n2222), .ZN(n2221) );
  NAND2_X1 U2801 ( .A1(n4402), .A2(REG2_REG_18__SCAN_IN), .ZN(n2222) );
  NOR2_X1 U2802 ( .A1(n2290), .A2(IR_REG_29__SCAN_IN), .ZN(n2819) );
  INV_X1 U2803 ( .A(IR_REG_0__SCAN_IN), .ZN(n2174) );
  OAI21_X1 U2804 ( .B1(n3604), .B2(n2093), .A(n3047), .ZN(n3019) );
  NAND2_X1 U2805 ( .A1(n3014), .A2(n3013), .ZN(n2093) );
  OAI21_X2 U2806 ( .B1(n3068), .B2(n3067), .A(n3626), .ZN(n3113) );
  OAI21_X2 U2807 ( .B1(n3155), .B2(n3130), .A(n3632), .ZN(n3175) );
  NAND2_X2 U2808 ( .A1(n4063), .A2(n3549), .ZN(n3994) );
  NAND2_X2 U2809 ( .A1(n4062), .A2(n3600), .ZN(n4063) );
  OR2_X2 U2810 ( .A1(n4076), .A2(n3606), .ZN(n4077) );
  OAI21_X2 U2811 ( .B1(n3207), .B2(n3653), .A(n3634), .ZN(n3264) );
  AND3_X2 U2812 ( .A1(n2179), .A2(n2140), .A3(n2064), .ZN(n2302) );
  NOR2_X2 U2813 ( .A1(n2253), .A2(n2320), .ZN(n2140) );
  NAND2_X2 U2814 ( .A1(n3614), .A2(n3013), .ZN(n3602) );
  NOR2_X2 U2815 ( .A1(n3844), .A2(n3845), .ZN(n3843) );
  OAI21_X2 U2816 ( .B1(n3883), .B2(n3673), .A(n3364), .ZN(n3844) );
  OR2_X2 U2817 ( .A1(n3900), .A2(n3674), .ZN(n3883) );
  AOI21_X1 U2818 ( .B1(n3958), .B2(n3672), .A(n3553), .ZN(n3900) );
  NAND4_X1 U2819 ( .A1(n2100), .A2(n2099), .A3(n2098), .A4(n2097), .ZN(n2253)
         );
  AND2_X1 U2820 ( .A1(n2104), .A2(n3109), .ZN(n2103) );
  NAND2_X1 U2821 ( .A1(n2106), .A2(n3107), .ZN(n2105) );
  NAND2_X1 U2822 ( .A1(n4015), .A2(n2111), .ZN(n2108) );
  NAND2_X1 U2823 ( .A1(n2108), .A2(n2109), .ZN(n3956) );
  NAND2_X1 U2824 ( .A1(n4015), .A2(n3336), .ZN(n4003) );
  OR2_X1 U2825 ( .A1(n3337), .A2(n2116), .ZN(n2115) );
  INV_X1 U2826 ( .A(n3336), .ZN(n2116) );
  OAI211_X1 U2827 ( .C1(n3825), .C2(n2126), .A(n2122), .B(n2117), .ZN(n4138)
         );
  OAI21_X1 U2828 ( .B1(n3270), .B2(n2129), .A(n2127), .ZN(n4093) );
  INV_X1 U2829 ( .A(n3599), .ZN(n2131) );
  INV_X1 U2830 ( .A(n3270), .ZN(n2132) );
  OAI21_X1 U2831 ( .B1(n3936), .B2(n2135), .A(n2133), .ZN(n3877) );
  INV_X1 U2832 ( .A(n3938), .ZN(n2137) );
  INV_X1 U2833 ( .A(n3936), .ZN(n2138) );
  NAND2_X1 U2834 ( .A1(n2140), .A2(n2139), .ZN(n2588) );
  OAI22_X1 U2835 ( .A1(n3956), .A2(n3340), .B1(n3339), .B2(n3942), .ZN(n3936)
         );
  NOR2_X1 U2836 ( .A1(n3223), .A2(n3222), .ZN(n3269) );
  AOI21_X1 U2837 ( .B1(n4100), .B2(n3704), .A(n3289), .ZN(n3290) );
  NAND2_X1 U2838 ( .A1(n3010), .A2(n3009), .ZN(n3044) );
  OAI22_X1 U2839 ( .A1(n3269), .A2(n3268), .B1(n3267), .B2(n3266), .ZN(n3270)
         );
  NAND2_X1 U2840 ( .A1(n2971), .A2(n2973), .ZN(n3614) );
  NAND2_X1 U2841 ( .A1(n2141), .A2(n2143), .ZN(n2597) );
  NAND2_X1 U2842 ( .A1(n3380), .A2(n2145), .ZN(n2141) );
  NOR2_X1 U2843 ( .A1(n2155), .A2(n2154), .ZN(n2153) );
  NAND2_X1 U2844 ( .A1(n3094), .A2(n3095), .ZN(n2159) );
  NAND2_X1 U2845 ( .A1(n2159), .A2(n2158), .ZN(n2474) );
  INV_X1 U2846 ( .A(n3430), .ZN(n2163) );
  NAND2_X1 U2847 ( .A1(n2171), .A2(n2169), .ZN(n3392) );
  NOR2_X2 U2848 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2272)
         );
  MUX2_X1 U2849 ( .A(n2174), .B(n2173), .S(n2433), .Z(n4384) );
  NAND2_X4 U2850 ( .A1(n2172), .A2(n2326), .ZN(n2433) );
  NOR2_X1 U2851 ( .A1(n2176), .A2(n2588), .ZN(n2300) );
  NAND2_X1 U2852 ( .A1(n2191), .A2(n2071), .ZN(U3258) );
  NAND3_X1 U2853 ( .A1(n2193), .A2(n4373), .A3(n2192), .ZN(n2191) );
  NAND2_X1 U2854 ( .A1(n4371), .A2(n4372), .ZN(n2192) );
  NOR2_X2 U2855 ( .A1(n2321), .A2(n2194), .ZN(n4276) );
  NAND3_X1 U2856 ( .A1(n2197), .A2(IR_REG_2__SCAN_IN), .A3(IR_REG_31__SCAN_IN), 
        .ZN(n2196) );
  NAND2_X1 U2857 ( .A1(n2914), .A2(REG1_REG_6__SCAN_IN), .ZN(n2198) );
  NAND2_X1 U2858 ( .A1(n2198), .A2(n2072), .ZN(n2894) );
  OAI22_X1 U2859 ( .A1(n2199), .A2(n2905), .B1(n2202), .B2(n2899), .ZN(n3777)
         );
  NAND2_X1 U2860 ( .A1(n4364), .A2(n2205), .ZN(n2204) );
  OAI211_X1 U2861 ( .C1(n2209), .C2(n2207), .A(n2206), .B(n2203), .ZN(U3259)
         );
  OAI211_X1 U2862 ( .C1(n4364), .C2(n2215), .A(n2204), .B(n4359), .ZN(n2203)
         );
  AND2_X1 U2863 ( .A1(n2216), .A2(n2218), .ZN(n2205) );
  INV_X1 U2864 ( .A(n2229), .ZN(n4325) );
  NAND2_X1 U2865 ( .A1(n2707), .A2(n2230), .ZN(n2234) );
  NAND2_X1 U2866 ( .A1(n2340), .A2(n3418), .ZN(n3013) );
  NAND2_X1 U2867 ( .A1(n2321), .A2(n2272), .ZN(n2397) );
  AOI21_X1 U2868 ( .B1(n3240), .B2(n2263), .A(n2254), .ZN(n3254) );
  INV_X1 U2869 ( .A(n3240), .ZN(n2260) );
  AND2_X1 U2870 ( .A1(n2302), .A2(n2286), .ZN(n2298) );
  NAND2_X1 U2871 ( .A1(n2302), .A2(n2269), .ZN(n2290) );
  NAND2_X1 U2872 ( .A1(n3161), .A2(n3160), .ZN(n3159) );
  NAND2_X1 U2873 ( .A1(n2801), .A2(n2325), .ZN(n2323) );
  NAND2_X1 U2874 ( .A1(n4130), .A2(n4124), .ZN(n4131) );
  NAND2_X1 U2875 ( .A1(n2433), .A2(DATAI_1_), .ZN(n2338) );
  NAND2_X1 U2876 ( .A1(n3868), .A2(n3851), .ZN(n3850) );
  AND2_X1 U2877 ( .A1(n2975), .A2(n2974), .ZN(n2976) );
  AOI21_X1 U2878 ( .B1(n4443), .B2(n4140), .A(n4139), .ZN(n4141) );
  MUX2_X1 U2879 ( .A(n4313), .B(n2517), .S(n2433), .Z(n3309) );
  INV_X1 U2880 ( .A(IR_REG_25__SCAN_IN), .ZN(n2286) );
  AND2_X1 U2881 ( .A1(n2345), .A2(n2344), .ZN(n2271) );
  AND2_X1 U2882 ( .A1(n2429), .A2(n2428), .ZN(n2273) );
  NAND2_X1 U2883 ( .A1(n3707), .A2(n3218), .ZN(n2274) );
  AND2_X1 U2884 ( .A1(n2808), .A2(n2807), .ZN(n2275) );
  AND2_X1 U2885 ( .A1(n2776), .A2(n2775), .ZN(n2276) );
  NOR2_X1 U2886 ( .A1(n3721), .A2(n2331), .ZN(n2277) );
  AND2_X1 U2887 ( .A1(n2053), .A2(REG0_REG_2__SCAN_IN), .ZN(n2278) );
  INV_X1 U2888 ( .A(n4105), .ZN(n3288) );
  INV_X1 U2889 ( .A(n3309), .ZN(n3287) );
  INV_X1 U2890 ( .A(n3241), .ZN(n2486) );
  AND2_X1 U2891 ( .A1(n3976), .A2(n3356), .ZN(n3665) );
  INV_X1 U2892 ( .A(IR_REG_26__SCAN_IN), .ZN(n2287) );
  INV_X1 U2893 ( .A(IR_REG_2__SCAN_IN), .ZN(n2280) );
  AND2_X1 U2894 ( .A1(n3393), .A2(n3394), .ZN(n2676) );
  INV_X1 U2895 ( .A(n2745), .ZN(n2374) );
  NAND2_X1 U2896 ( .A1(n3184), .A2(n3183), .ZN(n3215) );
  INV_X1 U2897 ( .A(IR_REG_14__SCAN_IN), .ZN(n2557) );
  AND2_X1 U2898 ( .A1(n2622), .A2(n2623), .ZN(n2621) );
  OAI22_X1 U2899 ( .A1(n2340), .A2(n2661), .B1(n2745), .B2(n2973), .ZN(n2356)
         );
  NOR2_X1 U2900 ( .A1(n2815), .A2(n2769), .ZN(n2311) );
  AND2_X1 U2901 ( .A1(n2366), .A2(REG3_REG_2__SCAN_IN), .ZN(n2293) );
  OR3_X1 U2902 ( .A1(n2462), .A2(IR_REG_7__SCAN_IN), .A3(IR_REG_8__SCAN_IN), 
        .ZN(n2465) );
  OR2_X1 U2903 ( .A1(n3822), .A2(n3821), .ZN(n3823) );
  OR2_X1 U2904 ( .A1(n3345), .A2(n3344), .ZN(n3346) );
  OR2_X1 U2905 ( .A1(n2629), .A2(n3481), .ZN(n2640) );
  AND2_X1 U2906 ( .A1(n3703), .A2(n3462), .ZN(n3333) );
  NAND2_X1 U2907 ( .A1(n3137), .A2(n3632), .ZN(n3184) );
  INV_X1 U2908 ( .A(n3966), .ZN(n3339) );
  OR2_X1 U2909 ( .A1(n3190), .A2(n3189), .ZN(n3219) );
  OR2_X1 U2910 ( .A1(n2666), .A2(n4633), .ZN(n2680) );
  OR2_X1 U2911 ( .A1(n2439), .A2(n2438), .ZN(n2456) );
  INV_X1 U2912 ( .A(n3960), .ZN(n3431) );
  AND2_X1 U2913 ( .A1(n2582), .A2(REG3_REG_17__SCAN_IN), .ZN(n2598) );
  OR2_X1 U2914 ( .A1(n2456), .A2(n2891), .ZN(n2476) );
  NOR2_X1 U2915 ( .A1(n2523), .A2(n3324), .ZN(n2538) );
  OR2_X1 U2916 ( .A1(n2551), .A2(n3516), .ZN(n2562) );
  AND2_X1 U2917 ( .A1(n2708), .A2(REG3_REG_26__SCAN_IN), .ZN(n2724) );
  NOR2_X1 U2918 ( .A1(n3785), .A2(n4304), .ZN(n4316) );
  INV_X1 U2919 ( .A(n4365), .ZN(n4366) );
  INV_X1 U2920 ( .A(n3699), .ZN(n3867) );
  NAND2_X1 U2921 ( .A1(n4085), .A2(n3354), .ZN(n4054) );
  INV_X1 U2922 ( .A(n3184), .ZN(n3629) );
  INV_X1 U2923 ( .A(n3009), .ZN(n3604) );
  INV_X1 U2924 ( .A(n3026), .ZN(n3028) );
  INV_X1 U2925 ( .A(n3265), .ZN(n3266) );
  AND2_X1 U2926 ( .A1(n2970), .A2(n3559), .ZN(n4065) );
  NAND2_X1 U2927 ( .A1(n2348), .A2(n4400), .ZN(n3024) );
  INV_X1 U2928 ( .A(n4045), .ZN(n3462) );
  AND3_X1 U2929 ( .A1(n3536), .A2(n3535), .A3(n3534), .ZN(n3561) );
  INV_X1 U2930 ( .A(n2366), .ZN(n2714) );
  NOR2_X1 U2931 ( .A1(n2466), .A2(n2501), .ZN(n3778) );
  AND2_X1 U2932 ( .A1(n3716), .A2(n2837), .ZN(n4359) );
  OR2_X1 U2933 ( .A1(n3217), .A2(n3629), .ZN(n4446) );
  AND2_X1 U2934 ( .A1(n3625), .A2(n3640), .ZN(n3591) );
  AOI21_X1 U2935 ( .B1(n3028), .B2(n4501), .A(n2825), .ZN(n3037) );
  NAND2_X1 U2936 ( .A1(n2433), .A2(DATAI_21_), .ZN(n3966) );
  AND2_X1 U2937 ( .A1(n4385), .A2(n2790), .ZN(n4460) );
  NAND2_X1 U2938 ( .A1(n2757), .A2(n2756), .ZN(n3026) );
  INV_X1 U2939 ( .A(n3428), .ZN(n3525) );
  NAND2_X1 U2940 ( .A1(n2731), .A2(n2730), .ZN(n3699) );
  INV_X1 U2941 ( .A(n4275), .ZN(n2848) );
  INV_X1 U2942 ( .A(n4373), .ZN(n4328) );
  INV_X1 U2943 ( .A(n4412), .ZN(n4313) );
  INV_X1 U2944 ( .A(n4005), .ZN(n4092) );
  INV_X1 U2945 ( .A(n4378), .ZN(n4088) );
  NAND2_X1 U2946 ( .A1(n4474), .A2(n4443), .ZN(n4206) );
  AND2_X2 U2947 ( .A1(n3038), .A2(n3037), .ZN(n4474) );
  NAND2_X1 U2948 ( .A1(n4463), .A2(n4443), .ZN(n4261) );
  INV_X1 U2949 ( .A(n4463), .ZN(n4461) );
  INV_X1 U2950 ( .A(n4399), .ZN(n4398) );
  INV_X1 U2951 ( .A(n2332), .ZN(n4263) );
  INV_X1 U2952 ( .A(n2790), .ZN(n4266) );
  INV_X1 U2953 ( .A(n3786), .ZN(n4411) );
  INV_X1 U2954 ( .A(n3709), .ZN(U4043) );
  NAND2_X1 U2955 ( .A1(n2319), .A2(n2280), .ZN(n2320) );
  NOR2_X1 U2956 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2288)
         );
  INV_X1 U2957 ( .A(IR_REG_29__SCAN_IN), .ZN(n2291) );
  NOR2_X1 U2958 ( .A1(n2278), .A2(n2293), .ZN(n2297) );
  INV_X1 U2959 ( .A(n2331), .ZN(n2294) );
  NOR2_X2 U2960 ( .A1(n2332), .A2(n2294), .ZN(n2343) );
  NAND2_X1 U2961 ( .A1(n2343), .A2(REG2_REG_2__SCAN_IN), .ZN(n2295) );
  INV_X1 U2962 ( .A(IR_REG_31__SCAN_IN), .ZN(n2820) );
  NOR2_X1 U2963 ( .A1(n2298), .A2(n2820), .ZN(n2299) );
  MUX2_X1 U2964 ( .A(n2820), .B(n2299), .S(IR_REG_26__SCAN_IN), .Z(n2301) );
  INV_X1 U2965 ( .A(n2298), .ZN(n2306) );
  NOR2_X1 U2966 ( .A1(n2302), .A2(n2820), .ZN(n2304) );
  NAND2_X1 U2967 ( .A1(n2307), .A2(IR_REG_31__SCAN_IN), .ZN(n2773) );
  NAND2_X1 U2968 ( .A1(n2773), .A2(n2772), .ZN(n2308) );
  NAND2_X1 U2969 ( .A1(n2312), .A2(IR_REG_31__SCAN_IN), .ZN(n2313) );
  MUX2_X1 U2970 ( .A(IR_REG_31__SCAN_IN), .B(n2313), .S(IR_REG_21__SCAN_IN), 
        .Z(n2314) );
  NAND2_X1 U2971 ( .A1(n2314), .A2(n2065), .ZN(n3579) );
  INV_X1 U2972 ( .A(IR_REG_19__SCAN_IN), .ZN(n2315) );
  NAND2_X1 U2973 ( .A1(n2328), .A2(n2315), .ZN(n2316) );
  NAND2_X1 U2974 ( .A1(n2316), .A2(IR_REG_31__SCAN_IN), .ZN(n2318) );
  INV_X1 U2975 ( .A(n2320), .ZN(n2321) );
  NAND2_X1 U2976 ( .A1(n2325), .A2(IR_REG_27__SCAN_IN), .ZN(n2326) );
  MUX2_X1 U2977 ( .A(n4276), .B(DATAI_2_), .S(n2433), .Z(n3034) );
  INV_X1 U2978 ( .A(n3034), .ZN(n3042) );
  NAND2_X1 U2979 ( .A1(n2065), .A2(IR_REG_31__SCAN_IN), .ZN(n2327) );
  NAND2_X1 U2980 ( .A1(n2790), .A2(n3579), .ZN(n4383) );
  INV_X1 U2981 ( .A(n4383), .ZN(n2330) );
  OAI22_X1 U2982 ( .A1(n3006), .A2(n2748), .B1(n3042), .B2(n2661), .ZN(n2361)
         );
  XNOR2_X1 U2983 ( .A(n2360), .B(n2361), .ZN(n2930) );
  NAND2_X1 U2984 ( .A1(n2366), .A2(REG3_REG_1__SCAN_IN), .ZN(n2336) );
  INV_X1 U2985 ( .A(REG1_REG_1__SCAN_IN), .ZN(n3721) );
  NAND2_X1 U2986 ( .A1(n2277), .A2(n2332), .ZN(n2334) );
  NAND2_X1 U2987 ( .A1(n2343), .A2(REG2_REG_1__SCAN_IN), .ZN(n2333) );
  NAND2_X1 U2988 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2337)
         );
  INV_X1 U2989 ( .A(n4277), .ZN(n2339) );
  XOR2_X1 U2990 ( .A(n2356), .B(n2734), .Z(n2341) );
  OAI22_X1 U2991 ( .A1(n2340), .A2(n2748), .B1(n2661), .B2(n2973), .ZN(n2357)
         );
  NAND2_X1 U2992 ( .A1(n2341), .A2(n2357), .ZN(n2932) );
  INV_X1 U2993 ( .A(n2932), .ZN(n2342) );
  NOR2_X1 U2994 ( .A1(n2930), .A2(n2342), .ZN(n2359) );
  INV_X1 U2995 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4464) );
  NAND2_X1 U2996 ( .A1(n2366), .A2(REG3_REG_0__SCAN_IN), .ZN(n2345) );
  NAND2_X1 U2997 ( .A1(n2343), .A2(REG2_REG_0__SCAN_IN), .ZN(n2344) );
  NAND2_X1 U2998 ( .A1(n2054), .A2(REG0_REG_0__SCAN_IN), .ZN(n2346) );
  INV_X1 U2999 ( .A(n2975), .ZN(n2347) );
  INV_X1 U3000 ( .A(n2348), .ZN(n2349) );
  AOI22_X1 U3001 ( .A1(n2974), .A2(n2051), .B1(IR_REG_0__SCAN_IN), .B2(n2349), 
        .ZN(n2350) );
  NAND2_X1 U3002 ( .A1(n2351), .A2(n2350), .ZN(n2922) );
  AND2_X1 U3003 ( .A1(n2974), .A2(n2374), .ZN(n2352) );
  OR2_X1 U3004 ( .A1(n2348), .A2(n4464), .ZN(n2353) );
  NAND2_X1 U3005 ( .A1(n2354), .A2(n2353), .ZN(n2923) );
  NAND2_X1 U3006 ( .A1(n2922), .A2(n2923), .ZN(n2921) );
  NAND2_X1 U3007 ( .A1(n2354), .A2(n2734), .ZN(n2355) );
  NAND2_X1 U3008 ( .A1(n2921), .A2(n2355), .ZN(n3415) );
  XNOR2_X1 U3009 ( .A(n2356), .B(n2734), .ZN(n2358) );
  XNOR2_X1 U3010 ( .A(n2358), .B(n2357), .ZN(n3416) );
  NAND2_X1 U3011 ( .A1(n3415), .A2(n3416), .ZN(n2931) );
  NAND2_X1 U3012 ( .A1(n2359), .A2(n2931), .ZN(n2933) );
  INV_X1 U3013 ( .A(n2360), .ZN(n2363) );
  INV_X1 U3014 ( .A(n2361), .ZN(n2362) );
  NAND2_X1 U3015 ( .A1(n2363), .A2(n2362), .ZN(n2364) );
  NAND2_X1 U3016 ( .A1(n2933), .A2(n2364), .ZN(n2939) );
  INV_X1 U3017 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2365) );
  INV_X1 U3018 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3088) );
  NAND2_X1 U3019 ( .A1(n2668), .A2(n3088), .ZN(n2369) );
  NAND2_X1 U3020 ( .A1(n2055), .A2(REG0_REG_3__SCAN_IN), .ZN(n2368) );
  NAND2_X1 U3021 ( .A1(n2343), .A2(REG2_REG_3__SCAN_IN), .ZN(n2367) );
  NAND2_X1 U3022 ( .A1(n3050), .A2(n2051), .ZN(n2376) );
  NAND2_X1 U3023 ( .A1(n2320), .A2(IR_REG_31__SCAN_IN), .ZN(n2372) );
  NAND2_X1 U3024 ( .A1(n2372), .A2(n2371), .ZN(n2388) );
  OR2_X1 U3025 ( .A1(n2372), .A2(n2371), .ZN(n2373) );
  MUX2_X1 U3026 ( .A(n4275), .B(DATAI_3_), .S(n2433), .Z(n3080) );
  NAND2_X1 U3027 ( .A1(n3080), .A2(n2374), .ZN(n2375) );
  AOI22_X1 U3028 ( .A1(n3050), .A2(n2737), .B1(n3080), .B2(n2051), .ZN(n2379)
         );
  XNOR2_X1 U3029 ( .A(n2378), .B(n2379), .ZN(n2940) );
  NAND2_X1 U3030 ( .A1(n2939), .A2(n2940), .ZN(n2382) );
  INV_X1 U3031 ( .A(n2378), .ZN(n2380) );
  NAND2_X1 U3032 ( .A1(n2380), .A2(n2379), .ZN(n2381) );
  NAND2_X1 U3033 ( .A1(n2056), .A2(REG0_REG_4__SCAN_IN), .ZN(n2387) );
  OAI21_X1 U3034 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        n2411), .ZN(n3057) );
  INV_X1 U3035 ( .A(n3057), .ZN(n2997) );
  NAND2_X1 U3036 ( .A1(n2668), .A2(n2997), .ZN(n2386) );
  NAND2_X1 U3037 ( .A1(n2343), .A2(REG2_REG_4__SCAN_IN), .ZN(n2385) );
  INV_X1 U3038 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2862) );
  OR2_X1 U3039 ( .A1(n3533), .A2(n2862), .ZN(n2384) );
  NAND2_X1 U3040 ( .A1(n2388), .A2(IR_REG_31__SCAN_IN), .ZN(n2389) );
  MUX2_X1 U3041 ( .A(n4274), .B(DATAI_4_), .S(n2433), .Z(n3064) );
  OAI22_X1 U3042 ( .A1(n3070), .A2(n2661), .B1(n2745), .B2(n3055), .ZN(n2390)
         );
  XNOR2_X1 U3043 ( .A(n2390), .B(n2746), .ZN(n2392) );
  OAI22_X1 U3044 ( .A1(n3070), .A2(n2748), .B1(n2661), .B2(n3055), .ZN(n2391)
         );
  XNOR2_X1 U3045 ( .A(n2392), .B(n2391), .ZN(n2994) );
  NAND2_X1 U3046 ( .A1(n2392), .A2(n2391), .ZN(n2946) );
  NAND2_X1 U3047 ( .A1(n2053), .A2(REG0_REG_5__SCAN_IN), .ZN(n2396) );
  XNOR2_X1 U3048 ( .A(n2411), .B(REG3_REG_5__SCAN_IN), .ZN(n3075) );
  NAND2_X1 U3049 ( .A1(n2668), .A2(n3075), .ZN(n2395) );
  NAND2_X1 U3050 ( .A1(n2343), .A2(REG2_REG_5__SCAN_IN), .ZN(n2394) );
  INV_X1 U3051 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2857) );
  OR2_X1 U3052 ( .A1(n3533), .A2(n2857), .ZN(n2393) );
  NAND2_X1 U3053 ( .A1(n2397), .A2(IR_REG_31__SCAN_IN), .ZN(n2398) );
  MUX2_X1 U3054 ( .A(IR_REG_31__SCAN_IN), .B(n2398), .S(IR_REG_5__SCAN_IN), 
        .Z(n2400) );
  INV_X1 U3055 ( .A(n2432), .ZN(n2399) );
  NAND2_X1 U3056 ( .A1(n2400), .A2(n2399), .ZN(n2871) );
  INV_X1 U3057 ( .A(DATAI_5_), .ZN(n2401) );
  MUX2_X1 U3058 ( .A(n2871), .B(n2401), .S(n2433), .Z(n3106) );
  OAI22_X1 U3059 ( .A1(n3115), .A2(n2661), .B1(n2745), .B2(n3106), .ZN(n2402)
         );
  XNOR2_X1 U3060 ( .A(n2402), .B(n2734), .ZN(n2405) );
  INV_X1 U3061 ( .A(n2405), .ZN(n2403) );
  OAI22_X1 U3062 ( .A1(n3115), .A2(n2748), .B1(n2661), .B2(n3106), .ZN(n2404)
         );
  NAND2_X1 U3063 ( .A1(n2403), .A2(n2404), .ZN(n2406) );
  XNOR2_X1 U3064 ( .A(n2405), .B(n2404), .ZN(n2948) );
  INV_X1 U3065 ( .A(n2406), .ZN(n2407) );
  INV_X1 U3066 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2408) );
  OR2_X1 U3067 ( .A1(n3533), .A2(n2408), .ZN(n2416) );
  NAND2_X1 U3068 ( .A1(n2056), .A2(REG0_REG_6__SCAN_IN), .ZN(n2415) );
  INV_X1 U3069 ( .A(n2411), .ZN(n2409) );
  AOI21_X1 U3070 ( .B1(n2409), .B2(REG3_REG_5__SCAN_IN), .A(
        REG3_REG_6__SCAN_IN), .ZN(n2412) );
  NAND2_X1 U3071 ( .A1(REG3_REG_5__SCAN_IN), .A2(REG3_REG_6__SCAN_IN), .ZN(
        n2410) );
  OR2_X1 U3072 ( .A1(n2412), .A2(n2423), .ZN(n3147) );
  INV_X1 U3073 ( .A(n3147), .ZN(n2962) );
  NAND2_X1 U3074 ( .A1(n2668), .A2(n2962), .ZN(n2414) );
  NAND2_X1 U3075 ( .A1(n2343), .A2(REG2_REG_6__SCAN_IN), .ZN(n2413) );
  NAND4_X1 U3076 ( .A1(n2416), .A2(n2415), .A3(n2414), .A4(n2413), .ZN(n3710)
         );
  NAND2_X1 U3077 ( .A1(n3710), .A2(n2737), .ZN(n2419) );
  OR2_X1 U3078 ( .A1(n2432), .A2(n2820), .ZN(n2417) );
  XNOR2_X1 U3079 ( .A(n2417), .B(IR_REG_6__SCAN_IN), .ZN(n4272) );
  MUX2_X1 U3080 ( .A(n4272), .B(DATAI_6_), .S(n2433), .Z(n3134) );
  NAND2_X1 U3081 ( .A1(n3134), .A2(n2051), .ZN(n2418) );
  NAND2_X1 U3082 ( .A1(n2419), .A2(n2418), .ZN(n2957) );
  NAND2_X1 U3083 ( .A1(n3710), .A2(n2051), .ZN(n2421) );
  NAND2_X1 U3084 ( .A1(n3134), .A2(n2374), .ZN(n2420) );
  NAND2_X1 U3085 ( .A1(n2421), .A2(n2420), .ZN(n2422) );
  XNOR2_X1 U3086 ( .A(n2422), .B(n2746), .ZN(n2956) );
  NAND2_X1 U3087 ( .A1(n2423), .A2(REG3_REG_7__SCAN_IN), .ZN(n2439) );
  OR2_X1 U3088 ( .A1(n2423), .A2(REG3_REG_7__SCAN_IN), .ZN(n2424) );
  AND2_X1 U3089 ( .A1(n2439), .A2(n2424), .ZN(n3162) );
  NAND2_X1 U3090 ( .A1(n2668), .A2(n3162), .ZN(n2426) );
  NAND2_X1 U3091 ( .A1(n2055), .A2(REG0_REG_7__SCAN_IN), .ZN(n2425) );
  INV_X1 U3092 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2427) );
  OR2_X1 U3093 ( .A1(n3533), .A2(n2427), .ZN(n2429) );
  NAND2_X1 U3094 ( .A1(n2343), .A2(REG2_REG_7__SCAN_IN), .ZN(n2428) );
  NAND2_X1 U3095 ( .A1(n2432), .A2(n2431), .ZN(n2462) );
  NAND2_X1 U3096 ( .A1(n2462), .A2(IR_REG_31__SCAN_IN), .ZN(n2447) );
  XNOR2_X1 U3097 ( .A(n2447), .B(IR_REG_7__SCAN_IN), .ZN(n4271) );
  MUX2_X1 U3098 ( .A(n4271), .B(DATAI_7_), .S(n2433), .Z(n3138) );
  OAI22_X1 U3099 ( .A1(n3129), .A2(n2661), .B1(n2745), .B2(n3160), .ZN(n2434)
         );
  XNOR2_X1 U3100 ( .A(n2434), .B(n2734), .ZN(n2435) );
  OAI22_X1 U3101 ( .A1(n3129), .A2(n2748), .B1(n2661), .B2(n3160), .ZN(n2436)
         );
  XNOR2_X1 U3102 ( .A(n2435), .B(n2436), .ZN(n3000) );
  INV_X1 U3103 ( .A(n2435), .ZN(n2437) );
  NAND2_X1 U3104 ( .A1(n2054), .A2(REG0_REG_8__SCAN_IN), .ZN(n2445) );
  NAND2_X1 U3105 ( .A1(n2439), .A2(n2438), .ZN(n2440) );
  AND2_X1 U3106 ( .A1(n2456), .A2(n2440), .ZN(n3141) );
  NAND2_X1 U3107 ( .A1(n2668), .A2(n3141), .ZN(n2444) );
  NAND2_X1 U3108 ( .A1(n2343), .A2(REG2_REG_8__SCAN_IN), .ZN(n2443) );
  INV_X1 U3109 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2441) );
  OR2_X1 U3110 ( .A1(n3533), .A2(n2441), .ZN(n2442) );
  INV_X1 U3111 ( .A(IR_REG_7__SCAN_IN), .ZN(n2446) );
  NAND2_X1 U3112 ( .A1(n2447), .A2(n2446), .ZN(n2448) );
  NAND2_X1 U3113 ( .A1(n2448), .A2(IR_REG_31__SCAN_IN), .ZN(n2450) );
  INV_X1 U3114 ( .A(IR_REG_8__SCAN_IN), .ZN(n2449) );
  XNOR2_X1 U3115 ( .A(n2450), .B(n2449), .ZN(n2908) );
  INV_X1 U3116 ( .A(DATAI_8_), .ZN(n2812) );
  MUX2_X1 U3117 ( .A(n2908), .B(n2812), .S(n2433), .Z(n3181) );
  OAI22_X1 U3118 ( .A1(n3182), .A2(n2661), .B1(n2745), .B2(n3181), .ZN(n2451)
         );
  XNOR2_X1 U3119 ( .A(n2451), .B(n2746), .ZN(n2452) );
  OAI22_X1 U3120 ( .A1(n3182), .A2(n2748), .B1(n2661), .B2(n3181), .ZN(n2453)
         );
  AND2_X1 U3121 ( .A1(n2452), .A2(n2453), .ZN(n3096) );
  INV_X1 U3122 ( .A(n2452), .ZN(n2455) );
  INV_X1 U3123 ( .A(n2453), .ZN(n2454) );
  NAND2_X1 U3124 ( .A1(n2455), .A2(n2454), .ZN(n3095) );
  INV_X1 U3125 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2898) );
  OR2_X1 U3126 ( .A1(n3533), .A2(n2898), .ZN(n2461) );
  NAND2_X1 U3127 ( .A1(n2053), .A2(REG0_REG_9__SCAN_IN), .ZN(n2460) );
  NAND2_X1 U3128 ( .A1(n2456), .A2(n2891), .ZN(n2457) );
  AND2_X1 U3129 ( .A1(n2476), .A2(n2457), .ZN(n3196) );
  NAND2_X1 U3130 ( .A1(n2668), .A2(n3196), .ZN(n2459) );
  NAND2_X1 U3131 ( .A1(n2343), .A2(REG2_REG_9__SCAN_IN), .ZN(n2458) );
  NAND4_X1 U3132 ( .A1(n2461), .A2(n2460), .A3(n2459), .A4(n2458), .ZN(n3707)
         );
  NAND2_X1 U3133 ( .A1(n3707), .A2(n2051), .ZN(n2468) );
  NAND2_X1 U3134 ( .A1(n2465), .A2(IR_REG_31__SCAN_IN), .ZN(n2463) );
  MUX2_X1 U3135 ( .A(IR_REG_31__SCAN_IN), .B(n2463), .S(IR_REG_9__SCAN_IN), 
        .Z(n2464) );
  INV_X1 U3136 ( .A(n2464), .ZN(n2466) );
  MUX2_X1 U3137 ( .A(n3778), .B(DATAI_9_), .S(n2433), .Z(n3218) );
  NAND2_X1 U3138 ( .A1(n3218), .A2(n2374), .ZN(n2467) );
  NAND2_X1 U3139 ( .A1(n2468), .A2(n2467), .ZN(n2469) );
  XNOR2_X1 U3140 ( .A(n2469), .B(n2746), .ZN(n2470) );
  AOI22_X1 U3141 ( .A1(n3707), .A2(n2737), .B1(n3218), .B2(n2051), .ZN(n2471)
         );
  XNOR2_X1 U3142 ( .A(n2470), .B(n2471), .ZN(n3169) );
  INV_X1 U3143 ( .A(n2470), .ZN(n2472) );
  NAND2_X1 U3144 ( .A1(n2472), .A2(n2471), .ZN(n2473) );
  NAND2_X1 U3145 ( .A1(n2474), .A2(n2473), .ZN(n3239) );
  INV_X1 U3146 ( .A(n3239), .ZN(n2487) );
  OR2_X1 U3147 ( .A1(n3533), .A2(n4287), .ZN(n2481) );
  NAND2_X1 U31480 ( .A1(n2056), .A2(REG0_REG_10__SCAN_IN), .ZN(n2480) );
  AND2_X1 U31490 ( .A1(n2476), .A2(n2475), .ZN(n2477) );
  NOR2_X1 U3150 ( .A1(n2493), .A2(n2477), .ZN(n3244) );
  NAND2_X1 U3151 ( .A1(n2668), .A2(n3244), .ZN(n2479) );
  NAND2_X1 U3152 ( .A1(n2343), .A2(REG2_REG_10__SCAN_IN), .ZN(n2478) );
  NAND4_X1 U3153 ( .A1(n2481), .A2(n2480), .A3(n2479), .A4(n2478), .ZN(n3706)
         );
  NAND2_X1 U3154 ( .A1(n3706), .A2(n2051), .ZN(n2484) );
  OR2_X1 U3155 ( .A1(n2501), .A2(n2820), .ZN(n2482) );
  XNOR2_X1 U3156 ( .A(n2482), .B(IR_REG_10__SCAN_IN), .ZN(n3779) );
  MUX2_X1 U3157 ( .A(n3779), .B(DATAI_10_), .S(n2433), .Z(n3265) );
  NAND2_X1 U3158 ( .A1(n3265), .A2(n2374), .ZN(n2483) );
  NAND2_X1 U3159 ( .A1(n2484), .A2(n2483), .ZN(n2485) );
  XNOR2_X1 U3160 ( .A(n2485), .B(n2734), .ZN(n2488) );
  AOI22_X1 U3161 ( .A1(n3706), .A2(n2737), .B1(n2051), .B2(n3265), .ZN(n2489)
         );
  XNOR2_X1 U3162 ( .A(n2488), .B(n2489), .ZN(n3241) );
  INV_X1 U3163 ( .A(n2488), .ZN(n2491) );
  INV_X1 U3164 ( .A(n2489), .ZN(n2490) );
  NAND2_X1 U3165 ( .A1(n2491), .A2(n2490), .ZN(n2492) );
  NAND2_X1 U3166 ( .A1(n2055), .A2(REG0_REG_11__SCAN_IN), .ZN(n2499) );
  OR2_X1 U3167 ( .A1(n2493), .A2(REG3_REG_11__SCAN_IN), .ZN(n2494) );
  NAND2_X1 U3168 ( .A1(n2493), .A2(REG3_REG_11__SCAN_IN), .ZN(n2508) );
  AND2_X1 U3169 ( .A1(n2494), .A2(n2508), .ZN(n3279) );
  NAND2_X1 U3170 ( .A1(n2668), .A2(n3279), .ZN(n2498) );
  NAND2_X1 U3171 ( .A1(n3531), .A2(REG2_REG_11__SCAN_IN), .ZN(n2497) );
  INV_X1 U3172 ( .A(REG1_REG_11__SCAN_IN), .ZN(n2495) );
  OR2_X1 U3173 ( .A1(n3533), .A2(n2495), .ZN(n2496) );
  INV_X1 U3174 ( .A(IR_REG_10__SCAN_IN), .ZN(n2500) );
  NAND2_X1 U3175 ( .A1(n2501), .A2(n2500), .ZN(n2502) );
  NAND2_X1 U3176 ( .A1(n2502), .A2(IR_REG_31__SCAN_IN), .ZN(n2504) );
  INV_X1 U3177 ( .A(IR_REG_11__SCAN_IN), .ZN(n2503) );
  NAND2_X1 U3178 ( .A1(n2504), .A2(n2503), .ZN(n2515) );
  OR2_X1 U3179 ( .A1(n2504), .A2(n2503), .ZN(n2505) );
  MUX2_X1 U3180 ( .A(n3783), .B(DATAI_11_), .S(n2433), .Z(n3284) );
  OAI22_X1 U3181 ( .A1(n3263), .A2(n2748), .B1(n2661), .B2(n3277), .ZN(n3230)
         );
  OAI22_X1 U3182 ( .A1(n3263), .A2(n2661), .B1(n2745), .B2(n3277), .ZN(n2506)
         );
  XNOR2_X1 U3183 ( .A(n2506), .B(n2746), .ZN(n3229) );
  NAND2_X1 U3184 ( .A1(n2054), .A2(REG0_REG_12__SCAN_IN), .ZN(n2514) );
  INV_X1 U3185 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2507) );
  NAND2_X1 U3186 ( .A1(n2508), .A2(n2507), .ZN(n2509) );
  AND2_X1 U3187 ( .A1(n2523), .A2(n2509), .ZN(n3315) );
  NAND2_X1 U3188 ( .A1(n2668), .A2(n3315), .ZN(n2513) );
  NAND2_X1 U3189 ( .A1(n2343), .A2(REG2_REG_12__SCAN_IN), .ZN(n2512) );
  INV_X1 U3190 ( .A(REG1_REG_12__SCAN_IN), .ZN(n2510) );
  OR2_X1 U3191 ( .A1(n3533), .A2(n2510), .ZN(n2511) );
  NAND2_X1 U3192 ( .A1(n2515), .A2(IR_REG_31__SCAN_IN), .ZN(n2516) );
  XNOR2_X1 U3193 ( .A(n2516), .B(IR_REG_12__SCAN_IN), .ZN(n4412) );
  INV_X1 U3194 ( .A(DATAI_12_), .ZN(n2517) );
  OAI22_X1 U3195 ( .A1(n4105), .A2(n2661), .B1(n2745), .B2(n3309), .ZN(n2518)
         );
  XNOR2_X1 U3196 ( .A(n2518), .B(n2746), .ZN(n2519) );
  OAI22_X1 U3197 ( .A1(n4105), .A2(n2748), .B1(n2661), .B2(n3309), .ZN(n2520)
         );
  AND2_X1 U3198 ( .A1(n2519), .A2(n2520), .ZN(n3256) );
  INV_X1 U3199 ( .A(n2519), .ZN(n2522) );
  INV_X1 U3200 ( .A(n2520), .ZN(n2521) );
  NAND2_X1 U3201 ( .A1(n2522), .A2(n2521), .ZN(n3255) );
  NAND2_X1 U3202 ( .A1(n2053), .A2(REG0_REG_13__SCAN_IN), .ZN(n2528) );
  AND2_X1 U3203 ( .A1(n2523), .A2(n3324), .ZN(n2524) );
  NOR2_X1 U3204 ( .A1(n2538), .A2(n2524), .ZN(n4114) );
  NAND2_X1 U3205 ( .A1(n2668), .A2(n4114), .ZN(n2527) );
  NAND2_X1 U3206 ( .A1(n3531), .A2(REG2_REG_13__SCAN_IN), .ZN(n2526) );
  INV_X1 U3207 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4201) );
  OR2_X1 U3208 ( .A1(n3533), .A2(n4201), .ZN(n2525) );
  OR2_X1 U3209 ( .A1(n2529), .A2(n2820), .ZN(n2530) );
  XNOR2_X1 U32100 ( .A(n2530), .B(IR_REG_13__SCAN_IN), .ZN(n3786) );
  INV_X1 U32110 ( .A(DATAI_13_), .ZN(n4410) );
  MUX2_X1 U32120 ( .A(n4411), .B(n4410), .S(n2433), .Z(n4112) );
  OAI22_X1 U32130 ( .A1(n3384), .A2(n2661), .B1(n2745), .B2(n4112), .ZN(n2531)
         );
  XNOR2_X1 U32140 ( .A(n2531), .B(n2734), .ZN(n3321) );
  NAND2_X1 U32150 ( .A1(n3320), .A2(n3321), .ZN(n2532) );
  OAI22_X1 U32160 ( .A1(n3384), .A2(n2748), .B1(n2661), .B2(n4112), .ZN(n3322)
         );
  NAND2_X1 U32170 ( .A1(n2532), .A2(n3322), .ZN(n2537) );
  OR2_X1 U32180 ( .A1(n3254), .A2(n3256), .ZN(n2535) );
  INV_X1 U32190 ( .A(n3321), .ZN(n2533) );
  AND2_X1 U32200 ( .A1(n2533), .A2(n3255), .ZN(n2534) );
  NAND2_X1 U32210 ( .A1(n2535), .A2(n2534), .ZN(n2536) );
  NAND2_X1 U32220 ( .A1(n2537), .A2(n2536), .ZN(n3380) );
  NAND2_X1 U32230 ( .A1(n2054), .A2(REG0_REG_14__SCAN_IN), .ZN(n2543) );
  NAND2_X1 U32240 ( .A1(n2538), .A2(REG3_REG_14__SCAN_IN), .ZN(n2551) );
  OR2_X1 U32250 ( .A1(n2538), .A2(REG3_REG_14__SCAN_IN), .ZN(n2539) );
  AND2_X1 U32260 ( .A1(n2551), .A2(n2539), .ZN(n3388) );
  NAND2_X1 U32270 ( .A1(n2668), .A2(n3388), .ZN(n2542) );
  NAND2_X1 U32280 ( .A1(n3531), .A2(REG2_REG_14__SCAN_IN), .ZN(n2541) );
  INV_X1 U32290 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4327) );
  OR2_X1 U32300 ( .A1(n3533), .A2(n4327), .ZN(n2540) );
  OR2_X1 U32310 ( .A1(n2544), .A2(n2820), .ZN(n2545) );
  XNOR2_X1 U32320 ( .A(n2545), .B(IR_REG_14__SCAN_IN), .ZN(n4334) );
  MUX2_X1 U32330 ( .A(n4334), .B(DATAI_14_), .S(n2433), .Z(n3331) );
  INV_X1 U32340 ( .A(n3331), .ZN(n3385) );
  OAI22_X1 U32350 ( .A1(n4083), .A2(n2661), .B1(n3385), .B2(n2745), .ZN(n2546)
         );
  XNOR2_X1 U32360 ( .A(n2546), .B(n2746), .ZN(n2547) );
  OAI22_X1 U32370 ( .A1(n4083), .A2(n2748), .B1(n3385), .B2(n2661), .ZN(n2548)
         );
  AND2_X1 U32380 ( .A1(n2547), .A2(n2548), .ZN(n3382) );
  INV_X1 U32390 ( .A(n2547), .ZN(n2550) );
  INV_X1 U32400 ( .A(n2548), .ZN(n2549) );
  NAND2_X1 U32410 ( .A1(n2550), .A2(n2549), .ZN(n3381) );
  NAND2_X1 U32420 ( .A1(n2056), .A2(REG0_REG_15__SCAN_IN), .ZN(n2556) );
  INV_X1 U32430 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3516) );
  NAND2_X1 U32440 ( .A1(n2551), .A2(n3516), .ZN(n2552) );
  AND2_X1 U32450 ( .A1(n2562), .A2(n2552), .ZN(n4086) );
  NAND2_X1 U32460 ( .A1(n2668), .A2(n4086), .ZN(n2555) );
  NAND2_X1 U32470 ( .A1(n3531), .A2(REG2_REG_15__SCAN_IN), .ZN(n2554) );
  INV_X1 U32480 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3788) );
  OR2_X1 U32490 ( .A1(n3533), .A2(n3788), .ZN(n2553) );
  NAND2_X1 U32500 ( .A1(n2544), .A2(n2557), .ZN(n2558) );
  NAND2_X1 U32510 ( .A1(n2558), .A2(IR_REG_31__SCAN_IN), .ZN(n2569) );
  XNOR2_X1 U32520 ( .A(n2569), .B(IR_REG_15__SCAN_IN), .ZN(n3789) );
  MUX2_X1 U32530 ( .A(n3789), .B(DATAI_15_), .S(n2433), .Z(n4084) );
  OAI22_X1 U32540 ( .A1(n3452), .A2(n2661), .B1(n2745), .B2(n3354), .ZN(n2559)
         );
  XNOR2_X1 U32550 ( .A(n2559), .B(n2734), .ZN(n2579) );
  INV_X1 U32560 ( .A(n2579), .ZN(n2560) );
  NAND2_X1 U32570 ( .A1(n2055), .A2(REG0_REG_16__SCAN_IN), .ZN(n2567) );
  INV_X1 U32580 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2561) );
  AND2_X1 U32590 ( .A1(n2562), .A2(n2561), .ZN(n2563) );
  NOR2_X1 U32600 ( .A1(n2582), .A2(n2563), .ZN(n4056) );
  NAND2_X1 U32610 ( .A1(n2668), .A2(n4056), .ZN(n2566) );
  NAND2_X1 U32620 ( .A1(n3531), .A2(REG2_REG_16__SCAN_IN), .ZN(n2565) );
  INV_X1 U32630 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4353) );
  OR2_X1 U32640 ( .A1(n3533), .A2(n4353), .ZN(n2564) );
  NAND2_X1 U32650 ( .A1(n2569), .A2(n2568), .ZN(n2570) );
  NAND2_X1 U32660 ( .A1(n2570), .A2(IR_REG_31__SCAN_IN), .ZN(n2571) );
  XNOR2_X1 U32670 ( .A(n2571), .B(n4502), .ZN(n4405) );
  INV_X1 U32680 ( .A(n4405), .ZN(n2572) );
  MUX2_X1 U32690 ( .A(n2572), .B(DATAI_16_), .S(n2433), .Z(n4055) );
  OAI22_X1 U32700 ( .A1(n3517), .A2(n2661), .B1(n4060), .B2(n2745), .ZN(n2573)
         );
  XNOR2_X1 U32710 ( .A(n2573), .B(n2734), .ZN(n2575) );
  OAI22_X1 U32720 ( .A1(n3517), .A2(n2748), .B1(n4060), .B2(n2661), .ZN(n2576)
         );
  INV_X1 U32730 ( .A(n2576), .ZN(n2574) );
  NAND2_X1 U32740 ( .A1(n2575), .A2(n2574), .ZN(n2581) );
  INV_X1 U32750 ( .A(n2575), .ZN(n2577) );
  NAND2_X1 U32760 ( .A1(n2577), .A2(n2576), .ZN(n2578) );
  AND2_X1 U32770 ( .A1(n2581), .A2(n2578), .ZN(n3451) );
  OAI22_X1 U32780 ( .A1(n3452), .A2(n2748), .B1(n2661), .B2(n3354), .ZN(n3515)
         );
  NAND2_X1 U32790 ( .A1(n2055), .A2(REG0_REG_17__SCAN_IN), .ZN(n2587) );
  NOR2_X1 U32800 ( .A1(n2582), .A2(REG3_REG_17__SCAN_IN), .ZN(n2583) );
  NOR2_X1 U32810 ( .A1(n2598), .A2(n2583), .ZN(n4046) );
  NAND2_X1 U32820 ( .A1(n2668), .A2(n4046), .ZN(n2586) );
  NAND2_X1 U32830 ( .A1(n3531), .A2(REG2_REG_17__SCAN_IN), .ZN(n2585) );
  INV_X1 U32840 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4648) );
  OR2_X1 U32850 ( .A1(n3533), .A2(n4648), .ZN(n2584) );
  NAND2_X1 U32860 ( .A1(n2588), .A2(IR_REG_31__SCAN_IN), .ZN(n2589) );
  MUX2_X1 U32870 ( .A(IR_REG_31__SCAN_IN), .B(n2589), .S(IR_REG_17__SCAN_IN), 
        .Z(n2591) );
  INV_X1 U32880 ( .A(n2590), .ZN(n2604) );
  NAND2_X1 U32890 ( .A1(n2591), .A2(n2604), .ZN(n3776) );
  INV_X1 U32900 ( .A(DATAI_17_), .ZN(n4512) );
  MUX2_X1 U32910 ( .A(n3776), .B(n4512), .S(n2433), .Z(n4045) );
  OAI22_X1 U32920 ( .A1(n4061), .A2(n2661), .B1(n2745), .B2(n4045), .ZN(n2592)
         );
  XNOR2_X1 U32930 ( .A(n2592), .B(n2746), .ZN(n2593) );
  OAI22_X1 U32940 ( .A1(n4061), .A2(n2748), .B1(n2661), .B2(n4045), .ZN(n2594)
         );
  NAND2_X1 U32950 ( .A1(n2593), .A2(n2594), .ZN(n3459) );
  INV_X1 U32960 ( .A(n2593), .ZN(n2596) );
  INV_X1 U32970 ( .A(n2594), .ZN(n2595) );
  NAND2_X1 U32980 ( .A1(n2596), .A2(n2595), .ZN(n3458) );
  NAND2_X1 U32990 ( .A1(n2597), .A2(n3458), .ZN(n3400) );
  NAND2_X1 U33000 ( .A1(n2053), .A2(REG0_REG_18__SCAN_IN), .ZN(n2603) );
  OR2_X1 U33010 ( .A1(n2598), .A2(REG3_REG_18__SCAN_IN), .ZN(n2599) );
  AND2_X1 U33020 ( .A1(n2609), .A2(n2599), .ZN(n4028) );
  NAND2_X1 U33030 ( .A1(n2668), .A2(n4028), .ZN(n2602) );
  NAND2_X1 U33040 ( .A1(n3531), .A2(REG2_REG_18__SCAN_IN), .ZN(n2601) );
  INV_X1 U33050 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3798) );
  OR2_X1 U33060 ( .A1(n3533), .A2(n3798), .ZN(n2600) );
  NAND2_X1 U33070 ( .A1(n2604), .A2(IR_REG_31__SCAN_IN), .ZN(n2605) );
  MUX2_X1 U33080 ( .A(IR_REG_31__SCAN_IN), .B(n2605), .S(IR_REG_18__SCAN_IN), 
        .Z(n2607) );
  AND2_X1 U33090 ( .A1(n2607), .A2(n2606), .ZN(n4402) );
  MUX2_X1 U33100 ( .A(n4402), .B(DATAI_18_), .S(n2433), .Z(n4025) );
  OAI22_X1 U33110 ( .A1(n4038), .A2(n2748), .B1(n2661), .B2(n3335), .ZN(n3496)
         );
  OAI22_X1 U33120 ( .A1(n4038), .A2(n2661), .B1(n2745), .B2(n3335), .ZN(n2608)
         );
  XNOR2_X1 U33130 ( .A(n2608), .B(n2746), .ZN(n3497) );
  INV_X1 U33140 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4179) );
  OR2_X1 U33150 ( .A1(n3533), .A2(n4179), .ZN(n2614) );
  NAND2_X1 U33160 ( .A1(n2054), .A2(REG0_REG_19__SCAN_IN), .ZN(n2613) );
  INV_X1 U33170 ( .A(REG3_REG_19__SCAN_IN), .ZN(n3409) );
  NAND2_X1 U33180 ( .A1(n2609), .A2(n3409), .ZN(n2610) );
  AND2_X1 U33190 ( .A1(n2629), .A2(n2610), .ZN(n4009) );
  NAND2_X1 U33200 ( .A1(n2668), .A2(n4009), .ZN(n2612) );
  NAND2_X1 U33210 ( .A1(n3531), .A2(REG2_REG_19__SCAN_IN), .ZN(n2611) );
  NAND2_X1 U33220 ( .A1(n4021), .A2(n2051), .ZN(n2616) );
  MUX2_X1 U33230 ( .A(n4269), .B(DATAI_19_), .S(n2433), .Z(n3411) );
  NAND2_X1 U33240 ( .A1(n3411), .A2(n2374), .ZN(n2615) );
  NAND2_X1 U33250 ( .A1(n2616), .A2(n2615), .ZN(n2617) );
  XNOR2_X1 U33260 ( .A(n2617), .B(n2746), .ZN(n2622) );
  NAND2_X1 U33270 ( .A1(n4021), .A2(n2737), .ZN(n2619) );
  NAND2_X1 U33280 ( .A1(n3411), .A2(n2051), .ZN(n2618) );
  NAND2_X1 U33290 ( .A1(n2619), .A2(n2618), .ZN(n2623) );
  AOI21_X1 U33300 ( .B1(n3496), .B2(n3497), .A(n2621), .ZN(n2620) );
  NAND2_X1 U33310 ( .A1(n3400), .A2(n2620), .ZN(n2628) );
  INV_X1 U33320 ( .A(n3497), .ZN(n3401) );
  INV_X1 U33330 ( .A(n3496), .ZN(n3402) );
  INV_X1 U33340 ( .A(n2621), .ZN(n3406) );
  NAND3_X1 U33350 ( .A1(n3401), .A2(n3402), .A3(n3406), .ZN(n2626) );
  INV_X1 U33360 ( .A(n2622), .ZN(n2625) );
  INV_X1 U33370 ( .A(n2623), .ZN(n2624) );
  NAND2_X1 U33380 ( .A1(n2625), .A2(n2624), .ZN(n3405) );
  NAND2_X1 U33390 ( .A1(n2628), .A2(n2627), .ZN(n3425) );
  NAND2_X1 U33400 ( .A1(n2056), .A2(REG0_REG_20__SCAN_IN), .ZN(n2634) );
  INV_X1 U33410 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3481) );
  NAND2_X1 U33420 ( .A1(n2629), .A2(n3481), .ZN(n2630) );
  NAND2_X1 U33430 ( .A1(n2640), .A2(n2630), .ZN(n3987) );
  INV_X1 U33440 ( .A(n3987), .ZN(n3484) );
  NAND2_X1 U33450 ( .A1(n2668), .A2(n3484), .ZN(n2633) );
  NAND2_X1 U33460 ( .A1(n3531), .A2(REG2_REG_20__SCAN_IN), .ZN(n2632) );
  INV_X1 U33470 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4174) );
  OR2_X1 U33480 ( .A1(n3533), .A2(n4174), .ZN(n2631) );
  OAI22_X1 U33490 ( .A1(n3999), .A2(n2661), .B1(n2745), .B2(n3974), .ZN(n2635)
         );
  XNOR2_X1 U33500 ( .A(n2635), .B(n2746), .ZN(n2636) );
  OAI22_X1 U33510 ( .A1(n3999), .A2(n2748), .B1(n2661), .B2(n3974), .ZN(n2637)
         );
  NAND2_X1 U33520 ( .A1(n2636), .A2(n2637), .ZN(n3477) );
  NAND2_X1 U3353 ( .A1(n3425), .A2(n3477), .ZN(n3476) );
  INV_X1 U33540 ( .A(n2636), .ZN(n2639) );
  INV_X1 U3355 ( .A(n2637), .ZN(n2638) );
  NAND2_X1 U3356 ( .A1(n2639), .A2(n2638), .ZN(n3479) );
  INV_X1 U3357 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4169) );
  OR2_X1 U3358 ( .A1(n3533), .A2(n4169), .ZN(n2645) );
  NAND2_X1 U3359 ( .A1(n2055), .A2(REG0_REG_21__SCAN_IN), .ZN(n2644) );
  INV_X1 U3360 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3432) );
  AND2_X1 U3361 ( .A1(n2640), .A2(n3432), .ZN(n2641) );
  NOR2_X1 U3362 ( .A1(n2655), .A2(n2641), .ZN(n3968) );
  NAND2_X1 U3363 ( .A1(n2668), .A2(n3968), .ZN(n2643) );
  NAND2_X1 U3364 ( .A1(n3531), .A2(REG2_REG_21__SCAN_IN), .ZN(n2642) );
  NAND2_X1 U3365 ( .A1(n3942), .A2(n2051), .ZN(n2647) );
  NAND2_X1 U3366 ( .A1(n2374), .A2(n3339), .ZN(n2646) );
  NAND2_X1 U3367 ( .A1(n2647), .A2(n2646), .ZN(n2648) );
  XNOR2_X1 U3368 ( .A(n2648), .B(n2734), .ZN(n2650) );
  NOR2_X1 U3369 ( .A1(n2661), .A2(n3966), .ZN(n2649) );
  AOI21_X1 U3370 ( .B1(n3942), .B2(n2737), .A(n2649), .ZN(n2651) );
  INV_X1 U3371 ( .A(n2650), .ZN(n2653) );
  INV_X1 U3372 ( .A(n2651), .ZN(n2652) );
  NAND2_X1 U3373 ( .A1(n2653), .A2(n2652), .ZN(n3424) );
  INV_X1 U3374 ( .A(REG1_REG_22__SCAN_IN), .ZN(n2654) );
  OR2_X1 U3375 ( .A1(n3533), .A2(n2654), .ZN(n2660) );
  NAND2_X1 U3376 ( .A1(n2053), .A2(REG0_REG_22__SCAN_IN), .ZN(n2659) );
  OR2_X1 U3377 ( .A1(n2655), .A2(REG3_REG_22__SCAN_IN), .ZN(n2656) );
  NAND2_X1 U3378 ( .A1(n2655), .A2(REG3_REG_22__SCAN_IN), .ZN(n2666) );
  AND2_X1 U3379 ( .A1(n2656), .A2(n2666), .ZN(n3948) );
  NAND2_X1 U3380 ( .A1(n2668), .A2(n3948), .ZN(n2658) );
  NAND2_X1 U3381 ( .A1(n3531), .A2(REG2_REG_22__SCAN_IN), .ZN(n2657) );
  NAND2_X1 U3382 ( .A1(n3960), .A2(n2051), .ZN(n2663) );
  NAND2_X1 U3383 ( .A1(n2374), .A2(n3951), .ZN(n2662) );
  NAND2_X1 U3384 ( .A1(n2663), .A2(n2662), .ZN(n2664) );
  XNOR2_X1 U3385 ( .A(n2664), .B(n2734), .ZN(n2675) );
  NOR2_X1 U3386 ( .A1(n2661), .A2(n3491), .ZN(n2665) );
  AOI21_X1 U3387 ( .B1(n3960), .B2(n2737), .A(n2665), .ZN(n2674) );
  XNOR2_X1 U3388 ( .A(n2675), .B(n2674), .ZN(n3489) );
  INV_X1 U3389 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4633) );
  NAND2_X1 U3390 ( .A1(n2666), .A2(n4633), .ZN(n2667) );
  AND2_X1 U3391 ( .A1(n2680), .A2(n2667), .ZN(n3931) );
  NAND2_X1 U3392 ( .A1(n3931), .A2(n2668), .ZN(n2672) );
  INV_X1 U3393 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4160) );
  OR2_X1 U3394 ( .A1(n3533), .A2(n4160), .ZN(n2671) );
  NAND2_X1 U3395 ( .A1(n2054), .A2(REG0_REG_23__SCAN_IN), .ZN(n2670) );
  NAND2_X1 U3396 ( .A1(n3531), .A2(REG2_REG_23__SCAN_IN), .ZN(n2669) );
  OAI22_X1 U3397 ( .A1(n3945), .A2(n2661), .B1(n2745), .B2(n3928), .ZN(n2673)
         );
  XNOR2_X1 U3398 ( .A(n2673), .B(n2734), .ZN(n2677) );
  OAI22_X1 U3399 ( .A1(n3945), .A2(n2748), .B1(n2661), .B2(n3928), .ZN(n2678)
         );
  XNOR2_X1 U3400 ( .A(n2677), .B(n2678), .ZN(n3393) );
  NAND2_X1 U3401 ( .A1(n2675), .A2(n2674), .ZN(n3394) );
  INV_X1 U3402 ( .A(n2677), .ZN(n2679) );
  NAND2_X1 U3403 ( .A1(n2679), .A2(n2678), .ZN(n2690) );
  INV_X1 U3404 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3471) );
  AND2_X1 U3405 ( .A1(n2680), .A2(n3471), .ZN(n2681) );
  OR2_X1 U3406 ( .A1(n2681), .A2(n2695), .ZN(n3470) );
  AOI22_X1 U3407 ( .A1(n2682), .A2(REG1_REG_24__SCAN_IN), .B1(n2054), .B2(
        REG0_REG_24__SCAN_IN), .ZN(n2684) );
  NAND2_X1 U3408 ( .A1(n2343), .A2(REG2_REG_24__SCAN_IN), .ZN(n2683) );
  NOR2_X1 U3409 ( .A1(n2661), .A2(n3903), .ZN(n2685) );
  AOI21_X1 U3410 ( .B1(n3700), .B2(n2737), .A(n2685), .ZN(n2691) );
  AND2_X1 U3411 ( .A1(n2690), .A2(n2691), .ZN(n2686) );
  NAND2_X1 U3412 ( .A1(n3700), .A2(n2051), .ZN(n2688) );
  NAND2_X1 U3413 ( .A1(n2374), .A2(n3908), .ZN(n2687) );
  NAND2_X1 U3414 ( .A1(n2688), .A2(n2687), .ZN(n2689) );
  XNOR2_X1 U3415 ( .A(n2689), .B(n2746), .ZN(n3469) );
  NAND2_X1 U3416 ( .A1(n3467), .A2(n3469), .ZN(n2694) );
  INV_X1 U3417 ( .A(n2691), .ZN(n2692) );
  NAND2_X1 U3418 ( .A1(n2693), .A2(n2692), .ZN(n3466) );
  NAND2_X1 U3419 ( .A1(n2694), .A2(n3466), .ZN(n3439) );
  NOR2_X1 U3420 ( .A1(n2695), .A2(REG3_REG_25__SCAN_IN), .ZN(n2696) );
  OR2_X1 U3421 ( .A1(n2708), .A2(n2696), .ZN(n3441) );
  AOI22_X1 U3422 ( .A1(n3531), .A2(REG2_REG_25__SCAN_IN), .B1(n2056), .B2(
        REG0_REG_25__SCAN_IN), .ZN(n2698) );
  INV_X1 U3423 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4153) );
  OR2_X1 U3424 ( .A1(n3533), .A2(n4153), .ZN(n2697) );
  NAND2_X1 U3425 ( .A1(n3905), .A2(n2051), .ZN(n2700) );
  NAND2_X1 U3426 ( .A1(n2374), .A2(n3342), .ZN(n2699) );
  NAND2_X1 U3427 ( .A1(n2700), .A2(n2699), .ZN(n2701) );
  XNOR2_X1 U3428 ( .A(n2701), .B(n2734), .ZN(n2703) );
  NOR2_X1 U3429 ( .A1(n2661), .A2(n3891), .ZN(n2702) );
  AOI21_X1 U3430 ( .B1(n3905), .B2(n2737), .A(n2702), .ZN(n2704) );
  NAND2_X1 U3431 ( .A1(n2703), .A2(n2704), .ZN(n3437) );
  INV_X1 U3432 ( .A(n2703), .ZN(n2706) );
  INV_X1 U3433 ( .A(n2704), .ZN(n2705) );
  NAND2_X1 U3434 ( .A1(n2706), .A2(n2705), .ZN(n3438) );
  NOR2_X1 U3435 ( .A1(n2708), .A2(REG3_REG_26__SCAN_IN), .ZN(n2709) );
  INV_X1 U3436 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4149) );
  NAND2_X1 U3437 ( .A1(n3531), .A2(REG2_REG_26__SCAN_IN), .ZN(n2711) );
  NAND2_X1 U3438 ( .A1(n2053), .A2(REG0_REG_26__SCAN_IN), .ZN(n2710) );
  OAI211_X1 U3439 ( .C1(n3533), .C2(n4149), .A(n2711), .B(n2710), .ZN(n2712)
         );
  INV_X1 U3440 ( .A(n2712), .ZN(n2713) );
  NAND2_X1 U3441 ( .A1(n3887), .A2(n2051), .ZN(n2716) );
  NAND2_X1 U3442 ( .A1(n2433), .A2(DATAI_26_), .ZN(n3870) );
  NAND2_X1 U3443 ( .A1(n2374), .A2(n3864), .ZN(n2715) );
  NAND2_X1 U3444 ( .A1(n2716), .A2(n2715), .ZN(n2717) );
  XNOR2_X1 U3445 ( .A(n2717), .B(n2746), .ZN(n2720) );
  NAND2_X1 U3446 ( .A1(n3887), .A2(n2737), .ZN(n2719) );
  NAND2_X1 U3447 ( .A1(n2051), .A2(n3864), .ZN(n2718) );
  NAND2_X1 U3448 ( .A1(n2719), .A2(n2718), .ZN(n2721) );
  AND2_X1 U3449 ( .A1(n2720), .A2(n2721), .ZN(n3505) );
  INV_X1 U3450 ( .A(n2720), .ZN(n2723) );
  INV_X1 U3451 ( .A(n2721), .ZN(n2722) );
  NAND2_X1 U3452 ( .A1(n2723), .A2(n2722), .ZN(n3504) );
  NAND2_X1 U3453 ( .A1(n2724), .A2(REG3_REG_27__SCAN_IN), .ZN(n2738) );
  OR2_X1 U3454 ( .A1(n2724), .A2(REG3_REG_27__SCAN_IN), .ZN(n2725) );
  NAND2_X1 U3455 ( .A1(n3852), .A2(n2668), .ZN(n2731) );
  INV_X1 U3456 ( .A(REG1_REG_27__SCAN_IN), .ZN(n2728) );
  NAND2_X1 U3457 ( .A1(n3531), .A2(REG2_REG_27__SCAN_IN), .ZN(n2727) );
  NAND2_X1 U34580 ( .A1(n2056), .A2(REG0_REG_27__SCAN_IN), .ZN(n2726) );
  OAI211_X1 U34590 ( .C1(n3533), .C2(n2728), .A(n2727), .B(n2726), .ZN(n2729)
         );
  INV_X1 U3460 ( .A(n2729), .ZN(n2730) );
  NAND2_X1 U3461 ( .A1(n3699), .A2(n2051), .ZN(n2733) );
  NAND2_X1 U3462 ( .A1(n2374), .A2(n3613), .ZN(n2732) );
  NAND2_X1 U3463 ( .A1(n2733), .A2(n2732), .ZN(n2735) );
  XNOR2_X1 U3464 ( .A(n2735), .B(n2734), .ZN(n2751) );
  AND2_X1 U3465 ( .A1(n2051), .A2(n3613), .ZN(n2736) );
  AOI21_X1 U3466 ( .B1(n3699), .B2(n2737), .A(n2736), .ZN(n2752) );
  XNOR2_X1 U34670 ( .A(n2751), .B(n2752), .ZN(n3373) );
  INV_X1 U3468 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2793) );
  NAND2_X1 U34690 ( .A1(n2738), .A2(n2793), .ZN(n2739) );
  NAND2_X1 U3470 ( .A1(n3833), .A2(n2668), .ZN(n2744) );
  INV_X1 U34710 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4546) );
  NAND2_X1 U3472 ( .A1(n2055), .A2(REG0_REG_28__SCAN_IN), .ZN(n2741) );
  NAND2_X1 U34730 ( .A1(n3531), .A2(REG2_REG_28__SCAN_IN), .ZN(n2740) );
  OAI211_X1 U3474 ( .C1(n4546), .C2(n3533), .A(n2741), .B(n2740), .ZN(n2742)
         );
  INV_X1 U34750 ( .A(n2742), .ZN(n2743) );
  INV_X1 U3476 ( .A(n3351), .ZN(n3821) );
  OAI22_X1 U34770 ( .A1(n3822), .A2(n2661), .B1(n3821), .B2(n2745), .ZN(n2747)
         );
  XNOR2_X1 U3478 ( .A(n2747), .B(n2746), .ZN(n2750) );
  OAI22_X1 U34790 ( .A1(n3822), .A2(n2748), .B1(n3821), .B2(n2661), .ZN(n2749)
         );
  XNOR2_X1 U3480 ( .A(n2750), .B(n2749), .ZN(n2781) );
  INV_X1 U34810 ( .A(n2781), .ZN(n2776) );
  INV_X1 U3482 ( .A(n2751), .ZN(n2754) );
  INV_X1 U34830 ( .A(n2752), .ZN(n2753) );
  NAND2_X1 U3484 ( .A1(n2754), .A2(n2753), .ZN(n2779) );
  NAND2_X1 U34850 ( .A1(n2815), .A2(B_REG_SCAN_IN), .ZN(n2755) );
  INV_X1 U3486 ( .A(n2769), .ZN(n4265) );
  MUX2_X1 U34870 ( .A(n2755), .B(B_REG_SCAN_IN), .S(n4265), .Z(n2757) );
  NOR4_X1 U3488 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_15__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2761) );
  NOR4_X1 U34890 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_7__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2760) );
  NOR4_X1 U3490 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2759) );
  NOR4_X1 U34910 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_22__SCAN_IN), .ZN(n2758) );
  AND4_X1 U3492 ( .A1(n2761), .A2(n2760), .A3(n2759), .A4(n2758), .ZN(n2767)
         );
  NOR2_X1 U34930 ( .A1(D_REG_8__SCAN_IN), .A2(D_REG_27__SCAN_IN), .ZN(n2765)
         );
  NOR4_X1 U3494 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2764) );
  NOR4_X1 U34950 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_2__SCAN_IN), .A3(
        D_REG_3__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n2763) );
  NOR4_X1 U3496 ( .A1(D_REG_9__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_26__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2762) );
  AND4_X1 U34970 ( .A1(n2765), .A2(n2764), .A3(n2763), .A4(n2762), .ZN(n2766)
         );
  NAND2_X1 U3498 ( .A1(n2767), .A2(n2766), .ZN(n3027) );
  INV_X1 U34990 ( .A(D_REG_1__SCAN_IN), .ZN(n2824) );
  NOR2_X1 U3500 ( .A1(n3027), .A2(n2824), .ZN(n2768) );
  INV_X1 U35010 ( .A(n2756), .ZN(n2770) );
  NAND2_X1 U3502 ( .A1(n2770), .A2(n2815), .ZN(n3025) );
  OAI21_X1 U35030 ( .B1(n3026), .B2(n2768), .A(n3025), .ZN(n2968) );
  INV_X1 U3504 ( .A(n2968), .ZN(n2771) );
  INV_X1 U35050 ( .A(D_REG_0__SCAN_IN), .ZN(n4501) );
  XNOR2_X1 U35060 ( .A(n2773), .B(n2772), .ZN(n2831) );
  INV_X1 U35070 ( .A(n4269), .ZN(n3807) );
  INV_X1 U35080 ( .A(n3579), .ZN(n4267) );
  NAND2_X1 U35090 ( .A1(n4266), .A2(n4267), .ZN(n2830) );
  OAI211_X1 U35100 ( .C1(n4383), .C2(n3807), .A(n4059), .B(n2830), .ZN(n2783)
         );
  NOR2_X1 U35110 ( .A1(n3024), .A2(n2783), .ZN(n2774) );
  AND2_X1 U35120 ( .A1(n2779), .A2(n3428), .ZN(n2775) );
  NAND2_X1 U35130 ( .A1(n2777), .A2(n2276), .ZN(n2810) );
  NAND3_X1 U35140 ( .A1(n2778), .A2(n3428), .A3(n2781), .ZN(n2809) );
  INV_X1 U35150 ( .A(n2779), .ZN(n2780) );
  NAND3_X1 U35160 ( .A1(n2781), .A2(n3428), .A3(n2780), .ZN(n2808) );
  NAND2_X1 U35170 ( .A1(n2783), .A2(n4059), .ZN(n2784) );
  NAND2_X1 U35180 ( .A1(n2800), .A2(n2784), .ZN(n2786) );
  AND2_X1 U35190 ( .A1(n3686), .A2(n3807), .ZN(n2785) );
  OR2_X1 U35200 ( .A1(n2830), .A2(n2785), .ZN(n3021) );
  NAND2_X1 U35210 ( .A1(n2786), .A2(n3021), .ZN(n2924) );
  NAND2_X1 U35220 ( .A1(n2348), .A2(n2831), .ZN(n2787) );
  OAI21_X1 U35230 ( .B1(n2924), .B2(n2787), .A(STATE_REG_SCAN_IN), .ZN(n2789)
         );
  INV_X1 U35240 ( .A(n4400), .ZN(n2811) );
  INV_X1 U35250 ( .A(n2799), .ZN(n3693) );
  NAND2_X1 U35260 ( .A1(n2800), .A2(n3693), .ZN(n2925) );
  NAND2_X2 U35270 ( .A1(n2789), .A2(n2925), .ZN(n3522) );
  NOR3_X1 U35280 ( .A1(n2800), .A2(n4059), .A3(n3024), .ZN(n2791) );
  AND2_X1 U35290 ( .A1(n3686), .A2(n4269), .ZN(n4385) );
  NAND2_X1 U35300 ( .A1(n4460), .A2(n3579), .ZN(n3022) );
  OAI22_X1 U35310 ( .A1(n2792), .A2(n3821), .B1(STATE_REG_SCAN_IN), .B2(n2793), 
        .ZN(n2806) );
  INV_X1 U35320 ( .A(n2794), .ZN(n3819) );
  INV_X1 U35330 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2797) );
  NAND2_X1 U35340 ( .A1(n2054), .A2(REG0_REG_29__SCAN_IN), .ZN(n2796) );
  NAND2_X1 U35350 ( .A1(n3531), .A2(REG2_REG_29__SCAN_IN), .ZN(n2795) );
  OAI211_X1 U35360 ( .C1(n2797), .C2(n3533), .A(n2796), .B(n2795), .ZN(n2798)
         );
  AOI21_X1 U35370 ( .B1(n3819), .B2(n2668), .A(n2798), .ZN(n3596) );
  NOR2_X1 U35380 ( .A1(n2800), .A2(n2799), .ZN(n2804) );
  NAND2_X1 U35390 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(
        n2802) );
  NAND2_X1 U35400 ( .A1(n2801), .A2(n2802), .ZN(n2803) );
  NAND2_X1 U35410 ( .A1(n2804), .A2(n4264), .ZN(n3519) );
  OAI22_X1 U35420 ( .A1(n3596), .A2(n3518), .B1(n3867), .B2(n3519), .ZN(n2805)
         );
  AOI211_X1 U35430 ( .C1(n3833), .C2(n3522), .A(n2806), .B(n2805), .ZN(n2807)
         );
  NAND3_X1 U35440 ( .A1(n2810), .A2(n2809), .A3(n2275), .ZN(U3217) );
  INV_X2 U35450 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  MUX2_X1 U35460 ( .A(n2812), .B(n2908), .S(STATE_REG_SCAN_IN), .Z(n2813) );
  INV_X1 U35470 ( .A(n2813), .ZN(U3344) );
  NAND2_X1 U35480 ( .A1(U3149), .A2(DATAI_25_), .ZN(n2814) );
  OAI21_X1 U35490 ( .B1(n2815), .B2(U3149), .A(n2814), .ZN(U3327) );
  INV_X1 U35500 ( .A(DATAI_26_), .ZN(n4611) );
  NAND2_X1 U35510 ( .A1(n2756), .A2(STATE_REG_SCAN_IN), .ZN(n2816) );
  OAI21_X1 U35520 ( .B1(STATE_REG_SCAN_IN), .B2(n4611), .A(n2816), .ZN(U3326)
         );
  INV_X1 U35530 ( .A(DATAI_27_), .ZN(n2818) );
  XNOR2_X1 U35540 ( .A(n2801), .B(IR_REG_27__SCAN_IN), .ZN(n3815) );
  NAND2_X1 U35550 ( .A1(n3815), .A2(STATE_REG_SCAN_IN), .ZN(n2817) );
  OAI21_X1 U35560 ( .B1(STATE_REG_SCAN_IN), .B2(n2818), .A(n2817), .ZN(U3325)
         );
  INV_X1 U35570 ( .A(DATAI_31_), .ZN(n4635) );
  INV_X1 U35580 ( .A(n2819), .ZN(n2821) );
  OR4_X1 U35590 ( .A1(n2821), .A2(IR_REG_30__SCAN_IN), .A3(n2820), .A4(U3149), 
        .ZN(n2822) );
  OAI21_X1 U35600 ( .B1(STATE_REG_SCAN_IN), .B2(n4635), .A(n2822), .ZN(U3321)
         );
  INV_X1 U35610 ( .A(n3024), .ZN(n2926) );
  INV_X1 U35620 ( .A(n3025), .ZN(n2823) );
  AOI22_X1 U35630 ( .A1(n4399), .A2(n2824), .B1(n2823), .B2(n4400), .ZN(U3459)
         );
  AOI22_X1 U35640 ( .A1(n4399), .A2(n4501), .B1(n2825), .B2(n4400), .ZN(U3458)
         );
  INV_X1 U35650 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n4618) );
  NAND2_X1 U35660 ( .A1(n2975), .A2(U4043), .ZN(n2826) );
  OAI21_X1 U35670 ( .B1(U4043), .B2(n4618), .A(n2826), .ZN(U3550) );
  INV_X1 U35680 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n4493) );
  NAND2_X1 U35690 ( .A1(n3050), .A2(U4043), .ZN(n2827) );
  OAI21_X1 U35700 ( .B1(U4043), .B2(n4493), .A(n2827), .ZN(U3553) );
  INV_X1 U35710 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n4650) );
  INV_X1 U35720 ( .A(n3182), .ZN(n3188) );
  NAND2_X1 U35730 ( .A1(n3188), .A2(U4043), .ZN(n2828) );
  OAI21_X1 U35740 ( .B1(U4043), .B2(n4650), .A(n2828), .ZN(U3558) );
  INV_X1 U35750 ( .A(n2831), .ZN(n2829) );
  NAND2_X1 U35760 ( .A1(n2829), .A2(STATE_REG_SCAN_IN), .ZN(n3696) );
  NAND2_X1 U35770 ( .A1(n3024), .A2(n3696), .ZN(n2843) );
  INV_X1 U35780 ( .A(n2830), .ZN(n2972) );
  NAND2_X1 U35790 ( .A1(n2972), .A2(n2831), .ZN(n2832) );
  AND2_X1 U35800 ( .A1(n2433), .A2(n2832), .ZN(n2844) );
  INV_X1 U35810 ( .A(n4335), .ZN(n4376) );
  INV_X1 U3582 ( .A(n3815), .ZN(n2837) );
  XNOR2_X1 U3583 ( .A(n4276), .B(REG1_REG_2__SCAN_IN), .ZN(n3739) );
  AND2_X1 U3584 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3724)
         );
  NAND2_X1 U3585 ( .A1(n4277), .A2(REG1_REG_1__SCAN_IN), .ZN(n2833) );
  OAI211_X1 U3586 ( .C1(n4277), .C2(REG1_REG_1__SCAN_IN), .A(n3724), .B(n2833), 
        .ZN(n3722) );
  NAND2_X1 U3587 ( .A1(n3722), .A2(n2833), .ZN(n3738) );
  INV_X1 U3588 ( .A(n3738), .ZN(n2834) );
  NAND2_X1 U3589 ( .A1(n4276), .A2(REG1_REG_2__SCAN_IN), .ZN(n2835) );
  NAND2_X1 U3590 ( .A1(n2836), .A2(n2835), .ZN(n2859) );
  XNOR2_X1 U3591 ( .A(n2859), .B(n2848), .ZN(n2858) );
  XOR2_X1 U3592 ( .A(n2858), .B(REG1_REG_3__SCAN_IN), .Z(n2842) );
  NOR2_X1 U3593 ( .A1(n2837), .A2(n3732), .ZN(n3692) );
  INV_X1 U3594 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2838) );
  MUX2_X1 U3595 ( .A(REG2_REG_2__SCAN_IN), .B(n2838), .S(n4276), .Z(n3743) );
  INV_X1 U3596 ( .A(REG2_REG_1__SCAN_IN), .ZN(n4606) );
  XNOR2_X1 U3597 ( .A(n4277), .B(n4606), .ZN(n3726) );
  AND2_X1 U3598 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3731)
         );
  NAND2_X1 U3599 ( .A1(n3726), .A2(n3731), .ZN(n3725) );
  NAND2_X1 U3600 ( .A1(n4277), .A2(REG2_REG_1__SCAN_IN), .ZN(n2839) );
  NAND2_X1 U3601 ( .A1(n3725), .A2(n2839), .ZN(n3742) );
  NAND2_X1 U3602 ( .A1(n3743), .A2(n3742), .ZN(n3741) );
  NAND2_X1 U3603 ( .A1(n4276), .A2(REG2_REG_2__SCAN_IN), .ZN(n2840) );
  NAND2_X1 U3604 ( .A1(n3741), .A2(n2840), .ZN(n2850) );
  XNOR2_X1 U3605 ( .A(n2850), .B(n2848), .ZN(n2849) );
  XOR2_X1 U3606 ( .A(REG2_REG_3__SCAN_IN), .B(n2849), .Z(n2841) );
  AOI22_X1 U3607 ( .A1(n4359), .A2(n2842), .B1(n4373), .B2(n2841), .ZN(n2847)
         );
  INV_X1 U3608 ( .A(n2843), .ZN(n2845) );
  AOI22_X1 U3609 ( .A1(n4351), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n2846) );
  OAI211_X1 U3610 ( .C1(n2848), .C2(n4376), .A(n2847), .B(n2846), .ZN(U3243)
         );
  NAND2_X1 U3611 ( .A1(n2850), .A2(n4275), .ZN(n2851) );
  AOI22_X1 U3612 ( .A1(n2853), .A2(REG2_REG_4__SCAN_IN), .B1(n4274), .B2(n2852), .ZN(n2856) );
  INV_X1 U3613 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2854) );
  MUX2_X1 U3614 ( .A(REG2_REG_5__SCAN_IN), .B(n2854), .S(n2871), .Z(n2855) );
  AOI211_X1 U3615 ( .C1(n2856), .C2(n2855), .A(n2878), .B(n4328), .ZN(n2870)
         );
  AND2_X1 U3616 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n2951) );
  AOI21_X1 U3617 ( .B1(n4351), .B2(ADDR_REG_5__SCAN_IN), .A(n2951), .ZN(n2868)
         );
  MUX2_X1 U3618 ( .A(n2857), .B(REG1_REG_5__SCAN_IN), .S(n2871), .Z(n2866) );
  NAND2_X1 U3619 ( .A1(n2858), .A2(REG1_REG_3__SCAN_IN), .ZN(n2861) );
  NAND2_X1 U3620 ( .A1(n2859), .A2(n4275), .ZN(n2860) );
  NAND2_X1 U3621 ( .A1(n2863), .A2(n4274), .ZN(n2864) );
  NAND2_X1 U3622 ( .A1(n2865), .A2(n2866), .ZN(n2873) );
  OAI211_X1 U3623 ( .C1(n2866), .C2(n2865), .A(n4359), .B(n2873), .ZN(n2867)
         );
  OAI211_X1 U3624 ( .C1(n4376), .C2(n2871), .A(n2868), .B(n2867), .ZN(n2869)
         );
  OR2_X1 U3625 ( .A1(n2870), .A2(n2869), .ZN(U3245) );
  NOR2_X1 U3626 ( .A1(n4351), .A2(U4043), .ZN(U3148) );
  MUX2_X1 U3627 ( .A(n2427), .B(REG1_REG_7__SCAN_IN), .S(n4271), .Z(n2876) );
  INV_X1 U3628 ( .A(n2871), .ZN(n4273) );
  NAND2_X1 U3629 ( .A1(n4273), .A2(REG1_REG_5__SCAN_IN), .ZN(n2872) );
  NAND2_X1 U3630 ( .A1(n2873), .A2(n2872), .ZN(n2874) );
  INV_X1 U3631 ( .A(n4272), .ZN(n2916) );
  NAND2_X1 U3632 ( .A1(n2874), .A2(n4272), .ZN(n2875) );
  XOR2_X1 U3633 ( .A(n2876), .B(n2892), .Z(n2884) );
  NAND2_X1 U3634 ( .A1(n4351), .A2(ADDR_REG_7__SCAN_IN), .ZN(n2877) );
  NAND2_X1 U3635 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3001) );
  NAND2_X1 U3636 ( .A1(n2877), .A2(n3001), .ZN(n2882) );
  INV_X1 U3637 ( .A(REG2_REG_7__SCAN_IN), .ZN(n4482) );
  MUX2_X1 U3638 ( .A(n4482), .B(REG2_REG_7__SCAN_IN), .S(n4271), .Z(n2879) );
  NOR2_X1 U3639 ( .A1(n2880), .A2(n2879), .ZN(n2885) );
  AOI211_X1 U3640 ( .C1(n2880), .C2(n2879), .A(n4328), .B(n2885), .ZN(n2881)
         );
  AOI211_X1 U3641 ( .C1(n4335), .C2(n4271), .A(n2882), .B(n2881), .ZN(n2883)
         );
  OAI21_X1 U3642 ( .B1(n4362), .B2(n2884), .A(n2883), .ZN(U3247) );
  INV_X1 U3643 ( .A(n3778), .ZN(n4666) );
  AOI21_X1 U3644 ( .B1(n4271), .B2(REG2_REG_7__SCAN_IN), .A(n2885), .ZN(n2886)
         );
  INV_X1 U3645 ( .A(n2908), .ZN(n2896) );
  XNOR2_X1 U3646 ( .A(n2886), .B(n2896), .ZN(n2903) );
  INV_X1 U3647 ( .A(n2886), .ZN(n2887) );
  AOI22_X1 U3648 ( .A1(n2903), .A2(REG2_REG_8__SCAN_IN), .B1(n2896), .B2(n2887), .ZN(n2889) );
  INV_X1 U3649 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3761) );
  MUX2_X1 U3650 ( .A(n3761), .B(REG2_REG_9__SCAN_IN), .S(n3778), .Z(n2888) );
  NOR2_X1 U3651 ( .A1(n2889), .A2(n2888), .ZN(n3759) );
  AOI211_X1 U3652 ( .C1(n2889), .C2(n2888), .A(n4328), .B(n3759), .ZN(n2890)
         );
  INV_X1 U3653 ( .A(n2890), .ZN(n2902) );
  NOR2_X1 U3654 ( .A1(STATE_REG_SCAN_IN), .A2(n2891), .ZN(n3171) );
  OR2_X1 U3655 ( .A1(n4271), .A2(REG1_REG_7__SCAN_IN), .ZN(n2893) );
  NAND2_X1 U3656 ( .A1(n2894), .A2(n2893), .ZN(n2895) );
  INV_X1 U3657 ( .A(n2895), .ZN(n2897) );
  MUX2_X1 U3658 ( .A(n2898), .B(REG1_REG_9__SCAN_IN), .S(n3778), .Z(n2899) );
  AOI211_X1 U3659 ( .C1(n2086), .C2(n2899), .A(n3777), .B(n4362), .ZN(n2900)
         );
  AOI211_X1 U3660 ( .C1(n4351), .C2(ADDR_REG_9__SCAN_IN), .A(n3171), .B(n2900), 
        .ZN(n2901) );
  OAI211_X1 U3661 ( .C1(n4376), .C2(n4666), .A(n2902), .B(n2901), .ZN(U3249)
         );
  XOR2_X1 U3662 ( .A(REG2_REG_8__SCAN_IN), .B(n2903), .Z(n2911) );
  AOI211_X1 U3663 ( .C1(n2441), .C2(n2905), .A(n4362), .B(n2904), .ZN(n2910)
         );
  NAND2_X1 U3664 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3099) );
  INV_X1 U3665 ( .A(n3099), .ZN(n2906) );
  AOI21_X1 U3666 ( .B1(n4351), .B2(ADDR_REG_8__SCAN_IN), .A(n2906), .ZN(n2907)
         );
  OAI21_X1 U3667 ( .B1(n4376), .B2(n2908), .A(n2907), .ZN(n2909) );
  AOI211_X1 U3668 ( .C1(n2911), .C2(n4373), .A(n2910), .B(n2909), .ZN(n2912)
         );
  INV_X1 U3669 ( .A(n2912), .ZN(U3248) );
  XNOR2_X1 U3670 ( .A(n2913), .B(REG2_REG_6__SCAN_IN), .ZN(n2920) );
  XOR2_X1 U3671 ( .A(REG1_REG_6__SCAN_IN), .B(n2914), .Z(n2918) );
  AND2_X1 U3672 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n2961) );
  AOI21_X1 U3673 ( .B1(n4351), .B2(ADDR_REG_6__SCAN_IN), .A(n2961), .ZN(n2915)
         );
  OAI21_X1 U3674 ( .B1(n4376), .B2(n2916), .A(n2915), .ZN(n2917) );
  AOI21_X1 U3675 ( .B1(n4359), .B2(n2918), .A(n2917), .ZN(n2919) );
  OAI21_X1 U3676 ( .B1(n2920), .B2(n4328), .A(n2919), .ZN(U3246) );
  OAI21_X1 U3677 ( .B1(n2923), .B2(n2922), .A(n2921), .ZN(n3735) );
  INV_X1 U3678 ( .A(n2924), .ZN(n2927) );
  NAND3_X1 U3679 ( .A1(n2927), .A2(n2926), .A3(n2925), .ZN(n3420) );
  OAI22_X1 U3680 ( .A1(n2792), .A2(n4384), .B1(n2340), .B2(n3518), .ZN(n2928)
         );
  AOI21_X1 U3681 ( .B1(REG3_REG_0__SCAN_IN), .B2(n3420), .A(n2928), .ZN(n2929)
         );
  OAI21_X1 U3682 ( .B1(n3525), .B2(n3735), .A(n2929), .ZN(U3229) );
  NAND2_X1 U3683 ( .A1(n2931), .A2(n2932), .ZN(n2935) );
  INV_X1 U3684 ( .A(n2933), .ZN(n2934) );
  AOI21_X1 U3685 ( .B1(n2930), .B2(n2935), .A(n2934), .ZN(n2938) );
  INV_X1 U3686 ( .A(n3519), .ZN(n3417) );
  AOI22_X1 U3687 ( .A1(n3521), .A2(n3034), .B1(n3417), .B2(n2971), .ZN(n2937)
         );
  INV_X1 U3688 ( .A(n3518), .ZN(n3419) );
  AOI22_X1 U3689 ( .A1(REG3_REG_2__SCAN_IN), .A2(n3420), .B1(n3419), .B2(n3050), .ZN(n2936) );
  OAI211_X1 U3690 ( .C1(n2938), .C2(n3525), .A(n2937), .B(n2936), .ZN(U3234)
         );
  XOR2_X1 U3691 ( .A(n2940), .B(n2939), .Z(n2944) );
  MUX2_X1 U3692 ( .A(U3149), .B(n3522), .S(n3088), .Z(n2942) );
  OAI22_X1 U3693 ( .A1(n2792), .A2(n3086), .B1(n3006), .B2(n3519), .ZN(n2941)
         );
  AOI211_X1 U3694 ( .C1(n3419), .C2(n3712), .A(n2942), .B(n2941), .ZN(n2943)
         );
  OAI21_X1 U3695 ( .B1(n2944), .B2(n3525), .A(n2943), .ZN(U3215) );
  INV_X1 U3696 ( .A(n3522), .ZN(n2955) );
  INV_X1 U3697 ( .A(n3075), .ZN(n2954) );
  OR2_X1 U3698 ( .A1(n2945), .A2(n2994), .ZN(n2992) );
  NAND2_X1 U3699 ( .A1(n2992), .A2(n2946), .ZN(n2949) );
  NAND2_X1 U3700 ( .A1(n2949), .A2(n2948), .ZN(n2947) );
  OAI211_X1 U3701 ( .C1(n2949), .C2(n2948), .A(n2947), .B(n3428), .ZN(n2953)
         );
  INV_X1 U3702 ( .A(n3710), .ZN(n3104) );
  OAI22_X1 U3703 ( .A1(n3070), .A2(n3519), .B1(n3518), .B2(n3104), .ZN(n2950)
         );
  AOI211_X1 U3704 ( .C1(n3108), .C2(n3521), .A(n2951), .B(n2950), .ZN(n2952)
         );
  OAI211_X1 U3705 ( .C1(n2955), .C2(n2954), .A(n2953), .B(n2952), .ZN(U3224)
         );
  XOR2_X1 U3706 ( .A(n2957), .B(n2956), .Z(n2958) );
  XNOR2_X1 U3707 ( .A(n2959), .B(n2958), .ZN(n2965) );
  OAI22_X1 U3708 ( .A1(n3115), .A2(n3519), .B1(n3518), .B2(n3129), .ZN(n2960)
         );
  AOI211_X1 U3709 ( .C1(n3134), .C2(n3521), .A(n2961), .B(n2960), .ZN(n2964)
         );
  NAND2_X1 U3710 ( .A1(n3522), .A2(n2962), .ZN(n2963) );
  OAI211_X1 U3711 ( .C1(n2965), .C2(n3525), .A(n2964), .B(n2963), .ZN(U3236)
         );
  INV_X1 U3712 ( .A(n3021), .ZN(n2966) );
  OR2_X1 U3713 ( .A1(n3024), .A2(n2966), .ZN(n2967) );
  OR2_X1 U3714 ( .A1(n2968), .A2(n2967), .ZN(n2969) );
  NAND2_X1 U3715 ( .A1(n2973), .A2(n4384), .ZN(n3033) );
  OAI21_X1 U3716 ( .B1(n4384), .B2(n2973), .A(n3033), .ZN(n4421) );
  NAND2_X1 U3717 ( .A1(n4266), .A2(n4269), .ZN(n2970) );
  OR2_X1 U3718 ( .A1(n3579), .A2(n3686), .ZN(n3559) );
  NAND2_X1 U3719 ( .A1(n2347), .A2(n2974), .ZN(n3567) );
  INV_X1 U3720 ( .A(n3567), .ZN(n3616) );
  XNOR2_X1 U3721 ( .A(n3602), .B(n3616), .ZN(n2983) );
  OAI22_X1 U3722 ( .A1(n3006), .A2(n4388), .B1(n4059), .B2(n2973), .ZN(n2981)
         );
  OR2_X1 U3723 ( .A1(n3602), .A2(n2976), .ZN(n2977) );
  NAND2_X1 U3724 ( .A1(n3008), .A2(n2977), .ZN(n4422) );
  XNOR2_X1 U3725 ( .A(n2978), .B(n4266), .ZN(n2979) );
  NAND2_X1 U3726 ( .A1(n2979), .A2(n3807), .ZN(n4109) );
  NOR2_X1 U3727 ( .A1(n4422), .A2(n4109), .ZN(n2980) );
  AOI211_X1 U3728 ( .C1(n4071), .C2(n2975), .A(n2981), .B(n2980), .ZN(n2982)
         );
  OAI21_X1 U3729 ( .B1(n4065), .B2(n2983), .A(n2982), .ZN(n4424) );
  NAND2_X1 U3730 ( .A1(n4424), .A2(n4118), .ZN(n2990) );
  INV_X1 U3731 ( .A(n4422), .ZN(n2988) );
  NAND2_X1 U3732 ( .A1(n2984), .A2(n4269), .ZN(n3062) );
  INV_X1 U3733 ( .A(n3062), .ZN(n2985) );
  NAND2_X1 U3734 ( .A1(n4118), .A2(n2985), .ZN(n4123) );
  INV_X1 U3735 ( .A(n4123), .ZN(n4393) );
  INV_X1 U3736 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2986) );
  OAI22_X1 U3737 ( .A1(n4118), .A2(n4606), .B1(n2986), .B2(n4115), .ZN(n2987)
         );
  AOI21_X1 U3738 ( .B1(n2988), .B2(n4393), .A(n2987), .ZN(n2989) );
  OAI211_X1 U3739 ( .C1(n4088), .C2(n4421), .A(n2990), .B(n2989), .ZN(U3289)
         );
  AOI22_X1 U3740 ( .A1(n3419), .A2(n3711), .B1(n3417), .B2(n3050), .ZN(n2991)
         );
  NAND2_X1 U3741 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3749) );
  OAI211_X1 U3742 ( .C1(n2792), .C2(n3055), .A(n2991), .B(n3749), .ZN(n2996)
         );
  INV_X1 U3743 ( .A(n2992), .ZN(n2993) );
  AOI211_X1 U3744 ( .C1(n2994), .C2(n2945), .A(n3525), .B(n2993), .ZN(n2995)
         );
  AOI211_X1 U3745 ( .C1(n2997), .C2(n3522), .A(n2996), .B(n2995), .ZN(n2998)
         );
  INV_X1 U3746 ( .A(n2998), .ZN(U3227) );
  XNOR2_X1 U3747 ( .A(n2999), .B(n3000), .ZN(n3005) );
  AOI22_X1 U3748 ( .A1(n3419), .A2(n3188), .B1(n3417), .B2(n3710), .ZN(n3002)
         );
  OAI211_X1 U3749 ( .C1(n2792), .C2(n3160), .A(n3002), .B(n3001), .ZN(n3003)
         );
  AOI21_X1 U3750 ( .B1(n3162), .B2(n3522), .A(n3003), .ZN(n3004) );
  OAI21_X1 U3751 ( .B1(n3005), .B2(n3525), .A(n3004), .ZN(U3210) );
  NAND2_X1 U3752 ( .A1(n3006), .A2(n3034), .ZN(n3617) );
  INV_X1 U3753 ( .A(n3006), .ZN(n3713) );
  NAND2_X1 U3754 ( .A1(n3713), .A2(n3042), .ZN(n3620) );
  NAND2_X1 U3755 ( .A1(n3617), .A2(n3620), .ZN(n3009) );
  NAND2_X1 U3756 ( .A1(n2971), .A2(n3418), .ZN(n3007) );
  NAND2_X1 U3757 ( .A1(n3008), .A2(n3007), .ZN(n3012) );
  INV_X1 U3758 ( .A(n3012), .ZN(n3010) );
  INV_X1 U3759 ( .A(n3044), .ZN(n3011) );
  AOI21_X1 U3760 ( .B1(n3604), .B2(n3012), .A(n3011), .ZN(n3016) );
  INV_X1 U3761 ( .A(n3016), .ZN(n4379) );
  OR2_X1 U3762 ( .A1(n3602), .A2(n3567), .ZN(n3014) );
  INV_X1 U3763 ( .A(n3050), .ZN(n3048) );
  AOI22_X1 U3764 ( .A1(n2971), .A2(n4071), .B1(n3034), .B2(n4135), .ZN(n3015)
         );
  OAI21_X1 U3765 ( .B1(n3048), .B2(n4388), .A(n3015), .ZN(n3018) );
  NOR2_X1 U3766 ( .A1(n3016), .A2(n4109), .ZN(n3017) );
  AOI211_X1 U3767 ( .C1(n4386), .C2(n3019), .A(n3018), .B(n3017), .ZN(n4382)
         );
  INV_X1 U3768 ( .A(n4382), .ZN(n3020) );
  AOI21_X1 U3769 ( .B1(n4460), .B2(n4379), .A(n3020), .ZN(n3041) );
  NAND2_X1 U3770 ( .A1(n3022), .A2(n3021), .ZN(n3023) );
  NOR2_X1 U3771 ( .A1(n3024), .A2(n3023), .ZN(n3031) );
  OAI21_X1 U3772 ( .B1(n3026), .B2(D_REG_1__SCAN_IN), .A(n3025), .ZN(n3030) );
  NAND2_X1 U3773 ( .A1(n3028), .A2(n3027), .ZN(n3029) );
  INV_X1 U3774 ( .A(n3037), .ZN(n3032) );
  AOI21_X1 U3775 ( .B1(n3034), .B2(n3033), .A(n3087), .ZN(n4377) );
  INV_X1 U3776 ( .A(n4261), .ZN(n3035) );
  AOI22_X1 U3777 ( .A1(n4377), .A2(n3035), .B1(n4461), .B2(REG0_REG_2__SCAN_IN), .ZN(n3036) );
  OAI21_X1 U3778 ( .B1(n3041), .B2(n4461), .A(n3036), .ZN(U3471) );
  INV_X1 U3779 ( .A(n4206), .ZN(n3039) );
  AOI22_X1 U3780 ( .A1(n4377), .A2(n3039), .B1(REG1_REG_2__SCAN_IN), .B2(n4472), .ZN(n3040) );
  OAI21_X1 U3781 ( .B1(n3041), .B2(n4472), .A(n3040), .ZN(U3520) );
  NAND2_X1 U3782 ( .A1(n3006), .A2(n3042), .ZN(n3043) );
  NAND2_X1 U3783 ( .A1(n3048), .A2(n3086), .ZN(n3045) );
  NAND2_X1 U3784 ( .A1(n3712), .A2(n3055), .ZN(n3626) );
  NAND2_X1 U3785 ( .A1(n3070), .A2(n3064), .ZN(n3623) );
  OR2_X1 U3786 ( .A1(n3111), .A2(n3105), .ZN(n3065) );
  NAND2_X1 U3787 ( .A1(n3111), .A2(n3105), .ZN(n3046) );
  AND2_X1 U3788 ( .A1(n3065), .A2(n3046), .ZN(n4435) );
  INV_X1 U3789 ( .A(n4435), .ZN(n3061) );
  NAND2_X1 U3790 ( .A1(n3047), .A2(n3617), .ZN(n3079) );
  NAND2_X1 U3791 ( .A1(n3048), .A2(n3080), .ZN(n3622) );
  NAND2_X1 U3792 ( .A1(n3050), .A2(n3086), .ZN(n3619) );
  NAND2_X1 U3793 ( .A1(n3079), .A2(n3603), .ZN(n3049) );
  XOR2_X1 U3794 ( .A(n3105), .B(n3068), .Z(n3054) );
  INV_X1 U3795 ( .A(n4109), .ZN(n4387) );
  AOI22_X1 U3796 ( .A1(n3050), .A2(n4071), .B1(n3064), .B2(n4135), .ZN(n3051)
         );
  OAI21_X1 U3797 ( .B1(n3115), .B2(n4388), .A(n3051), .ZN(n3052) );
  AOI21_X1 U3798 ( .B1(n4435), .B2(n4387), .A(n3052), .ZN(n3053) );
  OAI21_X1 U3799 ( .B1(n4065), .B2(n3054), .A(n3053), .ZN(n4433) );
  NAND2_X1 U3800 ( .A1(n3087), .A2(n3086), .ZN(n3085) );
  INV_X1 U3801 ( .A(n3085), .ZN(n3056) );
  OAI211_X1 U3802 ( .C1(n3056), .C2(n3055), .A(n4443), .B(n3073), .ZN(n4432)
         );
  OAI22_X1 U3803 ( .A1(n4432), .A2(n4269), .B1(n4115), .B2(n3057), .ZN(n3058)
         );
  OAI21_X1 U3804 ( .B1(n4433), .B2(n3058), .A(n4118), .ZN(n3060) );
  NAND2_X1 U3805 ( .A1(n4281), .A2(REG2_REG_4__SCAN_IN), .ZN(n3059) );
  OAI211_X1 U3806 ( .C1(n3061), .C2(n4123), .A(n3060), .B(n3059), .ZN(U3286)
         );
  NAND2_X1 U3807 ( .A1(n4109), .A2(n3062), .ZN(n3063) );
  AND2_X1 U3808 ( .A1(n3711), .A2(n3106), .ZN(n3112) );
  INV_X1 U3809 ( .A(n3112), .ZN(n3625) );
  NAND2_X1 U3810 ( .A1(n3115), .A2(n3108), .ZN(n3640) );
  NAND2_X1 U3811 ( .A1(n3712), .A2(n3064), .ZN(n3109) );
  NAND2_X1 U3812 ( .A1(n3065), .A2(n3109), .ZN(n3066) );
  XOR2_X1 U3813 ( .A(n3591), .B(n3066), .Z(n4439) );
  INV_X1 U3814 ( .A(n3623), .ZN(n3067) );
  XOR2_X1 U3815 ( .A(n3591), .B(n3113), .Z(n3072) );
  AOI22_X1 U3816 ( .A1(n3710), .A2(n4101), .B1(n4135), .B2(n3108), .ZN(n3069)
         );
  OAI21_X1 U3817 ( .B1(n3070), .B2(n4104), .A(n3069), .ZN(n3071) );
  AOI21_X1 U3818 ( .B1(n3072), .B2(n4386), .A(n3071), .ZN(n4437) );
  MUX2_X1 U3819 ( .A(n4437), .B(n2854), .S(n4281), .Z(n3077) );
  AND2_X1 U3820 ( .A1(n3073), .A2(n3108), .ZN(n3074) );
  NOR2_X1 U3821 ( .A1(n3119), .A2(n3074), .ZN(n4442) );
  AOI22_X1 U3822 ( .A1(n4442), .A2(n4378), .B1(n3075), .B2(n4392), .ZN(n3076)
         );
  OAI211_X1 U3823 ( .C1(n4092), .C2(n4439), .A(n3077), .B(n3076), .ZN(U3285)
         );
  XNOR2_X1 U3824 ( .A(n3078), .B(n3603), .ZN(n4428) );
  XNOR2_X1 U3825 ( .A(n3079), .B(n3603), .ZN(n3083) );
  AOI22_X1 U3826 ( .A1(n3712), .A2(n4101), .B1(n4135), .B2(n3080), .ZN(n3081)
         );
  OAI21_X1 U3827 ( .B1(n3006), .B2(n4104), .A(n3081), .ZN(n3082) );
  AOI21_X1 U3828 ( .B1(n3083), .B2(n4386), .A(n3082), .ZN(n3084) );
  OAI21_X1 U3829 ( .B1(n4428), .B2(n4109), .A(n3084), .ZN(n4430) );
  INV_X1 U3830 ( .A(n4430), .ZN(n3093) );
  INV_X2 U3831 ( .A(n4118), .ZN(n4281) );
  INV_X1 U3832 ( .A(n4428), .ZN(n3091) );
  OAI21_X1 U3833 ( .B1(n3087), .B2(n3086), .A(n3085), .ZN(n4426) );
  AOI22_X1 U3834 ( .A1(n4281), .A2(REG2_REG_3__SCAN_IN), .B1(n4392), .B2(n3088), .ZN(n3089) );
  OAI21_X1 U3835 ( .B1(n4088), .B2(n4426), .A(n3089), .ZN(n3090) );
  AOI21_X1 U3836 ( .B1(n3091), .B2(n4393), .A(n3090), .ZN(n3092) );
  OAI21_X1 U3837 ( .B1(n3093), .B2(n4281), .A(n3092), .ZN(U3287) );
  INV_X1 U3838 ( .A(n3095), .ZN(n3097) );
  NOR2_X1 U3839 ( .A1(n3097), .A2(n3096), .ZN(n3098) );
  XNOR2_X1 U3840 ( .A(n3094), .B(n3098), .ZN(n3103) );
  AOI22_X1 U3841 ( .A1(n3417), .A2(n3708), .B1(n3419), .B2(n3707), .ZN(n3100)
         );
  OAI211_X1 U3842 ( .C1(n2792), .C2(n3181), .A(n3100), .B(n3099), .ZN(n3101)
         );
  AOI21_X1 U3843 ( .B1(n3141), .B2(n3522), .A(n3101), .ZN(n3102) );
  OAI21_X1 U3844 ( .B1(n3103), .B2(n3525), .A(n3102), .ZN(U3218) );
  NAND2_X1 U3845 ( .A1(n3104), .A2(n3134), .ZN(n3628) );
  NAND2_X1 U3846 ( .A1(n3710), .A2(n3118), .ZN(n3638) );
  AND2_X1 U3847 ( .A1(n3628), .A2(n3638), .ZN(n3607) );
  AND2_X1 U3848 ( .A1(n3115), .A2(n3106), .ZN(n3110) );
  INV_X1 U3849 ( .A(n3110), .ZN(n3107) );
  XOR2_X1 U3850 ( .A(n3607), .B(n3136), .Z(n3149) );
  INV_X1 U3851 ( .A(n4460), .ZN(n4427) );
  INV_X1 U3852 ( .A(n4453), .ZN(n4438) );
  XNOR2_X1 U3853 ( .A(n3127), .B(n3607), .ZN(n3117) );
  AOI22_X1 U3854 ( .A1(n3708), .A2(n4101), .B1(n4135), .B2(n3134), .ZN(n3114)
         );
  OAI21_X1 U3855 ( .B1(n3115), .B2(n4104), .A(n3114), .ZN(n3116) );
  AOI21_X1 U3856 ( .B1(n3117), .B2(n4386), .A(n3116), .ZN(n3154) );
  OAI21_X1 U3857 ( .B1(n3149), .B2(n4438), .A(n3154), .ZN(n3125) );
  NOR2_X1 U3858 ( .A1(n3119), .A2(n3118), .ZN(n3120) );
  OR2_X1 U3859 ( .A1(n3161), .A2(n3120), .ZN(n3146) );
  INV_X1 U3860 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3121) );
  OAI22_X1 U3861 ( .A1(n3146), .A2(n4261), .B1(n4463), .B2(n3121), .ZN(n3122)
         );
  AOI21_X1 U3862 ( .B1(n3125), .B2(n4463), .A(n3122), .ZN(n3123) );
  INV_X1 U3863 ( .A(n3123), .ZN(U3479) );
  OAI22_X1 U3864 ( .A1(n3146), .A2(n4206), .B1(n4474), .B2(n2408), .ZN(n3124)
         );
  AOI21_X1 U3865 ( .B1(n3125), .B2(n4474), .A(n3124), .ZN(n3126) );
  INV_X1 U3866 ( .A(n3126), .ZN(U3524) );
  NAND2_X1 U3867 ( .A1(n3127), .A2(n3638), .ZN(n3128) );
  NAND2_X1 U3868 ( .A1(n3129), .A2(n3138), .ZN(n3137) );
  INV_X1 U3869 ( .A(n3137), .ZN(n3130) );
  NAND2_X1 U3870 ( .A1(n3708), .A2(n3160), .ZN(n3632) );
  NAND2_X1 U3871 ( .A1(n3182), .A2(n3187), .ZN(n3633) );
  NAND2_X1 U3872 ( .A1(n3188), .A2(n3181), .ZN(n3631) );
  AND2_X1 U3873 ( .A1(n3633), .A2(n3631), .ZN(n3587) );
  XNOR2_X1 U3874 ( .A(n3175), .B(n3587), .ZN(n3133) );
  INV_X1 U3875 ( .A(n3707), .ZN(n3214) );
  OAI22_X1 U3876 ( .A1(n3214), .A2(n4388), .B1(n4059), .B2(n3181), .ZN(n3131)
         );
  AOI21_X1 U3877 ( .B1(n4071), .B2(n3708), .A(n3131), .ZN(n3132) );
  OAI21_X1 U3878 ( .B1(n3133), .B2(n4065), .A(n3132), .ZN(n3200) );
  INV_X1 U3879 ( .A(n3200), .ZN(n3145) );
  AND2_X1 U3880 ( .A1(n3710), .A2(n3134), .ZN(n3135) );
  NAND2_X1 U3881 ( .A1(n3708), .A2(n3138), .ZN(n3185) );
  NAND2_X1 U3882 ( .A1(n4446), .A2(n3185), .ZN(n3139) );
  XNOR2_X1 U3883 ( .A(n3139), .B(n3587), .ZN(n3201) );
  NAND2_X1 U3884 ( .A1(n3159), .A2(n3187), .ZN(n3140) );
  AOI22_X1 U3885 ( .A1(n4281), .A2(REG2_REG_8__SCAN_IN), .B1(n3141), .B2(n4392), .ZN(n3142) );
  OAI21_X1 U3886 ( .B1(n3206), .B2(n4088), .A(n3142), .ZN(n3143) );
  AOI21_X1 U3887 ( .B1(n3201), .B2(n4005), .A(n3143), .ZN(n3144) );
  OAI21_X1 U3888 ( .B1(n3145), .B2(n4281), .A(n3144), .ZN(U3282) );
  INV_X1 U3889 ( .A(n3146), .ZN(n3152) );
  INV_X1 U3890 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3148) );
  OAI22_X1 U3891 ( .A1(n4118), .A2(n3148), .B1(n3147), .B2(n4115), .ZN(n3151)
         );
  NOR2_X1 U3892 ( .A1(n3149), .A2(n4092), .ZN(n3150) );
  AOI211_X1 U3893 ( .C1(n3152), .C2(n4378), .A(n3151), .B(n3150), .ZN(n3153)
         );
  OAI21_X1 U3894 ( .B1(n4281), .B2(n3154), .A(n3153), .ZN(U3284) );
  OAI22_X1 U3895 ( .A1(n3182), .A2(n4388), .B1(n3160), .B2(n4059), .ZN(n3158)
         );
  XOR2_X1 U3896 ( .A(n3629), .B(n3155), .Z(n3156) );
  NOR2_X1 U3897 ( .A1(n3156), .A2(n4065), .ZN(n3157) );
  AOI211_X1 U3898 ( .C1(n4071), .C2(n3710), .A(n3158), .B(n3157), .ZN(n4449)
         );
  OAI211_X1 U3899 ( .C1(n3161), .C2(n3160), .A(n4443), .B(n3159), .ZN(n4448)
         );
  INV_X1 U3900 ( .A(n4448), .ZN(n3165) );
  INV_X1 U3901 ( .A(n3162), .ZN(n3163) );
  OAI22_X1 U3902 ( .A1(n4118), .A2(n4482), .B1(n3163), .B2(n4115), .ZN(n3164)
         );
  AOI21_X1 U3903 ( .B1(n3165), .B2(n4027), .A(n3164), .ZN(n3167) );
  NAND2_X1 U3904 ( .A1(n3217), .A2(n3629), .ZN(n4445) );
  NAND3_X1 U3905 ( .A1(n4446), .A2(n4445), .A3(n4005), .ZN(n3166) );
  OAI211_X1 U3906 ( .C1(n4449), .C2(n4281), .A(n3167), .B(n3166), .ZN(U3283)
         );
  XOR2_X1 U3907 ( .A(n3168), .B(n3169), .Z(n3174) );
  INV_X1 U3908 ( .A(n3706), .ZN(n3267) );
  OAI22_X1 U3909 ( .A1(n3182), .A2(n3519), .B1(n3518), .B2(n3267), .ZN(n3170)
         );
  AOI211_X1 U3910 ( .C1(n3218), .C2(n3521), .A(n3171), .B(n3170), .ZN(n3173)
         );
  NAND2_X1 U3911 ( .A1(n3522), .A2(n3196), .ZN(n3172) );
  OAI211_X1 U3912 ( .C1(n3174), .C2(n3525), .A(n3173), .B(n3172), .ZN(U3228)
         );
  NAND2_X1 U3913 ( .A1(n3176), .A2(n3631), .ZN(n3207) );
  INV_X1 U3914 ( .A(n3218), .ZN(n3213) );
  AND2_X1 U3915 ( .A1(n3707), .A2(n3213), .ZN(n3653) );
  INV_X1 U3916 ( .A(n3653), .ZN(n3177) );
  NAND2_X1 U3917 ( .A1(n3214), .A2(n3218), .ZN(n3634) );
  NAND2_X1 U3918 ( .A1(n3177), .A2(n3634), .ZN(n3576) );
  XNOR2_X1 U3919 ( .A(n3207), .B(n3576), .ZN(n3180) );
  AOI22_X1 U3920 ( .A1(n3706), .A2(n4101), .B1(n4135), .B2(n3218), .ZN(n3178)
         );
  OAI21_X1 U3921 ( .B1(n3182), .B2(n4104), .A(n3178), .ZN(n3179) );
  AOI21_X1 U3922 ( .B1(n3180), .B2(n4386), .A(n3179), .ZN(n4450) );
  AND2_X1 U3923 ( .A1(n3182), .A2(n3181), .ZN(n3190) );
  OR2_X1 U3924 ( .A1(n3217), .A2(n3215), .ZN(n3191) );
  INV_X1 U3925 ( .A(n3185), .ZN(n3186) );
  AOI21_X1 U3926 ( .B1(n3188), .B2(n3187), .A(n3186), .ZN(n3189) );
  NAND2_X1 U3927 ( .A1(n3191), .A2(n3219), .ZN(n3192) );
  XOR2_X1 U3928 ( .A(n3576), .B(n3192), .Z(n4454) );
  INV_X1 U3929 ( .A(n3224), .ZN(n3194) );
  OAI21_X1 U3930 ( .B1(n3195), .B2(n3213), .A(n3194), .ZN(n4451) );
  AOI22_X1 U3931 ( .A1(n4281), .A2(REG2_REG_9__SCAN_IN), .B1(n3196), .B2(n4392), .ZN(n3197) );
  OAI21_X1 U3932 ( .B1(n4451), .B2(n4088), .A(n3197), .ZN(n3198) );
  AOI21_X1 U3933 ( .B1(n4454), .B2(n4005), .A(n3198), .ZN(n3199) );
  OAI21_X1 U3934 ( .B1(n4281), .B2(n4450), .A(n3199), .ZN(U3281) );
  INV_X1 U3935 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3202) );
  AOI21_X1 U3936 ( .B1(n3201), .B2(n4453), .A(n3200), .ZN(n3204) );
  MUX2_X1 U3937 ( .A(n3202), .B(n3204), .S(n4463), .Z(n3203) );
  OAI21_X1 U3938 ( .B1(n3206), .B2(n4261), .A(n3203), .ZN(U3483) );
  MUX2_X1 U3939 ( .A(n2441), .B(n3204), .S(n4474), .Z(n3205) );
  OAI21_X1 U3940 ( .B1(n3206), .B2(n4206), .A(n3205), .ZN(U3526) );
  NAND2_X1 U3941 ( .A1(n3267), .A2(n3265), .ZN(n3652) );
  NAND2_X1 U3942 ( .A1(n3706), .A2(n3266), .ZN(n3649) );
  NAND2_X1 U3943 ( .A1(n3652), .A2(n3649), .ZN(n3577) );
  INV_X1 U3944 ( .A(n3577), .ZN(n3208) );
  XNOR2_X1 U3945 ( .A(n3264), .B(n3208), .ZN(n3212) );
  NAND2_X1 U3946 ( .A1(n3265), .A2(n4135), .ZN(n3210) );
  NAND2_X1 U3947 ( .A1(n3707), .A2(n4071), .ZN(n3209) );
  OAI211_X1 U3948 ( .C1(n3263), .C2(n4388), .A(n3210), .B(n3209), .ZN(n3211)
         );
  AOI21_X1 U3949 ( .B1(n3212), .B2(n4386), .A(n3211), .ZN(n3248) );
  AND2_X1 U3950 ( .A1(n3214), .A2(n3213), .ZN(n3221) );
  NOR2_X1 U3951 ( .A1(n3217), .A2(n3216), .ZN(n3223) );
  AND2_X1 U3952 ( .A1(n2274), .A2(n3219), .ZN(n3220) );
  NOR2_X1 U3953 ( .A1(n3221), .A2(n3220), .ZN(n3222) );
  XNOR2_X1 U3954 ( .A(n3269), .B(n3577), .ZN(n3246) );
  NOR2_X1 U3955 ( .A1(n3224), .A2(n3266), .ZN(n3225) );
  OR2_X1 U3956 ( .A1(n3278), .A2(n3225), .ZN(n3253) );
  AOI22_X1 U3957 ( .A1(n4281), .A2(REG2_REG_10__SCAN_IN), .B1(n3244), .B2(
        n4392), .ZN(n3226) );
  OAI21_X1 U3958 ( .B1(n3253), .B2(n4088), .A(n3226), .ZN(n3227) );
  AOI21_X1 U3959 ( .B1(n3246), .B2(n4005), .A(n3227), .ZN(n3228) );
  OAI21_X1 U3960 ( .B1(n3248), .B2(n4281), .A(n3228), .ZN(U3280) );
  XOR2_X1 U3961 ( .A(n3230), .B(n3229), .Z(n3231) );
  XNOR2_X1 U3962 ( .A(n3232), .B(n3231), .ZN(n3237) );
  INV_X1 U3963 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3233) );
  NOR2_X1 U3964 ( .A1(STATE_REG_SCAN_IN), .A2(n3233), .ZN(n4297) );
  OAI22_X1 U3965 ( .A1(n4105), .A2(n3518), .B1(n3519), .B2(n3267), .ZN(n3234)
         );
  AOI211_X1 U3966 ( .C1(n3284), .C2(n3521), .A(n4297), .B(n3234), .ZN(n3236)
         );
  NAND2_X1 U3967 ( .A1(n3522), .A2(n3279), .ZN(n3235) );
  OAI211_X1 U3968 ( .C1(n3237), .C2(n3525), .A(n3236), .B(n3235), .ZN(U3233)
         );
  AOI22_X1 U3969 ( .A1(n3417), .A2(n3707), .B1(n3419), .B2(n3705), .ZN(n3238)
         );
  NAND2_X1 U3970 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4288) );
  OAI211_X1 U3971 ( .C1(n2792), .C2(n3266), .A(n3238), .B(n4288), .ZN(n3243)
         );
  AOI211_X1 U3972 ( .C1(n3241), .C2(n3239), .A(n3525), .B(n2260), .ZN(n3242)
         );
  AOI211_X1 U3973 ( .C1(n3244), .C2(n3522), .A(n3243), .B(n3242), .ZN(n3245)
         );
  INV_X1 U3974 ( .A(n3245), .ZN(U3214) );
  NAND2_X1 U3975 ( .A1(n3246), .A2(n4453), .ZN(n3247) );
  AND2_X1 U3976 ( .A1(n3248), .A2(n3247), .ZN(n3251) );
  INV_X1 U3977 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4287) );
  MUX2_X1 U3978 ( .A(n3251), .B(n4287), .S(n4472), .Z(n3249) );
  OAI21_X1 U3979 ( .B1(n3253), .B2(n4206), .A(n3249), .ZN(U3528) );
  INV_X1 U3980 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3250) );
  MUX2_X1 U3981 ( .A(n3251), .B(n3250), .S(n4461), .Z(n3252) );
  OAI21_X1 U3982 ( .B1(n3253), .B2(n4261), .A(n3252), .ZN(U3487) );
  INV_X1 U3983 ( .A(n3255), .ZN(n3257) );
  NOR2_X1 U3984 ( .A1(n3257), .A2(n3256), .ZN(n3258) );
  XNOR2_X1 U3985 ( .A(n3254), .B(n3258), .ZN(n3262) );
  OAI22_X1 U3986 ( .A1(n3263), .A2(n3519), .B1(n3518), .B2(n3384), .ZN(n3260)
         );
  NAND2_X1 U3987 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4306) );
  OAI21_X1 U3988 ( .B1(n2792), .B2(n3309), .A(n4306), .ZN(n3259) );
  AOI211_X1 U3989 ( .C1(n3315), .C2(n3522), .A(n3260), .B(n3259), .ZN(n3261)
         );
  OAI21_X1 U3990 ( .B1(n3262), .B2(n3525), .A(n3261), .ZN(U3221) );
  NAND2_X1 U3991 ( .A1(n3263), .A2(n3284), .ZN(n3305) );
  NAND2_X1 U3992 ( .A1(n3705), .A2(n3277), .ZN(n3307) );
  XOR2_X1 U3993 ( .A(n3599), .B(n3308), .Z(n3275) );
  OAI22_X1 U3994 ( .A1(n4105), .A2(n4388), .B1(n3277), .B2(n4059), .ZN(n3273)
         );
  NOR2_X1 U3995 ( .A1(n3706), .A2(n3265), .ZN(n3268) );
  NAND2_X1 U3996 ( .A1(n3270), .A2(n3599), .ZN(n3271) );
  AND2_X1 U3997 ( .A1(n3286), .A2(n3271), .ZN(n3276) );
  NOR2_X1 U3998 ( .A1(n3276), .A2(n4109), .ZN(n3272) );
  AOI211_X1 U3999 ( .C1(n4071), .C2(n3706), .A(n3273), .B(n3272), .ZN(n3274)
         );
  OAI21_X1 U4000 ( .B1(n4065), .B2(n3275), .A(n3274), .ZN(n4457) );
  INV_X1 U4001 ( .A(n4457), .ZN(n3283) );
  INV_X1 U4002 ( .A(n3276), .ZN(n4459) );
  OAI21_X1 U4003 ( .B1(n3278), .B2(n3277), .A(n3313), .ZN(n4456) );
  AOI22_X1 U4004 ( .A1(n4281), .A2(REG2_REG_11__SCAN_IN), .B1(n3279), .B2(
        n4392), .ZN(n3280) );
  OAI21_X1 U4005 ( .B1(n4456), .B2(n4088), .A(n3280), .ZN(n3281) );
  AOI21_X1 U4006 ( .B1(n4459), .B2(n4393), .A(n3281), .ZN(n3282) );
  OAI21_X1 U4007 ( .B1(n3283), .B2(n4281), .A(n3282), .ZN(U3279) );
  AOI21_X1 U4008 ( .B1(n3384), .B2(n4112), .A(n4093), .ZN(n3289) );
  NAND2_X1 U4009 ( .A1(n4083), .A2(n3331), .ZN(n3547) );
  NAND2_X1 U4010 ( .A1(n4102), .A2(n3385), .ZN(n3543) );
  NAND2_X1 U4011 ( .A1(n3547), .A2(n3543), .ZN(n3352) );
  NAND2_X1 U4012 ( .A1(n3290), .A2(n3352), .ZN(n3330) );
  OAI21_X1 U4013 ( .B1(n3290), .B2(n3352), .A(n3330), .ZN(n4196) );
  INV_X1 U4014 ( .A(n4196), .ZN(n3303) );
  NAND2_X1 U4015 ( .A1(n3288), .A2(n3309), .ZN(n4094) );
  NAND2_X1 U4016 ( .A1(n3704), .A2(n4112), .ZN(n3571) );
  NAND2_X1 U4017 ( .A1(n4094), .A2(n3571), .ZN(n3292) );
  INV_X1 U4018 ( .A(n3307), .ZN(n3650) );
  NOR2_X1 U4019 ( .A1(n3292), .A2(n3650), .ZN(n3291) );
  NAND2_X1 U4020 ( .A1(n3308), .A2(n3291), .ZN(n3294) );
  NAND2_X1 U4021 ( .A1(n4105), .A2(n3287), .ZN(n4096) );
  NAND2_X1 U4022 ( .A1(n3305), .A2(n4096), .ZN(n3293) );
  INV_X1 U4023 ( .A(n3292), .ZN(n3655) );
  NOR2_X1 U4024 ( .A1(n3704), .A2(n4112), .ZN(n3572) );
  AOI21_X1 U4025 ( .B1(n3293), .B2(n3655), .A(n3572), .ZN(n3661) );
  NAND2_X1 U4026 ( .A1(n3294), .A2(n3661), .ZN(n3548) );
  XNOR2_X1 U4027 ( .A(n3548), .B(n3352), .ZN(n3297) );
  OAI22_X1 U4028 ( .A1(n3452), .A2(n4388), .B1(n3385), .B2(n4059), .ZN(n3295)
         );
  AOI21_X1 U4029 ( .B1(n4071), .B2(n3704), .A(n3295), .ZN(n3296) );
  OAI21_X1 U4030 ( .B1(n3297), .B2(n4065), .A(n3296), .ZN(n4195) );
  INV_X1 U4031 ( .A(n4111), .ZN(n3299) );
  INV_X1 U4032 ( .A(n4085), .ZN(n3298) );
  OAI21_X1 U4033 ( .B1(n3299), .B2(n3385), .A(n3298), .ZN(n4253) );
  AOI22_X1 U4034 ( .A1(n4281), .A2(REG2_REG_14__SCAN_IN), .B1(n3388), .B2(
        n4392), .ZN(n3300) );
  OAI21_X1 U4035 ( .B1(n4253), .B2(n4088), .A(n3300), .ZN(n3301) );
  AOI21_X1 U4036 ( .B1(n4195), .B2(n4118), .A(n3301), .ZN(n3302) );
  OAI21_X1 U4037 ( .B1(n3303), .B2(n4092), .A(n3302), .ZN(U3276) );
  NAND2_X1 U4038 ( .A1(n4096), .A2(n4094), .ZN(n3578) );
  XNOR2_X1 U4039 ( .A(n3304), .B(n3578), .ZN(n4204) );
  INV_X1 U4040 ( .A(n4204), .ZN(n3319) );
  INV_X1 U4041 ( .A(n3305), .ZN(n3306) );
  AOI21_X1 U4042 ( .B1(n3308), .B2(n3307), .A(n3306), .ZN(n4097) );
  XOR2_X1 U40430 ( .A(n3578), .B(n4097), .Z(n3312) );
  OAI22_X1 U4044 ( .A1(n3384), .A2(n4388), .B1(n4059), .B2(n3309), .ZN(n3310)
         );
  AOI21_X1 U4045 ( .B1(n4071), .B2(n3705), .A(n3310), .ZN(n3311) );
  OAI21_X1 U4046 ( .B1(n3312), .B2(n4065), .A(n3311), .ZN(n4203) );
  NAND2_X1 U4047 ( .A1(n3313), .A2(n3287), .ZN(n3314) );
  NAND2_X1 U4048 ( .A1(n4110), .A2(n3314), .ZN(n4262) );
  AOI22_X1 U4049 ( .A1(n4281), .A2(REG2_REG_12__SCAN_IN), .B1(n3315), .B2(
        n4392), .ZN(n3316) );
  OAI21_X1 U4050 ( .B1(n4262), .B2(n4088), .A(n3316), .ZN(n3317) );
  AOI21_X1 U4051 ( .B1(n4203), .B2(n4118), .A(n3317), .ZN(n3318) );
  OAI21_X1 U4052 ( .B1(n3319), .B2(n4092), .A(n3318), .ZN(U3278) );
  XOR2_X1 U4053 ( .A(n3322), .B(n3321), .Z(n3323) );
  XNOR2_X1 U4054 ( .A(n3320), .B(n3323), .ZN(n3328) );
  NOR2_X1 U4055 ( .A1(STATE_REG_SCAN_IN), .A2(n3324), .ZN(n4317) );
  OAI22_X1 U4056 ( .A1(n4105), .A2(n3519), .B1(n3518), .B2(n4083), .ZN(n3325)
         );
  AOI211_X1 U4057 ( .C1(n4100), .C2(n3521), .A(n4317), .B(n3325), .ZN(n3327)
         );
  NAND2_X1 U4058 ( .A1(n3522), .A2(n4114), .ZN(n3326) );
  OAI211_X1 U4059 ( .C1(n3328), .C2(n3525), .A(n3327), .B(n3326), .ZN(U3231)
         );
  INV_X1 U4060 ( .A(n3850), .ZN(n3329) );
  OAI21_X1 U4061 ( .B1(n3329), .B2(n3821), .A(n3827), .ZN(n3835) );
  OR2_X1 U4062 ( .A1(n3835), .A2(n4206), .ZN(n3369) );
  NAND2_X1 U4063 ( .A1(n4070), .A2(n4084), .ZN(n3332) );
  NAND2_X1 U4064 ( .A1(n3517), .A2(n4055), .ZN(n3545) );
  INV_X1 U4065 ( .A(n3517), .ZN(n4080) );
  NAND2_X1 U4066 ( .A1(n4080), .A2(n4060), .ZN(n4035) );
  NAND2_X1 U4067 ( .A1(n3545), .A2(n4035), .ZN(n4066) );
  NAND2_X1 U4068 ( .A1(n4061), .A2(n4045), .ZN(n3334) );
  INV_X1 U4069 ( .A(n4061), .ZN(n3703) );
  NAND2_X1 U4070 ( .A1(n4038), .A2(n4025), .ZN(n3995) );
  NAND2_X1 U4071 ( .A1(n3702), .A2(n3335), .ZN(n3996) );
  NAND2_X1 U4072 ( .A1(n3995), .A2(n3996), .ZN(n4016) );
  NAND2_X1 U4073 ( .A1(n4017), .A2(n4016), .ZN(n4015) );
  NAND2_X1 U4074 ( .A1(n4021), .A2(n3411), .ZN(n3338) );
  NOR2_X1 U4075 ( .A1(n4021), .A2(n3411), .ZN(n3337) );
  INV_X1 U4076 ( .A(n3999), .ZN(n3961) );
  NOR2_X1 U4077 ( .A1(n3975), .A2(n3966), .ZN(n3340) );
  NAND2_X1 U4078 ( .A1(n3431), .A2(n3951), .ZN(n3921) );
  NAND2_X1 U4079 ( .A1(n3960), .A2(n3491), .ZN(n3361) );
  NAND2_X1 U4080 ( .A1(n3960), .A2(n3951), .ZN(n3341) );
  NOR2_X1 U4081 ( .A1(n3924), .A2(n3903), .ZN(n3878) );
  AND2_X1 U4082 ( .A1(n3905), .A2(n3342), .ZN(n3345) );
  OR2_X1 U4083 ( .A1(n3878), .A2(n3345), .ZN(n3347) );
  OR2_X1 U4084 ( .A1(n3905), .A2(n3342), .ZN(n3343) );
  NAND2_X1 U4085 ( .A1(n3924), .A2(n3903), .ZN(n3879) );
  AND2_X1 U4086 ( .A1(n3343), .A2(n3879), .ZN(n3344) );
  NAND2_X1 U4087 ( .A1(n3887), .A2(n3864), .ZN(n3349) );
  NOR2_X1 U4088 ( .A1(n3887), .A2(n3864), .ZN(n3348) );
  NAND2_X1 U4089 ( .A1(n3867), .A2(n3851), .ZN(n3350) );
  NOR2_X1 U4090 ( .A1(n3822), .A2(n3351), .ZN(n3811) );
  XNOR2_X1 U4091 ( .A(n3825), .B(n3820), .ZN(n3832) );
  INV_X1 U4092 ( .A(n3352), .ZN(n3590) );
  NAND2_X1 U4093 ( .A1(n3548), .A2(n3590), .ZN(n3353) );
  NAND2_X1 U4094 ( .A1(n3353), .A2(n3547), .ZN(n4076) );
  NAND2_X1 U4095 ( .A1(n3452), .A2(n4084), .ZN(n3546) );
  NAND2_X1 U4096 ( .A1(n4070), .A2(n3354), .ZN(n3544) );
  NAND2_X1 U4097 ( .A1(n3546), .A2(n3544), .ZN(n3606) );
  INV_X1 U4098 ( .A(n4066), .ZN(n3600) );
  NAND2_X1 U4099 ( .A1(n3703), .A2(n4045), .ZN(n3664) );
  AND2_X1 U4100 ( .A1(n4035), .A2(n3664), .ZN(n3549) );
  NAND2_X1 U4101 ( .A1(n4061), .A2(n3462), .ZN(n3993) );
  NAND2_X1 U4102 ( .A1(n3995), .A2(n3993), .ZN(n3355) );
  NAND2_X1 U4103 ( .A1(n4021), .A2(n4007), .ZN(n3568) );
  AND2_X1 U4104 ( .A1(n3996), .A2(n3568), .ZN(n3357) );
  NOR2_X1 U4105 ( .A1(n4021), .A2(n4007), .ZN(n3569) );
  AOI21_X1 U4106 ( .B1(n3355), .B2(n3357), .A(n3569), .ZN(n3976) );
  NAND2_X1 U4107 ( .A1(n3999), .A2(n3984), .ZN(n3356) );
  NAND2_X1 U4108 ( .A1(n3994), .A2(n3665), .ZN(n3359) );
  INV_X1 U4109 ( .A(n3357), .ZN(n3977) );
  AND2_X1 U4110 ( .A1(n3961), .A2(n3974), .ZN(n3358) );
  AOI21_X1 U4111 ( .B1(n3665), .B2(n3977), .A(n3358), .ZN(n3669) );
  INV_X1 U4112 ( .A(n3921), .ZN(n3360) );
  NOR2_X1 U4113 ( .A1(n3942), .A2(n3966), .ZN(n3918) );
  NOR2_X1 U4114 ( .A1(n3360), .A2(n3918), .ZN(n3672) );
  OR2_X1 U4115 ( .A1(n3945), .A2(n3363), .ZN(n3586) );
  AND2_X1 U4116 ( .A1(n3586), .A2(n3361), .ZN(n3676) );
  AND2_X1 U4117 ( .A1(n3942), .A2(n3966), .ZN(n3917) );
  NAND2_X1 U4118 ( .A1(n3921), .A2(n3917), .ZN(n3362) );
  NAND2_X1 U4119 ( .A1(n3676), .A2(n3362), .ZN(n3553) );
  OR2_X1 U4120 ( .A1(n3700), .A2(n3903), .ZN(n3585) );
  NAND2_X1 U4121 ( .A1(n3945), .A2(n3363), .ZN(n3898) );
  NAND2_X1 U4122 ( .A1(n3585), .A2(n3898), .ZN(n3674) );
  OR2_X1 U4123 ( .A1(n3887), .A2(n3870), .ZN(n3597) );
  OR2_X1 U4124 ( .A1(n3905), .A2(n3891), .ZN(n3858) );
  NAND2_X1 U4125 ( .A1(n3597), .A2(n3858), .ZN(n3673) );
  NAND2_X1 U4126 ( .A1(n3905), .A2(n3891), .ZN(n3566) );
  NAND2_X1 U4127 ( .A1(n3700), .A2(n3903), .ZN(n3882) );
  AND2_X1 U4128 ( .A1(n3566), .A2(n3882), .ZN(n3860) );
  NAND2_X1 U4129 ( .A1(n3887), .A2(n3870), .ZN(n3598) );
  OAI21_X1 U4130 ( .B1(n3673), .B2(n3860), .A(n3598), .ZN(n3678) );
  INV_X1 U4131 ( .A(n3678), .ZN(n3364) );
  XNOR2_X1 U4132 ( .A(n3699), .B(n3613), .ZN(n3840) );
  INV_X1 U4133 ( .A(n3840), .ZN(n3845) );
  NOR2_X1 U4134 ( .A1(n3699), .A2(n3851), .ZN(n3542) );
  NOR2_X2 U4135 ( .A1(n3843), .A2(n3542), .ZN(n3812) );
  XOR2_X1 U4136 ( .A(n3820), .B(n3812), .Z(n3367) );
  OAI22_X1 U4137 ( .A1(n3596), .A2(n4388), .B1(n4059), .B2(n3821), .ZN(n3365)
         );
  AOI21_X1 U4138 ( .B1(n4071), .B2(n3699), .A(n3365), .ZN(n3366) );
  OAI21_X1 U4139 ( .B1(n3367), .B2(n4065), .A(n3366), .ZN(n3837) );
  AOI21_X1 U4140 ( .B1(n3832), .B2(n4453), .A(n3837), .ZN(n3370) );
  MUX2_X1 U4141 ( .A(n4546), .B(n3370), .S(n4474), .Z(n3368) );
  NAND2_X1 U4142 ( .A1(n3369), .A2(n3368), .ZN(U3546) );
  INV_X1 U4143 ( .A(REG0_REG_28__SCAN_IN), .ZN(n3371) );
  MUX2_X1 U4144 ( .A(n3371), .B(n3370), .S(n4463), .Z(n3372) );
  OAI21_X1 U4145 ( .B1(n3835), .B2(n4261), .A(n3372), .ZN(U3514) );
  XNOR2_X1 U4146 ( .A(n3374), .B(n3373), .ZN(n3379) );
  INV_X1 U4147 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3375) );
  OAI22_X1 U4148 ( .A1(n2792), .A2(n3851), .B1(STATE_REG_SCAN_IN), .B2(n3375), 
        .ZN(n3377) );
  INV_X1 U4149 ( .A(n3887), .ZN(n3842) );
  OAI22_X1 U4150 ( .A1(n3822), .A2(n3518), .B1(n3842), .B2(n3519), .ZN(n3376)
         );
  AOI211_X1 U4151 ( .C1(n3852), .C2(n3522), .A(n3377), .B(n3376), .ZN(n3378)
         );
  OAI21_X1 U4152 ( .B1(n3379), .B2(n3525), .A(n3378), .ZN(U3211) );
  NOR2_X1 U4153 ( .A1(n2147), .A2(n3382), .ZN(n3383) );
  XNOR2_X1 U4154 ( .A(n3380), .B(n3383), .ZN(n3390) );
  OAI22_X1 U4155 ( .A1(n3452), .A2(n3518), .B1(n3519), .B2(n3384), .ZN(n3387)
         );
  NAND2_X1 U4156 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4336) );
  OAI21_X1 U4157 ( .B1(n2792), .B2(n3385), .A(n4336), .ZN(n3386) );
  AOI211_X1 U4158 ( .C1(n3388), .C2(n3522), .A(n3387), .B(n3386), .ZN(n3389)
         );
  OAI21_X1 U4159 ( .B1(n3390), .B2(n3525), .A(n3389), .ZN(U3212) );
  NAND2_X1 U4160 ( .A1(n3391), .A2(n3428), .ZN(n3399) );
  AOI21_X1 U4161 ( .B1(n3392), .B2(n3394), .A(n3393), .ZN(n3398) );
  OAI22_X1 U4162 ( .A1(n3924), .A2(n3518), .B1(n3519), .B2(n3431), .ZN(n3396)
         );
  OAI22_X1 U4163 ( .A1(n2792), .A2(n3928), .B1(STATE_REG_SCAN_IN), .B2(n4633), 
        .ZN(n3395) );
  AOI211_X1 U4164 ( .C1(n3931), .C2(n3522), .A(n3396), .B(n3395), .ZN(n3397)
         );
  OAI21_X1 U4165 ( .B1(n3399), .B2(n3398), .A(n3397), .ZN(U3213) );
  INV_X1 U4166 ( .A(n3400), .ZN(n3404) );
  AOI21_X1 U4167 ( .B1(n3400), .B2(n3402), .A(n3401), .ZN(n3403) );
  AOI21_X1 U4168 ( .B1(n3404), .B2(n3496), .A(n3403), .ZN(n3408) );
  NAND2_X1 U4169 ( .A1(n3406), .A2(n3405), .ZN(n3407) );
  XNOR2_X1 U4170 ( .A(n3408), .B(n3407), .ZN(n3414) );
  NOR2_X1 U4171 ( .A1(STATE_REG_SCAN_IN), .A2(n3409), .ZN(n3805) );
  OAI22_X1 U4172 ( .A1(n4038), .A2(n3519), .B1(n3518), .B2(n3999), .ZN(n3410)
         );
  AOI211_X1 U4173 ( .C1(n3411), .C2(n3521), .A(n3805), .B(n3410), .ZN(n3413)
         );
  NAND2_X1 U4174 ( .A1(n3522), .A2(n4009), .ZN(n3412) );
  OAI211_X1 U4175 ( .C1(n3414), .C2(n3525), .A(n3413), .B(n3412), .ZN(U3216)
         );
  OAI211_X1 U4176 ( .C1(n3416), .C2(n3415), .A(n2931), .B(n3428), .ZN(n3423)
         );
  AOI22_X1 U4177 ( .A1(n3521), .A2(n3418), .B1(n3417), .B2(n2975), .ZN(n3422)
         );
  AOI22_X1 U4178 ( .A1(REG3_REG_1__SCAN_IN), .A2(n3420), .B1(n3419), .B2(n3713), .ZN(n3421) );
  NAND3_X1 U4179 ( .A1(n3423), .A2(n3422), .A3(n3421), .ZN(U3219) );
  NAND2_X1 U4180 ( .A1(n2089), .A2(n3424), .ZN(n3429) );
  INV_X1 U4181 ( .A(n3479), .ZN(n3426) );
  OAI211_X1 U4182 ( .C1(n3425), .C2(n3426), .A(n3477), .B(n3429), .ZN(n3427)
         );
  OAI211_X1 U4183 ( .C1(n3430), .C2(n3429), .A(n3428), .B(n3427), .ZN(n3436)
         );
  OAI22_X1 U4184 ( .A1(n3999), .A2(n3519), .B1(n3518), .B2(n3431), .ZN(n3434)
         );
  OAI22_X1 U4185 ( .A1(n2792), .A2(n3966), .B1(STATE_REG_SCAN_IN), .B2(n3432), 
        .ZN(n3433) );
  AOI211_X1 U4186 ( .C1(n3968), .C2(n3522), .A(n3434), .B(n3433), .ZN(n3435)
         );
  NAND2_X1 U4187 ( .A1(n3436), .A2(n3435), .ZN(U3220) );
  NAND2_X1 U4188 ( .A1(n3438), .A2(n3437), .ZN(n3440) );
  XOR2_X1 U4189 ( .A(n3440), .B(n3439), .Z(n3446) );
  INV_X1 U4190 ( .A(n3441), .ZN(n3893) );
  INV_X1 U4191 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3442) );
  OAI22_X1 U4192 ( .A1(n2792), .A2(n3891), .B1(STATE_REG_SCAN_IN), .B2(n3442), 
        .ZN(n3444) );
  OAI22_X1 U4193 ( .A1(n3842), .A2(n3518), .B1(n3924), .B2(n3519), .ZN(n3443)
         );
  AOI211_X1 U4194 ( .C1(n3893), .C2(n3522), .A(n3444), .B(n3443), .ZN(n3445)
         );
  OAI21_X1 U4195 ( .B1(n3446), .B2(n3525), .A(n3445), .ZN(U3222) );
  INV_X1 U4196 ( .A(n3447), .ZN(n3449) );
  OAI21_X1 U4197 ( .B1(n3449), .B2(n3515), .A(n3448), .ZN(n3450) );
  XOR2_X1 U4198 ( .A(n3451), .B(n3450), .Z(n3456) );
  OAI22_X1 U4199 ( .A1(n4061), .A2(n3518), .B1(n3519), .B2(n3452), .ZN(n3454)
         );
  NAND2_X1 U4200 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4349) );
  OAI21_X1 U4201 ( .B1(n2792), .B2(n4060), .A(n4349), .ZN(n3453) );
  AOI211_X1 U4202 ( .C1(n4056), .C2(n3522), .A(n3454), .B(n3453), .ZN(n3455)
         );
  OAI21_X1 U4203 ( .B1(n3456), .B2(n3525), .A(n3455), .ZN(U3223) );
  NAND2_X1 U4204 ( .A1(n3459), .A2(n3458), .ZN(n3460) );
  XNOR2_X1 U4205 ( .A(n3457), .B(n3460), .ZN(n3465) );
  AND2_X1 U4206 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n3775) );
  OAI22_X1 U4207 ( .A1(n3517), .A2(n3519), .B1(n3518), .B2(n4038), .ZN(n3461)
         );
  AOI211_X1 U4208 ( .C1(n3462), .C2(n3521), .A(n3775), .B(n3461), .ZN(n3464)
         );
  NAND2_X1 U4209 ( .A1(n3522), .A2(n4046), .ZN(n3463) );
  OAI211_X1 U4210 ( .C1(n3465), .C2(n3525), .A(n3464), .B(n3463), .ZN(U3225)
         );
  NAND2_X1 U4211 ( .A1(n3466), .A2(n3467), .ZN(n3468) );
  XOR2_X1 U4212 ( .A(n3469), .B(n3468), .Z(n3475) );
  INV_X1 U4213 ( .A(n3470), .ZN(n3911) );
  OAI22_X1 U4214 ( .A1(n2792), .A2(n3903), .B1(STATE_REG_SCAN_IN), .B2(n3471), 
        .ZN(n3473) );
  INV_X1 U4215 ( .A(n3905), .ZN(n3509) );
  OAI22_X1 U4216 ( .A1(n3509), .A2(n3518), .B1(n3945), .B2(n3519), .ZN(n3472)
         );
  AOI211_X1 U4217 ( .C1(n3911), .C2(n3522), .A(n3473), .B(n3472), .ZN(n3474)
         );
  OAI21_X1 U4218 ( .B1(n3475), .B2(n3525), .A(n3474), .ZN(U3226) );
  INV_X1 U4219 ( .A(n3476), .ZN(n3480) );
  AOI21_X1 U4220 ( .B1(n3477), .B2(n3479), .A(n3425), .ZN(n3478) );
  AOI21_X1 U4221 ( .B1(n3480), .B2(n3479), .A(n3478), .ZN(n3486) );
  INV_X1 U4222 ( .A(n4021), .ZN(n3499) );
  OAI22_X1 U4223 ( .A1(n3499), .A2(n3519), .B1(n3518), .B2(n3975), .ZN(n3483)
         );
  OAI22_X1 U4224 ( .A1(n2792), .A2(n3974), .B1(STATE_REG_SCAN_IN), .B2(n3481), 
        .ZN(n3482) );
  AOI211_X1 U4225 ( .C1(n3484), .C2(n3522), .A(n3483), .B(n3482), .ZN(n3485)
         );
  OAI21_X1 U4226 ( .B1(n3486), .B2(n3525), .A(n3485), .ZN(U3230) );
  INV_X1 U4227 ( .A(n3392), .ZN(n3487) );
  AOI21_X1 U4228 ( .B1(n3489), .B2(n3488), .A(n3487), .ZN(n3495) );
  OAI22_X1 U4229 ( .A1(n3945), .A2(n3518), .B1(n3519), .B2(n3975), .ZN(n3493)
         );
  INV_X1 U4230 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3490) );
  OAI22_X1 U4231 ( .A1(n2792), .A2(n3491), .B1(STATE_REG_SCAN_IN), .B2(n3490), 
        .ZN(n3492) );
  AOI211_X1 U4232 ( .C1(n3948), .C2(n3522), .A(n3493), .B(n3492), .ZN(n3494)
         );
  OAI21_X1 U4233 ( .B1(n3495), .B2(n3525), .A(n3494), .ZN(U3232) );
  XNOR2_X1 U4234 ( .A(n3497), .B(n3496), .ZN(n3498) );
  XNOR2_X1 U4235 ( .A(n3400), .B(n3498), .ZN(n3503) );
  AND2_X1 U4236 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4365) );
  OAI22_X1 U4237 ( .A1(n3499), .A2(n3518), .B1(n3519), .B2(n4061), .ZN(n3500)
         );
  AOI211_X1 U4238 ( .C1(n4025), .C2(n3521), .A(n4365), .B(n3500), .ZN(n3502)
         );
  NAND2_X1 U4239 ( .A1(n3522), .A2(n4028), .ZN(n3501) );
  OAI211_X1 U4240 ( .C1(n3503), .C2(n3525), .A(n3502), .B(n3501), .ZN(U3235)
         );
  NOR2_X1 U4241 ( .A1(n2233), .A2(n3505), .ZN(n3506) );
  INV_X1 U4242 ( .A(n3507), .ZN(n3872) );
  INV_X1 U4243 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3508) );
  OAI22_X1 U4244 ( .A1(n2792), .A2(n3870), .B1(STATE_REG_SCAN_IN), .B2(n3508), 
        .ZN(n3511) );
  OAI22_X1 U4245 ( .A1(n3867), .A2(n3518), .B1(n3509), .B2(n3519), .ZN(n3510)
         );
  AOI211_X1 U4246 ( .C1(n3872), .C2(n3522), .A(n3511), .B(n3510), .ZN(n3512)
         );
  OAI21_X1 U4247 ( .B1(n3513), .B2(n3525), .A(n3512), .ZN(U3237) );
  NAND2_X1 U4248 ( .A1(n3447), .A2(n3448), .ZN(n3514) );
  XOR2_X1 U4249 ( .A(n3515), .B(n3514), .Z(n3526) );
  NOR2_X1 U4250 ( .A1(STATE_REG_SCAN_IN), .A2(n3516), .ZN(n4342) );
  OAI22_X1 U4251 ( .A1(n4083), .A2(n3519), .B1(n3518), .B2(n3517), .ZN(n3520)
         );
  AOI211_X1 U4252 ( .C1(n4084), .C2(n3521), .A(n4342), .B(n3520), .ZN(n3524)
         );
  NAND2_X1 U4253 ( .A1(n3522), .A2(n4086), .ZN(n3523) );
  OAI211_X1 U4254 ( .C1(n3526), .C2(n3525), .A(n3524), .B(n3523), .ZN(U3238)
         );
  NAND2_X1 U4255 ( .A1(n2433), .A2(DATAI_29_), .ZN(n3595) );
  NOR2_X1 U4256 ( .A1(n3596), .A2(n3828), .ZN(n3527) );
  OR2_X1 U4257 ( .A1(n3811), .A2(n3527), .ZN(n3677) );
  INV_X1 U4258 ( .A(n3677), .ZN(n3540) );
  OR2_X1 U4259 ( .A1(n3809), .A2(n3542), .ZN(n3539) );
  INV_X1 U4260 ( .A(n3596), .ZN(n3698) );
  INV_X1 U4261 ( .A(REG1_REG_30__SCAN_IN), .ZN(n3530) );
  NAND2_X1 U4262 ( .A1(n3531), .A2(REG2_REG_30__SCAN_IN), .ZN(n3529) );
  NAND2_X1 U4263 ( .A1(n2053), .A2(REG0_REG_30__SCAN_IN), .ZN(n3528) );
  OAI211_X1 U4264 ( .C1(n3533), .C2(n3530), .A(n3529), .B(n3528), .ZN(n3816)
         );
  NAND2_X1 U4265 ( .A1(n2433), .A2(DATAI_30_), .ZN(n4124) );
  OR2_X1 U4266 ( .A1(n3816), .A2(n4124), .ZN(n3538) );
  NAND2_X1 U4267 ( .A1(n3531), .A2(REG2_REG_31__SCAN_IN), .ZN(n3536) );
  NAND2_X1 U4268 ( .A1(n2055), .A2(REG0_REG_31__SCAN_IN), .ZN(n3535) );
  INV_X1 U4269 ( .A(REG1_REG_31__SCAN_IN), .ZN(n3532) );
  OR2_X1 U4270 ( .A1(n3533), .A2(n3532), .ZN(n3534) );
  INV_X1 U4271 ( .A(n3561), .ZN(n4127) );
  NAND2_X1 U4272 ( .A1(n2433), .A2(DATAI_31_), .ZN(n4125) );
  AND2_X1 U4273 ( .A1(n4127), .A2(n4125), .ZN(n3682) );
  INV_X1 U4274 ( .A(n3682), .ZN(n3537) );
  AND2_X1 U4275 ( .A1(n3538), .A2(n3537), .ZN(n3581) );
  OAI21_X1 U4276 ( .B1(n3698), .B2(n3595), .A(n3581), .ZN(n3541) );
  AOI21_X1 U4277 ( .B1(n3540), .B2(n3539), .A(n3541), .ZN(n3681) );
  NAND3_X1 U4278 ( .A1(n3840), .A2(n3540), .A3(n3598), .ZN(n3558) );
  NOR4_X1 U4279 ( .A1(n3809), .A2(n3542), .A3(n3673), .A4(n3541), .ZN(n3557)
         );
  NAND2_X1 U4280 ( .A1(n3544), .A2(n3543), .ZN(n3647) );
  AND2_X1 U4281 ( .A1(n3647), .A2(n3546), .ZN(n3660) );
  INV_X1 U4282 ( .A(n3660), .ZN(n3643) );
  INV_X1 U4283 ( .A(n3545), .ZN(n3662) );
  AOI21_X1 U4284 ( .B1(n3547), .B2(n3546), .A(n3660), .ZN(n3657) );
  AOI211_X1 U4285 ( .C1(n3548), .C2(n3643), .A(n3662), .B(n3657), .ZN(n3551)
         );
  INV_X1 U4286 ( .A(n3549), .ZN(n3550) );
  OAI21_X1 U4287 ( .B1(n3551), .B2(n3550), .A(n3665), .ZN(n3552) );
  NAND2_X1 U4288 ( .A1(n3552), .A2(n3669), .ZN(n3554) );
  AOI21_X1 U4289 ( .B1(n3672), .B2(n3554), .A(n3553), .ZN(n3555) );
  OAI21_X1 U4290 ( .B1(n3555), .B2(n3674), .A(n3860), .ZN(n3556) );
  AOI22_X1 U4291 ( .A1(n3681), .A2(n3558), .B1(n3557), .B2(n3556), .ZN(n3565)
         );
  NOR2_X1 U4292 ( .A1(n4127), .A2(n4124), .ZN(n3564) );
  INV_X1 U4293 ( .A(n3559), .ZN(n3563) );
  INV_X1 U4294 ( .A(n3816), .ZN(n3560) );
  INV_X1 U4295 ( .A(n4124), .ZN(n4136) );
  NOR2_X1 U4296 ( .A1(n3560), .A2(n4136), .ZN(n3575) );
  INV_X1 U4297 ( .A(n4125), .ZN(n4128) );
  OAI21_X1 U4298 ( .B1(n3575), .B2(n3561), .A(n4128), .ZN(n3562) );
  OAI211_X1 U4299 ( .C1(n3565), .C2(n3564), .A(n3563), .B(n3562), .ZN(n3690)
         );
  NAND2_X1 U4300 ( .A1(n3858), .A2(n3566), .ZN(n3885) );
  INV_X1 U4301 ( .A(n3885), .ZN(n3584) );
  NAND2_X1 U4302 ( .A1(n2975), .A2(n4384), .ZN(n3615) );
  AND2_X1 U4303 ( .A1(n3567), .A2(n3615), .ZN(n4391) );
  INV_X1 U4304 ( .A(n3568), .ZN(n3570) );
  OR2_X1 U4305 ( .A1(n3570), .A2(n3569), .ZN(n4004) );
  INV_X1 U4306 ( .A(n3571), .ZN(n3573) );
  OR2_X1 U4307 ( .A1(n3573), .A2(n3572), .ZN(n4099) );
  NOR2_X1 U4308 ( .A1(n4127), .A2(n4125), .ZN(n3574) );
  NOR2_X1 U4309 ( .A1(n3575), .A2(n3574), .ZN(n3683) );
  NOR3_X1 U4310 ( .A1(n3578), .A2(n3577), .A3(n3576), .ZN(n3580) );
  NAND4_X1 U4311 ( .A1(n3581), .A2(n3683), .A3(n3580), .A4(n3579), .ZN(n3582)
         );
  NOR3_X1 U4312 ( .A1(n4004), .A2(n4099), .A3(n3582), .ZN(n3583) );
  NAND3_X1 U4313 ( .A1(n3584), .A2(n4391), .A3(n3583), .ZN(n3594) );
  NAND2_X1 U4314 ( .A1(n3882), .A2(n3585), .ZN(n3902) );
  INV_X1 U4315 ( .A(n3902), .ZN(n3589) );
  NAND2_X1 U4316 ( .A1(n3586), .A2(n3898), .ZN(n3922) );
  INV_X1 U4317 ( .A(n3922), .ZN(n3588) );
  AND2_X1 U4318 ( .A1(n3993), .A2(n3664), .ZN(n4036) );
  NAND4_X1 U4319 ( .A1(n3589), .A2(n3588), .A3(n4036), .A4(n3587), .ZN(n3593)
         );
  INV_X1 U4320 ( .A(n4016), .ZN(n4019) );
  NAND4_X1 U4321 ( .A1(n4019), .A2(n3591), .A3(n3590), .A4(n3629), .ZN(n3592)
         );
  NOR4_X1 U4322 ( .A1(n3820), .A2(n3594), .A3(n3593), .A4(n3592), .ZN(n3612)
         );
  XNOR2_X1 U4323 ( .A(n3596), .B(n3595), .ZN(n3826) );
  NAND2_X1 U4324 ( .A1(n3598), .A2(n3597), .ZN(n3861) );
  INV_X1 U4325 ( .A(n3861), .ZN(n3601) );
  NAND3_X1 U4326 ( .A1(n3601), .A2(n3600), .A3(n3599), .ZN(n3610) );
  XNOR2_X1 U4327 ( .A(n3999), .B(n3984), .ZN(n3978) );
  INV_X1 U4328 ( .A(n3602), .ZN(n3605) );
  NAND4_X1 U4329 ( .A1(n3605), .A2(n3105), .A3(n3604), .A4(n3603), .ZN(n3609)
         );
  NOR2_X1 U4330 ( .A1(n3918), .A2(n3917), .ZN(n3957) );
  INV_X1 U4331 ( .A(n3606), .ZN(n4078) );
  NAND4_X1 U4332 ( .A1(n3957), .A2(n4078), .A3(n3938), .A4(n3607), .ZN(n3608)
         );
  NOR4_X1 U4333 ( .A1(n3610), .A2(n3978), .A3(n3609), .A4(n3608), .ZN(n3611)
         );
  NAND4_X1 U4334 ( .A1(n3612), .A2(n3826), .A3(n3840), .A4(n3611), .ZN(n3688)
         );
  NOR2_X1 U4335 ( .A1(n3867), .A2(n3613), .ZN(n3680) );
  OAI211_X1 U4336 ( .C1(n3616), .C2(n4267), .A(n3615), .B(n3614), .ZN(n3618)
         );
  NAND3_X1 U4337 ( .A1(n3618), .A2(n3617), .A3(n3013), .ZN(n3621) );
  NAND3_X1 U4338 ( .A1(n3621), .A2(n3620), .A3(n3619), .ZN(n3624) );
  NAND3_X1 U4339 ( .A1(n3624), .A2(n3623), .A3(n3622), .ZN(n3627) );
  NAND4_X1 U4340 ( .A1(n3627), .A2(n3626), .A3(n3625), .A4(n3638), .ZN(n3630)
         );
  NAND3_X1 U4341 ( .A1(n3630), .A2(n3629), .A3(n3628), .ZN(n3637) );
  AND2_X1 U4342 ( .A1(n3632), .A2(n3631), .ZN(n3639) );
  INV_X1 U4343 ( .A(n3633), .ZN(n3636) );
  INV_X1 U4344 ( .A(n3634), .ZN(n3635) );
  AOI211_X1 U4345 ( .C1(n3637), .C2(n3639), .A(n3636), .B(n3635), .ZN(n3648)
         );
  INV_X1 U4346 ( .A(n3638), .ZN(n3642) );
  INV_X1 U4347 ( .A(n3639), .ZN(n3641) );
  NOR3_X1 U4348 ( .A1(n3642), .A2(n3641), .A3(n3640), .ZN(n3645) );
  INV_X1 U4349 ( .A(n3652), .ZN(n3644) );
  OAI21_X1 U4350 ( .B1(n3645), .B2(n3644), .A(n3643), .ZN(n3646) );
  OAI21_X1 U4351 ( .B1(n3648), .B2(n3647), .A(n3646), .ZN(n3656) );
  INV_X1 U4352 ( .A(n3649), .ZN(n3651) );
  AOI211_X1 U4353 ( .C1(n3653), .C2(n3652), .A(n3651), .B(n3650), .ZN(n3654)
         );
  NAND3_X1 U4354 ( .A1(n3656), .A2(n3655), .A3(n3654), .ZN(n3659) );
  INV_X1 U4355 ( .A(n3657), .ZN(n3658) );
  OAI211_X1 U4356 ( .C1(n3661), .C2(n3660), .A(n3659), .B(n3658), .ZN(n3663)
         );
  AOI21_X1 U4357 ( .B1(n3663), .B2(n4035), .A(n3662), .ZN(n3667) );
  INV_X1 U4358 ( .A(n3664), .ZN(n3666) );
  OAI21_X1 U4359 ( .B1(n3667), .B2(n3666), .A(n3665), .ZN(n3670) );
  INV_X1 U4360 ( .A(n3917), .ZN(n3668) );
  NAND3_X1 U4361 ( .A1(n3670), .A2(n3669), .A3(n3668), .ZN(n3671) );
  NAND2_X1 U4362 ( .A1(n3672), .A2(n3671), .ZN(n3675) );
  AOI211_X1 U4363 ( .C1(n3676), .C2(n3675), .A(n3674), .B(n3673), .ZN(n3679)
         );
  NOR4_X1 U4364 ( .A1(n3680), .A2(n3679), .A3(n3678), .A4(n3677), .ZN(n3685)
         );
  INV_X1 U4365 ( .A(n3681), .ZN(n3684) );
  OAI22_X1 U4366 ( .A1(n3685), .A2(n3684), .B1(n3683), .B2(n3682), .ZN(n3687)
         );
  MUX2_X1 U4367 ( .A(n3688), .B(n3687), .S(n3686), .Z(n3689) );
  NAND2_X1 U4368 ( .A1(n3690), .A2(n3689), .ZN(n3691) );
  XNOR2_X1 U4369 ( .A(n3691), .B(n4269), .ZN(n3697) );
  NAND2_X1 U4370 ( .A1(n3693), .A2(n3692), .ZN(n3694) );
  OAI211_X1 U4371 ( .C1(n4266), .C2(n3696), .A(n3694), .B(B_REG_SCAN_IN), .ZN(
        n3695) );
  OAI21_X1 U4372 ( .B1(n3697), .B2(n3696), .A(n3695), .ZN(U3239) );
  MUX2_X1 U4373 ( .A(n4127), .B(DATAO_REG_31__SCAN_IN), .S(n3709), .Z(U3581)
         );
  MUX2_X1 U4374 ( .A(n3816), .B(DATAO_REG_30__SCAN_IN), .S(n3709), .Z(U3580)
         );
  MUX2_X1 U4375 ( .A(DATAO_REG_29__SCAN_IN), .B(n3698), .S(U4043), .Z(U3579)
         );
  INV_X1 U4376 ( .A(n3822), .ZN(n3849) );
  MUX2_X1 U4377 ( .A(DATAO_REG_28__SCAN_IN), .B(n3849), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4378 ( .A(n3699), .B(DATAO_REG_27__SCAN_IN), .S(n3709), .Z(U3577)
         );
  MUX2_X1 U4379 ( .A(n3887), .B(DATAO_REG_26__SCAN_IN), .S(n3709), .Z(U3576)
         );
  MUX2_X1 U4380 ( .A(n3905), .B(DATAO_REG_25__SCAN_IN), .S(n3709), .Z(U3575)
         );
  MUX2_X1 U4381 ( .A(n3700), .B(DATAO_REG_24__SCAN_IN), .S(n3709), .Z(U3574)
         );
  MUX2_X1 U4382 ( .A(DATAO_REG_23__SCAN_IN), .B(n3701), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U4383 ( .A(n3960), .B(DATAO_REG_22__SCAN_IN), .S(n3709), .Z(U3572)
         );
  MUX2_X1 U4384 ( .A(n3942), .B(DATAO_REG_21__SCAN_IN), .S(n3709), .Z(U3571)
         );
  MUX2_X1 U4385 ( .A(n3961), .B(DATAO_REG_20__SCAN_IN), .S(n3709), .Z(U3570)
         );
  MUX2_X1 U4386 ( .A(n4021), .B(DATAO_REG_19__SCAN_IN), .S(n3709), .Z(U3569)
         );
  MUX2_X1 U4387 ( .A(DATAO_REG_18__SCAN_IN), .B(n3702), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4388 ( .A(DATAO_REG_17__SCAN_IN), .B(n3703), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4389 ( .A(DATAO_REG_16__SCAN_IN), .B(n4080), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4390 ( .A(n4070), .B(DATAO_REG_15__SCAN_IN), .S(n3709), .Z(U3565)
         );
  MUX2_X1 U4391 ( .A(DATAO_REG_14__SCAN_IN), .B(n4102), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4392 ( .A(n3704), .B(DATAO_REG_13__SCAN_IN), .S(n3709), .Z(U3563)
         );
  MUX2_X1 U4393 ( .A(n3288), .B(DATAO_REG_12__SCAN_IN), .S(n3709), .Z(U3562)
         );
  MUX2_X1 U4394 ( .A(DATAO_REG_11__SCAN_IN), .B(n3705), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4395 ( .A(n3706), .B(DATAO_REG_10__SCAN_IN), .S(n3709), .Z(U3560)
         );
  MUX2_X1 U4396 ( .A(n3707), .B(DATAO_REG_9__SCAN_IN), .S(n3709), .Z(U3559) );
  MUX2_X1 U4397 ( .A(DATAO_REG_7__SCAN_IN), .B(n3708), .S(U4043), .Z(U3557) );
  MUX2_X1 U4398 ( .A(n3710), .B(DATAO_REG_6__SCAN_IN), .S(n3709), .Z(U3556) );
  MUX2_X1 U4399 ( .A(DATAO_REG_5__SCAN_IN), .B(n3711), .S(U4043), .Z(U3555) );
  MUX2_X1 U4400 ( .A(DATAO_REG_4__SCAN_IN), .B(n3712), .S(U4043), .Z(U3554) );
  MUX2_X1 U4401 ( .A(DATAO_REG_2__SCAN_IN), .B(n3713), .S(U4043), .Z(U3552) );
  MUX2_X1 U4402 ( .A(DATAO_REG_1__SCAN_IN), .B(n2971), .S(U4043), .Z(U3551) );
  NAND3_X1 U4403 ( .A1(n4359), .A2(IR_REG_0__SCAN_IN), .A3(n4464), .ZN(n3720)
         );
  NAND2_X1 U4404 ( .A1(n4351), .A2(ADDR_REG_0__SCAN_IN), .ZN(n3719) );
  NAND2_X1 U4405 ( .A1(U3149), .A2(REG3_REG_0__SCAN_IN), .ZN(n3718) );
  INV_X1 U4406 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4395) );
  AOI21_X1 U4407 ( .B1(n3815), .B2(n4395), .A(n3732), .ZN(n3737) );
  NOR2_X1 U4408 ( .A1(n3815), .A2(REG1_REG_0__SCAN_IN), .ZN(n3714) );
  OAI21_X1 U4409 ( .B1(IR_REG_0__SCAN_IN), .B2(n3714), .A(n3737), .ZN(n3715)
         );
  OAI211_X1 U4410 ( .C1(IR_REG_0__SCAN_IN), .C2(n3737), .A(n3716), .B(n3715), 
        .ZN(n3717) );
  NAND4_X1 U4411 ( .A1(n3720), .A2(n3719), .A3(n3718), .A4(n3717), .ZN(U3240)
         );
  AOI22_X1 U4412 ( .A1(n4351), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3730) );
  NAND2_X1 U4413 ( .A1(n4335), .A2(n4277), .ZN(n3729) );
  MUX2_X1 U4414 ( .A(REG1_REG_1__SCAN_IN), .B(n3721), .S(n4277), .Z(n3723) );
  OAI211_X1 U4415 ( .C1(n3724), .C2(n3723), .A(n4359), .B(n3722), .ZN(n3728)
         );
  OAI211_X1 U4416 ( .C1(n3726), .C2(n3731), .A(n4373), .B(n3725), .ZN(n3727)
         );
  NAND4_X1 U4417 ( .A1(n3730), .A2(n3729), .A3(n3728), .A4(n3727), .ZN(U3241)
         );
  INV_X1 U4418 ( .A(n3731), .ZN(n3733) );
  AOI21_X1 U4419 ( .B1(n3815), .B2(n3733), .A(n3732), .ZN(n3734) );
  OAI21_X1 U4420 ( .B1(n3735), .B2(n3815), .A(n3734), .ZN(n3736) );
  OAI211_X1 U4421 ( .C1(IR_REG_0__SCAN_IN), .C2(n3737), .A(n3736), .B(U4043), 
        .ZN(n3757) );
  AOI22_X1 U4422 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4351), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3746) );
  XNOR2_X1 U4423 ( .A(n3739), .B(n3738), .ZN(n3740) );
  AOI22_X1 U4424 ( .A1(n4276), .A2(n4335), .B1(n4359), .B2(n3740), .ZN(n3745)
         );
  OAI211_X1 U4425 ( .C1(n3743), .C2(n3742), .A(n4373), .B(n3741), .ZN(n3744)
         );
  NAND4_X1 U4426 ( .A1(n3757), .A2(n3746), .A3(n3745), .A4(n3744), .ZN(U3242)
         );
  NAND2_X1 U4427 ( .A1(n4351), .A2(ADDR_REG_4__SCAN_IN), .ZN(n3756) );
  XNOR2_X1 U4428 ( .A(n3747), .B(REG1_REG_4__SCAN_IN), .ZN(n3748) );
  NAND2_X1 U4429 ( .A1(n4359), .A2(n3748), .ZN(n3751) );
  NAND2_X1 U4430 ( .A1(n4335), .A2(n4274), .ZN(n3750) );
  AND3_X1 U4431 ( .A1(n3751), .A2(n3750), .A3(n3749), .ZN(n3755) );
  XNOR2_X1 U4432 ( .A(n3752), .B(REG2_REG_4__SCAN_IN), .ZN(n3753) );
  NAND2_X1 U4433 ( .A1(n4373), .A2(n3753), .ZN(n3754) );
  NAND4_X1 U4434 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(U3244)
         );
  INV_X1 U4435 ( .A(n3776), .ZN(n4270) );
  XNOR2_X1 U4436 ( .A(n3776), .B(REG2_REG_17__SCAN_IN), .ZN(n3773) );
  INV_X1 U4437 ( .A(n4334), .ZN(n4409) );
  NOR2_X1 U4438 ( .A1(n4117), .A2(n4411), .ZN(n4319) );
  NAND2_X1 U4439 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3783), .ZN(n3764) );
  INV_X1 U4440 ( .A(n3783), .ZN(n4414) );
  INV_X1 U4441 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3758) );
  AOI22_X1 U4442 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3783), .B1(n4414), .B2(
        n3758), .ZN(n4301) );
  INV_X1 U4443 ( .A(n3759), .ZN(n3760) );
  NAND2_X1 U4444 ( .A1(n3779), .A2(n3762), .ZN(n3763) );
  NAND2_X1 U4445 ( .A1(n4301), .A2(n4300), .ZN(n4299) );
  NAND2_X1 U4446 ( .A1(n3764), .A2(n4299), .ZN(n3765) );
  NAND2_X1 U4447 ( .A1(n4412), .A2(n3765), .ZN(n3766) );
  XNOR2_X1 U4448 ( .A(n3765), .B(n4313), .ZN(n4310) );
  NAND2_X1 U4449 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4310), .ZN(n4309) );
  NAND2_X1 U4450 ( .A1(n3766), .A2(n4309), .ZN(n4321) );
  OAI22_X1 U4451 ( .A1(n4319), .A2(n4321), .B1(REG2_REG_13__SCAN_IN), .B2(
        n3786), .ZN(n3767) );
  NOR2_X1 U4452 ( .A1(n4409), .A2(n3767), .ZN(n3768) );
  INV_X1 U4453 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4331) );
  XNOR2_X1 U4454 ( .A(n4409), .B(n3767), .ZN(n4330) );
  NOR2_X1 U4455 ( .A1(n4331), .A2(n4330), .ZN(n4329) );
  NOR2_X1 U4456 ( .A1(n3768), .A2(n4329), .ZN(n4344) );
  INV_X1 U4457 ( .A(n3789), .ZN(n4407) );
  INV_X1 U4458 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3769) );
  AOI22_X1 U4459 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4407), .B1(n3789), .B2(
        n3769), .ZN(n4345) );
  NOR2_X1 U4460 ( .A1(n4344), .A2(n4345), .ZN(n4343) );
  NAND2_X1 U4461 ( .A1(n3770), .A2(n4405), .ZN(n3771) );
  NAND2_X1 U4462 ( .A1(n3772), .A2(n3773), .ZN(n3802) );
  OAI21_X1 U4463 ( .B1(n3773), .B2(n3772), .A(n3802), .ZN(n3774) );
  AOI22_X1 U4464 ( .A1(n4270), .A2(n4335), .B1(n4373), .B2(n3774), .ZN(n3797)
         );
  AOI21_X1 U4465 ( .B1(n4351), .B2(ADDR_REG_17__SCAN_IN), .A(n3775), .ZN(n3796) );
  XNOR2_X1 U4466 ( .A(n3776), .B(REG1_REG_17__SCAN_IN), .ZN(n3793) );
  INV_X1 U4467 ( .A(n3779), .ZN(n4416) );
  NOR2_X1 U4468 ( .A1(n3780), .A2(n4416), .ZN(n3781) );
  NAND2_X1 U4469 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3783), .ZN(n3782) );
  OAI21_X1 U4470 ( .B1(REG1_REG_11__SCAN_IN), .B2(n3783), .A(n3782), .ZN(n4296) );
  NOR2_X1 U4471 ( .A1(n3784), .A2(n4313), .ZN(n3785) );
  XOR2_X1 U4472 ( .A(n3784), .B(n4412), .Z(n4305) );
  NOR2_X1 U4473 ( .A1(n2510), .A2(n4305), .ZN(n4304) );
  AOI22_X1 U4474 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4411), .B1(n3786), .B2(
        n4201), .ZN(n4315) );
  NOR2_X1 U4475 ( .A1(n4316), .A2(n4315), .ZN(n4314) );
  XNOR2_X1 U4476 ( .A(n4409), .B(n3787), .ZN(n4326) );
  AOI22_X1 U4477 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4407), .B1(n3789), .B2(
        n3788), .ZN(n4340) );
  NAND2_X1 U4478 ( .A1(n3790), .A2(n4405), .ZN(n3791) );
  XOR2_X1 U4479 ( .A(n4405), .B(n3790), .Z(n4354) );
  NAND2_X1 U4480 ( .A1(n4354), .A2(n4353), .ZN(n4352) );
  NAND2_X1 U4481 ( .A1(n3791), .A2(n4352), .ZN(n3792) );
  NAND2_X1 U4482 ( .A1(n3792), .A2(n3793), .ZN(n3799) );
  OAI21_X1 U4483 ( .B1(n3793), .B2(n3792), .A(n3799), .ZN(n3794) );
  NAND2_X1 U4484 ( .A1(n4359), .A2(n3794), .ZN(n3795) );
  NAND3_X1 U4485 ( .A1(n3797), .A2(n3796), .A3(n3795), .ZN(U3257) );
  INV_X1 U4486 ( .A(n4402), .ZN(n4375) );
  AOI22_X1 U4487 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4375), .B1(n4402), .B2(
        n3798), .ZN(n4363) );
  OAI21_X1 U4488 ( .B1(REG1_REG_17__SCAN_IN), .B2(n4270), .A(n3799), .ZN(n4364) );
  XNOR2_X1 U4489 ( .A(n4269), .B(REG1_REG_19__SCAN_IN), .ZN(n3800) );
  NAND2_X1 U4490 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4402), .ZN(n3801) );
  OAI21_X1 U4491 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4402), .A(n3801), .ZN(n4372) );
  OAI21_X1 U4492 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4270), .A(n3802), .ZN(n4371) );
  INV_X1 U4493 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3803) );
  MUX2_X1 U4494 ( .A(REG2_REG_19__SCAN_IN), .B(n3803), .S(n4269), .Z(n3804) );
  AOI21_X1 U4495 ( .B1(n4351), .B2(ADDR_REG_19__SCAN_IN), .A(n3805), .ZN(n3806) );
  OAI21_X1 U4496 ( .B1(n4376), .B2(n3807), .A(n3806), .ZN(n3808) );
  INV_X1 U4497 ( .A(n3809), .ZN(n3810) );
  OAI21_X1 U4498 ( .B1(n3812), .B2(n3811), .A(n3810), .ZN(n3813) );
  XNOR2_X1 U4499 ( .A(n3813), .B(n3826), .ZN(n3814) );
  NAND2_X1 U4500 ( .A1(n3814), .A2(n4386), .ZN(n3818) );
  AOI21_X1 U4501 ( .B1(n3815), .B2(B_REG_SCAN_IN), .A(n4388), .ZN(n4126) );
  AOI22_X1 U4502 ( .A1(n3816), .A2(n4126), .B1(n3828), .B2(n4135), .ZN(n3817)
         );
  OAI211_X1 U4503 ( .C1(n3822), .C2(n4104), .A(n3818), .B(n3817), .ZN(n4139)
         );
  AOI21_X1 U4504 ( .B1(n3819), .B2(n4392), .A(n4139), .ZN(n3831) );
  INV_X1 U4505 ( .A(n3820), .ZN(n3824) );
  NAND2_X1 U4506 ( .A1(n4138), .A2(n4005), .ZN(n3830) );
  AOI21_X1 U4507 ( .B1(n3828), .B2(n3827), .A(n4130), .ZN(n4140) );
  AOI22_X1 U4508 ( .A1(n4140), .A2(n4378), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4281), .ZN(n3829) );
  OAI211_X1 U4509 ( .C1(n4281), .C2(n3831), .A(n3830), .B(n3829), .ZN(U3354)
         );
  INV_X1 U4510 ( .A(n3832), .ZN(n3839) );
  AOI22_X1 U4511 ( .A1(n3833), .A2(n4392), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4281), .ZN(n3834) );
  OAI21_X1 U4512 ( .B1(n3835), .B2(n4088), .A(n3834), .ZN(n3836) );
  AOI21_X1 U4513 ( .B1(n3837), .B2(n4396), .A(n3836), .ZN(n3838) );
  OAI21_X1 U4514 ( .B1(n3839), .B2(n4092), .A(n3838), .ZN(U3262) );
  XNOR2_X1 U4515 ( .A(n3841), .B(n3840), .ZN(n4143) );
  OAI22_X1 U4516 ( .A1(n3842), .A2(n4104), .B1(n3851), .B2(n4059), .ZN(n3848)
         );
  AOI21_X1 U4517 ( .B1(n3845), .B2(n3844), .A(n3843), .ZN(n3846) );
  NOR2_X1 U4518 ( .A1(n3846), .A2(n4065), .ZN(n3847) );
  AOI211_X1 U4519 ( .C1(n4101), .C2(n3849), .A(n3848), .B(n3847), .ZN(n4144)
         );
  NOR2_X1 U4520 ( .A1(n4144), .A2(n4281), .ZN(n3855) );
  OAI21_X1 U4521 ( .B1(n3868), .B2(n3851), .A(n3850), .ZN(n4146) );
  AOI22_X1 U4522 ( .A1(n3852), .A2(n4392), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4281), .ZN(n3853) );
  OAI21_X1 U4523 ( .B1(n4146), .B2(n4088), .A(n3853), .ZN(n3854) );
  AOI211_X1 U4524 ( .C1(n4143), .C2(n4005), .A(n3855), .B(n3854), .ZN(n3856)
         );
  INV_X1 U4525 ( .A(n3856), .ZN(U3263) );
  XNOR2_X1 U4526 ( .A(n3857), .B(n3861), .ZN(n4148) );
  INV_X1 U4527 ( .A(n4148), .ZN(n3876) );
  INV_X1 U4528 ( .A(n3858), .ZN(n3859) );
  AOI21_X1 U4529 ( .B1(n3883), .B2(n3860), .A(n3859), .ZN(n3862) );
  XNOR2_X1 U4530 ( .A(n3862), .B(n3861), .ZN(n3863) );
  NAND2_X1 U4531 ( .A1(n3863), .A2(n4386), .ZN(n3866) );
  AOI22_X1 U4532 ( .A1(n3905), .A2(n4071), .B1(n3864), .B2(n4135), .ZN(n3865)
         );
  OAI211_X1 U4533 ( .C1(n3867), .C2(n4388), .A(n3866), .B(n3865), .ZN(n4147)
         );
  INV_X1 U4534 ( .A(n3890), .ZN(n3871) );
  INV_X1 U4535 ( .A(n3868), .ZN(n3869) );
  AOI22_X1 U4536 ( .A1(n3872), .A2(n4392), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4281), .ZN(n3873) );
  OAI21_X1 U4537 ( .B1(n4218), .B2(n4088), .A(n3873), .ZN(n3874) );
  AOI21_X1 U4538 ( .B1(n4147), .B2(n4396), .A(n3874), .ZN(n3875) );
  OAI21_X1 U4539 ( .B1(n3876), .B2(n4092), .A(n3875), .ZN(U3264) );
  OR2_X1 U4540 ( .A1(n3877), .A2(n3878), .ZN(n3880) );
  NAND2_X1 U4541 ( .A1(n3880), .A2(n3879), .ZN(n3881) );
  XNOR2_X1 U4542 ( .A(n3881), .B(n3885), .ZN(n4152) );
  INV_X1 U4543 ( .A(n4152), .ZN(n3897) );
  NAND2_X1 U4544 ( .A1(n3883), .A2(n3882), .ZN(n3884) );
  XOR2_X1 U4545 ( .A(n3885), .B(n3884), .Z(n3889) );
  OAI22_X1 U4546 ( .A1(n3924), .A2(n4104), .B1(n3891), .B2(n4059), .ZN(n3886)
         );
  AOI21_X1 U4547 ( .B1(n4101), .B2(n3887), .A(n3886), .ZN(n3888) );
  OAI21_X1 U4548 ( .B1(n3889), .B2(n4065), .A(n3888), .ZN(n4151) );
  INV_X1 U4549 ( .A(n3910), .ZN(n3892) );
  OAI21_X1 U4550 ( .B1(n3892), .B2(n3891), .A(n3890), .ZN(n4222) );
  AOI22_X1 U4551 ( .A1(n4281), .A2(REG2_REG_25__SCAN_IN), .B1(n3893), .B2(
        n4392), .ZN(n3894) );
  OAI21_X1 U4552 ( .B1(n4222), .B2(n4088), .A(n3894), .ZN(n3895) );
  AOI21_X1 U4553 ( .B1(n4151), .B2(n4118), .A(n3895), .ZN(n3896) );
  OAI21_X1 U4554 ( .B1(n3897), .B2(n4092), .A(n3896), .ZN(U3265) );
  XOR2_X1 U4555 ( .A(n3902), .B(n3877), .Z(n4156) );
  INV_X1 U4556 ( .A(n4156), .ZN(n3915) );
  INV_X1 U4557 ( .A(n3898), .ZN(n3899) );
  NOR2_X1 U4558 ( .A1(n3900), .A2(n3899), .ZN(n3901) );
  XOR2_X1 U4559 ( .A(n3902), .B(n3901), .Z(n3907) );
  OAI22_X1 U4560 ( .A1(n3945), .A2(n4104), .B1(n3903), .B2(n4059), .ZN(n3904)
         );
  AOI21_X1 U4561 ( .B1(n3905), .B2(n4101), .A(n3904), .ZN(n3906) );
  OAI21_X1 U4562 ( .B1(n3907), .B2(n4065), .A(n3906), .ZN(n4155) );
  NAND2_X1 U4563 ( .A1(n3930), .A2(n3908), .ZN(n3909) );
  NAND2_X1 U4564 ( .A1(n3910), .A2(n3909), .ZN(n4226) );
  AOI22_X1 U4565 ( .A1(n4281), .A2(REG2_REG_24__SCAN_IN), .B1(n3911), .B2(
        n4392), .ZN(n3912) );
  OAI21_X1 U4566 ( .B1(n4226), .B2(n4088), .A(n3912), .ZN(n3913) );
  AOI21_X1 U4567 ( .B1(n4155), .B2(n4118), .A(n3913), .ZN(n3914) );
  OAI21_X1 U4568 ( .B1(n3915), .B2(n4092), .A(n3914), .ZN(U3266) );
  XOR2_X1 U4569 ( .A(n3922), .B(n3916), .Z(n4159) );
  INV_X1 U4570 ( .A(n4159), .ZN(n3935) );
  OR2_X1 U4571 ( .A1(n3958), .A2(n3917), .ZN(n3920) );
  INV_X1 U4572 ( .A(n3918), .ZN(n3919) );
  NAND2_X1 U4573 ( .A1(n3920), .A2(n3919), .ZN(n3939) );
  NAND2_X1 U4574 ( .A1(n3939), .A2(n3938), .ZN(n3941) );
  NAND2_X1 U4575 ( .A1(n3941), .A2(n3921), .ZN(n3923) );
  XNOR2_X1 U4576 ( .A(n3923), .B(n3922), .ZN(n3927) );
  OAI22_X1 U4577 ( .A1(n3924), .A2(n4388), .B1(n4059), .B2(n3928), .ZN(n3925)
         );
  AOI21_X1 U4578 ( .B1(n4071), .B2(n3960), .A(n3925), .ZN(n3926) );
  OAI21_X1 U4579 ( .B1(n3927), .B2(n4065), .A(n3926), .ZN(n4158) );
  OR2_X1 U4580 ( .A1(n3949), .A2(n3928), .ZN(n3929) );
  NAND2_X1 U4581 ( .A1(n3930), .A2(n3929), .ZN(n4230) );
  AOI22_X1 U4582 ( .A1(n4281), .A2(REG2_REG_23__SCAN_IN), .B1(n3931), .B2(
        n4392), .ZN(n3932) );
  OAI21_X1 U4583 ( .B1(n4230), .B2(n4088), .A(n3932), .ZN(n3933) );
  AOI21_X1 U4584 ( .B1(n4158), .B2(n4396), .A(n3933), .ZN(n3934) );
  OAI21_X1 U4585 ( .B1(n3935), .B2(n4092), .A(n3934), .ZN(U3267) );
  OAI21_X1 U4586 ( .B1(n2138), .B2(n2137), .A(n3937), .ZN(n4166) );
  OR2_X1 U4587 ( .A1(n3939), .A2(n3938), .ZN(n3940) );
  NAND2_X1 U4588 ( .A1(n3941), .A2(n3940), .ZN(n3947) );
  NAND2_X1 U4589 ( .A1(n3951), .A2(n4135), .ZN(n3944) );
  NAND2_X1 U4590 ( .A1(n3942), .A2(n4071), .ZN(n3943) );
  OAI211_X1 U4591 ( .C1(n3945), .C2(n4388), .A(n3944), .B(n3943), .ZN(n3946)
         );
  AOI21_X1 U4592 ( .B1(n3947), .B2(n4386), .A(n3946), .ZN(n4165) );
  AOI22_X1 U4593 ( .A1(n4281), .A2(REG2_REG_22__SCAN_IN), .B1(n3948), .B2(
        n4392), .ZN(n3953) );
  INV_X1 U4594 ( .A(n3949), .ZN(n4163) );
  INV_X1 U4595 ( .A(n3950), .ZN(n3965) );
  NAND2_X1 U4596 ( .A1(n3965), .A2(n3951), .ZN(n4162) );
  NAND3_X1 U4597 ( .A1(n4163), .A2(n4378), .A3(n4162), .ZN(n3952) );
  OAI211_X1 U4598 ( .C1(n4165), .C2(n4281), .A(n3953), .B(n3952), .ZN(n3954)
         );
  INV_X1 U4599 ( .A(n3954), .ZN(n3955) );
  OAI21_X1 U4600 ( .B1(n4166), .B2(n4092), .A(n3955), .ZN(U3268) );
  XNOR2_X1 U4601 ( .A(n3956), .B(n3957), .ZN(n4168) );
  INV_X1 U4602 ( .A(n4168), .ZN(n3972) );
  XNOR2_X1 U4603 ( .A(n3958), .B(n3957), .ZN(n3964) );
  NOR2_X1 U4604 ( .A1(n3966), .A2(n4059), .ZN(n3959) );
  AOI21_X1 U4605 ( .B1(n3960), .B2(n4101), .A(n3959), .ZN(n3963) );
  NAND2_X1 U4606 ( .A1(n3961), .A2(n4071), .ZN(n3962) );
  OAI211_X1 U4607 ( .C1(n3964), .C2(n4065), .A(n3963), .B(n3962), .ZN(n4167)
         );
  INV_X1 U4608 ( .A(n3986), .ZN(n3967) );
  OAI21_X1 U4609 ( .B1(n3967), .B2(n3966), .A(n3965), .ZN(n4235) );
  AOI22_X1 U4610 ( .A1(n4281), .A2(REG2_REG_21__SCAN_IN), .B1(n3968), .B2(
        n4392), .ZN(n3969) );
  OAI21_X1 U4611 ( .B1(n4235), .B2(n4088), .A(n3969), .ZN(n3970) );
  AOI21_X1 U4612 ( .B1(n4167), .B2(n4118), .A(n3970), .ZN(n3971) );
  OAI21_X1 U4613 ( .B1(n3972), .B2(n4092), .A(n3971), .ZN(U3269) );
  XNOR2_X1 U4614 ( .A(n3973), .B(n3978), .ZN(n4171) );
  OAI22_X1 U4615 ( .A1(n3975), .A2(n4388), .B1(n4059), .B2(n3974), .ZN(n3982)
         );
  OAI21_X1 U4616 ( .B1(n3994), .B2(n3977), .A(n3976), .ZN(n3979) );
  XNOR2_X1 U4617 ( .A(n3979), .B(n3978), .ZN(n3980) );
  NOR2_X1 U4618 ( .A1(n3980), .A2(n4065), .ZN(n3981) );
  AOI211_X1 U4619 ( .C1(n4071), .C2(n4021), .A(n3982), .B(n3981), .ZN(n3983)
         );
  OAI21_X1 U4620 ( .B1(n4171), .B2(n4109), .A(n3983), .ZN(n4172) );
  NAND2_X1 U4621 ( .A1(n4172), .A2(n4396), .ZN(n3992) );
  NAND2_X1 U4622 ( .A1(n4006), .A2(n3984), .ZN(n3985) );
  NAND2_X1 U4623 ( .A1(n3986), .A2(n3985), .ZN(n4238) );
  INV_X1 U4624 ( .A(n4238), .ZN(n3990) );
  INV_X1 U4625 ( .A(REG2_REG_20__SCAN_IN), .ZN(n3988) );
  OAI22_X1 U4626 ( .A1(n4118), .A2(n3988), .B1(n3987), .B2(n4115), .ZN(n3989)
         );
  AOI21_X1 U4627 ( .B1(n3990), .B2(n4378), .A(n3989), .ZN(n3991) );
  OAI211_X1 U4628 ( .C1(n4171), .C2(n4123), .A(n3992), .B(n3991), .ZN(U3270)
         );
  NAND2_X1 U4629 ( .A1(n3994), .A2(n3993), .ZN(n4020) );
  INV_X1 U4630 ( .A(n3995), .ZN(n3997) );
  OAI21_X1 U4631 ( .B1(n4020), .B2(n3997), .A(n3996), .ZN(n3998) );
  XNOR2_X1 U4632 ( .A(n3998), .B(n4004), .ZN(n4002) );
  NOR2_X1 U4633 ( .A1(n4038), .A2(n4104), .ZN(n4001) );
  OAI22_X1 U4634 ( .A1(n3999), .A2(n4388), .B1(n4059), .B2(n4007), .ZN(n4000)
         );
  AOI211_X1 U4635 ( .C1(n4002), .C2(n4386), .A(n4001), .B(n4000), .ZN(n4176)
         );
  XNOR2_X1 U4636 ( .A(n4003), .B(n4004), .ZN(n4178) );
  NAND2_X1 U4637 ( .A1(n4178), .A2(n4005), .ZN(n4014) );
  OAI21_X1 U4638 ( .B1(n4008), .B2(n4007), .A(n4006), .ZN(n4242) );
  INV_X1 U4639 ( .A(n4242), .ZN(n4012) );
  INV_X1 U4640 ( .A(n4009), .ZN(n4010) );
  OAI22_X1 U4641 ( .A1(n4118), .A2(n3803), .B1(n4010), .B2(n4115), .ZN(n4011)
         );
  AOI21_X1 U4642 ( .B1(n4012), .B2(n4378), .A(n4011), .ZN(n4013) );
  OAI211_X1 U4643 ( .C1(n4281), .C2(n4176), .A(n4014), .B(n4013), .ZN(U3271)
         );
  OAI21_X1 U4644 ( .B1(n4017), .B2(n4016), .A(n4015), .ZN(n4018) );
  INV_X1 U4645 ( .A(n4018), .ZN(n4183) );
  XNOR2_X1 U4646 ( .A(n4020), .B(n4019), .ZN(n4024) );
  AOI22_X1 U4647 ( .A1(n4021), .A2(n4101), .B1(n4025), .B2(n4135), .ZN(n4022)
         );
  OAI21_X1 U4648 ( .B1(n4061), .B2(n4104), .A(n4022), .ZN(n4023) );
  AOI21_X1 U4649 ( .B1(n4024), .B2(n4386), .A(n4023), .ZN(n4182) );
  INV_X1 U4650 ( .A(n4182), .ZN(n4032) );
  XNOR2_X1 U4651 ( .A(n4043), .B(n4025), .ZN(n4026) );
  NAND2_X1 U4652 ( .A1(n4026), .A2(n4443), .ZN(n4181) );
  INV_X1 U4653 ( .A(n4027), .ZN(n4030) );
  AOI22_X1 U4654 ( .A1(n4281), .A2(REG2_REG_18__SCAN_IN), .B1(n4028), .B2(
        n4392), .ZN(n4029) );
  OAI21_X1 U4655 ( .B1(n4181), .B2(n4030), .A(n4029), .ZN(n4031) );
  AOI21_X1 U4656 ( .B1(n4032), .B2(n4396), .A(n4031), .ZN(n4033) );
  OAI21_X1 U4657 ( .B1(n4183), .B2(n4092), .A(n4033), .ZN(U3272) );
  XNOR2_X1 U4658 ( .A(n4034), .B(n4036), .ZN(n4185) );
  INV_X1 U4659 ( .A(n4185), .ZN(n4050) );
  NAND2_X1 U4660 ( .A1(n4063), .A2(n4035), .ZN(n4037) );
  XNOR2_X1 U4661 ( .A(n4037), .B(n4036), .ZN(n4041) );
  OAI22_X1 U4662 ( .A1(n4038), .A2(n4388), .B1(n4059), .B2(n4045), .ZN(n4039)
         );
  AOI21_X1 U4663 ( .B1(n4071), .B2(n4080), .A(n4039), .ZN(n4040) );
  OAI21_X1 U4664 ( .B1(n4041), .B2(n4065), .A(n4040), .ZN(n4184) );
  INV_X1 U4665 ( .A(n4042), .ZN(n4053) );
  INV_X1 U4666 ( .A(n4043), .ZN(n4044) );
  OAI21_X1 U4667 ( .B1(n4053), .B2(n4045), .A(n4044), .ZN(n4247) );
  AOI22_X1 U4668 ( .A1(n4281), .A2(REG2_REG_17__SCAN_IN), .B1(n4046), .B2(
        n4392), .ZN(n4047) );
  OAI21_X1 U4669 ( .B1(n4247), .B2(n4088), .A(n4047), .ZN(n4048) );
  AOI21_X1 U4670 ( .B1(n4184), .B2(n4396), .A(n4048), .ZN(n4049) );
  OAI21_X1 U4671 ( .B1(n4050), .B2(n4092), .A(n4049), .ZN(U3273) );
  OAI21_X1 U4672 ( .B1(n4052), .B2(n4066), .A(n4051), .ZN(n4190) );
  AOI21_X1 U4673 ( .B1(n4055), .B2(n4054), .A(n4053), .ZN(n4187) );
  INV_X1 U4674 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4058) );
  INV_X1 U4675 ( .A(n4056), .ZN(n4057) );
  OAI22_X1 U4676 ( .A1(n4118), .A2(n4058), .B1(n4057), .B2(n4115), .ZN(n4073)
         );
  OAI22_X1 U4677 ( .A1(n4061), .A2(n4388), .B1(n4060), .B2(n4059), .ZN(n4069)
         );
  INV_X1 U4678 ( .A(n4062), .ZN(n4067) );
  INV_X1 U4679 ( .A(n4063), .ZN(n4064) );
  AOI211_X1 U4680 ( .C1(n4067), .C2(n4066), .A(n4065), .B(n4064), .ZN(n4068)
         );
  AOI211_X1 U4681 ( .C1(n4071), .C2(n4070), .A(n4069), .B(n4068), .ZN(n4189)
         );
  NOR2_X1 U4682 ( .A1(n4189), .A2(n4281), .ZN(n4072) );
  AOI211_X1 U4683 ( .C1(n4187), .C2(n4378), .A(n4073), .B(n4072), .ZN(n4074)
         );
  OAI21_X1 U4684 ( .B1(n4092), .B2(n4190), .A(n4074), .ZN(U3274) );
  XNOR2_X1 U4685 ( .A(n4075), .B(n4078), .ZN(n4194) );
  INV_X1 U4686 ( .A(n4076), .ZN(n4079) );
  OAI211_X1 U4687 ( .C1(n4079), .C2(n4078), .A(n4386), .B(n4077), .ZN(n4082)
         );
  AOI22_X1 U4688 ( .A1(n4080), .A2(n4101), .B1(n4135), .B2(n4084), .ZN(n4081)
         );
  OAI211_X1 U4689 ( .C1(n4083), .C2(n4104), .A(n4082), .B(n4081), .ZN(n4191)
         );
  XNOR2_X1 U4690 ( .A(n4085), .B(n4084), .ZN(n4192) );
  INV_X1 U4691 ( .A(n4192), .ZN(n4089) );
  AOI22_X1 U4692 ( .A1(n4281), .A2(REG2_REG_15__SCAN_IN), .B1(n4086), .B2(
        n4392), .ZN(n4087) );
  OAI21_X1 U4693 ( .B1(n4089), .B2(n4088), .A(n4087), .ZN(n4090) );
  AOI21_X1 U4694 ( .B1(n4191), .B2(n4396), .A(n4090), .ZN(n4091) );
  OAI21_X1 U4695 ( .B1(n4194), .B2(n4092), .A(n4091), .ZN(U3275) );
  XOR2_X1 U4696 ( .A(n4099), .B(n4093), .Z(n4198) );
  INV_X1 U4697 ( .A(n4094), .ZN(n4095) );
  AOI21_X1 U4698 ( .B1(n4097), .B2(n4096), .A(n4095), .ZN(n4098) );
  XOR2_X1 U4699 ( .A(n4099), .B(n4098), .Z(n4107) );
  AOI22_X1 U4700 ( .A1(n4102), .A2(n4101), .B1(n4135), .B2(n4100), .ZN(n4103)
         );
  OAI21_X1 U4701 ( .B1(n4105), .B2(n4104), .A(n4103), .ZN(n4106) );
  AOI21_X1 U4702 ( .B1(n4107), .B2(n4386), .A(n4106), .ZN(n4108) );
  OAI21_X1 U4703 ( .B1(n4198), .B2(n4109), .A(n4108), .ZN(n4199) );
  NAND2_X1 U4704 ( .A1(n4199), .A2(n4396), .ZN(n4122) );
  INV_X1 U4705 ( .A(n4110), .ZN(n4113) );
  OAI21_X1 U4706 ( .B1(n4113), .B2(n4112), .A(n4111), .ZN(n4257) );
  INV_X1 U4707 ( .A(n4257), .ZN(n4120) );
  INV_X1 U4708 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4117) );
  INV_X1 U4709 ( .A(n4114), .ZN(n4116) );
  OAI22_X1 U4710 ( .A1(n4118), .A2(n4117), .B1(n4116), .B2(n4115), .ZN(n4119)
         );
  AOI21_X1 U4711 ( .B1(n4120), .B2(n4378), .A(n4119), .ZN(n4121) );
  OAI211_X1 U4712 ( .C1(n4198), .C2(n4123), .A(n4122), .B(n4121), .ZN(U3277)
         );
  AND2_X1 U4713 ( .A1(n4127), .A2(n4126), .ZN(n4134) );
  AOI21_X1 U4714 ( .B1(n4128), .B2(n4135), .A(n4134), .ZN(n4280) );
  MUX2_X1 U4715 ( .A(n3532), .B(n4280), .S(n4474), .Z(n4129) );
  OAI21_X1 U4716 ( .B1(n4209), .B2(n4206), .A(n4129), .ZN(U3549) );
  INV_X1 U4717 ( .A(n4130), .ZN(n4133) );
  INV_X1 U4718 ( .A(n4131), .ZN(n4132) );
  INV_X1 U4719 ( .A(n4282), .ZN(n4212) );
  AOI21_X1 U4720 ( .B1(n4136), .B2(n4135), .A(n4134), .ZN(n4284) );
  MUX2_X1 U4721 ( .A(n3530), .B(n4284), .S(n4474), .Z(n4137) );
  OAI21_X1 U4722 ( .B1(n4212), .B2(n4206), .A(n4137), .ZN(U3548) );
  NAND2_X1 U4723 ( .A1(n4138), .A2(n4453), .ZN(n4142) );
  NAND2_X1 U4724 ( .A1(n4142), .A2(n4141), .ZN(n4213) );
  MUX2_X1 U4725 ( .A(REG1_REG_29__SCAN_IN), .B(n4213), .S(n4474), .Z(U3547) );
  INV_X1 U4726 ( .A(n4443), .ZN(n4455) );
  NAND2_X1 U4727 ( .A1(n4143), .A2(n4453), .ZN(n4145) );
  OAI211_X1 U4728 ( .C1(n4455), .C2(n4146), .A(n4145), .B(n4144), .ZN(n4214)
         );
  MUX2_X1 U4729 ( .A(REG1_REG_27__SCAN_IN), .B(n4214), .S(n4474), .Z(U3545) );
  AOI21_X1 U4730 ( .B1(n4148), .B2(n4453), .A(n4147), .ZN(n4215) );
  MUX2_X1 U4731 ( .A(n4149), .B(n4215), .S(n4474), .Z(n4150) );
  OAI21_X1 U4732 ( .B1(n4206), .B2(n4218), .A(n4150), .ZN(U3544) );
  AOI21_X1 U4733 ( .B1(n4152), .B2(n4453), .A(n4151), .ZN(n4219) );
  MUX2_X1 U4734 ( .A(n4153), .B(n4219), .S(n4474), .Z(n4154) );
  OAI21_X1 U4735 ( .B1(n4206), .B2(n4222), .A(n4154), .ZN(U3543) );
  INV_X1 U4736 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4589) );
  AOI21_X1 U4737 ( .B1(n4156), .B2(n4453), .A(n4155), .ZN(n4223) );
  MUX2_X1 U4738 ( .A(n4589), .B(n4223), .S(n4474), .Z(n4157) );
  OAI21_X1 U4739 ( .B1(n4206), .B2(n4226), .A(n4157), .ZN(U3542) );
  AOI21_X1 U4740 ( .B1(n4159), .B2(n4453), .A(n4158), .ZN(n4227) );
  MUX2_X1 U4741 ( .A(n4160), .B(n4227), .S(n4474), .Z(n4161) );
  OAI21_X1 U4742 ( .B1(n4206), .B2(n4230), .A(n4161), .ZN(U3541) );
  NAND3_X1 U4743 ( .A1(n4163), .A2(n4443), .A3(n4162), .ZN(n4164) );
  OAI211_X1 U4744 ( .C1(n4166), .C2(n4438), .A(n4165), .B(n4164), .ZN(n4231)
         );
  MUX2_X1 U4745 ( .A(REG1_REG_22__SCAN_IN), .B(n4231), .S(n4474), .Z(U3540) );
  AOI21_X1 U4746 ( .B1(n4168), .B2(n4453), .A(n4167), .ZN(n4232) );
  MUX2_X1 U4747 ( .A(n4169), .B(n4232), .S(n4474), .Z(n4170) );
  OAI21_X1 U4748 ( .B1(n4206), .B2(n4235), .A(n4170), .ZN(U3539) );
  INV_X1 U4749 ( .A(n4171), .ZN(n4173) );
  AOI21_X1 U4750 ( .B1(n4460), .B2(n4173), .A(n4172), .ZN(n4236) );
  MUX2_X1 U4751 ( .A(n4174), .B(n4236), .S(n4474), .Z(n4175) );
  OAI21_X1 U4752 ( .B1(n4206), .B2(n4238), .A(n4175), .ZN(U3538) );
  INV_X1 U4753 ( .A(n4176), .ZN(n4177) );
  AOI21_X1 U4754 ( .B1(n4178), .B2(n4453), .A(n4177), .ZN(n4239) );
  MUX2_X1 U4755 ( .A(n4179), .B(n4239), .S(n4474), .Z(n4180) );
  OAI21_X1 U4756 ( .B1(n4206), .B2(n4242), .A(n4180), .ZN(U3537) );
  OAI211_X1 U4757 ( .C1(n4183), .C2(n4438), .A(n4182), .B(n4181), .ZN(n4243)
         );
  MUX2_X1 U4758 ( .A(REG1_REG_18__SCAN_IN), .B(n4243), .S(n4474), .Z(U3536) );
  AOI21_X1 U4759 ( .B1(n4185), .B2(n4453), .A(n4184), .ZN(n4244) );
  MUX2_X1 U4760 ( .A(n4648), .B(n4244), .S(n4474), .Z(n4186) );
  OAI21_X1 U4761 ( .B1(n4206), .B2(n4247), .A(n4186), .ZN(U3535) );
  NAND2_X1 U4762 ( .A1(n4187), .A2(n4443), .ZN(n4188) );
  OAI211_X1 U4763 ( .C1(n4190), .C2(n4438), .A(n4189), .B(n4188), .ZN(n4248)
         );
  MUX2_X1 U4764 ( .A(REG1_REG_16__SCAN_IN), .B(n4248), .S(n4474), .Z(U3534) );
  AOI21_X1 U4765 ( .B1(n4443), .B2(n4192), .A(n4191), .ZN(n4193) );
  OAI21_X1 U4766 ( .B1(n4194), .B2(n4438), .A(n4193), .ZN(n4249) );
  MUX2_X1 U4767 ( .A(REG1_REG_15__SCAN_IN), .B(n4249), .S(n4474), .Z(U3533) );
  AOI21_X1 U4768 ( .B1(n4196), .B2(n4453), .A(n4195), .ZN(n4250) );
  MUX2_X1 U4769 ( .A(n4327), .B(n4250), .S(n4474), .Z(n4197) );
  OAI21_X1 U4770 ( .B1(n4206), .B2(n4253), .A(n4197), .ZN(U3532) );
  INV_X1 U4771 ( .A(n4198), .ZN(n4200) );
  AOI21_X1 U4772 ( .B1(n4460), .B2(n4200), .A(n4199), .ZN(n4254) );
  MUX2_X1 U4773 ( .A(n4201), .B(n4254), .S(n4474), .Z(n4202) );
  OAI21_X1 U4774 ( .B1(n4206), .B2(n4257), .A(n4202), .ZN(U3531) );
  AOI21_X1 U4775 ( .B1(n4453), .B2(n4204), .A(n4203), .ZN(n4258) );
  MUX2_X1 U4776 ( .A(n2510), .B(n4258), .S(n4474), .Z(n4205) );
  OAI21_X1 U4777 ( .B1(n4262), .B2(n4206), .A(n4205), .ZN(U3530) );
  INV_X1 U4778 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4207) );
  MUX2_X1 U4779 ( .A(n4207), .B(n4280), .S(n4463), .Z(n4208) );
  OAI21_X1 U4780 ( .B1(n4209), .B2(n4261), .A(n4208), .ZN(U3517) );
  INV_X1 U4781 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4210) );
  MUX2_X1 U4782 ( .A(n4210), .B(n4284), .S(n4463), .Z(n4211) );
  OAI21_X1 U4783 ( .B1(n4212), .B2(n4261), .A(n4211), .ZN(U3516) );
  MUX2_X1 U4784 ( .A(REG0_REG_29__SCAN_IN), .B(n4213), .S(n4463), .Z(U3515) );
  MUX2_X1 U4785 ( .A(REG0_REG_27__SCAN_IN), .B(n4214), .S(n4463), .Z(U3513) );
  INV_X1 U4786 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4216) );
  MUX2_X1 U4787 ( .A(n4216), .B(n4215), .S(n4463), .Z(n4217) );
  OAI21_X1 U4788 ( .B1(n4218), .B2(n4261), .A(n4217), .ZN(U3512) );
  INV_X1 U4789 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4220) );
  MUX2_X1 U4790 ( .A(n4220), .B(n4219), .S(n4463), .Z(n4221) );
  OAI21_X1 U4791 ( .B1(n4222), .B2(n4261), .A(n4221), .ZN(U3511) );
  INV_X1 U4792 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4224) );
  MUX2_X1 U4793 ( .A(n4224), .B(n4223), .S(n4463), .Z(n4225) );
  OAI21_X1 U4794 ( .B1(n4226), .B2(n4261), .A(n4225), .ZN(U3510) );
  INV_X1 U4795 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4228) );
  MUX2_X1 U4796 ( .A(n4228), .B(n4227), .S(n4463), .Z(n4229) );
  OAI21_X1 U4797 ( .B1(n4230), .B2(n4261), .A(n4229), .ZN(U3509) );
  MUX2_X1 U4798 ( .A(REG0_REG_22__SCAN_IN), .B(n4231), .S(n4463), .Z(U3508) );
  INV_X1 U4799 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4233) );
  MUX2_X1 U4800 ( .A(n4233), .B(n4232), .S(n4463), .Z(n4234) );
  OAI21_X1 U4801 ( .B1(n4235), .B2(n4261), .A(n4234), .ZN(U3507) );
  INV_X1 U4802 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4620) );
  MUX2_X1 U4803 ( .A(n4620), .B(n4236), .S(n4463), .Z(n4237) );
  OAI21_X1 U4804 ( .B1(n4238), .B2(n4261), .A(n4237), .ZN(U3506) );
  INV_X1 U4805 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4240) );
  MUX2_X1 U4806 ( .A(n4240), .B(n4239), .S(n4463), .Z(n4241) );
  OAI21_X1 U4807 ( .B1(n4242), .B2(n4261), .A(n4241), .ZN(U3505) );
  MUX2_X1 U4808 ( .A(REG0_REG_18__SCAN_IN), .B(n4243), .S(n4463), .Z(U3503) );
  INV_X1 U4809 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4245) );
  MUX2_X1 U4810 ( .A(n4245), .B(n4244), .S(n4463), .Z(n4246) );
  OAI21_X1 U4811 ( .B1(n4247), .B2(n4261), .A(n4246), .ZN(U3501) );
  MUX2_X1 U4812 ( .A(REG0_REG_16__SCAN_IN), .B(n4248), .S(n4463), .Z(U3499) );
  MUX2_X1 U4813 ( .A(REG0_REG_15__SCAN_IN), .B(n4249), .S(n4463), .Z(U3497) );
  INV_X1 U4814 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4251) );
  MUX2_X1 U4815 ( .A(n4251), .B(n4250), .S(n4463), .Z(n4252) );
  OAI21_X1 U4816 ( .B1(n4253), .B2(n4261), .A(n4252), .ZN(U3495) );
  INV_X1 U4817 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4255) );
  MUX2_X1 U4818 ( .A(n4255), .B(n4254), .S(n4463), .Z(n4256) );
  OAI21_X1 U4819 ( .B1(n4257), .B2(n4261), .A(n4256), .ZN(U3493) );
  INV_X1 U4820 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4259) );
  MUX2_X1 U4821 ( .A(n4259), .B(n4258), .S(n4463), .Z(n4260) );
  OAI21_X1 U4822 ( .B1(n4262), .B2(n4261), .A(n4260), .ZN(U3491) );
  MUX2_X1 U4823 ( .A(n4263), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U4824 ( .A(n2294), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U4825 ( .A(DATAI_28_), .B(n4264), .S(STATE_REG_SCAN_IN), .Z(U3324)
         );
  MUX2_X1 U4826 ( .A(DATAI_24_), .B(n4265), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U4827 ( .A(DATAI_22_), .B(n4266), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U4828 ( .A(DATAI_21_), .B(n4267), .S(STATE_REG_SCAN_IN), .Z(U3331)
         );
  MUX2_X1 U4829 ( .A(DATAI_20_), .B(n4268), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4830 ( .A(DATAI_19_), .B(n4269), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U4831 ( .A(DATAI_17_), .B(n4270), .S(STATE_REG_SCAN_IN), .Z(U3335)
         );
  MUX2_X1 U4832 ( .A(DATAI_7_), .B(n4271), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U4833 ( .A(n4272), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U4834 ( .A(n4273), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U4835 ( .A(DATAI_4_), .B(n4274), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4836 ( .A(n4275), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4837 ( .A(DATAI_2_), .B(n4276), .S(STATE_REG_SCAN_IN), .Z(U3350) );
  MUX2_X1 U4838 ( .A(n4277), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U4839 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(STATE_REG_SCAN_IN), 
        .Z(U3352) );
  AOI22_X1 U4840 ( .A1(n4278), .A2(n4378), .B1(n4281), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n4279) );
  OAI21_X1 U4841 ( .B1(n4281), .B2(n4280), .A(n4279), .ZN(U3260) );
  AOI22_X1 U4842 ( .A1(n4282), .A2(n4378), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4281), .ZN(n4283) );
  OAI21_X1 U4843 ( .B1(n4281), .B2(n4284), .A(n4283), .ZN(U3261) );
  AOI211_X1 U4844 ( .C1(n4287), .C2(n4286), .A(n4285), .B(n4362), .ZN(n4290)
         );
  INV_X1 U4845 ( .A(n4288), .ZN(n4289) );
  AOI211_X1 U4846 ( .C1(n4351), .C2(ADDR_REG_10__SCAN_IN), .A(n4290), .B(n4289), .ZN(n4294) );
  OAI211_X1 U4847 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4292), .A(n4373), .B(n4291), .ZN(n4293) );
  OAI211_X1 U4848 ( .C1(n4376), .C2(n4416), .A(n4294), .B(n4293), .ZN(U3250)
         );
  AOI211_X1 U4849 ( .C1(n2085), .C2(n4296), .A(n4295), .B(n4362), .ZN(n4298)
         );
  AOI211_X1 U4850 ( .C1(n4351), .C2(ADDR_REG_11__SCAN_IN), .A(n4298), .B(n4297), .ZN(n4303) );
  OAI211_X1 U4851 ( .C1(n4301), .C2(n4300), .A(n4373), .B(n4299), .ZN(n4302)
         );
  OAI211_X1 U4852 ( .C1(n4376), .C2(n4414), .A(n4303), .B(n4302), .ZN(U3251)
         );
  AOI211_X1 U4853 ( .C1(n2510), .C2(n4305), .A(n4304), .B(n4362), .ZN(n4308)
         );
  INV_X1 U4854 ( .A(n4306), .ZN(n4307) );
  AOI211_X1 U4855 ( .C1(n4351), .C2(ADDR_REG_12__SCAN_IN), .A(n4308), .B(n4307), .ZN(n4312) );
  OAI211_X1 U4856 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4310), .A(n4373), .B(n4309), .ZN(n4311) );
  OAI211_X1 U4857 ( .C1(n4376), .C2(n4313), .A(n4312), .B(n4311), .ZN(U3252)
         );
  AOI211_X1 U4858 ( .C1(n4316), .C2(n4315), .A(n4314), .B(n4362), .ZN(n4318)
         );
  AOI211_X1 U4859 ( .C1(n4351), .C2(ADDR_REG_13__SCAN_IN), .A(n4318), .B(n4317), .ZN(n4324) );
  AOI21_X1 U4860 ( .B1(n4117), .B2(n4411), .A(n4319), .ZN(n4322) );
  AOI21_X1 U4861 ( .B1(n4322), .B2(n4321), .A(n4328), .ZN(n4320) );
  OAI21_X1 U4862 ( .B1(n4322), .B2(n4321), .A(n4320), .ZN(n4323) );
  OAI211_X1 U4863 ( .C1(n4376), .C2(n4411), .A(n4324), .B(n4323), .ZN(U3253)
         );
  NAND2_X1 U4864 ( .A1(ADDR_REG_14__SCAN_IN), .A2(n4351), .ZN(n4338) );
  AOI211_X1 U4865 ( .C1(n4327), .C2(n4326), .A(n4325), .B(n4362), .ZN(n4333)
         );
  AOI211_X1 U4866 ( .C1(n4331), .C2(n4330), .A(n4329), .B(n4328), .ZN(n4332)
         );
  AOI211_X1 U4867 ( .C1(n4335), .C2(n4334), .A(n4333), .B(n4332), .ZN(n4337)
         );
  NAND3_X1 U4868 ( .A1(n4338), .A2(n4337), .A3(n4336), .ZN(U3254) );
  AOI211_X1 U4869 ( .C1(n2073), .C2(n4340), .A(n4339), .B(n4362), .ZN(n4341)
         );
  AOI211_X1 U4870 ( .C1(n4351), .C2(ADDR_REG_15__SCAN_IN), .A(n4342), .B(n4341), .ZN(n4348) );
  AOI21_X1 U4871 ( .B1(n4345), .B2(n4344), .A(n4343), .ZN(n4346) );
  NAND2_X1 U4872 ( .A1(n4373), .A2(n4346), .ZN(n4347) );
  OAI211_X1 U4873 ( .C1(n4376), .C2(n4407), .A(n4348), .B(n4347), .ZN(U3255)
         );
  INV_X1 U4874 ( .A(n4349), .ZN(n4350) );
  AOI21_X1 U4875 ( .B1(n4351), .B2(ADDR_REG_16__SCAN_IN), .A(n4350), .ZN(n4361) );
  OAI21_X1 U4876 ( .B1(n4354), .B2(n4353), .A(n4352), .ZN(n4358) );
  OAI21_X1 U4877 ( .B1(n4356), .B2(n4058), .A(n4355), .ZN(n4357) );
  AOI22_X1 U4878 ( .A1(n4359), .A2(n4358), .B1(n4373), .B2(n4357), .ZN(n4360)
         );
  OAI211_X1 U4879 ( .C1(n4405), .C2(n4376), .A(n4361), .B(n4360), .ZN(U3256)
         );
  NAND2_X1 U4880 ( .A1(n4351), .A2(ADDR_REG_18__SCAN_IN), .ZN(n4367) );
  NAND2_X1 U4881 ( .A1(n4367), .A2(n4366), .ZN(n4368) );
  AOI22_X1 U4882 ( .A1(REG2_REG_2__SCAN_IN), .A2(n4281), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4392), .ZN(n4381) );
  AOI22_X1 U4883 ( .A1(n4379), .A2(n4393), .B1(n4378), .B2(n4377), .ZN(n4380)
         );
  OAI211_X1 U4884 ( .C1(n4281), .C2(n4382), .A(n4381), .B(n4380), .ZN(U3288)
         );
  NOR2_X1 U4885 ( .A1(n4384), .A2(n4383), .ZN(n4418) );
  INV_X1 U4886 ( .A(n4385), .ZN(n4390) );
  NOR2_X1 U4887 ( .A1(n4387), .A2(n4386), .ZN(n4389) );
  OAI22_X1 U4888 ( .A1(n4391), .A2(n4389), .B1(n2340), .B2(n4388), .ZN(n4417)
         );
  AOI21_X1 U4889 ( .B1(n4418), .B2(n4390), .A(n4417), .ZN(n4397) );
  INV_X1 U4890 ( .A(n4391), .ZN(n4419) );
  AOI22_X1 U4891 ( .A1(n4419), .A2(n4393), .B1(REG3_REG_0__SCAN_IN), .B2(n4392), .ZN(n4394) );
  OAI221_X1 U4892 ( .B1(n4281), .B2(n4397), .C1(n4396), .C2(n4395), .A(n4394), 
        .ZN(U3290) );
  AND2_X1 U4893 ( .A1(D_REG_31__SCAN_IN), .A2(n4399), .ZN(U3291) );
  AND2_X1 U4894 ( .A1(D_REG_30__SCAN_IN), .A2(n4399), .ZN(U3292) );
  AND2_X1 U4895 ( .A1(D_REG_29__SCAN_IN), .A2(n4399), .ZN(U3293) );
  AND2_X1 U4896 ( .A1(D_REG_28__SCAN_IN), .A2(n4399), .ZN(U3294) );
  INV_X1 U4897 ( .A(D_REG_27__SCAN_IN), .ZN(n4499) );
  NOR2_X1 U4898 ( .A1(n4398), .A2(n4499), .ZN(U3295) );
  INV_X1 U4899 ( .A(D_REG_26__SCAN_IN), .ZN(n4605) );
  NOR2_X1 U4900 ( .A1(n4398), .A2(n4605), .ZN(U3296) );
  INV_X1 U4901 ( .A(D_REG_25__SCAN_IN), .ZN(n4631) );
  NOR2_X1 U4902 ( .A1(n4398), .A2(n4631), .ZN(U3297) );
  AND2_X1 U4903 ( .A1(D_REG_24__SCAN_IN), .A2(n4399), .ZN(U3298) );
  AND2_X1 U4904 ( .A1(D_REG_23__SCAN_IN), .A2(n4399), .ZN(U3299) );
  AND2_X1 U4905 ( .A1(D_REG_22__SCAN_IN), .A2(n4399), .ZN(U3300) );
  AND2_X1 U4906 ( .A1(D_REG_21__SCAN_IN), .A2(n4399), .ZN(U3301) );
  AND2_X1 U4907 ( .A1(D_REG_20__SCAN_IN), .A2(n4399), .ZN(U3302) );
  AND2_X1 U4908 ( .A1(D_REG_19__SCAN_IN), .A2(n4399), .ZN(U3303) );
  INV_X1 U4909 ( .A(D_REG_18__SCAN_IN), .ZN(n4630) );
  NOR2_X1 U4910 ( .A1(n4398), .A2(n4630), .ZN(U3304) );
  AND2_X1 U4911 ( .A1(D_REG_17__SCAN_IN), .A2(n4399), .ZN(U3305) );
  AND2_X1 U4912 ( .A1(D_REG_16__SCAN_IN), .A2(n4399), .ZN(U3306) );
  AND2_X1 U4913 ( .A1(D_REG_15__SCAN_IN), .A2(n4399), .ZN(U3307) );
  AND2_X1 U4914 ( .A1(D_REG_14__SCAN_IN), .A2(n4399), .ZN(U3308) );
  AND2_X1 U4915 ( .A1(D_REG_13__SCAN_IN), .A2(n4399), .ZN(U3309) );
  INV_X1 U4916 ( .A(D_REG_12__SCAN_IN), .ZN(n4515) );
  NOR2_X1 U4917 ( .A1(n4398), .A2(n4515), .ZN(U3310) );
  INV_X1 U4918 ( .A(D_REG_11__SCAN_IN), .ZN(n4621) );
  NOR2_X1 U4919 ( .A1(n4398), .A2(n4621), .ZN(U3311) );
  AND2_X1 U4920 ( .A1(D_REG_10__SCAN_IN), .A2(n4399), .ZN(U3312) );
  INV_X1 U4921 ( .A(D_REG_9__SCAN_IN), .ZN(n4476) );
  NOR2_X1 U4922 ( .A1(n4398), .A2(n4476), .ZN(U3313) );
  INV_X1 U4923 ( .A(D_REG_8__SCAN_IN), .ZN(n4477) );
  NOR2_X1 U4924 ( .A1(n4398), .A2(n4477), .ZN(U3314) );
  AND2_X1 U4925 ( .A1(D_REG_7__SCAN_IN), .A2(n4399), .ZN(U3315) );
  AND2_X1 U4926 ( .A1(D_REG_6__SCAN_IN), .A2(n4399), .ZN(U3316) );
  INV_X1 U4927 ( .A(D_REG_5__SCAN_IN), .ZN(n4514) );
  NOR2_X1 U4928 ( .A1(n4398), .A2(n4514), .ZN(U3317) );
  AND2_X1 U4929 ( .A1(D_REG_4__SCAN_IN), .A2(n4399), .ZN(U3318) );
  AND2_X1 U4930 ( .A1(D_REG_3__SCAN_IN), .A2(n4399), .ZN(U3319) );
  AND2_X1 U4931 ( .A1(D_REG_2__SCAN_IN), .A2(n4399), .ZN(U3320) );
  INV_X1 U4932 ( .A(DATAI_23_), .ZN(n4401) );
  AOI21_X1 U4933 ( .B1(U3149), .B2(n4401), .A(n4400), .ZN(U3329) );
  OAI22_X1 U4934 ( .A1(U3149), .A2(n4402), .B1(DATAI_18_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4403) );
  INV_X1 U4935 ( .A(n4403), .ZN(U3334) );
  INV_X1 U4936 ( .A(DATAI_16_), .ZN(n4404) );
  AOI22_X1 U4937 ( .A1(STATE_REG_SCAN_IN), .A2(n4405), .B1(n4404), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U4938 ( .A(DATAI_15_), .ZN(n4406) );
  AOI22_X1 U4939 ( .A1(STATE_REG_SCAN_IN), .A2(n4407), .B1(n4406), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U4940 ( .A(DATAI_14_), .ZN(n4408) );
  AOI22_X1 U4941 ( .A1(STATE_REG_SCAN_IN), .A2(n4409), .B1(n4408), .B2(U3149), 
        .ZN(U3338) );
  AOI22_X1 U4942 ( .A1(STATE_REG_SCAN_IN), .A2(n4411), .B1(n4410), .B2(U3149), 
        .ZN(U3339) );
  OAI22_X1 U4943 ( .A1(U3149), .A2(n4412), .B1(DATAI_12_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4413) );
  INV_X1 U4944 ( .A(n4413), .ZN(U3340) );
  INV_X1 U4945 ( .A(DATAI_11_), .ZN(n4511) );
  AOI22_X1 U4946 ( .A1(STATE_REG_SCAN_IN), .A2(n4414), .B1(n4511), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U4947 ( .A(DATAI_10_), .ZN(n4415) );
  AOI22_X1 U4948 ( .A1(STATE_REG_SCAN_IN), .A2(n4416), .B1(n4415), .B2(U3149), 
        .ZN(U3342) );
  AOI211_X1 U4949 ( .C1(n4460), .C2(n4419), .A(n4418), .B(n4417), .ZN(n4465)
         );
  INV_X1 U4950 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4420) );
  AOI22_X1 U4951 ( .A1(n4463), .A2(n4465), .B1(n4420), .B2(n4461), .ZN(U3467)
         );
  OAI22_X1 U4952 ( .A1(n4422), .A2(n4427), .B1(n4455), .B2(n4421), .ZN(n4423)
         );
  NOR2_X1 U4953 ( .A1(n4424), .A2(n4423), .ZN(n4466) );
  INV_X1 U4954 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4425) );
  AOI22_X1 U4955 ( .A1(n4463), .A2(n4466), .B1(n4425), .B2(n4461), .ZN(U3469)
         );
  OAI22_X1 U4956 ( .A1(n4428), .A2(n4427), .B1(n4455), .B2(n4426), .ZN(n4429)
         );
  NOR2_X1 U4957 ( .A1(n4430), .A2(n4429), .ZN(n4467) );
  INV_X1 U4958 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4431) );
  AOI22_X1 U4959 ( .A1(n4463), .A2(n4467), .B1(n4431), .B2(n4461), .ZN(U3473)
         );
  INV_X1 U4960 ( .A(n4432), .ZN(n4434) );
  AOI211_X1 U4961 ( .C1(n4435), .C2(n4460), .A(n4434), .B(n4433), .ZN(n4468)
         );
  INV_X1 U4962 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4436) );
  AOI22_X1 U4963 ( .A1(n4463), .A2(n4468), .B1(n4436), .B2(n4461), .ZN(U3475)
         );
  INV_X1 U4964 ( .A(n4437), .ZN(n4441) );
  NOR2_X1 U4965 ( .A1(n4439), .A2(n4438), .ZN(n4440) );
  AOI211_X1 U4966 ( .C1(n4443), .C2(n4442), .A(n4441), .B(n4440), .ZN(n4469)
         );
  INV_X1 U4967 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4444) );
  AOI22_X1 U4968 ( .A1(n4463), .A2(n4469), .B1(n4444), .B2(n4461), .ZN(U3477)
         );
  NAND3_X1 U4969 ( .A1(n4446), .A2(n4445), .A3(n4453), .ZN(n4447) );
  AND3_X1 U4970 ( .A1(n4449), .A2(n4448), .A3(n4447), .ZN(n4470) );
  INV_X1 U4971 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4636) );
  AOI22_X1 U4972 ( .A1(n4463), .A2(n4470), .B1(n4636), .B2(n4461), .ZN(U3481)
         );
  OAI21_X1 U4973 ( .B1(n4455), .B2(n4451), .A(n4450), .ZN(n4452) );
  AOI21_X1 U4974 ( .B1(n4454), .B2(n4453), .A(n4452), .ZN(n4471) );
  INV_X1 U4975 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4489) );
  AOI22_X1 U4976 ( .A1(n4463), .A2(n4471), .B1(n4489), .B2(n4461), .ZN(U3485)
         );
  NOR2_X1 U4977 ( .A1(n4456), .A2(n4455), .ZN(n4458) );
  AOI211_X1 U4978 ( .C1(n4460), .C2(n4459), .A(n4458), .B(n4457), .ZN(n4473)
         );
  INV_X1 U4979 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4462) );
  AOI22_X1 U4980 ( .A1(n4463), .A2(n4473), .B1(n4462), .B2(n4461), .ZN(U3489)
         );
  AOI22_X1 U4981 ( .A1(n4474), .A2(n4465), .B1(n4464), .B2(n4472), .ZN(U3518)
         );
  AOI22_X1 U4982 ( .A1(n4474), .A2(n4466), .B1(n3721), .B2(n4472), .ZN(U3519)
         );
  AOI22_X1 U4983 ( .A1(n4474), .A2(n4467), .B1(n2365), .B2(n4472), .ZN(U3521)
         );
  AOI22_X1 U4984 ( .A1(n4474), .A2(n4468), .B1(n2862), .B2(n4472), .ZN(U3522)
         );
  AOI22_X1 U4985 ( .A1(n4474), .A2(n4469), .B1(n2857), .B2(n4472), .ZN(U3523)
         );
  AOI22_X1 U4986 ( .A1(n4474), .A2(n4470), .B1(n2427), .B2(n4472), .ZN(U3525)
         );
  AOI22_X1 U4987 ( .A1(n4474), .A2(n4471), .B1(n2898), .B2(n4472), .ZN(U3527)
         );
  AOI22_X1 U4988 ( .A1(n4474), .A2(n4473), .B1(n2495), .B2(n4472), .ZN(U3529)
         );
  AOI22_X1 U4989 ( .A1(n4477), .A2(keyinput93), .B1(keyinput115), .B2(n4476), 
        .ZN(n4475) );
  OAI221_X1 U4990 ( .B1(n4477), .B2(keyinput93), .C1(n4476), .C2(keyinput115), 
        .A(n4475), .ZN(n4486) );
  AOI22_X1 U4991 ( .A1(n4650), .A2(keyinput75), .B1(n4618), .B2(keyinput124), 
        .ZN(n4478) );
  OAI221_X1 U4992 ( .B1(n4650), .B2(keyinput75), .C1(n4618), .C2(keyinput124), 
        .A(n4478), .ZN(n4485) );
  INV_X1 U4993 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n4645) );
  AOI22_X1 U4994 ( .A1(n4645), .A2(keyinput74), .B1(n4633), .B2(keyinput84), 
        .ZN(n4479) );
  OAI221_X1 U4995 ( .B1(n4645), .B2(keyinput74), .C1(n4633), .C2(keyinput84), 
        .A(n4479), .ZN(n4484) );
  INV_X1 U4996 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n4481) );
  AOI22_X1 U4997 ( .A1(n4482), .A2(keyinput82), .B1(keyinput67), .B2(n4481), 
        .ZN(n4480) );
  OAI221_X1 U4998 ( .B1(n4482), .B2(keyinput82), .C1(n4481), .C2(keyinput67), 
        .A(n4480), .ZN(n4483) );
  NOR4_X1 U4999 ( .A1(n4486), .A2(n4485), .A3(n4484), .A4(n4483), .ZN(n4526)
         );
  AOI22_X1 U5000 ( .A1(n4620), .A2(keyinput120), .B1(keyinput72), .B2(n4636), 
        .ZN(n4487) );
  OAI221_X1 U5001 ( .B1(n4620), .B2(keyinput120), .C1(n4636), .C2(keyinput72), 
        .A(n4487), .ZN(n4497) );
  AOI22_X1 U5002 ( .A1(n4489), .A2(keyinput127), .B1(n4648), .B2(keyinput87), 
        .ZN(n4488) );
  OAI221_X1 U5003 ( .B1(n4489), .B2(keyinput127), .C1(n4648), .C2(keyinput87), 
        .A(n4488), .ZN(n4496) );
  XNOR2_X1 U5004 ( .A(REG1_REG_2__SCAN_IN), .B(keyinput69), .ZN(n4492) );
  XNOR2_X1 U5005 ( .A(REG0_REG_18__SCAN_IN), .B(keyinput125), .ZN(n4491) );
  XNOR2_X1 U5006 ( .A(REG2_REG_1__SCAN_IN), .B(keyinput99), .ZN(n4490) );
  NAND3_X1 U5007 ( .A1(n4492), .A2(n4491), .A3(n4490), .ZN(n4495) );
  XNOR2_X1 U5008 ( .A(n4493), .B(keyinput101), .ZN(n4494) );
  NOR4_X1 U5009 ( .A1(n4497), .A2(n4496), .A3(n4495), .A4(n4494), .ZN(n4525)
         );
  AOI22_X1 U5010 ( .A1(n4621), .A2(keyinput114), .B1(n4499), .B2(keyinput89), 
        .ZN(n4498) );
  OAI221_X1 U5011 ( .B1(n4621), .B2(keyinput114), .C1(n4499), .C2(keyinput89), 
        .A(n4498), .ZN(n4509) );
  AOI22_X1 U5012 ( .A1(n4502), .A2(keyinput79), .B1(keyinput78), .B2(n4501), 
        .ZN(n4500) );
  OAI221_X1 U5013 ( .B1(n4502), .B2(keyinput79), .C1(n4501), .C2(keyinput78), 
        .A(n4500), .ZN(n4508) );
  XNOR2_X1 U5014 ( .A(n4631), .B(keyinput109), .ZN(n4507) );
  XNOR2_X1 U5015 ( .A(IR_REG_28__SCAN_IN), .B(keyinput107), .ZN(n4505) );
  XNOR2_X1 U5016 ( .A(IR_REG_17__SCAN_IN), .B(keyinput71), .ZN(n4504) );
  XNOR2_X1 U5017 ( .A(IR_REG_22__SCAN_IN), .B(keyinput70), .ZN(n4503) );
  NAND3_X1 U5018 ( .A1(n4505), .A2(n4504), .A3(n4503), .ZN(n4506) );
  NOR4_X1 U5019 ( .A1(n4509), .A2(n4508), .A3(n4507), .A4(n4506), .ZN(n4524)
         );
  AOI22_X1 U5020 ( .A1(n4512), .A2(keyinput106), .B1(keyinput112), .B2(n4511), 
        .ZN(n4510) );
  OAI221_X1 U5021 ( .B1(n4512), .B2(keyinput106), .C1(n4511), .C2(keyinput112), 
        .A(n4510), .ZN(n4522) );
  AOI22_X1 U5022 ( .A1(n4515), .A2(keyinput80), .B1(n4514), .B2(keyinput68), 
        .ZN(n4513) );
  OAI221_X1 U5023 ( .B1(n4515), .B2(keyinput80), .C1(n4514), .C2(keyinput68), 
        .A(n4513), .ZN(n4521) );
  XNOR2_X1 U5024 ( .A(IR_REG_0__SCAN_IN), .B(keyinput103), .ZN(n4519) );
  XNOR2_X1 U5025 ( .A(IR_REG_1__SCAN_IN), .B(keyinput111), .ZN(n4518) );
  XNOR2_X1 U5026 ( .A(IR_REG_6__SCAN_IN), .B(keyinput86), .ZN(n4517) );
  XNOR2_X1 U5027 ( .A(IR_REG_3__SCAN_IN), .B(keyinput94), .ZN(n4516) );
  NAND4_X1 U5028 ( .A1(n4519), .A2(n4518), .A3(n4517), .A4(n4516), .ZN(n4520)
         );
  NOR3_X1 U5029 ( .A1(n4522), .A2(n4521), .A3(n4520), .ZN(n4523) );
  AND4_X1 U5030 ( .A1(n4526), .A2(n4525), .A3(n4524), .A4(n4523), .ZN(n4665)
         );
  OAI22_X1 U5031 ( .A1(REG2_REG_20__SCAN_IN), .A2(keyinput97), .B1(
        REG2_REG_12__SCAN_IN), .B2(keyinput83), .ZN(n4527) );
  AOI221_X1 U5032 ( .B1(REG2_REG_20__SCAN_IN), .B2(keyinput97), .C1(keyinput83), .C2(REG2_REG_12__SCAN_IN), .A(n4527), .ZN(n4534) );
  OAI22_X1 U5033 ( .A1(REG2_REG_24__SCAN_IN), .A2(keyinput91), .B1(keyinput76), 
        .B2(DATAO_REG_24__SCAN_IN), .ZN(n4528) );
  AOI221_X1 U5034 ( .B1(REG2_REG_24__SCAN_IN), .B2(keyinput91), .C1(
        DATAO_REG_24__SCAN_IN), .C2(keyinput76), .A(n4528), .ZN(n4533) );
  OAI22_X1 U5035 ( .A1(REG3_REG_4__SCAN_IN), .A2(keyinput85), .B1(keyinput81), 
        .B2(REG3_REG_0__SCAN_IN), .ZN(n4529) );
  AOI221_X1 U5036 ( .B1(REG3_REG_4__SCAN_IN), .B2(keyinput85), .C1(
        REG3_REG_0__SCAN_IN), .C2(keyinput81), .A(n4529), .ZN(n4532) );
  OAI22_X1 U5037 ( .A1(ADDR_REG_9__SCAN_IN), .A2(keyinput90), .B1(keyinput116), 
        .B2(ADDR_REG_8__SCAN_IN), .ZN(n4530) );
  AOI221_X1 U5038 ( .B1(ADDR_REG_9__SCAN_IN), .B2(keyinput90), .C1(
        ADDR_REG_8__SCAN_IN), .C2(keyinput116), .A(n4530), .ZN(n4531) );
  NAND4_X1 U5039 ( .A1(n4534), .A2(n4533), .A3(n4532), .A4(n4531), .ZN(n4563)
         );
  OAI22_X1 U5040 ( .A1(REG2_REG_5__SCAN_IN), .A2(keyinput123), .B1(
        REG1_REG_31__SCAN_IN), .B2(keyinput104), .ZN(n4535) );
  AOI221_X1 U5041 ( .B1(REG2_REG_5__SCAN_IN), .B2(keyinput123), .C1(
        keyinput104), .C2(REG1_REG_31__SCAN_IN), .A(n4535), .ZN(n4542) );
  OAI22_X1 U5042 ( .A1(REG1_REG_25__SCAN_IN), .A2(keyinput113), .B1(
        REG1_REG_18__SCAN_IN), .B2(keyinput118), .ZN(n4536) );
  AOI221_X1 U5043 ( .B1(REG1_REG_25__SCAN_IN), .B2(keyinput113), .C1(
        keyinput118), .C2(REG1_REG_18__SCAN_IN), .A(n4536), .ZN(n4541) );
  OAI22_X1 U5044 ( .A1(ADDR_REG_2__SCAN_IN), .A2(keyinput66), .B1(
        DATAO_REG_16__SCAN_IN), .B2(keyinput96), .ZN(n4537) );
  AOI221_X1 U5045 ( .B1(ADDR_REG_2__SCAN_IN), .B2(keyinput66), .C1(keyinput96), 
        .C2(DATAO_REG_16__SCAN_IN), .A(n4537), .ZN(n4540) );
  OAI22_X1 U5046 ( .A1(REG0_REG_26__SCAN_IN), .A2(keyinput100), .B1(
        REG0_REG_22__SCAN_IN), .B2(keyinput122), .ZN(n4538) );
  AOI221_X1 U5047 ( .B1(REG0_REG_26__SCAN_IN), .B2(keyinput100), .C1(
        keyinput122), .C2(REG0_REG_22__SCAN_IN), .A(n4538), .ZN(n4539) );
  NAND4_X1 U5048 ( .A1(n4542), .A2(n4541), .A3(n4540), .A4(n4539), .ZN(n4562)
         );
  OAI22_X1 U5049 ( .A1(IR_REG_20__SCAN_IN), .A2(keyinput110), .B1(
        IR_REG_8__SCAN_IN), .B2(keyinput73), .ZN(n4543) );
  AOI221_X1 U5050 ( .B1(IR_REG_20__SCAN_IN), .B2(keyinput110), .C1(keyinput73), 
        .C2(IR_REG_8__SCAN_IN), .A(n4543), .ZN(n4551) );
  OAI22_X1 U5051 ( .A1(D_REG_26__SCAN_IN), .A2(keyinput95), .B1(keyinput92), 
        .B2(REG0_REG_2__SCAN_IN), .ZN(n4544) );
  AOI221_X1 U5052 ( .B1(D_REG_26__SCAN_IN), .B2(keyinput95), .C1(
        REG0_REG_2__SCAN_IN), .C2(keyinput92), .A(n4544), .ZN(n4550) );
  OAI22_X1 U5053 ( .A1(n4546), .A2(keyinput102), .B1(n2838), .B2(keyinput105), 
        .ZN(n4545) );
  AOI221_X1 U5054 ( .B1(n4546), .B2(keyinput102), .C1(keyinput105), .C2(n2838), 
        .A(n4545), .ZN(n4549) );
  OAI22_X1 U5055 ( .A1(n4589), .A2(keyinput108), .B1(keyinput88), .B2(
        IR_REG_31__SCAN_IN), .ZN(n4547) );
  AOI221_X1 U5056 ( .B1(n4589), .B2(keyinput108), .C1(IR_REG_31__SCAN_IN), 
        .C2(keyinput88), .A(n4547), .ZN(n4548) );
  NAND4_X1 U5057 ( .A1(n4551), .A2(n4550), .A3(n4549), .A4(n4548), .ZN(n4561)
         );
  OAI22_X1 U5058 ( .A1(DATAI_26_), .A2(keyinput98), .B1(keyinput65), .B2(
        DATAI_31_), .ZN(n4552) );
  AOI221_X1 U5059 ( .B1(DATAI_26_), .B2(keyinput98), .C1(DATAI_31_), .C2(
        keyinput65), .A(n4552), .ZN(n4559) );
  OAI22_X1 U5060 ( .A1(REG3_REG_3__SCAN_IN), .A2(keyinput119), .B1(DATAI_23_), 
        .B2(keyinput64), .ZN(n4553) );
  AOI221_X1 U5061 ( .B1(REG3_REG_3__SCAN_IN), .B2(keyinput119), .C1(keyinput64), .C2(DATAI_23_), .A(n4553), .ZN(n4558) );
  OAI22_X1 U5062 ( .A1(D_REG_18__SCAN_IN), .A2(keyinput121), .B1(keyinput126), 
        .B2(DATAI_9_), .ZN(n4554) );
  AOI221_X1 U5063 ( .B1(D_REG_18__SCAN_IN), .B2(keyinput121), .C1(DATAI_9_), 
        .C2(keyinput126), .A(n4554), .ZN(n4557) );
  OAI22_X1 U5064 ( .A1(REG3_REG_14__SCAN_IN), .A2(keyinput77), .B1(DATAI_0_), 
        .B2(keyinput117), .ZN(n4555) );
  AOI221_X1 U5065 ( .B1(REG3_REG_14__SCAN_IN), .B2(keyinput77), .C1(
        keyinput117), .C2(DATAI_0_), .A(n4555), .ZN(n4556) );
  NAND4_X1 U5066 ( .A1(n4559), .A2(n4558), .A3(n4557), .A4(n4556), .ZN(n4560)
         );
  NOR4_X1 U5067 ( .A1(n4563), .A2(n4562), .A3(n4561), .A4(n4560), .ZN(n4664)
         );
  AOI22_X1 U5068 ( .A1(REG2_REG_2__SCAN_IN), .A2(keyinput41), .B1(
        REG1_REG_2__SCAN_IN), .B2(keyinput5), .ZN(n4564) );
  OAI221_X1 U5069 ( .B1(REG2_REG_2__SCAN_IN), .B2(keyinput41), .C1(
        REG1_REG_2__SCAN_IN), .C2(keyinput5), .A(n4564), .ZN(n4571) );
  AOI22_X1 U5070 ( .A1(REG2_REG_20__SCAN_IN), .A2(keyinput33), .B1(
        REG1_REG_25__SCAN_IN), .B2(keyinput49), .ZN(n4565) );
  OAI221_X1 U5071 ( .B1(REG2_REG_20__SCAN_IN), .B2(keyinput33), .C1(
        REG1_REG_25__SCAN_IN), .C2(keyinput49), .A(n4565), .ZN(n4570) );
  AOI22_X1 U5072 ( .A1(D_REG_8__SCAN_IN), .A2(keyinput29), .B1(
        IR_REG_8__SCAN_IN), .B2(keyinput9), .ZN(n4566) );
  OAI221_X1 U5073 ( .B1(D_REG_8__SCAN_IN), .B2(keyinput29), .C1(
        IR_REG_8__SCAN_IN), .C2(keyinput9), .A(n4566), .ZN(n4569) );
  AOI22_X1 U5074 ( .A1(DATAO_REG_3__SCAN_IN), .A2(keyinput37), .B1(
        D_REG_27__SCAN_IN), .B2(keyinput25), .ZN(n4567) );
  OAI221_X1 U5075 ( .B1(DATAO_REG_3__SCAN_IN), .B2(keyinput37), .C1(
        D_REG_27__SCAN_IN), .C2(keyinput25), .A(n4567), .ZN(n4568) );
  NOR4_X1 U5076 ( .A1(n4571), .A2(n4570), .A3(n4569), .A4(n4568), .ZN(n4602)
         );
  AOI22_X1 U5077 ( .A1(ADDR_REG_8__SCAN_IN), .A2(keyinput52), .B1(
        REG0_REG_26__SCAN_IN), .B2(keyinput36), .ZN(n4572) );
  OAI221_X1 U5078 ( .B1(ADDR_REG_8__SCAN_IN), .B2(keyinput52), .C1(
        REG0_REG_26__SCAN_IN), .C2(keyinput36), .A(n4572), .ZN(n4579) );
  AOI22_X1 U5079 ( .A1(DATAI_11_), .A2(keyinput48), .B1(REG3_REG_14__SCAN_IN), 
        .B2(keyinput13), .ZN(n4573) );
  OAI221_X1 U5080 ( .B1(DATAI_11_), .B2(keyinput48), .C1(REG3_REG_14__SCAN_IN), 
        .C2(keyinput13), .A(n4573), .ZN(n4578) );
  AOI22_X1 U5081 ( .A1(D_REG_12__SCAN_IN), .A2(keyinput16), .B1(
        D_REG_5__SCAN_IN), .B2(keyinput4), .ZN(n4574) );
  OAI221_X1 U5082 ( .B1(D_REG_12__SCAN_IN), .B2(keyinput16), .C1(
        D_REG_5__SCAN_IN), .C2(keyinput4), .A(n4574), .ZN(n4577) );
  AOI22_X1 U5083 ( .A1(DATAO_REG_24__SCAN_IN), .A2(keyinput12), .B1(
        DATAO_REG_16__SCAN_IN), .B2(keyinput32), .ZN(n4575) );
  OAI221_X1 U5084 ( .B1(DATAO_REG_24__SCAN_IN), .B2(keyinput12), .C1(
        DATAO_REG_16__SCAN_IN), .C2(keyinput32), .A(n4575), .ZN(n4576) );
  NOR4_X1 U5085 ( .A1(n4579), .A2(n4578), .A3(n4577), .A4(n4576), .ZN(n4601)
         );
  AOI22_X1 U5086 ( .A1(REG0_REG_22__SCAN_IN), .A2(keyinput58), .B1(
        REG1_REG_28__SCAN_IN), .B2(keyinput38), .ZN(n4580) );
  OAI221_X1 U5087 ( .B1(REG0_REG_22__SCAN_IN), .B2(keyinput58), .C1(
        REG1_REG_28__SCAN_IN), .C2(keyinput38), .A(n4580), .ZN(n4587) );
  AOI22_X1 U5088 ( .A1(REG2_REG_7__SCAN_IN), .A2(keyinput18), .B1(
        IR_REG_6__SCAN_IN), .B2(keyinput22), .ZN(n4581) );
  OAI221_X1 U5089 ( .B1(REG2_REG_7__SCAN_IN), .B2(keyinput18), .C1(
        IR_REG_6__SCAN_IN), .C2(keyinput22), .A(n4581), .ZN(n4586) );
  AOI22_X1 U5090 ( .A1(ADDR_REG_2__SCAN_IN), .A2(keyinput2), .B1(
        D_REG_0__SCAN_IN), .B2(keyinput14), .ZN(n4582) );
  OAI221_X1 U5091 ( .B1(ADDR_REG_2__SCAN_IN), .B2(keyinput2), .C1(
        D_REG_0__SCAN_IN), .C2(keyinput14), .A(n4582), .ZN(n4585) );
  AOI22_X1 U5092 ( .A1(ADDR_REG_3__SCAN_IN), .A2(keyinput3), .B1(DATAI_23_), 
        .B2(keyinput0), .ZN(n4583) );
  OAI221_X1 U5093 ( .B1(ADDR_REG_3__SCAN_IN), .B2(keyinput3), .C1(DATAI_23_), 
        .C2(keyinput0), .A(n4583), .ZN(n4584) );
  NOR4_X1 U5094 ( .A1(n4587), .A2(n4586), .A3(n4585), .A4(n4584), .ZN(n4600)
         );
  INV_X1 U5095 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4590) );
  AOI22_X1 U5096 ( .A1(n4590), .A2(keyinput28), .B1(keyinput44), .B2(n4589), 
        .ZN(n4588) );
  OAI221_X1 U5097 ( .B1(n4590), .B2(keyinput28), .C1(n4589), .C2(keyinput44), 
        .A(n4588), .ZN(n4598) );
  AOI22_X1 U5098 ( .A1(REG2_REG_5__SCAN_IN), .A2(keyinput59), .B1(
        IR_REG_0__SCAN_IN), .B2(keyinput39), .ZN(n4591) );
  OAI221_X1 U5099 ( .B1(REG2_REG_5__SCAN_IN), .B2(keyinput59), .C1(
        IR_REG_0__SCAN_IN), .C2(keyinput39), .A(n4591), .ZN(n4597) );
  AOI22_X1 U5100 ( .A1(REG0_REG_9__SCAN_IN), .A2(keyinput63), .B1(
        IR_REG_16__SCAN_IN), .B2(keyinput15), .ZN(n4592) );
  OAI221_X1 U5101 ( .B1(REG0_REG_9__SCAN_IN), .B2(keyinput63), .C1(
        IR_REG_16__SCAN_IN), .C2(keyinput15), .A(n4592), .ZN(n4596) );
  XOR2_X1 U5102 ( .A(D_REG_9__SCAN_IN), .B(keyinput51), .Z(n4594) );
  XNOR2_X1 U5103 ( .A(IR_REG_31__SCAN_IN), .B(keyinput24), .ZN(n4593) );
  NAND2_X1 U5104 ( .A1(n4594), .A2(n4593), .ZN(n4595) );
  NOR4_X1 U5105 ( .A1(n4598), .A2(n4597), .A3(n4596), .A4(n4595), .ZN(n4599)
         );
  NAND4_X1 U5106 ( .A1(n4602), .A2(n4601), .A3(n4600), .A4(n4599), .ZN(n4663)
         );
  INV_X1 U5107 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4604) );
  AOI22_X1 U5108 ( .A1(n4605), .A2(keyinput31), .B1(keyinput27), .B2(n4604), 
        .ZN(n4603) );
  OAI221_X1 U5109 ( .B1(n4605), .B2(keyinput31), .C1(n4604), .C2(keyinput27), 
        .A(n4603), .ZN(n4615) );
  XNOR2_X1 U5110 ( .A(n4606), .B(keyinput35), .ZN(n4614) );
  XNOR2_X1 U5111 ( .A(DATAI_17_), .B(keyinput42), .ZN(n4610) );
  XNOR2_X1 U5112 ( .A(IR_REG_28__SCAN_IN), .B(keyinput43), .ZN(n4609) );
  XNOR2_X1 U5113 ( .A(IR_REG_3__SCAN_IN), .B(keyinput30), .ZN(n4608) );
  XNOR2_X1 U5114 ( .A(IR_REG_1__SCAN_IN), .B(keyinput47), .ZN(n4607) );
  NAND4_X1 U5115 ( .A1(n4610), .A2(n4609), .A3(n4608), .A4(n4607), .ZN(n4613)
         );
  XNOR2_X1 U5116 ( .A(keyinput34), .B(n4611), .ZN(n4612) );
  NOR4_X1 U5117 ( .A1(n4615), .A2(n4614), .A3(n4613), .A4(n4612), .ZN(n4661)
         );
  INV_X1 U5118 ( .A(DATAI_9_), .ZN(n4617) );
  AOI22_X1 U5119 ( .A1(n4618), .A2(keyinput60), .B1(n4617), .B2(keyinput62), 
        .ZN(n4616) );
  OAI221_X1 U5120 ( .B1(n4618), .B2(keyinput60), .C1(n4617), .C2(keyinput62), 
        .A(n4616), .ZN(n4628) );
  AOI22_X1 U5121 ( .A1(n3532), .A2(keyinput40), .B1(n4620), .B2(keyinput56), 
        .ZN(n4619) );
  OAI221_X1 U5122 ( .B1(n3532), .B2(keyinput40), .C1(n4620), .C2(keyinput56), 
        .A(n4619), .ZN(n4627) );
  XNOR2_X1 U5123 ( .A(n4621), .B(keyinput50), .ZN(n4626) );
  XNOR2_X1 U5124 ( .A(REG1_REG_18__SCAN_IN), .B(keyinput54), .ZN(n4624) );
  XNOR2_X1 U5125 ( .A(IR_REG_20__SCAN_IN), .B(keyinput46), .ZN(n4623) );
  XNOR2_X1 U5126 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput55), .ZN(n4622) );
  NAND3_X1 U5127 ( .A1(n4624), .A2(n4623), .A3(n4622), .ZN(n4625) );
  NOR4_X1 U5128 ( .A1(n4628), .A2(n4627), .A3(n4626), .A4(n4625), .ZN(n4660)
         );
  AOI22_X1 U5129 ( .A1(n4631), .A2(keyinput45), .B1(keyinput57), .B2(n4630), 
        .ZN(n4629) );
  OAI221_X1 U5130 ( .B1(n4631), .B2(keyinput45), .C1(n4630), .C2(keyinput57), 
        .A(n4629), .ZN(n4643) );
  INV_X1 U5131 ( .A(REG0_REG_18__SCAN_IN), .ZN(n4634) );
  AOI22_X1 U5132 ( .A1(n4634), .A2(keyinput61), .B1(n4633), .B2(keyinput20), 
        .ZN(n4632) );
  OAI221_X1 U5133 ( .B1(n4634), .B2(keyinput61), .C1(n4633), .C2(keyinput20), 
        .A(n4632), .ZN(n4642) );
  XNOR2_X1 U5134 ( .A(n4635), .B(keyinput1), .ZN(n4641) );
  XOR2_X1 U5135 ( .A(n4636), .B(keyinput8), .Z(n4639) );
  XNOR2_X1 U5136 ( .A(DATAI_0_), .B(keyinput53), .ZN(n4638) );
  XNOR2_X1 U5137 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput21), .ZN(n4637) );
  NAND3_X1 U5138 ( .A1(n4639), .A2(n4638), .A3(n4637), .ZN(n4640) );
  NOR4_X1 U5139 ( .A1(n4643), .A2(n4642), .A3(n4641), .A4(n4640), .ZN(n4659)
         );
  INV_X1 U5140 ( .A(REG2_REG_12__SCAN_IN), .ZN(n4646) );
  AOI22_X1 U5141 ( .A1(n4646), .A2(keyinput19), .B1(keyinput10), .B2(n4645), 
        .ZN(n4644) );
  OAI221_X1 U5142 ( .B1(n4646), .B2(keyinput19), .C1(n4645), .C2(keyinput10), 
        .A(n4644), .ZN(n4657) );
  INV_X1 U5143 ( .A(ADDR_REG_9__SCAN_IN), .ZN(n4649) );
  AOI22_X1 U5144 ( .A1(n4649), .A2(keyinput26), .B1(n4648), .B2(keyinput23), 
        .ZN(n4647) );
  OAI221_X1 U5145 ( .B1(n4649), .B2(keyinput26), .C1(n4648), .C2(keyinput23), 
        .A(n4647), .ZN(n4656) );
  XNOR2_X1 U5146 ( .A(n4650), .B(keyinput11), .ZN(n4655) );
  XNOR2_X1 U5147 ( .A(IR_REG_22__SCAN_IN), .B(keyinput6), .ZN(n4653) );
  XNOR2_X1 U5148 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput17), .ZN(n4652) );
  XNOR2_X1 U5149 ( .A(IR_REG_17__SCAN_IN), .B(keyinput7), .ZN(n4651) );
  NAND3_X1 U5150 ( .A1(n4653), .A2(n4652), .A3(n4651), .ZN(n4654) );
  NOR4_X1 U5151 ( .A1(n4657), .A2(n4656), .A3(n4655), .A4(n4654), .ZN(n4658)
         );
  NAND4_X1 U5152 ( .A1(n4661), .A2(n4660), .A3(n4659), .A4(n4658), .ZN(n4662)
         );
  AOI211_X1 U5153 ( .C1(n4665), .C2(n4664), .A(n4663), .B(n4662), .ZN(n4669)
         );
  NAND2_X1 U5154 ( .A1(n4666), .A2(STATE_REG_SCAN_IN), .ZN(n4667) );
  OAI21_X1 U5155 ( .B1(DATAI_9_), .B2(STATE_REG_SCAN_IN), .A(n4667), .ZN(n4668) );
  XNOR2_X1 U5156 ( .A(n4669), .B(n4668), .ZN(U3343) );
  CLKBUF_X1 U2331 ( .A(n2343), .Z(n3531) );
  CLKBUF_X1 U2387 ( .A(n4396), .Z(n4118) );
endmodule

