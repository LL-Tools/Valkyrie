

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884;

  CLKBUF_X2 U2374 ( .A(n2408), .Z(n2416) );
  INV_X2 U2375 ( .A(IR_REG_0__SCAN_IN), .ZN(n4428) );
  NAND2_X1 U2376 ( .A1(n3594), .A2(n3139), .ZN(n2968) );
  INV_X1 U2377 ( .A(n2132), .ZN(n2952) );
  INV_X1 U2378 ( .A(n3594), .ZN(n3627) );
  INV_X2 U2380 ( .A(IR_REG_31__SCAN_IN), .ZN(n2194) );
  INV_X2 U2381 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND2_X1 U2383 ( .A1(n2949), .A2(n2768), .ZN(n3628) );
  OAI21_X2 U2384 ( .B1(n4209), .B2(n3880), .A(n3881), .ZN(n4186) );
  AOI21_X2 U2385 ( .B1(n4223), .B2(n2599), .A(n2598), .ZN(n4209) );
  OAI21_X2 U2386 ( .B1(n3229), .B2(n2280), .A(n2279), .ZN(n3319) );
  OAI21_X1 U2387 ( .B1(n3166), .B2(n3165), .A(n3164), .ZN(n3229) );
  BUF_X1 U2388 ( .A(n2968), .Z(n3631) );
  OR2_X1 U2389 ( .A1(n2946), .A2(n2403), .ZN(n3891) );
  INV_X2 U2390 ( .A(n3604), .ZN(n3630) );
  NAND2_X1 U2391 ( .A1(n2403), .A2(n3005), .ZN(n3055) );
  NAND2_X1 U2392 ( .A1(n2381), .A2(n4409), .ZN(n2393) );
  AND2_X1 U2393 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2360)
         );
  NAND2_X1 U2394 ( .A1(n3661), .A2(n3575), .ZN(n3664) );
  NAND2_X1 U2395 ( .A1(n2311), .A2(n2167), .ZN(n2317) );
  NAND2_X1 U2396 ( .A1(n2351), .A2(n2350), .ZN(n4245) );
  NAND2_X1 U2397 ( .A1(n3449), .A2(n2568), .ZN(n3485) );
  OR2_X2 U2398 ( .A1(n3338), .A2(n3706), .ZN(n2201) );
  CLKBUF_X1 U2399 ( .A(n3798), .Z(n3746) );
  AOI21_X1 U2400 ( .B1(n2286), .B2(n2287), .A(n2284), .ZN(n2283) );
  NAND2_X1 U2401 ( .A1(n2896), .A2(n2266), .ZN(n4008) );
  NOR2_X2 U2402 ( .A1(n2933), .A2(n4539), .ZN(n2934) );
  NAND2_X2 U2403 ( .A1(n2993), .A2(n4239), .ZN(n4421) );
  NAND2_X1 U2404 ( .A1(n3891), .A2(n3889), .ZN(n2320) );
  AND2_X1 U2405 ( .A1(n3904), .A2(n3907), .ZN(n2363) );
  INV_X2 U2406 ( .A(n2968), .ZN(n2945) );
  INV_X1 U2407 ( .A(n3194), .ZN(n3984) );
  NAND4_X1 U2408 ( .A1(n2420), .A2(n2419), .A3(n2418), .A4(n2417), .ZN(n3150)
         );
  AND2_X1 U2409 ( .A1(n2439), .A2(n2438), .ZN(n3194) );
  NAND4_X1 U2410 ( .A1(n2413), .A2(n2412), .A3(n2411), .A4(n2410), .ZN(n3027)
         );
  AND2_X2 U2411 ( .A1(n2769), .A2(n2997), .ZN(n3604) );
  INV_X1 U2412 ( .A(n3004), .ZN(n3005) );
  INV_X1 U2413 ( .A(n2768), .ZN(n2997) );
  AND2_X1 U2414 ( .A1(n2740), .A2(n2739), .ZN(n2741) );
  INV_X1 U2415 ( .A(n3077), .ZN(n3062) );
  NAND2_X1 U2416 ( .A1(n2729), .A2(n2728), .ZN(n3624) );
  INV_X1 U2417 ( .A(n2745), .ZN(n4410) );
  AND2_X1 U2418 ( .A1(n2383), .A2(n2382), .ZN(n2408) );
  XNOR2_X1 U2419 ( .A(n2721), .B(IR_REG_26__SCAN_IN), .ZN(n2739) );
  NAND2_X1 U2420 ( .A1(n2380), .A2(n2379), .ZN(n2382) );
  XNOR2_X1 U2421 ( .A(n2674), .B(n2730), .ZN(n2928) );
  NAND2_X1 U2422 ( .A1(n2662), .A2(IR_REG_31__SCAN_IN), .ZN(n2663) );
  AND2_X1 U2423 ( .A1(n2662), .A2(n2597), .ZN(n4412) );
  MUX2_X1 U2424 ( .A(IR_REG_31__SCAN_IN), .B(n2378), .S(IR_REG_29__SCAN_IN), 
        .Z(n2380) );
  NAND2_X1 U2425 ( .A1(n2724), .A2(IR_REG_31__SCAN_IN), .ZN(n2721) );
  NAND2_X1 U2426 ( .A1(n2723), .A2(IR_REG_25__SCAN_IN), .ZN(n2729) );
  OAI21_X1 U2427 ( .B1(n2667), .B2(IR_REG_18__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2596) );
  OR2_X1 U2428 ( .A1(n2722), .A2(n2189), .ZN(n2188) );
  AND2_X1 U2429 ( .A1(n2486), .A2(n2303), .ZN(n2302) );
  OR2_X1 U2430 ( .A1(IR_REG_18__SCAN_IN), .A2(n2666), .ZN(n2669) );
  NAND3_X1 U2431 ( .A1(n2185), .A2(n2184), .A3(n2183), .ZN(n2830) );
  AND2_X1 U2432 ( .A1(n2365), .A2(n2462), .ZN(n2486) );
  AND4_X1 U2433 ( .A1(n2373), .A2(n2372), .A3(n2371), .A4(n2730), .ZN(n2374)
         );
  AND4_X1 U2434 ( .A1(n2367), .A2(n2369), .A3(n2368), .A4(n2553), .ZN(n2370)
         );
  AND2_X1 U2435 ( .A1(n2366), .A2(n2304), .ZN(n2303) );
  NOR2_X1 U2436 ( .A1(n2360), .A2(n2194), .ZN(n2190) );
  NOR2_X1 U2437 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2358)
         );
  NOR2_X1 U2438 ( .A1(IR_REG_2__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2206)
         );
  INV_X1 U2439 ( .A(IR_REG_15__SCAN_IN), .ZN(n2553) );
  NOR2_X1 U2440 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2368)
         );
  NOR2_X1 U2441 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2369)
         );
  NOR2_X1 U2442 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2367)
         );
  NOR2_X1 U2443 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2365)
         );
  INV_X1 U2444 ( .A(IR_REG_9__SCAN_IN), .ZN(n2366) );
  INV_X1 U2445 ( .A(IR_REG_19__SCAN_IN), .ZN(n2665) );
  INV_X1 U2446 ( .A(IR_REG_20__SCAN_IN), .ZN(n2664) );
  INV_X1 U2447 ( .A(IR_REG_22__SCAN_IN), .ZN(n2730) );
  OR2_X1 U2448 ( .A1(n2766), .A2(n4587), .ZN(n2222) );
  INV_X1 U2449 ( .A(n2947), .ZN(n2971) );
  NOR2_X2 U2450 ( .A1(n3055), .A2(n3056), .ZN(n3054) );
  AND2_X1 U2451 ( .A1(n2769), .A2(n2997), .ZN(n2134) );
  AND2_X2 U2452 ( .A1(n2381), .A2(n2382), .ZN(n2409) );
  OR2_X2 U2453 ( .A1(n2381), .A2(n2382), .ZN(n2406) );
  INV_X1 U2454 ( .A(n2393), .ZN(n2135) );
  NOR2_X2 U2455 ( .A1(n4355), .A2(n4343), .ZN(n4258) );
  NOR2_X2 U2456 ( .A1(n4159), .A2(n2204), .ZN(n4120) );
  OR2_X2 U2457 ( .A1(n4176), .A2(n4155), .ZN(n4159) );
  INV_X1 U2458 ( .A(n2968), .ZN(n2136) );
  NOR2_X2 U2459 ( .A1(n4270), .A2(n4271), .ZN(n4269) );
  BUF_X4 U2460 ( .A(n2541), .Z(n2137) );
  BUF_X4 U2461 ( .A(n2541), .Z(n2138) );
  NAND3_X2 U2462 ( .A1(n2188), .A2(n2187), .A3(n2186), .ZN(n2541) );
  AOI21_X1 U2463 ( .B1(n2362), .B2(n2300), .A(n2299), .ZN(n2298) );
  INV_X1 U2464 ( .A(n3613), .ZN(n2299) );
  AND2_X1 U2465 ( .A1(n3511), .A2(n2296), .ZN(n2295) );
  NAND2_X1 U2466 ( .A1(n3227), .A2(n3228), .ZN(n2286) );
  INV_X1 U2467 ( .A(n2335), .ZN(n2334) );
  NAND2_X1 U2468 ( .A1(n4119), .A2(n4105), .ZN(n2339) );
  INV_X1 U2469 ( .A(n2240), .ZN(n2239) );
  NOR2_X1 U2470 ( .A1(n2346), .A2(n2343), .ZN(n2342) );
  INV_X1 U2471 ( .A(n2468), .ZN(n2343) );
  INV_X1 U2472 ( .A(n2347), .ZN(n2346) );
  OR2_X1 U2473 ( .A1(n3027), .A2(n2976), .ZN(n3892) );
  OR2_X1 U2474 ( .A1(n4290), .A2(n4348), .ZN(n2224) );
  NOR2_X1 U2475 ( .A1(n3228), .A2(n3227), .ZN(n2287) );
  AND2_X1 U2476 ( .A1(n3594), .A2(n3004), .ZN(n2772) );
  NOR2_X1 U2477 ( .A1(n2836), .A2(n2837), .ZN(n2852) );
  XNOR2_X1 U2478 ( .A(n2897), .B(n2901), .ZN(n2855) );
  XNOR2_X1 U2479 ( .A(n3996), .B(n4558), .ZN(n4496) );
  NOR2_X1 U2480 ( .A1(n4517), .A2(REG1_REG_16__SCAN_IN), .ZN(n4516) );
  NOR2_X1 U2481 ( .A1(n2258), .A2(n4529), .ZN(n4528) );
  CLKBUF_X1 U2482 ( .A(n2406), .Z(n2872) );
  AND2_X1 U2483 ( .A1(n4101), .A2(n4115), .ZN(n2340) );
  NAND2_X1 U2484 ( .A1(n3485), .A2(n2162), .ZN(n2351) );
  AND2_X1 U2485 ( .A1(n2928), .A2(n2745), .ZN(n3003) );
  AND2_X1 U2486 ( .A1(n2677), .A2(n2234), .ZN(n2359) );
  AND2_X1 U2487 ( .A1(n2374), .A2(n2391), .ZN(n2234) );
  INV_X1 U2488 ( .A(IR_REG_17__SCAN_IN), .ZN(n2233) );
  AND2_X1 U2489 ( .A1(n3065), .A2(n3064), .ZN(n3066) );
  AOI21_X1 U2490 ( .B1(n4026), .B2(n2270), .A(n4043), .ZN(n2269) );
  INV_X1 U2491 ( .A(n2221), .ZN(n2217) );
  INV_X1 U2492 ( .A(n3832), .ZN(n2216) );
  INV_X1 U2493 ( .A(n2314), .ZN(n2313) );
  OAI21_X1 U2494 ( .B1(n2156), .B2(n2315), .A(n3583), .ZN(n2314) );
  NAND2_X1 U2495 ( .A1(n2289), .A2(n2288), .ZN(n3531) );
  AOI21_X1 U2496 ( .B1(n2290), .B2(n2294), .A(n2169), .ZN(n2288) );
  AND2_X1 U2497 ( .A1(n2293), .A2(n2291), .ZN(n2290) );
  NAND2_X1 U2498 ( .A1(n4509), .A2(n4023), .ZN(n4025) );
  INV_X1 U2499 ( .A(n2333), .ZN(n2332) );
  OAI21_X1 U2500 ( .B1(n2336), .B2(n2334), .A(n2644), .ZN(n2333) );
  NAND2_X1 U2501 ( .A1(n4281), .A2(n2643), .ZN(n2644) );
  AND2_X1 U2502 ( .A1(n2166), .A2(n3931), .ZN(n2244) );
  INV_X1 U2503 ( .A(n2190), .ZN(n2189) );
  INV_X1 U2504 ( .A(n2193), .ZN(n2192) );
  OAI21_X1 U2505 ( .B1(n2389), .B2(n2194), .A(n2392), .ZN(n2193) );
  INV_X1 U2506 ( .A(IR_REG_27__SCAN_IN), .ZN(n2390) );
  NOR2_X1 U2507 ( .A1(n2348), .A2(n2491), .ZN(n2347) );
  INV_X1 U2508 ( .A(n2477), .ZN(n2348) );
  NAND2_X1 U2509 ( .A1(n2446), .A2(n2328), .ZN(n2325) );
  AND2_X1 U2510 ( .A1(n3120), .A2(n2426), .ZN(n2356) );
  AND2_X1 U2511 ( .A1(n3437), .A2(n2157), .ZN(n2354) );
  NAND2_X1 U2512 ( .A1(n2671), .A2(n2359), .ZN(n2681) );
  INV_X1 U2513 ( .A(IR_REG_25__SCAN_IN), .ZN(n2725) );
  INV_X1 U2514 ( .A(IR_REG_23__SCAN_IN), .ZN(n2744) );
  NAND2_X1 U2515 ( .A1(n2306), .A2(n2161), .ZN(n3683) );
  INV_X1 U2516 ( .A(n2362), .ZN(n2296) );
  OR2_X1 U2517 ( .A1(n2514), .A2(n4631), .ZN(n2525) );
  AND2_X1 U2518 ( .A1(n2492), .A2(REG3_REG_10__SCAN_IN), .ZN(n2502) );
  OR2_X1 U2519 ( .A1(n2525), .A2(n3615), .ZN(n2543) );
  INV_X1 U2520 ( .A(IR_REG_1__SCAN_IN), .ZN(n2273) );
  XNOR2_X1 U2521 ( .A(n2830), .B(n2272), .ZN(n2820) );
  INV_X1 U2522 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2272) );
  NAND2_X1 U2523 ( .A1(n2181), .A2(n2180), .ZN(n2179) );
  NOR2_X1 U2524 ( .A1(n2851), .A2(n2842), .ZN(n2271) );
  NOR2_X1 U2525 ( .A1(n2885), .A2(n2163), .ZN(n2897) );
  NAND2_X1 U2526 ( .A1(n2264), .A2(n2263), .ZN(n4009) );
  OAI21_X1 U2527 ( .B1(n4008), .B2(REG1_REG_7__SCAN_IN), .A(n2265), .ZN(n2264)
         );
  NAND2_X1 U2528 ( .A1(n4441), .A2(n4011), .ZN(n4012) );
  NAND2_X1 U2529 ( .A1(n4462), .A2(n4015), .ZN(n4017) );
  NAND2_X1 U2530 ( .A1(n4489), .A2(n4019), .ZN(n4021) );
  NAND2_X1 U2531 ( .A1(n2262), .A2(n2261), .ZN(n3996) );
  NAND2_X1 U2532 ( .A1(n4559), .A2(n4748), .ZN(n2261) );
  OR2_X1 U2533 ( .A1(n4485), .A2(n2168), .ZN(n2262) );
  NOR2_X1 U2534 ( .A1(n4496), .A2(n4497), .ZN(n4495) );
  XNOR2_X1 U2535 ( .A(n4025), .B(n4024), .ZN(n4517) );
  NOR2_X1 U2536 ( .A1(n4504), .A2(n2246), .ZN(n3999) );
  AND2_X1 U2537 ( .A1(n4003), .A2(REG2_REG_15__SCAN_IN), .ZN(n2246) );
  INV_X1 U2538 ( .A(n2219), .ZN(n2218) );
  OAI21_X1 U2539 ( .B1(n4086), .B2(n2220), .A(n2711), .ZN(n2219) );
  NAND2_X1 U2540 ( .A1(n2710), .A2(n2709), .ZN(n2220) );
  NOR2_X1 U2541 ( .A1(n4086), .A2(n3834), .ZN(n2221) );
  NOR2_X1 U2542 ( .A1(n4113), .A2(n3846), .ZN(n4096) );
  AND2_X1 U2543 ( .A1(n2339), .A2(n2635), .ZN(n2336) );
  NAND2_X1 U2544 ( .A1(n2152), .A2(n2339), .ZN(n2335) );
  NOR2_X1 U2545 ( .A1(n2613), .A2(n4805), .ZN(n2617) );
  AND2_X1 U2546 ( .A1(n2588), .A2(n2577), .ZN(n2350) );
  INV_X1 U2547 ( .A(n4248), .ZN(n2588) );
  NOR2_X1 U2548 ( .A1(n2238), .A2(n2159), .ZN(n2237) );
  NAND2_X1 U2549 ( .A1(n2227), .A2(n2231), .ZN(n2226) );
  AOI21_X1 U2550 ( .B1(n2231), .B2(n2230), .A(n2229), .ZN(n2228) );
  INV_X1 U2551 ( .A(n3906), .ZN(n2229) );
  INV_X1 U2552 ( .A(n3907), .ZN(n2230) );
  NAND2_X1 U2553 ( .A1(n3144), .A2(n2468), .ZN(n3304) );
  INV_X1 U2554 ( .A(n2446), .ZN(n2327) );
  OR2_X1 U2555 ( .A1(n3121), .A2(n2685), .ZN(n2686) );
  NAND2_X1 U2556 ( .A1(n2742), .A2(n2816), .ZN(n2988) );
  NAND2_X1 U2557 ( .A1(n2720), .A2(n2223), .ZN(n4063) );
  AND2_X1 U2558 ( .A1(n2224), .A2(n2719), .ZN(n2223) );
  XNOR2_X1 U2559 ( .A(n2173), .B(n2172), .ZN(n4060) );
  INV_X1 U2560 ( .A(n3878), .ZN(n2172) );
  INV_X1 U2561 ( .A(n2661), .ZN(n2173) );
  NAND2_X1 U2562 ( .A1(n4072), .A2(n2762), .ZN(n4270) );
  INV_X1 U2563 ( .A(n4342), .ZN(n4273) );
  NAND2_X1 U2564 ( .A1(n2713), .A2(n3844), .ZN(n4254) );
  INV_X1 U2565 ( .A(n2976), .ZN(n3056) );
  NAND2_X1 U2566 ( .A1(n2676), .A2(n3003), .ZN(n3139) );
  NAND2_X1 U2567 ( .A1(n2722), .A2(n2725), .ZN(n2724) );
  INV_X1 U2568 ( .A(n2724), .ZN(n2727) );
  AND2_X1 U2569 ( .A1(n2194), .A2(n2725), .ZN(n2726) );
  INV_X1 U2570 ( .A(IR_REG_2__SCAN_IN), .ZN(n4825) );
  NOR2_X1 U2571 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2398)
         );
  CLKBUF_X1 U2572 ( .A(n2769), .Z(n2742) );
  INV_X1 U2573 ( .A(n4322), .ZN(n4194) );
  OR2_X1 U2574 ( .A1(n2285), .A2(n2147), .ZN(n2280) );
  OR2_X1 U2575 ( .A1(n2283), .A2(n2147), .ZN(n2279) );
  NAND2_X1 U2576 ( .A1(n2951), .A2(n2952), .ZN(n2953) );
  AND2_X1 U2577 ( .A1(n2472), .A2(n2471), .ZN(n3327) );
  INV_X1 U2578 ( .A(n2934), .ZN(n3729) );
  OAI21_X1 U2579 ( .B1(n3718), .B2(n2393), .A(n2634), .ZN(n4101) );
  INV_X1 U2580 ( .A(n3327), .ZN(n3983) );
  OR2_X1 U2581 ( .A1(n2406), .A2(n2405), .ZN(n2413) );
  OR2_X1 U2582 ( .A1(n2855), .A2(n3090), .ZN(n2896) );
  XNOR2_X1 U2583 ( .A(n4017), .B(n4560), .ZN(n4480) );
  NAND2_X1 U2584 ( .A1(n4480), .A2(REG1_REG_12__SCAN_IN), .ZN(n4479) );
  XNOR2_X1 U2585 ( .A(n3999), .B(n4024), .ZN(n4515) );
  NAND2_X1 U2586 ( .A1(n4515), .A2(n3460), .ZN(n4514) );
  OAI21_X1 U2587 ( .B1(n4528), .B2(n2256), .A(n2255), .ZN(n2254) );
  AOI21_X1 U2588 ( .B1(n4531), .B2(ADDR_REG_18__SCAN_IN), .A(n4530), .ZN(n2255) );
  INV_X1 U2589 ( .A(n2257), .ZN(n2256) );
  NAND2_X1 U2590 ( .A1(n2268), .A2(n2142), .ZN(n4532) );
  NAND2_X1 U2591 ( .A1(n4425), .A2(n2938), .ZN(n4538) );
  AND2_X1 U2592 ( .A1(n4425), .A2(n2790), .ZN(n4533) );
  NOR2_X1 U2593 ( .A1(n4063), .A2(n2199), .ZN(n2198) );
  NOR2_X1 U2594 ( .A1(n4061), .A2(n4239), .ZN(n2199) );
  OR2_X1 U2595 ( .A1(n4421), .A2(n4065), .ZN(n2195) );
  OR2_X1 U2596 ( .A1(n2988), .A2(n2932), .ZN(n4239) );
  OR2_X1 U2597 ( .A1(n4261), .A2(n3139), .ZN(n4238) );
  AOI21_X1 U2598 ( .B1(n4060), .B2(n4582), .A(n4063), .ZN(n2766) );
  NAND2_X1 U2599 ( .A1(n4270), .A2(n2200), .ZN(n4062) );
  OR2_X1 U2600 ( .A1(n4072), .A2(n2762), .ZN(n2200) );
  INV_X1 U2601 ( .A(IR_REG_29__SCAN_IN), .ZN(n2376) );
  INV_X1 U2602 ( .A(n3651), .ZN(n2291) );
  NAND2_X1 U2603 ( .A1(n2946), .A2(n2403), .ZN(n3889) );
  CLKBUF_X1 U2604 ( .A(n3604), .Z(n3553) );
  INV_X1 U2605 ( .A(n3692), .ZN(n2316) );
  OR2_X1 U2606 ( .A1(n2623), .A2(n3755), .ZN(n2629) );
  NAND2_X1 U2607 ( .A1(n4038), .A2(n2259), .ZN(n2258) );
  NAND2_X1 U2608 ( .A1(n4037), .A2(n2260), .ZN(n2259) );
  INV_X1 U2609 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2260) );
  AND2_X1 U2610 ( .A1(n4203), .A2(n2701), .ZN(n3940) );
  NAND2_X1 U2611 ( .A1(n2245), .A2(n2242), .ZN(n4204) );
  NOR2_X1 U2612 ( .A1(n2698), .A2(n2243), .ZN(n2242) );
  INV_X1 U2613 ( .A(n2244), .ZN(n2243) );
  NOR2_X1 U2614 ( .A1(n3927), .A2(n2239), .ZN(n2238) );
  AND2_X1 U2615 ( .A1(n2241), .A2(n3868), .ZN(n2240) );
  OR2_X1 U2616 ( .A1(n3150), .A2(n3062), .ZN(n3897) );
  AOI21_X1 U2617 ( .B1(n4096), .B2(n2215), .A(n2214), .ZN(n2712) );
  NOR2_X1 U2618 ( .A1(n2217), .A2(n2216), .ZN(n2215) );
  OAI21_X1 U2619 ( .B1(n2218), .B2(n2216), .A(n2654), .ZN(n2214) );
  NOR2_X1 U2620 ( .A1(n3440), .A2(n3520), .ZN(n2205) );
  OR2_X1 U2621 ( .A1(n2813), .A2(n2756), .ZN(n2924) );
  INV_X1 U2622 ( .A(IR_REG_28__SCAN_IN), .ZN(n2391) );
  INV_X1 U2623 ( .A(IR_REG_5__SCAN_IN), .ZN(n2304) );
  OR2_X1 U2624 ( .A1(n2550), .A2(IR_REG_14__SCAN_IN), .ZN(n2551) );
  INV_X1 U2625 ( .A(IR_REG_7__SCAN_IN), .ZN(n2464) );
  AOI22_X1 U2626 ( .A1(n2295), .A2(n3703), .B1(n2298), .B2(n2140), .ZN(n2293)
         );
  NOR2_X1 U2627 ( .A1(n2295), .A2(n2298), .ZN(n2294) );
  NAND2_X1 U2628 ( .A1(n3780), .A2(n3781), .ZN(n2307) );
  NAND2_X1 U2629 ( .A1(n2310), .A2(n2309), .ZN(n2308) );
  INV_X1 U2630 ( .A(n3781), .ZN(n2309) );
  INV_X1 U2631 ( .A(n3780), .ZN(n2310) );
  INV_X1 U2632 ( .A(n3259), .ZN(n2284) );
  INV_X1 U2633 ( .A(n2286), .ZN(n2285) );
  INV_X1 U2634 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4631) );
  NAND2_X1 U2635 ( .A1(n3664), .A2(n3581), .ZN(n3750) );
  AND2_X1 U2636 ( .A1(n3583), .A2(n3584), .ZN(n3581) );
  OAI21_X1 U2637 ( .B1(n3697), .B2(n2312), .A(n2313), .ZN(n3586) );
  NAND2_X1 U2638 ( .A1(n3575), .A2(n2167), .ZN(n2312) );
  INV_X1 U2639 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2478) );
  NAND2_X1 U2640 ( .A1(n3319), .A2(n3318), .ZN(n3321) );
  NAND2_X1 U2641 ( .A1(n2775), .A2(REG1_REG_0__SCAN_IN), .ZN(n2776) );
  NOR2_X1 U2642 ( .A1(n2742), .A2(n4428), .ZN(n2770) );
  AND2_X1 U2643 ( .A1(n2138), .A2(DATAI_20_), .ZN(n4216) );
  OR2_X1 U2644 ( .A1(n2570), .A2(n2569), .ZN(n2579) );
  INV_X1 U2645 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2578) );
  NOR2_X1 U2646 ( .A1(n2543), .A2(n2364), .ZN(n2558) );
  OR2_X1 U2647 ( .A1(n2928), .A2(n4412), .ZN(n2949) );
  XNOR2_X1 U2648 ( .A(n2851), .B(n2842), .ZN(n2836) );
  NOR2_X1 U2649 ( .A1(n2253), .A2(n2252), .ZN(n2251) );
  INV_X1 U2650 ( .A(n2849), .ZN(n2253) );
  NAND2_X1 U2651 ( .A1(n2250), .A2(n2849), .ZN(n2247) );
  INV_X1 U2652 ( .A(n2848), .ZN(n2250) );
  NAND2_X1 U2653 ( .A1(n4435), .A2(n4010), .ZN(n4443) );
  NAND2_X1 U2654 ( .A1(n4458), .A2(n4014), .ZN(n4464) );
  INV_X1 U2655 ( .A(n4028), .ZN(n2270) );
  AOI21_X1 U2656 ( .B1(n2258), .B2(n4529), .A(n4527), .ZN(n2257) );
  AOI21_X1 U2657 ( .B1(n2332), .B2(n2334), .A(n2164), .ZN(n2330) );
  AOI21_X1 U2658 ( .B1(n4184), .B2(n2707), .A(n2706), .ZN(n4129) );
  INV_X1 U2659 ( .A(n4160), .ZN(n4155) );
  OR2_X1 U2660 ( .A1(n2606), .A2(n3698), .ZN(n2613) );
  INV_X1 U2661 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4805) );
  INV_X1 U2662 ( .A(n4151), .ZN(n4170) );
  NAND2_X1 U2663 ( .A1(n2600), .A2(REG3_REG_20__SCAN_IN), .ZN(n2606) );
  AND2_X1 U2664 ( .A1(n2590), .A2(REG3_REG_19__SCAN_IN), .ZN(n2600) );
  NAND2_X1 U2665 ( .A1(n4245), .A2(n2589), .ZN(n4223) );
  NAND2_X1 U2666 ( .A1(n2245), .A2(n2244), .ZN(n4225) );
  AOI21_X1 U2667 ( .B1(n2354), .B2(n2139), .A(n2160), .ZN(n2353) );
  AOI22_X1 U2668 ( .A1(n2192), .A2(n2194), .B1(n2190), .B2(n2375), .ZN(n2186)
         );
  NAND2_X1 U2669 ( .A1(n2722), .A2(n2192), .ZN(n2187) );
  NAND2_X1 U2670 ( .A1(n2236), .A2(n2240), .ZN(n3435) );
  NAND2_X1 U2671 ( .A1(n3334), .A2(n3927), .ZN(n2236) );
  AOI21_X1 U2672 ( .B1(n2347), .B2(n2345), .A(n2149), .ZN(n2344) );
  INV_X1 U2673 ( .A(n2476), .ZN(n2345) );
  NAND2_X1 U2674 ( .A1(n2689), .A2(n3909), .ZN(n3216) );
  NAND2_X1 U2675 ( .A1(n2226), .A2(n2141), .ZN(n2689) );
  OR2_X1 U2676 ( .A1(n2469), .A2(n4633), .ZN(n2479) );
  INV_X1 U2677 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4633) );
  OR2_X1 U2678 ( .A1(n2454), .A2(n2327), .ZN(n2326) );
  INV_X1 U2679 ( .A(n2324), .ZN(n2323) );
  OAI22_X1 U2680 ( .A1(n2454), .A2(n2325), .B1(n3239), .B2(n3167), .ZN(n2324)
         );
  NOR2_X1 U2681 ( .A1(n2447), .A2(n2857), .ZN(n2455) );
  NAND2_X1 U2682 ( .A1(n2455), .A2(REG3_REG_7__SCAN_IN), .ZN(n2469) );
  INV_X1 U2683 ( .A(n3236), .ZN(n3231) );
  NAND2_X1 U2684 ( .A1(n2687), .A2(n3903), .ZN(n3135) );
  NAND2_X1 U2685 ( .A1(n2209), .A2(n2143), .ZN(n2687) );
  AOI21_X1 U2686 ( .B1(n3914), .B2(n2212), .A(n2211), .ZN(n2210) );
  INV_X1 U2687 ( .A(n3901), .ZN(n2212) );
  INV_X1 U2688 ( .A(n3900), .ZN(n2211) );
  NAND2_X1 U2689 ( .A1(n2207), .A2(n3914), .ZN(n2209) );
  INV_X1 U2690 ( .A(n2686), .ZN(n2207) );
  AND2_X1 U2691 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2436) );
  NAND2_X1 U2692 ( .A1(n2357), .A2(n2426), .ZN(n3124) );
  NAND2_X1 U2693 ( .A1(n2176), .A2(n2404), .ZN(n3045) );
  NAND2_X1 U2694 ( .A1(n3892), .A2(n3895), .ZN(n3044) );
  OAI21_X1 U2695 ( .B1(n3888), .B2(n2320), .A(n3891), .ZN(n3047) );
  INV_X1 U2696 ( .A(n2320), .ZN(n3860) );
  AND2_X1 U2697 ( .A1(n2924), .A2(n2923), .ZN(n2992) );
  NOR2_X1 U2698 ( .A1(n2144), .A2(n4277), .ZN(n4072) );
  AND2_X1 U2699 ( .A1(n2653), .A2(n2652), .ZN(n4290) );
  NAND2_X1 U2700 ( .A1(n4120), .A2(n4105), .ZN(n4104) );
  NAND2_X1 U2701 ( .A1(n4140), .A2(n4122), .ZN(n2204) );
  NOR2_X1 U2702 ( .A1(n4159), .A2(n4302), .ZN(n4135) );
  INV_X1 U2703 ( .A(n4348), .ZN(n4303) );
  NAND2_X1 U2704 ( .A1(n4189), .A2(n4177), .ZN(n4176) );
  NAND2_X1 U2705 ( .A1(n2137), .A2(DATAI_22_), .ZN(n4177) );
  NOR2_X1 U2706 ( .A1(n4235), .A2(n4216), .ZN(n4215) );
  AND2_X1 U2707 ( .A1(n4215), .A2(n4195), .ZN(n4189) );
  NAND2_X1 U2708 ( .A1(n4258), .A2(n4257), .ZN(n4256) );
  OR2_X1 U2709 ( .A1(n4256), .A2(n3686), .ZN(n4235) );
  NAND2_X1 U2710 ( .A1(n2205), .A2(n2567), .ZN(n4355) );
  INV_X1 U2711 ( .A(n2205), .ZN(n3457) );
  NAND2_X1 U2712 ( .A1(n3441), .A2(n3515), .ZN(n3440) );
  NAND2_X1 U2713 ( .A1(n2355), .A2(n2354), .ZN(n3433) );
  AND2_X1 U2714 ( .A1(n2355), .A2(n2157), .ZN(n3434) );
  OR2_X1 U2715 ( .A1(n3366), .A2(n2139), .ZN(n2355) );
  NOR2_X1 U2716 ( .A1(n2201), .A2(n3494), .ZN(n3441) );
  NAND2_X1 U2717 ( .A1(n3217), .A2(n2158), .ZN(n3338) );
  INV_X1 U2718 ( .A(n4254), .ZN(n4233) );
  NAND2_X1 U2719 ( .A1(n3217), .A2(n3397), .ZN(n3289) );
  INV_X1 U2720 ( .A(n3671), .ZN(n3397) );
  AND2_X1 U2721 ( .A1(n3300), .A2(n3328), .ZN(n3217) );
  OR2_X1 U2722 ( .A1(n3140), .A2(n3231), .ZN(n3299) );
  NOR2_X1 U2723 ( .A1(n3299), .A2(n3306), .ZN(n3300) );
  INV_X1 U2724 ( .A(n3167), .ZN(n3193) );
  NAND2_X1 U2725 ( .A1(n3119), .A2(n3123), .ZN(n3118) );
  NOR2_X1 U2726 ( .A1(n3118), .A2(n3108), .ZN(n3085) );
  INV_X1 U2727 ( .A(n3176), .ZN(n3108) );
  AND2_X1 U2728 ( .A1(n3003), .A2(n4411), .ZN(n4342) );
  INV_X1 U2729 ( .A(n4307), .ZN(n4344) );
  INV_X1 U2730 ( .A(n3139), .ZN(n4354) );
  INV_X1 U2731 ( .A(n2990), .ZN(n2925) );
  INV_X1 U2732 ( .A(n4579), .ZN(n4565) );
  INV_X1 U2733 ( .A(n2739), .ZN(n2759) );
  NAND2_X1 U2734 ( .A1(n2733), .A2(IR_REG_31__SCAN_IN), .ZN(n2735) );
  XNOR2_X1 U2735 ( .A(n2743), .B(n2744), .ZN(n3069) );
  NAND2_X1 U2736 ( .A1(n2672), .A2(n2673), .ZN(n2745) );
  INV_X1 U2737 ( .A(n2440), .ZN(n2301) );
  AND2_X1 U2738 ( .A1(n2302), .A2(n2370), .ZN(n2235) );
  INV_X1 U2739 ( .A(IR_REG_11__SCAN_IN), .ZN(n2510) );
  AND2_X1 U2740 ( .A1(n2486), .A2(n2366), .ZN(n2305) );
  INV_X1 U2741 ( .A(IR_REG_4__SCAN_IN), .ZN(n4826) );
  INV_X1 U2742 ( .A(IR_REG_3__SCAN_IN), .ZN(n2422) );
  INV_X1 U2743 ( .A(n2281), .ZN(n3260) );
  AOI21_X1 U2744 ( .B1(n3229), .B2(n2282), .A(n2285), .ZN(n2281) );
  INV_X1 U2745 ( .A(n2287), .ZN(n2282) );
  AOI21_X1 U2746 ( .B1(n3788), .B2(n3790), .A(n3789), .ZN(n3626) );
  NAND2_X1 U2747 ( .A1(n2292), .A2(n2293), .ZN(n3653) );
  OR2_X1 U2748 ( .A1(n3510), .A2(n2294), .ZN(n2292) );
  NAND2_X1 U2749 ( .A1(n2138), .A2(DATAI_23_), .ZN(n4160) );
  INV_X1 U2750 ( .A(n3670), .ZN(n3708) );
  NAND2_X1 U2751 ( .A1(n2138), .A2(DATAI_25_), .ZN(n4122) );
  INV_X1 U2752 ( .A(n2276), .ZN(n2275) );
  NAND2_X1 U2753 ( .A1(n3155), .A2(n3107), .ZN(n3113) );
  OR2_X1 U2754 ( .A1(n2959), .A2(n2939), .ZN(n3795) );
  NAND2_X1 U2755 ( .A1(n3510), .A2(n3509), .ZN(n2297) );
  NAND2_X1 U2756 ( .A1(n2317), .A2(n3692), .ZN(n3772) );
  NAND2_X1 U2757 ( .A1(n2971), .A2(n2970), .ZN(n2972) );
  INV_X1 U2758 ( .A(n2969), .ZN(n2970) );
  AOI21_X1 U2759 ( .B1(n3740), .B2(n3737), .A(n3736), .ZN(n3783) );
  NAND2_X1 U2760 ( .A1(n2137), .A2(DATAI_26_), .ZN(n4105) );
  OR2_X1 U2761 ( .A1(n2959), .A2(n2937), .ZN(n3800) );
  INV_X1 U2762 ( .A(n3800), .ZN(n3805) );
  INV_X1 U2763 ( .A(n3795), .ZN(n3811) );
  INV_X1 U2764 ( .A(n4412), .ZN(n4050) );
  OAI211_X1 U2765 ( .C1(n2872), .C2(n4314), .A(n2620), .B(n2619), .ZN(n4304)
         );
  OAI211_X1 U2766 ( .C1(n2393), .C2(n4178), .A(n2616), .B(n2615), .ZN(n4322)
         );
  NAND4_X1 U2767 ( .A1(n2611), .A2(n2610), .A3(n2609), .A4(n2608), .ZN(n4206)
         );
  NAND4_X1 U2768 ( .A1(n2497), .A2(n2496), .A3(n2495), .A4(n2494), .ZN(n3399)
         );
  CLKBUF_X2 U2769 ( .A(U4043), .Z(n3985) );
  NAND2_X1 U2770 ( .A1(n2194), .A2(n2273), .ZN(n2183) );
  AOI21_X1 U2771 ( .B1(n2182), .B2(n2853), .A(n2913), .ZN(n2887) );
  NAND2_X1 U2772 ( .A1(n2909), .A2(REG2_REG_4__SCAN_IN), .ZN(n2249) );
  NAND2_X1 U2773 ( .A1(n2444), .A2(n2443), .ZN(n2891) );
  NAND2_X1 U2774 ( .A1(n2267), .A2(n2854), .ZN(n2266) );
  INV_X1 U2775 ( .A(n4600), .ZN(n4439) );
  XNOR2_X1 U2776 ( .A(n4009), .B(n4439), .ZN(n4436) );
  NAND2_X1 U2777 ( .A1(n4436), .A2(REG1_REG_8__SCAN_IN), .ZN(n4435) );
  XNOR2_X1 U2778 ( .A(n4012), .B(n4561), .ZN(n4459) );
  NAND2_X1 U2779 ( .A1(n4459), .A2(REG1_REG_10__SCAN_IN), .ZN(n4458) );
  NAND2_X1 U2780 ( .A1(n4479), .A2(n4018), .ZN(n4490) );
  NAND2_X1 U2781 ( .A1(n4500), .A2(n4022), .ZN(n4510) );
  NAND2_X1 U2782 ( .A1(n4510), .A2(n4511), .ZN(n4509) );
  NOR2_X1 U2783 ( .A1(n3997), .A2(n4495), .ZN(n4506) );
  AND2_X1 U2784 ( .A1(n2795), .A2(n2794), .ZN(n4531) );
  AND2_X1 U2785 ( .A1(n4425), .A2(n3966), .ZN(n4522) );
  NOR2_X1 U2786 ( .A1(n4029), .A2(n4028), .ZN(n4042) );
  NOR2_X1 U2787 ( .A1(n4516), .A2(n4026), .ZN(n4029) );
  NAND2_X1 U2788 ( .A1(n4000), .A2(n4514), .ZN(n4001) );
  INV_X1 U2789 ( .A(n4522), .ZN(n4527) );
  NAND2_X1 U2790 ( .A1(n2213), .A2(n2218), .ZN(n4066) );
  NAND2_X1 U2791 ( .A1(n4096), .A2(n2221), .ZN(n2213) );
  OAI21_X1 U2792 ( .B1(n4096), .B2(n2710), .A(n2709), .ZN(n4083) );
  INV_X1 U2793 ( .A(n4287), .ZN(n4119) );
  NAND2_X1 U2794 ( .A1(n2331), .A2(n2335), .ZN(n4085) );
  INV_X1 U2795 ( .A(n2340), .ZN(n2337) );
  NAND2_X1 U2796 ( .A1(n4111), .A2(n2635), .ZN(n2338) );
  NAND2_X1 U2797 ( .A1(n2351), .A2(n2577), .ZN(n4247) );
  NAND2_X1 U2798 ( .A1(n2245), .A2(n3931), .ZN(n3483) );
  NAND4_X1 U2799 ( .A1(n2519), .A2(n2518), .A3(n2517), .A4(n2516), .ZN(n3981)
         );
  NAND2_X1 U2800 ( .A1(n2226), .A2(n2228), .ZN(n3211) );
  NAND2_X1 U2801 ( .A1(n2349), .A2(n2477), .ZN(n3204) );
  NAND2_X1 U2802 ( .A1(n3304), .A2(n2476), .ZN(n2349) );
  AND2_X1 U2803 ( .A1(n4421), .A2(n3147), .ZN(n4188) );
  INV_X1 U2804 ( .A(n2322), .ZN(n3080) );
  AOI21_X1 U2805 ( .B1(n3013), .B2(n2445), .A(n2327), .ZN(n2322) );
  NAND2_X1 U2806 ( .A1(n2686), .A2(n3901), .ZN(n3015) );
  INV_X1 U2807 ( .A(n4238), .ZN(n4543) );
  INV_X1 U2808 ( .A(n4239), .ZN(n4539) );
  OR2_X1 U2809 ( .A1(n2765), .A2(n2990), .ZN(n4596) );
  INV_X2 U2810 ( .A(n4596), .ZN(n4599) );
  NAND2_X1 U2811 ( .A1(n3024), .A2(n2202), .ZN(n3039) );
  INV_X1 U2812 ( .A(n3119), .ZN(n2202) );
  INV_X1 U2813 ( .A(n4551), .ZN(n2816) );
  NAND2_X1 U2814 ( .A1(n2379), .A2(IR_REG_31__SCAN_IN), .ZN(n2377) );
  NAND2_X1 U2815 ( .A1(n2191), .A2(IR_REG_31__SCAN_IN), .ZN(n2718) );
  NAND2_X1 U2816 ( .A1(n2722), .A2(n2389), .ZN(n2191) );
  NOR2_X1 U2817 ( .A1(n2727), .A2(n2726), .ZN(n2728) );
  OAI21_X1 U2818 ( .B1(n2511), .B2(n2510), .A(n2520), .ZN(n4470) );
  OR2_X1 U2819 ( .A1(n2398), .A2(n2194), .ZN(n2414) );
  INV_X1 U2820 ( .A(n2254), .ZN(n4536) );
  NAND2_X1 U2821 ( .A1(n2196), .A2(n2148), .ZN(U3354) );
  NAND2_X1 U2822 ( .A1(n2197), .A2(n4421), .ZN(n2196) );
  OAI21_X1 U2823 ( .B1(n4062), .B2(n4238), .A(n2198), .ZN(n2197) );
  OR2_X1 U2824 ( .A1(n4062), .A2(n4338), .ZN(n2763) );
  INV_X4 U2825 ( .A(n2406), .ZN(n2457) );
  NOR2_X1 U2826 ( .A1(n3980), .A2(n3494), .ZN(n2139) );
  OR2_X1 U2827 ( .A1(n3703), .A2(n3511), .ZN(n2140) );
  AND2_X1 U2828 ( .A1(n2228), .A2(n2225), .ZN(n2141) );
  AND2_X1 U2829 ( .A1(n2269), .A2(n4534), .ZN(n2142) );
  AND2_X1 U2830 ( .A1(n2210), .A2(n2208), .ZN(n2143) );
  NOR2_X1 U2831 ( .A1(n2834), .A2(n2150), .ZN(n2851) );
  OAI21_X1 U2832 ( .B1(n2137), .B2(n4428), .A(n2402), .ZN(n3004) );
  INV_X1 U2833 ( .A(n3575), .ZN(n2315) );
  INV_X1 U2834 ( .A(n3511), .ZN(n2300) );
  OR2_X1 U2835 ( .A1(n4104), .A2(n4286), .ZN(n2144) );
  NOR2_X1 U2836 ( .A1(n2440), .A2(IR_REG_5__SCAN_IN), .ZN(n2442) );
  INV_X1 U2837 ( .A(n2393), .ZN(n2581) );
  INV_X1 U2838 ( .A(n2393), .ZN(n2407) );
  INV_X1 U2839 ( .A(n2912), .ZN(n2182) );
  AND2_X1 U2840 ( .A1(n3897), .A2(n3894), .ZN(n2145) );
  NAND4_X1 U2841 ( .A1(n2431), .A2(n2430), .A3(n2429), .A4(n2428), .ZN(n3099)
         );
  AND2_X1 U2842 ( .A1(n2432), .A2(n2424), .ZN(n4416) );
  NOR2_X1 U2843 ( .A1(IR_REG_25__SCAN_IN), .A2(IR_REG_26__SCAN_IN), .ZN(n2389)
         );
  BUF_X1 U2844 ( .A(n2948), .Z(n2946) );
  NAND4_X1 U2845 ( .A1(n2397), .A2(n2396), .A3(n2395), .A4(n2394), .ZN(n2948)
         );
  AND2_X1 U2846 ( .A1(n4287), .A2(n4100), .ZN(n2146) );
  NOR2_X1 U2847 ( .A1(n3258), .A2(n3257), .ZN(n2147) );
  NAND3_X1 U2848 ( .A1(n2358), .A2(n2206), .A3(n4428), .ZN(n2440) );
  XNOR2_X1 U2849 ( .A(n2377), .B(IR_REG_30__SCAN_IN), .ZN(n2381) );
  INV_X1 U2850 ( .A(n3123), .ZN(n3151) );
  NAND2_X1 U2851 ( .A1(n2398), .A2(n4825), .ZN(n2421) );
  AND2_X1 U2852 ( .A1(n4064), .A2(n2195), .ZN(n2148) );
  AND2_X1 U2853 ( .A1(n3673), .A2(n3328), .ZN(n2149) );
  AND2_X1 U2854 ( .A1(n2835), .A2(REG1_REG_2__SCAN_IN), .ZN(n2150) );
  AND2_X1 U2855 ( .A1(n2268), .A2(n2269), .ZN(n2151) );
  OR2_X1 U2856 ( .A1(n2146), .A2(n2340), .ZN(n2152) );
  AND2_X1 U2857 ( .A1(n2338), .A2(n2337), .ZN(n2153) );
  INV_X1 U2858 ( .A(n3107), .ZN(n2277) );
  AND2_X1 U2859 ( .A1(n3400), .A2(n3392), .ZN(n2154) );
  AND2_X1 U2860 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2155)
         );
  NAND2_X1 U2861 ( .A1(n2442), .A2(n2305), .ZN(n2489) );
  INV_X1 U2862 ( .A(n3915), .ZN(n2208) );
  NAND2_X1 U2863 ( .A1(n3675), .A2(n3404), .ZN(n3498) );
  AND2_X1 U2864 ( .A1(n2297), .A2(n2296), .ZN(n3612) );
  NOR2_X1 U2865 ( .A1(n3773), .A2(n2316), .ZN(n2156) );
  NAND2_X1 U2866 ( .A1(n3980), .A2(n3494), .ZN(n2157) );
  NAND2_X1 U2867 ( .A1(n2306), .A2(n2307), .ZN(n3682) );
  INV_X1 U2868 ( .A(n3703), .ZN(n3509) );
  AND2_X1 U2869 ( .A1(n3397), .A2(n3409), .ZN(n2158) );
  INV_X1 U2870 ( .A(n2567), .ZN(n3728) );
  OR2_X1 U2871 ( .A1(n3866), .A2(n2695), .ZN(n2159) );
  AND2_X1 U2872 ( .A1(n3808), .A2(n3515), .ZN(n2160) );
  AND2_X1 U2873 ( .A1(n3548), .A2(n2307), .ZN(n2161) );
  NAND2_X1 U2874 ( .A1(n4250), .A2(n3742), .ZN(n2162) );
  AND2_X1 U2875 ( .A1(n4415), .A2(REG1_REG_5__SCAN_IN), .ZN(n2163) );
  AND2_X1 U2876 ( .A1(n4290), .A2(n4277), .ZN(n3836) );
  INV_X1 U2877 ( .A(n2321), .ZN(n3888) );
  AND2_X1 U2878 ( .A1(n2960), .A2(n3004), .ZN(n2321) );
  NOR2_X1 U2879 ( .A1(n4281), .A2(n2643), .ZN(n2164) );
  OR2_X1 U2880 ( .A1(n2891), .A2(n2850), .ZN(n2165) );
  NAND2_X1 U2881 ( .A1(n3976), .A2(n3742), .ZN(n2166) );
  NAND2_X1 U2882 ( .A1(n2732), .A2(IR_REG_31__SCAN_IN), .ZN(n2743) );
  INV_X1 U2883 ( .A(n4020), .ZN(n4558) );
  XNOR2_X1 U2884 ( .A(n2735), .B(n2734), .ZN(n2738) );
  INV_X1 U2885 ( .A(n3917), .ZN(n2225) );
  NAND2_X1 U2886 ( .A1(n3393), .A2(n3392), .ZN(n3674) );
  NAND2_X1 U2887 ( .A1(n2278), .A2(n3103), .ZN(n3155) );
  NAND2_X1 U2888 ( .A1(n2235), .A2(n2301), .ZN(n2574) );
  NAND2_X1 U2889 ( .A1(n3564), .A2(n3565), .ZN(n2167) );
  AND2_X1 U2890 ( .A1(n2535), .A2(n2550), .ZN(n4483) );
  AND2_X1 U2891 ( .A1(n4483), .A2(REG2_REG_13__SCAN_IN), .ZN(n2168) );
  INV_X2 U2892 ( .A(n4587), .ZN(n4589) );
  AND2_X1 U2893 ( .A1(n3518), .A2(n3517), .ZN(n2169) );
  INV_X1 U2894 ( .A(n4140), .ZN(n4302) );
  INV_X1 U2895 ( .A(n2742), .ZN(n2775) );
  INV_X1 U2896 ( .A(n2445), .ZN(n2328) );
  AND2_X1 U2897 ( .A1(n2249), .A2(n2848), .ZN(n2170) );
  OR2_X1 U2898 ( .A1(n4589), .A2(n4716), .ZN(n2171) );
  INV_X1 U2899 ( .A(n4414), .ZN(n2265) );
  INV_X1 U2900 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2252) );
  NAND4_X1 U2901 ( .A1(n2401), .A2(n2175), .A3(n2174), .A4(n2400), .ZN(n2773)
         );
  NAND2_X1 U2902 ( .A1(n2409), .A2(REG2_REG_0__SCAN_IN), .ZN(n2174) );
  NAND2_X1 U2903 ( .A1(n2407), .A2(REG3_REG_0__SCAN_IN), .ZN(n2175) );
  NAND2_X1 U2904 ( .A1(n2318), .A2(n2176), .ZN(n2996) );
  NAND2_X1 U2905 ( .A1(n2876), .A2(n2320), .ZN(n2176) );
  NAND3_X1 U2906 ( .A1(n2671), .A2(n2359), .A3(n2376), .ZN(n2379) );
  NAND2_X1 U2907 ( .A1(n2181), .A2(n2177), .ZN(n2853) );
  INV_X1 U2908 ( .A(n2271), .ZN(n2177) );
  NAND2_X1 U2909 ( .A1(n2179), .A2(n2178), .ZN(n2914) );
  OAI21_X1 U2910 ( .B1(n2852), .B2(n2271), .A(n2182), .ZN(n2178) );
  NOR2_X1 U2911 ( .A1(n2271), .A2(n2182), .ZN(n2180) );
  INV_X1 U2912 ( .A(n2852), .ZN(n2181) );
  NOR2_X1 U2913 ( .A1(n2820), .A2(n2821), .ZN(n2819) );
  INV_X1 U2914 ( .A(n2398), .ZN(n2184) );
  NAND2_X1 U2915 ( .A1(n2155), .A2(IR_REG_0__SCAN_IN), .ZN(n2185) );
  INV_X1 U2916 ( .A(n2201), .ZN(n3367) );
  AND2_X2 U2917 ( .A1(n3062), .A2(n3054), .ZN(n3119) );
  INV_X2 U2918 ( .A(n2203), .ZN(n2671) );
  NAND4_X1 U2919 ( .A1(n2302), .A2(n2301), .A3(n2370), .A4(n2233), .ZN(n2203)
         );
  NAND2_X1 U2920 ( .A1(n2209), .A2(n2210), .ZN(n3081) );
  NAND3_X1 U2921 ( .A1(n2222), .A2(n2767), .A3(n2171), .ZN(U3515) );
  INV_X1 U2922 ( .A(n3135), .ZN(n2227) );
  OAI21_X1 U2923 ( .B1(n3135), .B2(n2688), .A(n3907), .ZN(n3305) );
  AOI21_X1 U2924 ( .B1(n2688), .B2(n3907), .A(n2232), .ZN(n2231) );
  INV_X1 U2925 ( .A(n3908), .ZN(n2232) );
  OAI21_X1 U2926 ( .B1(n3334), .B2(n2239), .A(n2237), .ZN(n2696) );
  OAI21_X1 U2927 ( .B1(n3334), .B2(n2692), .A(n3927), .ZN(n3821) );
  NAND2_X1 U2928 ( .A1(n3927), .A2(n2692), .ZN(n2241) );
  NAND2_X1 U2929 ( .A1(n3452), .A2(n3869), .ZN(n2245) );
  NAND2_X1 U2930 ( .A1(n2909), .A2(n2251), .ZN(n2248) );
  NAND3_X1 U2931 ( .A1(n2247), .A2(n2165), .A3(n2248), .ZN(n2900) );
  NAND2_X1 U2932 ( .A1(n2247), .A2(n2248), .ZN(n2888) );
  NAND2_X1 U2933 ( .A1(n4008), .A2(REG1_REG_7__SCAN_IN), .ZN(n2263) );
  INV_X1 U2934 ( .A(n2897), .ZN(n2267) );
  NAND2_X1 U2935 ( .A1(n4516), .A2(n2270), .ZN(n2268) );
  INV_X1 U2936 ( .A(n3154), .ZN(n2278) );
  NAND2_X1 U2937 ( .A1(n2275), .A2(n2274), .ZN(n3164) );
  NAND2_X1 U2938 ( .A1(n3154), .A2(n3107), .ZN(n2274) );
  OAI21_X1 U2939 ( .B1(n3103), .B2(n2277), .A(n3112), .ZN(n2276) );
  NAND2_X1 U2940 ( .A1(n3510), .A2(n2290), .ZN(n2289) );
  NAND2_X1 U2941 ( .A1(n3393), .A2(n2154), .ZN(n3675) );
  NAND2_X1 U2942 ( .A1(n3783), .A2(n2308), .ZN(n2306) );
  INV_X1 U2943 ( .A(n3697), .ZN(n2311) );
  NAND2_X1 U2944 ( .A1(n2317), .A2(n2156), .ZN(n3661) );
  AND2_X2 U2945 ( .A1(n2671), .A2(n2374), .ZN(n2722) );
  NAND2_X1 U2946 ( .A1(n2319), .A2(n3860), .ZN(n2318) );
  INV_X1 U2947 ( .A(n2876), .ZN(n2319) );
  XNOR2_X1 U2948 ( .A(n2321), .B(n3860), .ZN(n2880) );
  OAI21_X1 U2949 ( .B1(n3013), .B2(n2326), .A(n2323), .ZN(n3145) );
  INV_X1 U2950 ( .A(n3145), .ZN(n2467) );
  NAND2_X1 U2951 ( .A1(n4111), .A2(n2332), .ZN(n2329) );
  NAND2_X1 U2952 ( .A1(n2329), .A2(n2330), .ZN(n4070) );
  NAND2_X1 U2953 ( .A1(n4111), .A2(n2336), .ZN(n2331) );
  NAND2_X1 U2954 ( .A1(n3144), .A2(n2342), .ZN(n2341) );
  NAND2_X1 U2955 ( .A1(n2341), .A2(n2344), .ZN(n3222) );
  NAND2_X1 U2956 ( .A1(n3366), .A2(n2354), .ZN(n2352) );
  NAND2_X1 U2957 ( .A1(n2352), .A2(n2353), .ZN(n3422) );
  NAND2_X1 U2958 ( .A1(n3025), .A2(n2425), .ZN(n2357) );
  NAND2_X1 U2959 ( .A1(n2357), .A2(n2356), .ZN(n3126) );
  NAND2_X1 U2960 ( .A1(n2541), .A2(DATAI_0_), .ZN(n2402) );
  OAI21_X1 U2961 ( .B1(n2968), .B2(n2960), .A(n2771), .ZN(n2778) );
  OAI21_X1 U2962 ( .B1(n3498), .B2(n3497), .A(n3496), .ZN(n3499) );
  AOI21_X2 U2963 ( .B1(n3717), .B2(n3713), .A(n3715), .ZN(n3788) );
  OAI22_X1 U2964 ( .A1(n3097), .A2(n3096), .B1(n3095), .B2(n3094), .ZN(n3154)
         );
  NAND2_X1 U2965 ( .A1(n4589), .A2(n4354), .ZN(n4406) );
  OR2_X1 U2966 ( .A1(n4194), .A2(n4177), .ZN(n2361) );
  AND2_X1 U2967 ( .A1(n2138), .A2(DATAI_27_), .ZN(n4286) );
  AND2_X1 U2968 ( .A1(n3508), .A2(n3507), .ZN(n2362) );
  AOI21_X1 U2969 ( .B1(n2773), .B2(n3604), .A(n2772), .ZN(n2951) );
  NOR2_X1 U2970 ( .A1(n2974), .A2(n2975), .ZN(n3067) );
  NAND2_X1 U2971 ( .A1(n2777), .A2(n2778), .ZN(n2954) );
  AND2_X1 U2972 ( .A1(n2388), .A2(n2387), .ZN(n4281) );
  INV_X1 U2973 ( .A(n3389), .ZN(n3390) );
  INV_X1 U2974 ( .A(n3388), .ZN(n3391) );
  NAND2_X1 U2975 ( .A1(n3391), .A2(n3390), .ZN(n3392) );
  INV_X1 U2976 ( .A(n4286), .ZN(n2643) );
  INV_X1 U2977 ( .A(IR_REG_24__SCAN_IN), .ZN(n2734) );
  INV_X1 U2978 ( .A(n3624), .ZN(n2740) );
  INV_X1 U2979 ( .A(n3677), .ZN(n3400) );
  AOI21_X1 U2980 ( .B1(n3004), .B2(n3604), .A(n2770), .ZN(n2771) );
  INV_X1 U2981 ( .A(IR_REG_6__SCAN_IN), .ZN(n2462) );
  INV_X1 U2982 ( .A(n3685), .ZN(n3548) );
  INV_X1 U2983 ( .A(n3105), .ZN(n3106) );
  INV_X1 U2984 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2569) );
  NOR2_X1 U2985 ( .A1(n2629), .A2(n3719), .ZN(n2636) );
  INV_X1 U2986 ( .A(n2409), .ZN(n2505) );
  AND2_X1 U2987 ( .A1(n4281), .A2(n4286), .ZN(n3835) );
  AND2_X1 U2988 ( .A1(n4158), .A2(n4140), .ZN(n2627) );
  AND2_X1 U2989 ( .A1(n4304), .A2(n4155), .ZN(n2621) );
  INV_X1 U2990 ( .A(n2363), .ZN(n2466) );
  INV_X1 U2991 ( .A(n3742), .ZN(n4343) );
  NAND2_X1 U2992 ( .A1(n2636), .A2(REG3_REG_26__SCAN_IN), .ZN(n2646) );
  NAND2_X1 U2993 ( .A1(n2558), .A2(REG3_REG_16__SCAN_IN), .ZN(n2570) );
  NAND2_X1 U2994 ( .A1(n3104), .A2(n3106), .ZN(n3107) );
  NOR2_X1 U2995 ( .A1(n2579), .A2(n2578), .ZN(n2590) );
  OR2_X1 U2996 ( .A1(n2959), .A2(n2958), .ZN(n3807) );
  NOR2_X1 U2997 ( .A1(n3630), .A2(n2929), .ZN(n3967) );
  OR2_X1 U2998 ( .A1(n3793), .A2(n2393), .ZN(n2642) );
  INV_X1 U2999 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2857) );
  INV_X1 U3000 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3615) );
  OR3_X1 U3001 ( .A1(n2646), .A2(n3607), .A3(n2645), .ZN(n4061) );
  OR2_X1 U3002 ( .A1(n3951), .A2(n3835), .ZN(n4086) );
  AND2_X1 U3003 ( .A1(n4149), .A2(n2704), .ZN(n4151) );
  INV_X1 U3004 ( .A(n4345), .ZN(n3741) );
  OR2_X1 U3005 ( .A1(n2813), .A2(D_REG_1__SCAN_IN), .ZN(n2989) );
  OR2_X1 U3006 ( .A1(n2813), .A2(D_REG_0__SCAN_IN), .ZN(n2760) );
  AND2_X1 U3007 ( .A1(n2137), .A2(DATAI_28_), .ZN(n4277) );
  INV_X1 U3008 ( .A(n3494), .ZN(n3617) );
  INV_X1 U3009 ( .A(n3302), .ZN(n3306) );
  OR2_X1 U3010 ( .A1(n2938), .A2(n2922), .ZN(n4348) );
  NAND2_X1 U3011 ( .A1(n2675), .A2(n4050), .ZN(n4210) );
  OR2_X1 U3012 ( .A1(n2534), .A2(IR_REG_13__SCAN_IN), .ZN(n2550) );
  OR2_X1 U3013 ( .A1(n2463), .A2(n2194), .ZN(n2465) );
  AOI21_X1 U3014 ( .B1(n3529), .B2(n3528), .A(n3533), .ZN(n3727) );
  NAND2_X1 U3015 ( .A1(n2436), .A2(REG3_REG_5__SCAN_IN), .ZN(n2447) );
  NOR2_X1 U3016 ( .A1(n2479), .A2(n2478), .ZN(n2492) );
  NAND2_X1 U3017 ( .A1(n2502), .A2(REG3_REG_11__SCAN_IN), .ZN(n2514) );
  INV_X1 U3018 ( .A(n3807), .ZN(n3744) );
  OAI21_X1 U3019 ( .B1(n3073), .B2(U3149), .A(n3072), .ZN(n3798) );
  NAND2_X1 U3020 ( .A1(n2642), .A2(n2641), .ZN(n4287) );
  AND2_X1 U3021 ( .A1(n2573), .A2(n2572), .ZN(n4250) );
  NAND2_X1 U3022 ( .A1(n4490), .A2(n4491), .ZN(n4489) );
  AND2_X1 U3023 ( .A1(n2795), .A2(n2793), .ZN(n4425) );
  AND2_X1 U3024 ( .A1(n4226), .A2(n4227), .ZN(n4248) );
  NAND2_X1 U3025 ( .A1(n2760), .A2(n2814), .ZN(n2990) );
  NAND2_X1 U3026 ( .A1(n2137), .A2(DATAI_24_), .ZN(n4140) );
  NAND2_X1 U3027 ( .A1(n2137), .A2(DATAI_21_), .ZN(n4195) );
  INV_X1 U3028 ( .A(n3322), .ZN(n3328) );
  NAND2_X1 U3029 ( .A1(n4210), .A2(n4565), .ZN(n4582) );
  AND2_X1 U3030 ( .A1(n3007), .A2(n2928), .ZN(n4579) );
  NAND2_X1 U3031 ( .A1(n2739), .A2(n2737), .ZN(n2813) );
  INV_X1 U3032 ( .A(n2928), .ZN(n3969) );
  AND2_X1 U3033 ( .A1(n2555), .A2(n2564), .ZN(n4003) );
  OAI21_X1 U3034 ( .B1(n2465), .B2(n2464), .A(n2473), .ZN(n4414) );
  NAND2_X1 U3035 ( .A1(n3069), .A2(STATE_REG_SCAN_IN), .ZN(n4551) );
  INV_X1 U3036 ( .A(n4290), .ZN(n3973) );
  OAI211_X1 U3037 ( .C1(n2872), .C2(n4730), .A(n2626), .B(n2625), .ZN(n4116)
         );
  INV_X1 U3038 ( .A(n4250), .ZN(n3976) );
  INV_X1 U3039 ( .A(n4533), .ZN(n4518) );
  INV_X1 U3040 ( .A(n4553), .ZN(n4537) );
  INV_X1 U3041 ( .A(n4188), .ZN(n4265) );
  NAND2_X1 U3042 ( .A1(n4599), .A2(n4354), .ZN(n4338) );
  OR2_X1 U3043 ( .A1(n4062), .A2(n4406), .ZN(n2767) );
  AND3_X1 U3044 ( .A1(n4586), .A2(n4585), .A3(n4584), .ZN(n4598) );
  OR2_X1 U3045 ( .A1(n2765), .A2(n2925), .ZN(n4587) );
  INV_X1 U3046 ( .A(n4549), .ZN(n4550) );
  NAND2_X1 U3047 ( .A1(n2813), .A2(n2930), .ZN(n4549) );
  INV_X1 U3048 ( .A(n4024), .ZN(n4555) );
  NOR2_X1 U3049 ( .A1(n2742), .A2(n4551), .ZN(U4043) );
  INV_X1 U3050 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2761) );
  NAND2_X1 U3051 ( .A1(REG3_REG_14__SCAN_IN), .A2(REG3_REG_15__SCAN_IN), .ZN(
        n2364) );
  INV_X1 U3052 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3698) );
  NAND2_X1 U3053 ( .A1(n2617), .A2(REG3_REG_23__SCAN_IN), .ZN(n2623) );
  INV_X1 U3054 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3755) );
  INV_X1 U3055 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3719) );
  XNOR2_X1 U3056 ( .A(n2646), .B(REG3_REG_27__SCAN_IN), .ZN(n4088) );
  NOR2_X1 U3057 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2373)
         );
  NOR2_X1 U3058 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_21__SCAN_IN), .ZN(n2372)
         );
  NOR2_X1 U3059 ( .A1(IR_REG_23__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2371)
         );
  INV_X1 U3060 ( .A(n2389), .ZN(n2375) );
  NOR2_X1 U3061 ( .A1(IR_REG_27__SCAN_IN), .A2(n2375), .ZN(n2677) );
  NAND2_X1 U3062 ( .A1(n2681), .A2(IR_REG_31__SCAN_IN), .ZN(n2378) );
  INV_X1 U3063 ( .A(n2382), .ZN(n4409) );
  NAND2_X1 U3064 ( .A1(n4088), .A2(n2135), .ZN(n2388) );
  INV_X1 U3065 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4293) );
  INV_X2 U3066 ( .A(n2505), .ZN(n2648) );
  NAND2_X1 U3067 ( .A1(n2648), .A2(REG2_REG_27__SCAN_IN), .ZN(n2385) );
  INV_X1 U3068 ( .A(n2381), .ZN(n2383) );
  NAND2_X1 U3069 ( .A1(n2416), .A2(REG0_REG_27__SCAN_IN), .ZN(n2384) );
  OAI211_X1 U3070 ( .C1(n4293), .C2(n2872), .A(n2385), .B(n2384), .ZN(n2386)
         );
  INV_X1 U3071 ( .A(n2386), .ZN(n2387) );
  NAND2_X1 U3072 ( .A1(n2391), .A2(n2390), .ZN(n2392) );
  NAND2_X1 U3073 ( .A1(n2407), .A2(REG3_REG_1__SCAN_IN), .ZN(n2397) );
  NAND2_X1 U3074 ( .A1(n2457), .A2(REG1_REG_1__SCAN_IN), .ZN(n2396) );
  NAND2_X1 U3075 ( .A1(n2408), .A2(REG0_REG_1__SCAN_IN), .ZN(n2395) );
  NAND2_X1 U3076 ( .A1(n2409), .A2(REG2_REG_1__SCAN_IN), .ZN(n2394) );
  INV_X1 U3077 ( .A(DATAI_1_), .ZN(n2399) );
  MUX2_X1 U3078 ( .A(n2830), .B(n2399), .S(n2541), .Z(n2403) );
  NAND2_X1 U3079 ( .A1(n2457), .A2(REG1_REG_0__SCAN_IN), .ZN(n2401) );
  NAND2_X1 U3080 ( .A1(n2408), .A2(REG0_REG_0__SCAN_IN), .ZN(n2400) );
  INV_X1 U3081 ( .A(n2773), .ZN(n2960) );
  AND2_X1 U3082 ( .A1(n2773), .A2(n3004), .ZN(n2876) );
  INV_X1 U3083 ( .A(n2403), .ZN(n2962) );
  NAND2_X1 U3084 ( .A1(n2946), .A2(n2962), .ZN(n2404) );
  INV_X1 U3085 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2405) );
  NAND2_X1 U3086 ( .A1(n2407), .A2(REG3_REG_2__SCAN_IN), .ZN(n2412) );
  NAND2_X1 U3087 ( .A1(n2408), .A2(REG0_REG_2__SCAN_IN), .ZN(n2411) );
  NAND2_X1 U3088 ( .A1(n2409), .A2(REG2_REG_2__SCAN_IN), .ZN(n2410) );
  XNOR2_X2 U3089 ( .A(n2414), .B(n4825), .ZN(n2831) );
  INV_X1 U3090 ( .A(DATAI_2_), .ZN(n2415) );
  MUX2_X1 U3091 ( .A(n2831), .B(n2415), .S(n2138), .Z(n2976) );
  NAND2_X1 U3092 ( .A1(n3027), .A2(n2976), .ZN(n3895) );
  INV_X1 U3093 ( .A(n3044), .ZN(n2683) );
  OAI22_X1 U3094 ( .A1(n3045), .A2(n2683), .B1(n3056), .B2(n3027), .ZN(n3025)
         );
  INV_X1 U3095 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3074) );
  NAND2_X1 U3096 ( .A1(n2581), .A2(n3074), .ZN(n2420) );
  NAND2_X1 U3097 ( .A1(n2457), .A2(REG1_REG_3__SCAN_IN), .ZN(n2419) );
  NAND2_X1 U3098 ( .A1(n2416), .A2(REG0_REG_3__SCAN_IN), .ZN(n2418) );
  NAND2_X1 U3099 ( .A1(n2409), .A2(REG2_REG_3__SCAN_IN), .ZN(n2417) );
  NAND2_X1 U3100 ( .A1(n2421), .A2(IR_REG_31__SCAN_IN), .ZN(n2423) );
  NAND2_X1 U3101 ( .A1(n2423), .A2(n2422), .ZN(n2432) );
  OR2_X1 U3102 ( .A1(n2423), .A2(n2422), .ZN(n2424) );
  MUX2_X1 U3103 ( .A(n4416), .B(DATAI_3_), .S(n2138), .Z(n3077) );
  NAND2_X1 U3104 ( .A1(n3150), .A2(n3077), .ZN(n2425) );
  INV_X1 U3105 ( .A(n3150), .ZN(n3063) );
  NAND2_X1 U3106 ( .A1(n3063), .A2(n3062), .ZN(n2426) );
  NOR2_X1 U3107 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2427) );
  NOR2_X1 U3108 ( .A1(n2436), .A2(n2427), .ZN(n3160) );
  NAND2_X1 U3109 ( .A1(n2135), .A2(n3160), .ZN(n2431) );
  NAND2_X1 U3110 ( .A1(n2457), .A2(REG1_REG_4__SCAN_IN), .ZN(n2430) );
  NAND2_X1 U3111 ( .A1(n2409), .A2(REG2_REG_4__SCAN_IN), .ZN(n2429) );
  NAND2_X1 U3112 ( .A1(n2416), .A2(REG0_REG_4__SCAN_IN), .ZN(n2428) );
  NAND2_X1 U3113 ( .A1(n2432), .A2(IR_REG_31__SCAN_IN), .ZN(n2433) );
  XNOR2_X1 U3114 ( .A(n2433), .B(n4826), .ZN(n2912) );
  INV_X1 U3115 ( .A(DATAI_4_), .ZN(n2434) );
  MUX2_X1 U3116 ( .A(n2912), .B(n2434), .S(n2138), .Z(n3123) );
  OR2_X1 U3117 ( .A1(n3099), .A2(n3123), .ZN(n3898) );
  NAND2_X1 U3118 ( .A1(n3099), .A2(n3123), .ZN(n3901) );
  NAND2_X1 U3119 ( .A1(n3898), .A2(n3901), .ZN(n3120) );
  INV_X1 U3120 ( .A(n3120), .ZN(n3863) );
  NAND2_X1 U3121 ( .A1(n3099), .A2(n3151), .ZN(n2435) );
  NAND2_X1 U3122 ( .A1(n3126), .A2(n2435), .ZN(n3013) );
  AOI22_X1 U3123 ( .A1(n2457), .A2(REG1_REG_5__SCAN_IN), .B1(n2416), .B2(
        REG0_REG_5__SCAN_IN), .ZN(n2439) );
  OAI21_X1 U3124 ( .B1(n2436), .B2(REG3_REG_5__SCAN_IN), .A(n2447), .ZN(n3179)
         );
  INV_X1 U3125 ( .A(n3179), .ZN(n2437) );
  AOI22_X1 U3126 ( .A1(n2581), .A2(n2437), .B1(n2648), .B2(REG2_REG_5__SCAN_IN), .ZN(n2438) );
  NAND2_X1 U3127 ( .A1(n2440), .A2(IR_REG_31__SCAN_IN), .ZN(n2441) );
  MUX2_X1 U3128 ( .A(IR_REG_31__SCAN_IN), .B(n2441), .S(IR_REG_5__SCAN_IN), 
        .Z(n2444) );
  INV_X1 U3129 ( .A(n2442), .ZN(n2443) );
  INV_X1 U3130 ( .A(DATAI_5_), .ZN(n4624) );
  MUX2_X1 U3131 ( .A(n2891), .B(n4624), .S(n2137), .Z(n3176) );
  NAND2_X1 U3132 ( .A1(n3194), .A2(n3176), .ZN(n2445) );
  NAND2_X1 U3133 ( .A1(n3984), .A2(n3108), .ZN(n2446) );
  AND2_X1 U3134 ( .A1(n2447), .A2(n2857), .ZN(n2448) );
  NOR2_X1 U3135 ( .A1(n2455), .A2(n2448), .ZN(n3189) );
  NAND2_X1 U3136 ( .A1(n2581), .A2(n3189), .ZN(n2452) );
  NAND2_X1 U3137 ( .A1(n2457), .A2(REG1_REG_6__SCAN_IN), .ZN(n2451) );
  NAND2_X1 U3138 ( .A1(n2648), .A2(REG2_REG_6__SCAN_IN), .ZN(n2450) );
  NAND2_X1 U3139 ( .A1(n2416), .A2(REG0_REG_6__SCAN_IN), .ZN(n2449) );
  NAND4_X1 U3140 ( .A1(n2452), .A2(n2451), .A3(n2450), .A4(n2449), .ZN(n3239)
         );
  OR2_X1 U3141 ( .A1(n2442), .A2(n2194), .ZN(n2453) );
  XNOR2_X1 U3142 ( .A(n2453), .B(IR_REG_6__SCAN_IN), .ZN(n2854) );
  MUX2_X1 U3143 ( .A(n2854), .B(DATAI_6_), .S(n2137), .Z(n3167) );
  AND2_X1 U3144 ( .A1(n3239), .A2(n3167), .ZN(n2454) );
  OR2_X1 U3145 ( .A1(n2455), .A2(REG3_REG_7__SCAN_IN), .ZN(n2456) );
  AND2_X1 U3146 ( .A1(n2469), .A2(n2456), .ZN(n3240) );
  NAND2_X1 U3147 ( .A1(n2581), .A2(n3240), .ZN(n2461) );
  NAND2_X1 U31480 ( .A1(n2457), .A2(REG1_REG_7__SCAN_IN), .ZN(n2460) );
  NAND2_X1 U31490 ( .A1(n2648), .A2(REG2_REG_7__SCAN_IN), .ZN(n2459) );
  NAND2_X1 U3150 ( .A1(n2416), .A2(REG0_REG_7__SCAN_IN), .ZN(n2458) );
  NAND4_X1 U3151 ( .A1(n2461), .A2(n2460), .A3(n2459), .A4(n2458), .ZN(n3307)
         );
  AND2_X1 U3152 ( .A1(n2442), .A2(n2462), .ZN(n2463) );
  NAND2_X1 U3153 ( .A1(n2465), .A2(n2464), .ZN(n2473) );
  INV_X1 U3154 ( .A(DATAI_7_), .ZN(n4625) );
  MUX2_X1 U3155 ( .A(n4414), .B(n4625), .S(n2138), .Z(n3236) );
  OR2_X1 U3156 ( .A1(n3307), .A2(n3236), .ZN(n3904) );
  NAND2_X1 U3157 ( .A1(n3307), .A2(n3236), .ZN(n3907) );
  NAND2_X1 U3158 ( .A1(n2467), .A2(n2466), .ZN(n3144) );
  NAND2_X1 U3159 ( .A1(n3307), .A2(n3231), .ZN(n2468) );
  AOI22_X1 U3160 ( .A1(n2457), .A2(REG1_REG_8__SCAN_IN), .B1(n2416), .B2(
        REG0_REG_8__SCAN_IN), .ZN(n2472) );
  NAND2_X1 U3161 ( .A1(n2469), .A2(n4633), .ZN(n2470) );
  AND2_X1 U3162 ( .A1(n2479), .A2(n2470), .ZN(n4540) );
  AOI22_X1 U3163 ( .A1(n2581), .A2(n4540), .B1(n2648), .B2(REG2_REG_8__SCAN_IN), .ZN(n2471) );
  NAND2_X1 U3164 ( .A1(n2473), .A2(IR_REG_31__SCAN_IN), .ZN(n2474) );
  XNOR2_X1 U3165 ( .A(n2474), .B(IR_REG_8__SCAN_IN), .ZN(n4600) );
  INV_X1 U3166 ( .A(DATAI_8_), .ZN(n2475) );
  MUX2_X1 U3167 ( .A(n4439), .B(n2475), .S(n2137), .Z(n3302) );
  NAND2_X1 U3168 ( .A1(n3327), .A2(n3302), .ZN(n2476) );
  NAND2_X1 U3169 ( .A1(n3983), .A2(n3306), .ZN(n2477) );
  AND2_X1 U3170 ( .A1(n2479), .A2(n2478), .ZN(n2480) );
  OR2_X1 U3171 ( .A1(n2480), .A2(n2492), .ZN(n3332) );
  INV_X1 U3172 ( .A(n3332), .ZN(n2481) );
  NAND2_X1 U3173 ( .A1(n2581), .A2(n2481), .ZN(n2485) );
  NAND2_X1 U3174 ( .A1(n2457), .A2(REG1_REG_9__SCAN_IN), .ZN(n2484) );
  NAND2_X1 U3175 ( .A1(n2416), .A2(REG0_REG_9__SCAN_IN), .ZN(n2483) );
  NAND2_X1 U3176 ( .A1(n2648), .A2(REG2_REG_9__SCAN_IN), .ZN(n2482) );
  NAND4_X1 U3177 ( .A1(n2485), .A2(n2484), .A3(n2483), .A4(n2482), .ZN(n3982)
         );
  NAND2_X1 U3178 ( .A1(n2442), .A2(n2486), .ZN(n2487) );
  NAND2_X1 U3179 ( .A1(n2487), .A2(IR_REG_31__SCAN_IN), .ZN(n2488) );
  MUX2_X1 U3180 ( .A(IR_REG_31__SCAN_IN), .B(n2488), .S(IR_REG_9__SCAN_IN), 
        .Z(n2490) );
  AND2_X1 U3181 ( .A1(n2490), .A2(n2489), .ZN(n4440) );
  MUX2_X1 U3182 ( .A(n4440), .B(DATAI_9_), .S(n2138), .Z(n3322) );
  AND2_X1 U3183 ( .A1(n3982), .A2(n3322), .ZN(n2491) );
  INV_X1 U3184 ( .A(n3982), .ZN(n3673) );
  NAND2_X1 U3185 ( .A1(n2457), .A2(REG1_REG_10__SCAN_IN), .ZN(n2497) );
  NOR2_X1 U3186 ( .A1(n2492), .A2(REG3_REG_10__SCAN_IN), .ZN(n2493) );
  NOR2_X1 U3187 ( .A1(n2502), .A2(n2493), .ZN(n3680) );
  NAND2_X1 U3188 ( .A1(n2581), .A2(n3680), .ZN(n2496) );
  NAND2_X1 U3189 ( .A1(n2416), .A2(REG0_REG_10__SCAN_IN), .ZN(n2495) );
  NAND2_X1 U3190 ( .A1(n2648), .A2(REG2_REG_10__SCAN_IN), .ZN(n2494) );
  NAND2_X1 U3191 ( .A1(n2489), .A2(IR_REG_31__SCAN_IN), .ZN(n2498) );
  XNOR2_X1 U3192 ( .A(n2498), .B(IR_REG_10__SCAN_IN), .ZN(n4013) );
  MUX2_X1 U3193 ( .A(n4013), .B(DATAI_10_), .S(n2138), .Z(n3671) );
  NOR2_X1 U3194 ( .A1(n3399), .A2(n3671), .ZN(n2499) );
  NAND2_X1 U3195 ( .A1(n3399), .A2(n3671), .ZN(n2500) );
  OAI21_X1 U3196 ( .B1(n3222), .B2(n2499), .A(n2500), .ZN(n2501) );
  INV_X1 U3197 ( .A(n2501), .ZN(n3287) );
  OR2_X1 U3198 ( .A1(n2502), .A2(REG3_REG_11__SCAN_IN), .ZN(n2503) );
  NAND2_X1 U3199 ( .A1(n2514), .A2(n2503), .ZN(n3413) );
  INV_X1 U3200 ( .A(n3413), .ZN(n2504) );
  NAND2_X1 U3201 ( .A1(n2135), .A2(n2504), .ZN(n2509) );
  NAND2_X1 U3202 ( .A1(n2457), .A2(REG1_REG_11__SCAN_IN), .ZN(n2508) );
  NAND2_X1 U3203 ( .A1(n2648), .A2(REG2_REG_11__SCAN_IN), .ZN(n2507) );
  NAND2_X1 U3204 ( .A1(n2416), .A2(REG0_REG_11__SCAN_IN), .ZN(n2506) );
  NAND4_X1 U3205 ( .A1(n2509), .A2(n2508), .A3(n2507), .A4(n2506), .ZN(n3670)
         );
  NOR2_X1 U3206 ( .A1(n2489), .A2(IR_REG_10__SCAN_IN), .ZN(n2532) );
  OR2_X1 U3207 ( .A1(n2532), .A2(n2194), .ZN(n2511) );
  NAND2_X1 U3208 ( .A1(n2511), .A2(n2510), .ZN(n2520) );
  INV_X1 U3209 ( .A(DATAI_11_), .ZN(n2512) );
  MUX2_X1 U32100 ( .A(n4470), .B(n2512), .S(n2138), .Z(n3409) );
  OR2_X1 U32110 ( .A1(n3670), .A2(n3409), .ZN(n3333) );
  NAND2_X1 U32120 ( .A1(n3670), .A2(n3409), .ZN(n3924) );
  NAND2_X1 U32130 ( .A1(n3333), .A2(n3924), .ZN(n3854) );
  NAND2_X1 U32140 ( .A1(n3287), .A2(n3854), .ZN(n3286) );
  NAND2_X1 U32150 ( .A1(n3708), .A2(n3409), .ZN(n2513) );
  NAND2_X1 U32160 ( .A1(n3286), .A2(n2513), .ZN(n3337) );
  NAND2_X1 U32170 ( .A1(n2514), .A2(n4631), .ZN(n2515) );
  AND2_X1 U32180 ( .A1(n2525), .A2(n2515), .ZN(n3710) );
  NAND2_X1 U32190 ( .A1(n2581), .A2(n3710), .ZN(n2519) );
  NAND2_X1 U32200 ( .A1(n2457), .A2(REG1_REG_12__SCAN_IN), .ZN(n2518) );
  NAND2_X1 U32210 ( .A1(n2648), .A2(REG2_REG_12__SCAN_IN), .ZN(n2517) );
  NAND2_X1 U32220 ( .A1(n2416), .A2(REG0_REG_12__SCAN_IN), .ZN(n2516) );
  NAND2_X1 U32230 ( .A1(n2520), .A2(IR_REG_31__SCAN_IN), .ZN(n2521) );
  XNOR2_X1 U32240 ( .A(n2521), .B(IR_REG_12__SCAN_IN), .ZN(n4016) );
  MUX2_X1 U32250 ( .A(n4016), .B(DATAI_12_), .S(n2138), .Z(n3706) );
  NAND2_X1 U32260 ( .A1(n3981), .A2(n3706), .ZN(n2522) );
  NAND2_X1 U32270 ( .A1(n3337), .A2(n2522), .ZN(n2524) );
  OR2_X1 U32280 ( .A1(n3981), .A2(n3706), .ZN(n2523) );
  NAND2_X1 U32290 ( .A1(n2524), .A2(n2523), .ZN(n3366) );
  NAND2_X1 U32300 ( .A1(n2525), .A2(n3615), .ZN(n2526) );
  AND2_X1 U32310 ( .A1(n2543), .A2(n2526), .ZN(n3619) );
  NAND2_X1 U32320 ( .A1(n2135), .A2(n3619), .ZN(n2530) );
  NAND2_X1 U32330 ( .A1(n2457), .A2(REG1_REG_13__SCAN_IN), .ZN(n2529) );
  NAND2_X1 U32340 ( .A1(n2648), .A2(REG2_REG_13__SCAN_IN), .ZN(n2528) );
  NAND2_X1 U32350 ( .A1(n2416), .A2(REG0_REG_13__SCAN_IN), .ZN(n2527) );
  NAND4_X1 U32360 ( .A1(n2530), .A2(n2529), .A3(n2528), .A4(n2527), .ZN(n3980)
         );
  NOR2_X1 U32370 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U32380 ( .A1(n2532), .A2(n2531), .ZN(n2534) );
  NAND2_X1 U32390 ( .A1(n2534), .A2(IR_REG_31__SCAN_IN), .ZN(n2533) );
  MUX2_X1 U32400 ( .A(IR_REG_31__SCAN_IN), .B(n2533), .S(IR_REG_13__SCAN_IN), 
        .Z(n2535) );
  MUX2_X1 U32410 ( .A(n4483), .B(DATAI_13_), .S(n2137), .Z(n3494) );
  NAND2_X1 U32420 ( .A1(n2457), .A2(REG1_REG_14__SCAN_IN), .ZN(n2539) );
  XNOR2_X1 U32430 ( .A(n2543), .B(REG3_REG_14__SCAN_IN), .ZN(n3658) );
  NAND2_X1 U32440 ( .A1(n2581), .A2(n3658), .ZN(n2538) );
  NAND2_X1 U32450 ( .A1(n2416), .A2(REG0_REG_14__SCAN_IN), .ZN(n2537) );
  NAND2_X1 U32460 ( .A1(n2648), .A2(REG2_REG_14__SCAN_IN), .ZN(n2536) );
  NAND4_X1 U32470 ( .A1(n2539), .A2(n2538), .A3(n2537), .A4(n2536), .ZN(n3979)
         );
  NAND2_X1 U32480 ( .A1(n2550), .A2(IR_REG_31__SCAN_IN), .ZN(n2540) );
  XNOR2_X1 U32490 ( .A(n2540), .B(IR_REG_14__SCAN_IN), .ZN(n4020) );
  INV_X1 U32500 ( .A(DATAI_14_), .ZN(n2542) );
  MUX2_X1 U32510 ( .A(n4558), .B(n2542), .S(n2137), .Z(n3515) );
  OR2_X1 U32520 ( .A1(n3979), .A2(n3515), .ZN(n3817) );
  NAND2_X1 U32530 ( .A1(n3979), .A2(n3515), .ZN(n3818) );
  NAND2_X1 U32540 ( .A1(n3817), .A2(n3818), .ZN(n3437) );
  INV_X1 U32550 ( .A(n3979), .ZN(n3808) );
  INV_X1 U32560 ( .A(n2543), .ZN(n2544) );
  AOI21_X1 U32570 ( .B1(n2544), .B2(REG3_REG_14__SCAN_IN), .A(
        REG3_REG_15__SCAN_IN), .ZN(n2545) );
  OR2_X1 U32580 ( .A1(n2545), .A2(n2558), .ZN(n3814) );
  INV_X1 U32590 ( .A(n3814), .ZN(n3428) );
  NAND2_X1 U32600 ( .A1(n2135), .A2(n3428), .ZN(n2549) );
  NAND2_X1 U32610 ( .A1(n2457), .A2(REG1_REG_15__SCAN_IN), .ZN(n2548) );
  NAND2_X1 U32620 ( .A1(n2648), .A2(REG2_REG_15__SCAN_IN), .ZN(n2547) );
  NAND2_X1 U32630 ( .A1(n2416), .A2(REG0_REG_15__SCAN_IN), .ZN(n2546) );
  NAND4_X1 U32640 ( .A1(n2549), .A2(n2548), .A3(n2547), .A4(n2546), .ZN(n3978)
         );
  NAND2_X1 U32650 ( .A1(n2551), .A2(IR_REG_31__SCAN_IN), .ZN(n2554) );
  INV_X1 U32660 ( .A(n2554), .ZN(n2552) );
  NAND2_X1 U32670 ( .A1(n2552), .A2(IR_REG_15__SCAN_IN), .ZN(n2555) );
  NAND2_X1 U32680 ( .A1(n2554), .A2(n2553), .ZN(n2564) );
  MUX2_X1 U32690 ( .A(n4003), .B(DATAI_15_), .S(n2137), .Z(n3520) );
  NAND2_X1 U32700 ( .A1(n3978), .A2(n3520), .ZN(n2557) );
  NOR2_X1 U32710 ( .A1(n3978), .A2(n3520), .ZN(n2556) );
  AOI21_X1 U32720 ( .B1(n3422), .B2(n2557), .A(n2556), .ZN(n3450) );
  OR2_X1 U32730 ( .A1(n2558), .A2(REG3_REG_16__SCAN_IN), .ZN(n2559) );
  AND2_X1 U32740 ( .A1(n2559), .A2(n2570), .ZN(n3733) );
  NAND2_X1 U32750 ( .A1(n2581), .A2(n3733), .ZN(n2563) );
  NAND2_X1 U32760 ( .A1(n2457), .A2(REG1_REG_16__SCAN_IN), .ZN(n2562) );
  NAND2_X1 U32770 ( .A1(n2409), .A2(REG2_REG_16__SCAN_IN), .ZN(n2561) );
  NAND2_X1 U32780 ( .A1(n2416), .A2(REG0_REG_16__SCAN_IN), .ZN(n2560) );
  NAND4_X1 U32790 ( .A1(n2563), .A2(n2562), .A3(n2561), .A4(n2560), .ZN(n3977)
         );
  NAND2_X1 U32800 ( .A1(n2564), .A2(IR_REG_31__SCAN_IN), .ZN(n2565) );
  XNOR2_X1 U32810 ( .A(n2565), .B(IR_REG_16__SCAN_IN), .ZN(n4024) );
  INV_X1 U32820 ( .A(DATAI_16_), .ZN(n2566) );
  MUX2_X1 U32830 ( .A(n4555), .B(n2566), .S(n2138), .Z(n2567) );
  OR2_X1 U32840 ( .A1(n3977), .A2(n2567), .ZN(n3935) );
  NAND2_X1 U32850 ( .A1(n3977), .A2(n2567), .ZN(n3931) );
  NAND2_X1 U32860 ( .A1(n3935), .A2(n3931), .ZN(n3451) );
  NAND2_X1 U32870 ( .A1(n3450), .A2(n3451), .ZN(n3449) );
  NAND2_X1 U32880 ( .A1(n3977), .A2(n3728), .ZN(n2568) );
  AOI22_X1 U32890 ( .A1(n2457), .A2(REG1_REG_17__SCAN_IN), .B1(n2416), .B2(
        REG0_REG_17__SCAN_IN), .ZN(n2573) );
  NAND2_X1 U32900 ( .A1(n2570), .A2(n2569), .ZN(n2571) );
  AND2_X1 U32910 ( .A1(n2579), .A2(n2571), .ZN(n3745) );
  AOI22_X1 U32920 ( .A1(n2135), .A2(n3745), .B1(n2648), .B2(
        REG2_REG_17__SCAN_IN), .ZN(n2572) );
  NAND2_X1 U32930 ( .A1(n2574), .A2(IR_REG_31__SCAN_IN), .ZN(n2575) );
  MUX2_X1 U32940 ( .A(IR_REG_31__SCAN_IN), .B(n2575), .S(IR_REG_17__SCAN_IN), 
        .Z(n2576) );
  INV_X1 U32950 ( .A(n2671), .ZN(n2667) );
  NAND2_X1 U32960 ( .A1(n2576), .A2(n2667), .ZN(n4037) );
  INV_X1 U32970 ( .A(DATAI_17_), .ZN(n4617) );
  MUX2_X1 U32980 ( .A(n4037), .B(n4617), .S(n2137), .Z(n3742) );
  NAND2_X1 U32990 ( .A1(n3976), .A2(n4343), .ZN(n2577) );
  NAND2_X1 U33000 ( .A1(n2457), .A2(REG1_REG_18__SCAN_IN), .ZN(n2585) );
  AND2_X1 U33010 ( .A1(n2579), .A2(n2578), .ZN(n2580) );
  NOR2_X1 U33020 ( .A1(n2590), .A2(n2580), .ZN(n4259) );
  NAND2_X1 U33030 ( .A1(n2581), .A2(n4259), .ZN(n2584) );
  NAND2_X1 U33040 ( .A1(n2416), .A2(REG0_REG_18__SCAN_IN), .ZN(n2583) );
  NAND2_X1 U33050 ( .A1(n2648), .A2(REG2_REG_18__SCAN_IN), .ZN(n2582) );
  NAND4_X1 U33060 ( .A1(n2585), .A2(n2584), .A3(n2583), .A4(n2582), .ZN(n4345)
         );
  OR2_X1 U33070 ( .A1(n2671), .A2(n2194), .ZN(n2586) );
  XNOR2_X1 U33080 ( .A(n2586), .B(IR_REG_18__SCAN_IN), .ZN(n4553) );
  INV_X1 U33090 ( .A(DATAI_18_), .ZN(n2587) );
  MUX2_X1 U33100 ( .A(n4537), .B(n2587), .S(n2137), .Z(n4257) );
  OR2_X1 U33110 ( .A1(n4345), .A2(n4257), .ZN(n4226) );
  NAND2_X1 U33120 ( .A1(n4345), .A2(n4257), .ZN(n4227) );
  NAND2_X1 U33130 ( .A1(n3741), .A2(n4257), .ZN(n2589) );
  NOR2_X1 U33140 ( .A1(n2590), .A2(REG3_REG_19__SCAN_IN), .ZN(n2591) );
  OR2_X1 U33150 ( .A1(n2600), .A2(n2591), .ZN(n4240) );
  INV_X1 U33160 ( .A(n4240), .ZN(n3689) );
  NAND2_X1 U33170 ( .A1(n2581), .A2(n3689), .ZN(n2595) );
  NAND2_X1 U33180 ( .A1(n2457), .A2(REG1_REG_19__SCAN_IN), .ZN(n2594) );
  NAND2_X1 U33190 ( .A1(n2648), .A2(REG2_REG_19__SCAN_IN), .ZN(n2593) );
  NAND2_X1 U33200 ( .A1(n2416), .A2(REG0_REG_19__SCAN_IN), .ZN(n2592) );
  NAND4_X1 U33210 ( .A1(n2595), .A2(n2594), .A3(n2593), .A4(n2592), .ZN(n3975)
         );
  NAND2_X1 U33220 ( .A1(n2596), .A2(n2665), .ZN(n2662) );
  OR2_X1 U33230 ( .A1(n2596), .A2(n2665), .ZN(n2597) );
  MUX2_X1 U33240 ( .A(n4412), .B(DATAI_19_), .S(n2138), .Z(n3686) );
  NAND2_X1 U33250 ( .A1(n3975), .A2(n3686), .ZN(n2599) );
  NOR2_X1 U33260 ( .A1(n3975), .A2(n3686), .ZN(n2598) );
  OR2_X1 U33270 ( .A1(n2600), .A2(REG3_REG_20__SCAN_IN), .ZN(n2601) );
  AND2_X1 U33280 ( .A1(n2606), .A2(n2601), .ZN(n4214) );
  NAND2_X1 U33290 ( .A1(n2581), .A2(n4214), .ZN(n2605) );
  NAND2_X1 U33300 ( .A1(n2457), .A2(REG1_REG_20__SCAN_IN), .ZN(n2604) );
  NAND2_X1 U33310 ( .A1(n2416), .A2(REG0_REG_20__SCAN_IN), .ZN(n2603) );
  NAND2_X1 U33320 ( .A1(n2648), .A2(REG2_REG_20__SCAN_IN), .ZN(n2602) );
  NAND4_X1 U33330 ( .A1(n2605), .A2(n2604), .A3(n2603), .A4(n2602), .ZN(n3974)
         );
  AND2_X1 U33340 ( .A1(n3974), .A2(n4216), .ZN(n3880) );
  OR2_X1 U33350 ( .A1(n3974), .A2(n4216), .ZN(n3881) );
  NAND2_X1 U33360 ( .A1(n2606), .A2(n3698), .ZN(n2607) );
  AND2_X1 U33370 ( .A1(n2613), .A2(n2607), .ZN(n4191) );
  NAND2_X1 U33380 ( .A1(n2135), .A2(n4191), .ZN(n2611) );
  NAND2_X1 U33390 ( .A1(n2457), .A2(REG1_REG_21__SCAN_IN), .ZN(n2610) );
  NAND2_X1 U33400 ( .A1(n2648), .A2(REG2_REG_21__SCAN_IN), .ZN(n2609) );
  NAND2_X1 U33410 ( .A1(n2416), .A2(REG0_REG_21__SCAN_IN), .ZN(n2608) );
  INV_X1 U33420 ( .A(n4195), .ZN(n4321) );
  NAND2_X1 U33430 ( .A1(n4206), .A2(n4321), .ZN(n2612) );
  INV_X1 U33440 ( .A(n4206), .ZN(n3774) );
  AOI22_X1 U33450 ( .A1(n4186), .A2(n2612), .B1(n3774), .B2(n4195), .ZN(n4169)
         );
  AND2_X1 U33460 ( .A1(n2613), .A2(n4805), .ZN(n2614) );
  OR2_X1 U33470 ( .A1(n2614), .A2(n2617), .ZN(n4178) );
  AOI22_X1 U33480 ( .A1(n2457), .A2(REG1_REG_22__SCAN_IN), .B1(n2416), .B2(
        REG0_REG_22__SCAN_IN), .ZN(n2616) );
  NAND2_X1 U33490 ( .A1(n2648), .A2(REG2_REG_22__SCAN_IN), .ZN(n2615) );
  OR2_X1 U33500 ( .A1(n4322), .A2(n4177), .ZN(n4149) );
  NAND2_X1 U33510 ( .A1(n4322), .A2(n4177), .ZN(n2704) );
  NAND2_X1 U33520 ( .A1(n4169), .A2(n4170), .ZN(n4168) );
  NAND2_X1 U3353 ( .A1(n4168), .A2(n2361), .ZN(n4146) );
  INV_X1 U33540 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4314) );
  OR2_X1 U3355 ( .A1(n2617), .A2(REG3_REG_23__SCAN_IN), .ZN(n2618) );
  NAND2_X1 U3356 ( .A1(n2623), .A2(n2618), .ZN(n4162) );
  OR2_X1 U3357 ( .A1(n4162), .A2(n2393), .ZN(n2620) );
  AOI22_X1 U3358 ( .A1(n2648), .A2(REG2_REG_23__SCAN_IN), .B1(n2416), .B2(
        REG0_REG_23__SCAN_IN), .ZN(n2619) );
  INV_X1 U3359 ( .A(n4304), .ZN(n4172) );
  NAND2_X1 U3360 ( .A1(n4172), .A2(n4160), .ZN(n2622) );
  AOI21_X2 U3361 ( .B1(n4146), .B2(n2622), .A(n2621), .ZN(n4134) );
  INV_X1 U3362 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4730) );
  NAND2_X1 U3363 ( .A1(n2623), .A2(n3755), .ZN(n2624) );
  NAND2_X1 U3364 ( .A1(n2629), .A2(n2624), .ZN(n3754) );
  OR2_X1 U3365 ( .A1(n3754), .A2(n2393), .ZN(n2626) );
  AOI22_X1 U3366 ( .A1(n2648), .A2(REG2_REG_24__SCAN_IN), .B1(n2416), .B2(
        REG0_REG_24__SCAN_IN), .ZN(n2625) );
  NAND2_X1 U3367 ( .A1(n4116), .A2(n4302), .ZN(n2628) );
  INV_X1 U3368 ( .A(n4116), .ZN(n4158) );
  AOI21_X2 U3369 ( .B1(n4134), .B2(n2628), .A(n2627), .ZN(n4111) );
  AND2_X1 U3370 ( .A1(n2629), .A2(n3719), .ZN(n2630) );
  OR2_X1 U3371 ( .A1(n2636), .A2(n2630), .ZN(n3718) );
  INV_X1 U3372 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4300) );
  NAND2_X1 U3373 ( .A1(n2648), .A2(REG2_REG_25__SCAN_IN), .ZN(n2632) );
  NAND2_X1 U3374 ( .A1(n2416), .A2(REG0_REG_25__SCAN_IN), .ZN(n2631) );
  OAI211_X1 U3375 ( .C1(n4300), .C2(n2872), .A(n2632), .B(n2631), .ZN(n2633)
         );
  INV_X1 U3376 ( .A(n2633), .ZN(n2634) );
  INV_X1 U3377 ( .A(n4101), .ZN(n4308) );
  NAND2_X1 U3378 ( .A1(n4308), .A2(n4122), .ZN(n2635) );
  INV_X1 U3379 ( .A(n4122), .ZN(n4115) );
  OR2_X1 U3380 ( .A1(n2636), .A2(REG3_REG_26__SCAN_IN), .ZN(n2637) );
  NAND2_X1 U3381 ( .A1(n2646), .A2(n2637), .ZN(n3793) );
  INV_X1 U3382 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4732) );
  NAND2_X1 U3383 ( .A1(n2648), .A2(REG2_REG_26__SCAN_IN), .ZN(n2639) );
  NAND2_X1 U3384 ( .A1(n2408), .A2(REG0_REG_26__SCAN_IN), .ZN(n2638) );
  OAI211_X1 U3385 ( .C1(n4732), .C2(n2872), .A(n2639), .B(n2638), .ZN(n2640)
         );
  INV_X1 U3386 ( .A(n2640), .ZN(n2641) );
  INV_X1 U3387 ( .A(n4105), .ZN(n4100) );
  INV_X1 U3388 ( .A(n4281), .ZN(n3642) );
  INV_X1 U3389 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3607) );
  INV_X1 U3390 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2645) );
  OAI21_X1 U3391 ( .B1(n2646), .B2(n3607), .A(n2645), .ZN(n2647) );
  NAND2_X1 U3392 ( .A1(n2647), .A2(n4061), .ZN(n4073) );
  OR2_X1 U3393 ( .A1(n4073), .A2(n2393), .ZN(n2653) );
  INV_X1 U3394 ( .A(REG1_REG_28__SCAN_IN), .ZN(n4284) );
  NAND2_X1 U3395 ( .A1(n2648), .A2(REG2_REG_28__SCAN_IN), .ZN(n2650) );
  NAND2_X1 U3396 ( .A1(n2416), .A2(REG0_REG_28__SCAN_IN), .ZN(n2649) );
  OAI211_X1 U3397 ( .C1(n4284), .C2(n2872), .A(n2650), .B(n2649), .ZN(n2651)
         );
  INV_X1 U3398 ( .A(n2651), .ZN(n2652) );
  INV_X1 U3399 ( .A(n3836), .ZN(n2654) );
  INV_X1 U3400 ( .A(n4277), .ZN(n4077) );
  NAND2_X1 U3401 ( .A1(n3973), .A2(n4077), .ZN(n3832) );
  NAND2_X1 U3402 ( .A1(n2654), .A2(n3832), .ZN(n4068) );
  AOI22_X1 U3403 ( .A1(n4070), .A2(n4068), .B1(n4277), .B2(n3973), .ZN(n2661)
         );
  INV_X1 U3404 ( .A(n4061), .ZN(n2655) );
  NAND2_X1 U3405 ( .A1(n2655), .A2(n2581), .ZN(n2660) );
  NAND2_X1 U3406 ( .A1(n2648), .A2(REG2_REG_29__SCAN_IN), .ZN(n2657) );
  NAND2_X1 U3407 ( .A1(n2408), .A2(REG0_REG_29__SCAN_IN), .ZN(n2656) );
  OAI211_X1 U3408 ( .C1(n2761), .C2(n2872), .A(n2657), .B(n2656), .ZN(n2658)
         );
  INV_X1 U3409 ( .A(n2658), .ZN(n2659) );
  NAND2_X1 U3410 ( .A1(n2660), .A2(n2659), .ZN(n4278) );
  NAND2_X1 U3411 ( .A1(n2138), .A2(DATAI_29_), .ZN(n2762) );
  XNOR2_X1 U3412 ( .A(n4278), .B(n2762), .ZN(n3878) );
  XNOR2_X2 U3413 ( .A(n2663), .B(n2664), .ZN(n2676) );
  NAND2_X1 U3414 ( .A1(n2665), .A2(n2664), .ZN(n2666) );
  OAI21_X1 U3415 ( .B1(n2667), .B2(n2669), .A(IR_REG_31__SCAN_IN), .ZN(n2668)
         );
  MUX2_X1 U3416 ( .A(IR_REG_31__SCAN_IN), .B(n2668), .S(IR_REG_21__SCAN_IN), 
        .Z(n2672) );
  NOR2_X1 U3417 ( .A1(n2669), .A2(IR_REG_21__SCAN_IN), .ZN(n2670) );
  AND2_X1 U3418 ( .A1(n2671), .A2(n2670), .ZN(n2731) );
  INV_X1 U3419 ( .A(n2731), .ZN(n2673) );
  NAND2_X2 U3420 ( .A1(n2676), .A2(n4410), .ZN(n2768) );
  NAND2_X1 U3421 ( .A1(n2673), .A2(IR_REG_31__SCAN_IN), .ZN(n2674) );
  XNOR2_X1 U3422 ( .A(n2768), .B(n3969), .ZN(n2675) );
  AND2_X1 U3423 ( .A1(n2676), .A2(n4412), .ZN(n3007) );
  AND2_X1 U3424 ( .A1(n2722), .A2(n2677), .ZN(n2678) );
  NOR2_X1 U3425 ( .A1(n2678), .A2(n2194), .ZN(n2679) );
  MUX2_X1 U3426 ( .A(n2194), .B(n2679), .S(IR_REG_28__SCAN_IN), .Z(n2680) );
  INV_X1 U3427 ( .A(n2680), .ZN(n2682) );
  NAND2_X1 U3428 ( .A1(n2682), .A2(n2681), .ZN(n2938) );
  AND2_X1 U3429 ( .A1(n4410), .A2(n3969), .ZN(n2782) );
  INV_X1 U3430 ( .A(n2782), .ZN(n2922) );
  NAND2_X1 U3431 ( .A1(n3047), .A2(n2683), .ZN(n3046) );
  NAND2_X1 U3432 ( .A1(n3046), .A2(n3892), .ZN(n3026) );
  NAND2_X1 U3433 ( .A1(n3150), .A2(n3062), .ZN(n3894) );
  NAND2_X1 U3434 ( .A1(n3026), .A2(n2145), .ZN(n2684) );
  NAND2_X1 U3435 ( .A1(n2684), .A2(n3897), .ZN(n3121) );
  INV_X1 U3436 ( .A(n3898), .ZN(n2685) );
  OR2_X1 U3437 ( .A1(n3984), .A2(n3176), .ZN(n3914) );
  NAND2_X1 U3438 ( .A1(n3984), .A2(n3176), .ZN(n3900) );
  AND2_X1 U3439 ( .A1(n3239), .A2(n3193), .ZN(n3915) );
  OR2_X1 U3440 ( .A1(n3239), .A2(n3193), .ZN(n3903) );
  INV_X1 U3441 ( .A(n3904), .ZN(n2688) );
  OR2_X1 U3442 ( .A1(n3983), .A2(n3302), .ZN(n3908) );
  NAND2_X1 U3443 ( .A1(n3983), .A2(n3302), .ZN(n3906) );
  AND2_X1 U3444 ( .A1(n3982), .A2(n3328), .ZN(n3917) );
  OR2_X1 U3445 ( .A1(n3982), .A2(n3328), .ZN(n3909) );
  NAND2_X1 U3446 ( .A1(n3399), .A2(n3397), .ZN(n3923) );
  NAND2_X1 U3447 ( .A1(n3216), .A2(n3923), .ZN(n2690) );
  OR2_X1 U3448 ( .A1(n3399), .A2(n3397), .ZN(n3918) );
  NAND2_X1 U3449 ( .A1(n2690), .A2(n3918), .ZN(n3285) );
  NAND2_X1 U3450 ( .A1(n3285), .A2(n3924), .ZN(n3334) );
  INV_X1 U3451 ( .A(n3706), .ZN(n3505) );
  NAND2_X1 U3452 ( .A1(n3981), .A2(n3505), .ZN(n3359) );
  NAND2_X1 U3453 ( .A1(n3980), .A2(n3617), .ZN(n2691) );
  NAND2_X1 U3454 ( .A1(n3359), .A2(n2691), .ZN(n2692) );
  INV_X1 U3455 ( .A(n2692), .ZN(n3925) );
  OR2_X1 U3456 ( .A1(n3981), .A2(n3505), .ZN(n3358) );
  NAND2_X1 U3457 ( .A1(n3333), .A2(n3358), .ZN(n2694) );
  NOR2_X1 U34580 ( .A1(n3980), .A2(n3617), .ZN(n2693) );
  AOI21_X1 U34590 ( .B1(n3925), .B2(n2694), .A(n2693), .ZN(n3927) );
  INV_X1 U3460 ( .A(n3437), .ZN(n3868) );
  INV_X1 U3461 ( .A(n3520), .ZN(n3809) );
  OR2_X1 U3462 ( .A1(n3978), .A2(n3809), .ZN(n3820) );
  NAND2_X1 U3463 ( .A1(n3978), .A2(n3809), .ZN(n3819) );
  NAND2_X1 U3464 ( .A1(n3820), .A2(n3819), .ZN(n3866) );
  INV_X1 U3465 ( .A(n3817), .ZN(n2695) );
  NAND2_X1 U3466 ( .A1(n2696), .A2(n3819), .ZN(n3452) );
  INV_X1 U34670 ( .A(n3451), .ZN(n3869) );
  INV_X1 U3468 ( .A(n3686), .ZN(n4236) );
  NAND2_X1 U34690 ( .A1(n3975), .A2(n4236), .ZN(n2697) );
  NAND2_X1 U3470 ( .A1(n4227), .A2(n2697), .ZN(n2698) );
  INV_X1 U34710 ( .A(n2698), .ZN(n3936) );
  OR2_X1 U3472 ( .A1(n3976), .A2(n3742), .ZN(n4224) );
  NAND2_X1 U34730 ( .A1(n4226), .A2(n4224), .ZN(n2700) );
  NOR2_X1 U3474 ( .A1(n3975), .A2(n4236), .ZN(n2699) );
  AOI21_X1 U34750 ( .B1(n3936), .B2(n2700), .A(n2699), .ZN(n4203) );
  INV_X1 U3476 ( .A(n3974), .ZN(n4325) );
  NAND2_X1 U34770 ( .A1(n4325), .A2(n4216), .ZN(n2701) );
  NAND2_X1 U3478 ( .A1(n4204), .A2(n3940), .ZN(n2702) );
  INV_X1 U34790 ( .A(n4216), .ZN(n3766) );
  NAND2_X1 U3480 ( .A1(n3974), .A2(n3766), .ZN(n3824) );
  NAND2_X1 U34810 ( .A1(n2702), .A2(n3824), .ZN(n4184) );
  OR2_X1 U3482 ( .A1(n4206), .A2(n4195), .ZN(n4147) );
  NAND2_X1 U34830 ( .A1(n4149), .A2(n4147), .ZN(n3942) );
  INV_X1 U3484 ( .A(n3942), .ZN(n2707) );
  AND2_X1 U34850 ( .A1(n4206), .A2(n4195), .ZN(n4148) );
  AND2_X1 U3486 ( .A1(n4149), .A2(n4148), .ZN(n2705) );
  NAND2_X1 U34870 ( .A1(n4304), .A2(n4160), .ZN(n2703) );
  NAND2_X1 U3488 ( .A1(n2704), .A2(n2703), .ZN(n3945) );
  NOR2_X1 U34890 ( .A1(n2705), .A2(n3945), .ZN(n3826) );
  INV_X1 U3490 ( .A(n3826), .ZN(n2706) );
  NOR2_X1 U34910 ( .A1(n4116), .A2(n4140), .ZN(n3883) );
  NOR2_X1 U3492 ( .A1(n4304), .A2(n4160), .ZN(n4128) );
  NOR2_X1 U34930 ( .A1(n3883), .A2(n4128), .ZN(n3944) );
  INV_X1 U3494 ( .A(n3944), .ZN(n2708) );
  NAND2_X1 U34950 ( .A1(n4116), .A2(n4140), .ZN(n3816) );
  OAI21_X1 U3496 ( .B1(n4129), .B2(n2708), .A(n3816), .ZN(n4113) );
  AND2_X1 U34970 ( .A1(n4101), .A2(n4122), .ZN(n3846) );
  OR2_X1 U3498 ( .A1(n4101), .A2(n4122), .ZN(n3847) );
  INV_X1 U34990 ( .A(n3847), .ZN(n4095) );
  AOI21_X1 U3500 ( .B1(n4119), .B2(n4100), .A(n4095), .ZN(n3953) );
  INV_X1 U35010 ( .A(n3953), .ZN(n2710) );
  AND2_X1 U3502 ( .A1(n4287), .A2(n4105), .ZN(n3834) );
  INV_X1 U35030 ( .A(n3834), .ZN(n2709) );
  NOR2_X1 U3504 ( .A1(n4281), .A2(n4286), .ZN(n3951) );
  INV_X1 U35050 ( .A(n3835), .ZN(n2711) );
  XNOR2_X1 U35060 ( .A(n2712), .B(n3878), .ZN(n2714) );
  NAND2_X1 U35070 ( .A1(n3969), .A2(n4412), .ZN(n2713) );
  INV_X1 U35080 ( .A(n2676), .ZN(n4411) );
  NAND2_X1 U35090 ( .A1(n4410), .A2(n4411), .ZN(n3844) );
  NAND2_X1 U35100 ( .A1(n2714), .A2(n4254), .ZN(n2720) );
  INV_X1 U35110 ( .A(REG1_REG_30__SCAN_IN), .ZN(n2717) );
  NAND2_X1 U35120 ( .A1(n2409), .A2(REG2_REG_30__SCAN_IN), .ZN(n2716) );
  NAND2_X1 U35130 ( .A1(n2416), .A2(REG0_REG_30__SCAN_IN), .ZN(n2715) );
  OAI211_X1 U35140 ( .C1(n2872), .C2(n2717), .A(n2716), .B(n2715), .ZN(n3843)
         );
  XNOR2_X1 U35150 ( .A(n2718), .B(IR_REG_27__SCAN_IN), .ZN(n4423) );
  NAND2_X1 U35160 ( .A1(n2938), .A2(n2782), .ZN(n4307) );
  AOI21_X1 U35170 ( .B1(B_REG_SCAN_IN), .B2(n4423), .A(n4307), .ZN(n4055) );
  INV_X1 U35180 ( .A(n2762), .ZN(n3833) );
  AOI22_X1 U35190 ( .A1(n3843), .A2(n4055), .B1(n4342), .B2(n3833), .ZN(n2719)
         );
  NOR2_X1 U35200 ( .A1(n2722), .A2(n2194), .ZN(n2723) );
  NAND2_X1 U35210 ( .A1(n3624), .A2(B_REG_SCAN_IN), .ZN(n2736) );
  NAND2_X1 U35220 ( .A1(n2731), .A2(n2730), .ZN(n2732) );
  NAND2_X1 U35230 ( .A1(n2743), .A2(n2744), .ZN(n2733) );
  INV_X1 U35240 ( .A(n2738), .ZN(n2810) );
  MUX2_X1 U35250 ( .A(n2736), .B(B_REG_SCAN_IN), .S(n2810), .Z(n2737) );
  NAND2_X1 U35260 ( .A1(n3624), .A2(n2759), .ZN(n2923) );
  NAND2_X1 U35270 ( .A1(n2989), .A2(n2923), .ZN(n2758) );
  NAND2_X2 U35280 ( .A1(n2810), .A2(n2741), .ZN(n2769) );
  NAND2_X1 U35290 ( .A1(n4579), .A2(n2745), .ZN(n2932) );
  NAND2_X1 U35300 ( .A1(n2676), .A2(n4050), .ZN(n2920) );
  NAND2_X1 U35310 ( .A1(n2782), .A2(n2920), .ZN(n2986) );
  NAND2_X1 U35320 ( .A1(n2932), .A2(n2986), .ZN(n2746) );
  NOR2_X1 U35330 ( .A1(n2988), .A2(n2746), .ZN(n2757) );
  NOR3_X1 U35340 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_29__SCAN_IN), .ZN(n4865) );
  NOR3_X1 U35350 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .ZN(n2749) );
  NOR4_X1 U35360 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_17__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2748) );
  NOR4_X1 U35370 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2747) );
  NAND4_X1 U35380 ( .A1(n4865), .A2(n2749), .A3(n2748), .A4(n2747), .ZN(n2755)
         );
  NOR4_X1 U35390 ( .A1(D_REG_8__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n2753) );
  NOR4_X1 U35400 ( .A1(D_REG_3__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2752) );
  NOR4_X1 U35410 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2751) );
  NOR4_X1 U35420 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2750) );
  NAND4_X1 U35430 ( .A1(n2753), .A2(n2752), .A3(n2751), .A4(n2750), .ZN(n2754)
         );
  NOR2_X1 U35440 ( .A1(n2755), .A2(n2754), .ZN(n2756) );
  NAND3_X1 U35450 ( .A1(n2758), .A2(n2757), .A3(n2924), .ZN(n2765) );
  NAND2_X1 U35460 ( .A1(n2738), .A2(n2759), .ZN(n2814) );
  MUX2_X1 U35470 ( .A(n2761), .B(n2766), .S(n4599), .Z(n2764) );
  NAND2_X1 U35480 ( .A1(n3085), .A2(n3193), .ZN(n3140) );
  INV_X1 U35490 ( .A(n3409), .ZN(n3288) );
  NAND2_X1 U35500 ( .A1(n2764), .A2(n2763), .ZN(U3547) );
  AND2_X4 U35510 ( .A1(n2769), .A2(n2768), .ZN(n3594) );
  INV_X1 U35520 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2774) );
  NAND2_X1 U35530 ( .A1(n2951), .A2(n2776), .ZN(n2777) );
  OAI21_X1 U35540 ( .B1(n2778), .B2(n2777), .A(n2954), .ZN(n2940) );
  INV_X1 U35550 ( .A(n2938), .ZN(n2957) );
  INV_X1 U35560 ( .A(n4423), .ZN(n2790) );
  NAND3_X1 U35570 ( .A1(n2940), .A2(n2957), .A3(n2790), .ZN(n2781) );
  NOR2_X1 U35580 ( .A1(n2938), .A2(n2790), .ZN(n3966) );
  AND2_X1 U35590 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n2824) );
  INV_X1 U35600 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3012) );
  AND2_X1 U35610 ( .A1(n4423), .A2(n3012), .ZN(n2779) );
  OR2_X1 U35620 ( .A1(n2938), .A2(n2779), .ZN(n4424) );
  AOI22_X1 U35630 ( .A1(n3966), .A2(n2824), .B1(n4424), .B2(n4428), .ZN(n2780)
         );
  NAND3_X1 U35640 ( .A1(n2781), .A2(n3985), .A3(n2780), .ZN(n2918) );
  INV_X1 U35650 ( .A(n2918), .ZN(n2800) );
  OR2_X1 U35660 ( .A1(n3069), .A2(U3149), .ZN(n3971) );
  NAND2_X1 U35670 ( .A1(n2988), .A2(n3971), .ZN(n2795) );
  NAND2_X1 U35680 ( .A1(n2782), .A2(n3069), .ZN(n2783) );
  AND2_X1 U35690 ( .A1(n2783), .A2(n2137), .ZN(n2793) );
  INV_X1 U35700 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2784) );
  MUX2_X1 U35710 ( .A(n2784), .B(REG2_REG_1__SCAN_IN), .S(n2830), .Z(n2823) );
  NAND2_X1 U35720 ( .A1(n2823), .A2(n2824), .ZN(n2822) );
  INV_X1 U35730 ( .A(n2830), .ZN(n4417) );
  NAND2_X1 U35740 ( .A1(n4417), .A2(REG2_REG_1__SCAN_IN), .ZN(n2788) );
  NAND2_X1 U35750 ( .A1(n2822), .A2(n2788), .ZN(n2786) );
  INV_X1 U35760 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3053) );
  MUX2_X1 U35770 ( .A(n3053), .B(REG2_REG_2__SCAN_IN), .S(n2831), .Z(n2785) );
  NAND2_X1 U35780 ( .A1(n2786), .A2(n2785), .ZN(n2833) );
  MUX2_X1 U35790 ( .A(REG2_REG_2__SCAN_IN), .B(n3053), .S(n2831), .Z(n2787) );
  NAND3_X1 U35800 ( .A1(n2822), .A2(n2788), .A3(n2787), .ZN(n2789) );
  AND3_X1 U35810 ( .A1(n4522), .A2(n2833), .A3(n2789), .ZN(n2799) );
  NAND2_X1 U3582 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n2821) );
  AOI21_X1 U3583 ( .B1(REG1_REG_1__SCAN_IN), .B2(n4417), .A(n2819), .ZN(n2792)
         );
  XOR2_X1 U3584 ( .A(REG1_REG_2__SCAN_IN), .B(n2831), .Z(n2791) );
  NOR2_X1 U3585 ( .A1(n2792), .A2(n2791), .ZN(n2834) );
  AOI211_X1 U3586 ( .C1(n2792), .C2(n2791), .A(n2834), .B(n4518), .ZN(n2798)
         );
  INV_X1 U3587 ( .A(n2793), .ZN(n2794) );
  AOI22_X1 U3588 ( .A1(n4531), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n2796) );
  OAI21_X1 U3589 ( .B1(n4538), .B2(n2831), .A(n2796), .ZN(n2797) );
  OR4_X1 U3590 ( .A1(n2800), .A2(n2799), .A3(n2798), .A4(n2797), .ZN(U3242) );
  MUX2_X1 U3591 ( .A(n2434), .B(n2912), .S(STATE_REG_SCAN_IN), .Z(n2801) );
  INV_X1 U3592 ( .A(n2801), .ZN(U3348) );
  MUX2_X1 U3593 ( .A(n2831), .B(n2415), .S(U3149), .Z(n2802) );
  INV_X1 U3594 ( .A(n2802), .ZN(U3350) );
  INV_X1 U3595 ( .A(n2854), .ZN(n2901) );
  INV_X1 U3596 ( .A(DATAI_6_), .ZN(n2803) );
  MUX2_X1 U3597 ( .A(n2901), .B(n2803), .S(U3149), .Z(n2804) );
  INV_X1 U3598 ( .A(n2804), .ZN(U3346) );
  MUX2_X1 U3599 ( .A(n4470), .B(n2512), .S(U3149), .Z(n2805) );
  INV_X1 U3600 ( .A(n2805), .ZN(U3341) );
  INV_X1 U3601 ( .A(DATAI_22_), .ZN(n4611) );
  NAND2_X1 U3602 ( .A1(n3969), .A2(STATE_REG_SCAN_IN), .ZN(n2806) );
  OAI21_X1 U3603 ( .B1(STATE_REG_SCAN_IN), .B2(n4611), .A(n2806), .ZN(U3330)
         );
  INV_X1 U3604 ( .A(DATAI_26_), .ZN(n4608) );
  NAND2_X1 U3605 ( .A1(n2739), .A2(STATE_REG_SCAN_IN), .ZN(n2807) );
  OAI21_X1 U3606 ( .B1(STATE_REG_SCAN_IN), .B2(n4608), .A(n2807), .ZN(U3326)
         );
  INV_X1 U3607 ( .A(DATAI_27_), .ZN(n4605) );
  NAND2_X1 U3608 ( .A1(n4423), .A2(STATE_REG_SCAN_IN), .ZN(n2808) );
  OAI21_X1 U3609 ( .B1(STATE_REG_SCAN_IN), .B2(n4605), .A(n2808), .ZN(U3325)
         );
  INV_X1 U3610 ( .A(DATAI_31_), .ZN(n4602) );
  OR4_X1 U3611 ( .A1(n2379), .A2(IR_REG_30__SCAN_IN), .A3(U3149), .A4(n2194), 
        .ZN(n2809) );
  OAI21_X1 U3612 ( .B1(STATE_REG_SCAN_IN), .B2(n4602), .A(n2809), .ZN(U3321)
         );
  INV_X1 U3613 ( .A(DATAI_24_), .ZN(n4861) );
  NAND2_X1 U3614 ( .A1(n2810), .A2(STATE_REG_SCAN_IN), .ZN(n2811) );
  OAI21_X1 U3615 ( .B1(STATE_REG_SCAN_IN), .B2(n4861), .A(n2811), .ZN(U3328)
         );
  INV_X1 U3616 ( .A(DATAI_28_), .ZN(n4606) );
  NAND2_X1 U3617 ( .A1(n2957), .A2(STATE_REG_SCAN_IN), .ZN(n2812) );
  OAI21_X1 U3618 ( .B1(STATE_REG_SCAN_IN), .B2(n4606), .A(n2812), .ZN(U3324)
         );
  INV_X1 U3619 ( .A(n2988), .ZN(n2930) );
  INV_X1 U3620 ( .A(D_REG_0__SCAN_IN), .ZN(n4666) );
  INV_X1 U3621 ( .A(n2814), .ZN(n2815) );
  AOI22_X1 U3622 ( .A1(n4549), .A2(n4666), .B1(n2815), .B2(n2816), .ZN(U3458)
         );
  INV_X1 U3623 ( .A(D_REG_1__SCAN_IN), .ZN(n2818) );
  INV_X1 U3624 ( .A(n2923), .ZN(n2817) );
  AOI22_X1 U3625 ( .A1(n4549), .A2(n2818), .B1(n2817), .B2(n2816), .ZN(U3459)
         );
  NOR2_X1 U3626 ( .A1(n4531), .A2(U4043), .ZN(U3148) );
  AOI211_X1 U3627 ( .C1(n2821), .C2(n2820), .A(n2819), .B(n4518), .ZN(n2827)
         );
  OAI211_X1 U3628 ( .C1(n2824), .C2(n2823), .A(n4522), .B(n2822), .ZN(n2825)
         );
  INV_X1 U3629 ( .A(n2825), .ZN(n2826) );
  NOR2_X1 U3630 ( .A1(n2827), .A2(n2826), .ZN(n2829) );
  AOI22_X1 U3631 ( .A1(n4531), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n2828) );
  OAI211_X1 U3632 ( .C1(n2830), .C2(n4538), .A(n2829), .B(n2828), .ZN(U3241)
         );
  INV_X1 U3633 ( .A(n4416), .ZN(n2842) );
  INV_X1 U3634 ( .A(n2831), .ZN(n2835) );
  NAND2_X1 U3635 ( .A1(n2835), .A2(REG2_REG_2__SCAN_IN), .ZN(n2832) );
  NAND2_X1 U3636 ( .A1(n2833), .A2(n2832), .ZN(n2844) );
  XNOR2_X1 U3637 ( .A(n2844), .B(n2842), .ZN(n2843) );
  XOR2_X1 U3638 ( .A(REG2_REG_3__SCAN_IN), .B(n2843), .Z(n2839) );
  INV_X1 U3639 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2837) );
  AOI211_X1 U3640 ( .C1(n2837), .C2(n2836), .A(n2852), .B(n4518), .ZN(n2838)
         );
  AOI21_X1 U3641 ( .B1(n4522), .B2(n2839), .A(n2838), .ZN(n2841) );
  AOI22_X1 U3642 ( .A1(n4531), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n2840) );
  OAI211_X1 U3643 ( .C1(n2842), .C2(n4538), .A(n2841), .B(n2840), .ZN(U3243)
         );
  NAND2_X1 U3644 ( .A1(n2843), .A2(REG2_REG_3__SCAN_IN), .ZN(n2846) );
  NAND2_X1 U3645 ( .A1(n2844), .A2(n4416), .ZN(n2845) );
  NAND2_X1 U3646 ( .A1(n2846), .A2(n2845), .ZN(n2847) );
  XNOR2_X1 U3647 ( .A(n2847), .B(n2912), .ZN(n2909) );
  NAND2_X1 U3648 ( .A1(n2847), .A2(n2182), .ZN(n2848) );
  INV_X1 U3649 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2850) );
  MUX2_X1 U3650 ( .A(n2850), .B(REG2_REG_5__SCAN_IN), .S(n2891), .Z(n2849) );
  XNOR2_X1 U3651 ( .A(n2900), .B(n2854), .ZN(n2903) );
  XOR2_X1 U3652 ( .A(REG2_REG_6__SCAN_IN), .B(n2903), .Z(n2861) );
  INV_X1 U3653 ( .A(n2891), .ZN(n4415) );
  INV_X1 U3654 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4718) );
  NOR2_X1 U3655 ( .A1(n2914), .A2(n4718), .ZN(n2913) );
  XOR2_X1 U3656 ( .A(REG1_REG_5__SCAN_IN), .B(n2891), .Z(n2886) );
  NOR2_X1 U3657 ( .A1(n2887), .A2(n2886), .ZN(n2885) );
  INV_X1 U3658 ( .A(n2855), .ZN(n2856) );
  INV_X1 U3659 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3090) );
  OAI211_X1 U3660 ( .C1(REG1_REG_6__SCAN_IN), .C2(n2856), .A(n2896), .B(n4533), 
        .ZN(n2860) );
  NOR2_X1 U3661 ( .A1(STATE_REG_SCAN_IN), .A2(n2857), .ZN(n3171) );
  NOR2_X1 U3662 ( .A1(n4538), .A2(n2901), .ZN(n2858) );
  AOI211_X1 U3663 ( .C1(n4531), .C2(ADDR_REG_6__SCAN_IN), .A(n3171), .B(n2858), 
        .ZN(n2859) );
  OAI211_X1 U3664 ( .C1(n2861), .C2(n4527), .A(n2860), .B(n2859), .ZN(U3246)
         );
  INV_X1 U3665 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n4789) );
  NAND2_X1 U3666 ( .A1(n4345), .A2(U4043), .ZN(n2862) );
  OAI21_X1 U3667 ( .B1(U4043), .B2(n4789), .A(n2862), .ZN(U3568) );
  INV_X1 U3668 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n4828) );
  NAND2_X1 U3669 ( .A1(n4322), .A2(U4043), .ZN(n2863) );
  OAI21_X1 U3670 ( .B1(U4043), .B2(n4828), .A(n2863), .ZN(U3572) );
  INV_X1 U3671 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n4807) );
  NAND2_X1 U3672 ( .A1(n3843), .A2(n3985), .ZN(n2864) );
  OAI21_X1 U3673 ( .B1(n3985), .B2(n4807), .A(n2864), .ZN(U3580) );
  INV_X1 U3674 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n4830) );
  NAND2_X1 U3675 ( .A1(n3670), .A2(n3985), .ZN(n2865) );
  OAI21_X1 U3676 ( .B1(U4043), .B2(n4830), .A(n2865), .ZN(U3561) );
  INV_X1 U3677 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n4787) );
  NAND2_X1 U3678 ( .A1(n3399), .A2(n3985), .ZN(n2866) );
  OAI21_X1 U3679 ( .B1(U4043), .B2(n4787), .A(n2866), .ZN(U3560) );
  INV_X1 U3680 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n4829) );
  NAND2_X1 U3681 ( .A1(n3307), .A2(n3985), .ZN(n2867) );
  OAI21_X1 U3682 ( .B1(n3985), .B2(n4829), .A(n2867), .ZN(U3557) );
  INV_X1 U3683 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n4833) );
  NAND2_X1 U3684 ( .A1(n3150), .A2(n3985), .ZN(n2868) );
  OAI21_X1 U3685 ( .B1(n3985), .B2(n4833), .A(n2868), .ZN(U3553) );
  INV_X1 U3686 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n4832) );
  NAND2_X1 U3687 ( .A1(n3027), .A2(n3985), .ZN(n2869) );
  OAI21_X1 U3688 ( .B1(n3985), .B2(n4832), .A(n2869), .ZN(U3552) );
  INV_X1 U3689 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n4801) );
  INV_X1 U3690 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4266) );
  NAND2_X1 U3691 ( .A1(n2648), .A2(REG2_REG_31__SCAN_IN), .ZN(n2871) );
  NAND2_X1 U3692 ( .A1(n2416), .A2(REG0_REG_31__SCAN_IN), .ZN(n2870) );
  OAI211_X1 U3693 ( .C1(n2872), .C2(n4266), .A(n2871), .B(n2870), .ZN(n4056)
         );
  NAND2_X1 U3694 ( .A1(n4056), .A2(n3985), .ZN(n2873) );
  OAI21_X1 U3695 ( .B1(n3985), .B2(n4801), .A(n2873), .ZN(U3581) );
  INV_X1 U3696 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n4831) );
  NAND2_X1 U3697 ( .A1(n3239), .A2(n3985), .ZN(n2874) );
  OAI21_X1 U3698 ( .B1(n3985), .B2(n4831), .A(n2874), .ZN(U3556) );
  INV_X1 U3699 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n4834) );
  NAND2_X1 U3700 ( .A1(n2773), .A2(n3985), .ZN(n2875) );
  OAI21_X1 U3701 ( .B1(U4043), .B2(n4834), .A(n2875), .ZN(U3550) );
  NAND2_X1 U3702 ( .A1(n2773), .A2(n4303), .ZN(n2878) );
  NAND2_X1 U3703 ( .A1(n3027), .A2(n4344), .ZN(n2877) );
  OAI211_X1 U3704 ( .C1(n4273), .C2(n2403), .A(n2878), .B(n2877), .ZN(n2879)
         );
  INV_X1 U3705 ( .A(n2879), .ZN(n2882) );
  NAND2_X1 U3706 ( .A1(n2880), .A2(n4254), .ZN(n2881) );
  OAI211_X1 U3707 ( .C1(n2996), .C2(n4210), .A(n2882), .B(n2881), .ZN(n2994)
         );
  OAI21_X1 U3708 ( .B1(n3005), .B2(n2403), .A(n3055), .ZN(n3002) );
  OAI22_X1 U3709 ( .A1(n2996), .A2(n4565), .B1(n3139), .B2(n3002), .ZN(n2883)
         );
  NOR2_X1 U3710 ( .A1(n2994), .A2(n2883), .ZN(n4569) );
  NAND2_X1 U3711 ( .A1(n4596), .A2(REG1_REG_1__SCAN_IN), .ZN(n2884) );
  OAI21_X1 U3712 ( .B1(n4569), .B2(n4596), .A(n2884), .ZN(U3519) );
  AOI211_X1 U3713 ( .C1(n2887), .C2(n2886), .A(n4518), .B(n2885), .ZN(n2894)
         );
  MUX2_X1 U3714 ( .A(REG2_REG_5__SCAN_IN), .B(n2850), .S(n2891), .Z(n2889) );
  AOI211_X1 U3715 ( .C1(n2170), .C2(n2889), .A(n2888), .B(n4527), .ZN(n2893)
         );
  AND2_X1 U3716 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3115) );
  AOI21_X1 U3717 ( .B1(n4531), .B2(ADDR_REG_5__SCAN_IN), .A(n3115), .ZN(n2890)
         );
  OAI21_X1 U3718 ( .B1(n4538), .B2(n2891), .A(n2890), .ZN(n2892) );
  OR3_X1 U3719 ( .A1(n2894), .A2(n2893), .A3(n2892), .ZN(U3245) );
  INV_X1 U3720 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n4792) );
  NAND2_X1 U3721 ( .A1(n4304), .A2(U4043), .ZN(n2895) );
  OAI21_X1 U3722 ( .B1(n3985), .B2(n4792), .A(n2895), .ZN(U3573) );
  INV_X1 U3723 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4597) );
  MUX2_X1 U3724 ( .A(n4597), .B(REG1_REG_7__SCAN_IN), .S(n4414), .Z(n2898) );
  XNOR2_X1 U3725 ( .A(n4008), .B(n2898), .ZN(n2908) );
  AND2_X1 U3726 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3238) );
  NOR2_X1 U3727 ( .A1(n4538), .A2(n4414), .ZN(n2899) );
  AOI211_X1 U3728 ( .C1(n4531), .C2(ADDR_REG_7__SCAN_IN), .A(n3238), .B(n2899), 
        .ZN(n2907) );
  INV_X1 U3729 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3987) );
  MUX2_X1 U3730 ( .A(n3987), .B(REG2_REG_7__SCAN_IN), .S(n4414), .Z(n2905) );
  INV_X1 U3731 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3191) );
  INV_X1 U3732 ( .A(n2900), .ZN(n2902) );
  OAI22_X1 U3733 ( .A1(n2903), .A2(n3191), .B1(n2902), .B2(n2901), .ZN(n2904)
         );
  NAND2_X1 U3734 ( .A1(n2904), .A2(n2905), .ZN(n3986) );
  OAI211_X1 U3735 ( .C1(n2905), .C2(n2904), .A(n4522), .B(n3986), .ZN(n2906)
         );
  OAI211_X1 U3736 ( .C1(n2908), .C2(n4518), .A(n2907), .B(n2906), .ZN(U3247)
         );
  XOR2_X1 U3737 ( .A(REG2_REG_4__SCAN_IN), .B(n2909), .Z(n2917) );
  NAND2_X1 U3738 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3152) );
  INV_X1 U3739 ( .A(n3152), .ZN(n2910) );
  AOI21_X1 U3740 ( .B1(n4531), .B2(ADDR_REG_4__SCAN_IN), .A(n2910), .ZN(n2911)
         );
  OAI21_X1 U3741 ( .B1(n4538), .B2(n2912), .A(n2911), .ZN(n2916) );
  AOI211_X1 U3742 ( .C1(n4718), .C2(n2914), .A(n4518), .B(n2913), .ZN(n2915)
         );
  AOI211_X1 U3743 ( .C1(n4522), .C2(n2917), .A(n2916), .B(n2915), .ZN(n2919)
         );
  NAND2_X1 U3744 ( .A1(n2919), .A2(n2918), .ZN(U3244) );
  NAND2_X1 U3745 ( .A1(n3003), .A2(n2920), .ZN(n2921) );
  AND2_X1 U3746 ( .A1(n2922), .A2(n2921), .ZN(n2935) );
  NAND3_X1 U3747 ( .A1(n2925), .A2(n2992), .A3(n2989), .ZN(n2959) );
  OAI21_X1 U3748 ( .B1(n2935), .B2(n4342), .A(n2959), .ZN(n2926) );
  NAND2_X1 U3749 ( .A1(n2926), .A2(n2986), .ZN(n3071) );
  INV_X1 U3750 ( .A(n3071), .ZN(n2931) );
  INV_X1 U3751 ( .A(n3604), .ZN(n2927) );
  OR2_X1 U3752 ( .A1(n2949), .A2(n4551), .ZN(n2929) );
  NAND2_X1 U3753 ( .A1(n2959), .A2(n3967), .ZN(n3072) );
  NAND3_X1 U3754 ( .A1(n2931), .A2(n2930), .A3(n3072), .ZN(n2979) );
  INV_X1 U3755 ( .A(n2979), .ZN(n2966) );
  INV_X1 U3756 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2943) );
  NOR3_X1 U3757 ( .A1(n2959), .A2(n2988), .A3(n4273), .ZN(n2933) );
  INV_X1 U3758 ( .A(n2935), .ZN(n2936) );
  OR2_X1 U3759 ( .A1(n2988), .A2(n2936), .ZN(n2937) );
  INV_X1 U3760 ( .A(n2946), .ZN(n3049) );
  NAND2_X1 U3761 ( .A1(n3967), .A2(n2938), .ZN(n2939) );
  OAI22_X1 U3762 ( .A1(n2940), .A2(n3800), .B1(n3049), .B2(n3795), .ZN(n2941)
         );
  AOI21_X1 U3763 ( .B1(n3004), .B2(n3729), .A(n2941), .ZN(n2942) );
  OAI21_X1 U3764 ( .B1(n2966), .B2(n2943), .A(n2942), .ZN(U3229) );
  INV_X1 U3765 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2965) );
  NOR2_X1 U3766 ( .A1(n2927), .A2(n2403), .ZN(n2944) );
  AOI21_X1 U3767 ( .B1(n2946), .B2(n2136), .A(n2944), .ZN(n2947) );
  AOI22_X1 U3768 ( .A1(n2948), .A2(n2134), .B1(n2962), .B2(n3594), .ZN(n2950)
         );
  XNOR2_X1 U3769 ( .A(n2950), .B(n3628), .ZN(n2969) );
  XNOR2_X1 U3770 ( .A(n2971), .B(n2969), .ZN(n2955) );
  NAND2_X1 U3771 ( .A1(n2954), .A2(n2953), .ZN(n2956) );
  NAND2_X1 U3772 ( .A1(n2956), .A2(n2955), .ZN(n2973) );
  OAI211_X1 U3773 ( .C1(n2955), .C2(n2956), .A(n2973), .B(n3805), .ZN(n2964)
         );
  NAND2_X1 U3774 ( .A1(n3967), .A2(n2957), .ZN(n2958) );
  INV_X1 U3775 ( .A(n3027), .ZN(n3068) );
  OAI22_X1 U3776 ( .A1(n2960), .A2(n3807), .B1(n3795), .B2(n3068), .ZN(n2961)
         );
  AOI21_X1 U3777 ( .B1(n3729), .B2(n2962), .A(n2961), .ZN(n2963) );
  OAI211_X1 U3778 ( .C1(n2966), .C2(n2965), .A(n2964), .B(n2963), .ZN(U3219)
         );
  AOI22_X1 U3779 ( .A1(n3027), .A2(n3604), .B1(n3594), .B2(n3056), .ZN(n2967)
         );
  XNOR2_X1 U3780 ( .A(n2967), .B(n2133), .ZN(n3065) );
  AOI22_X1 U3781 ( .A1(n3027), .A2(n2945), .B1(n3604), .B2(n3056), .ZN(n3064)
         );
  XNOR2_X1 U3782 ( .A(n3065), .B(n3064), .ZN(n2975) );
  NAND2_X1 U3783 ( .A1(n2973), .A2(n2972), .ZN(n2974) );
  AOI21_X1 U3784 ( .B1(n2975), .B2(n2974), .A(n3067), .ZN(n2981) );
  OAI22_X1 U3785 ( .A1(n3063), .A2(n3795), .B1(n3807), .B2(n3049), .ZN(n2978)
         );
  NOR2_X1 U3786 ( .A1(n2934), .A2(n2976), .ZN(n2977) );
  AOI211_X1 U3787 ( .C1(REG3_REG_2__SCAN_IN), .C2(n2979), .A(n2978), .B(n2977), 
        .ZN(n2980) );
  OAI21_X1 U3788 ( .B1(n2981), .B2(n3800), .A(n2980), .ZN(U3234) );
  INV_X1 U3789 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n4795) );
  NAND2_X1 U3790 ( .A1(n4287), .A2(n3985), .ZN(n2982) );
  OAI21_X1 U3791 ( .B1(n3985), .B2(n4795), .A(n2982), .ZN(U3576) );
  INV_X1 U3792 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n4794) );
  NAND2_X1 U3793 ( .A1(n3642), .A2(n3985), .ZN(n2983) );
  OAI21_X1 U3794 ( .B1(n3985), .B2(n4794), .A(n2983), .ZN(U3577) );
  INV_X1 U3795 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n4808) );
  NAND2_X1 U3796 ( .A1(n4278), .A2(n3985), .ZN(n2984) );
  OAI21_X1 U3797 ( .B1(n3985), .B2(n4808), .A(n2984), .ZN(U3579) );
  INV_X1 U3798 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n4791) );
  NAND2_X1 U3799 ( .A1(n4101), .A2(U4043), .ZN(n2985) );
  OAI21_X1 U3800 ( .B1(n3985), .B2(n4791), .A(n2985), .ZN(U3575) );
  INV_X1 U3801 ( .A(n2986), .ZN(n2987) );
  NOR2_X1 U3802 ( .A1(n2988), .A2(n2987), .ZN(n2991) );
  NAND4_X1 U3803 ( .A1(n2992), .A2(n2991), .A3(n2990), .A4(n2989), .ZN(n2993)
         );
  NAND2_X1 U3804 ( .A1(n4421), .A2(n4050), .ZN(n4261) );
  MUX2_X1 U3805 ( .A(n2994), .B(REG2_REG_1__SCAN_IN), .S(n4222), .Z(n2995) );
  INV_X1 U3806 ( .A(n2995), .ZN(n3001) );
  INV_X1 U3807 ( .A(n2996), .ZN(n2999) );
  NAND2_X1 U3808 ( .A1(n2997), .A2(n4412), .ZN(n3146) );
  INV_X1 U3809 ( .A(n3146), .ZN(n2998) );
  NAND2_X1 U3810 ( .A1(n4421), .A2(n2998), .ZN(n4219) );
  INV_X1 U3811 ( .A(n4219), .ZN(n4544) );
  AOI22_X1 U3812 ( .A1(n2999), .A2(n4544), .B1(REG3_REG_1__SCAN_IN), .B2(n4539), .ZN(n3000) );
  OAI211_X1 U3813 ( .C1(n4238), .C2(n3002), .A(n3001), .B(n3000), .ZN(U3289)
         );
  NAND2_X1 U3814 ( .A1(n3004), .A2(n3003), .ZN(n4563) );
  NAND2_X1 U3815 ( .A1(n2773), .A2(n3005), .ZN(n3890) );
  NAND2_X1 U3816 ( .A1(n3888), .A2(n3890), .ZN(n3009) );
  INV_X1 U3817 ( .A(n3009), .ZN(n4566) );
  AOI21_X1 U3818 ( .B1(n4233), .B2(n4210), .A(n4566), .ZN(n3006) );
  AOI21_X1 U3819 ( .B1(n4344), .B2(n2946), .A(n3006), .ZN(n4564) );
  OAI21_X1 U3820 ( .B1(n3007), .B2(n4563), .A(n4564), .ZN(n3008) );
  AOI22_X1 U3821 ( .A1(n3008), .A2(n4421), .B1(REG3_REG_0__SCAN_IN), .B2(n4539), .ZN(n3011) );
  NAND2_X1 U3822 ( .A1(n4544), .A2(n3009), .ZN(n3010) );
  OAI211_X1 U3823 ( .C1(n4421), .C2(n3012), .A(n3011), .B(n3010), .ZN(U3290)
         );
  NAND2_X1 U3824 ( .A1(n3914), .A2(n3900), .ZN(n3014) );
  INV_X1 U3825 ( .A(n3014), .ZN(n3857) );
  XNOR2_X1 U3826 ( .A(n3013), .B(n3857), .ZN(n3175) );
  INV_X1 U3827 ( .A(n3099), .ZN(n3177) );
  XNOR2_X1 U3828 ( .A(n3015), .B(n3014), .ZN(n3016) );
  NAND2_X1 U3829 ( .A1(n3016), .A2(n4254), .ZN(n3183) );
  AOI22_X1 U3830 ( .A1(n3239), .A2(n4344), .B1(n4342), .B2(n3108), .ZN(n3017)
         );
  OAI211_X1 U3831 ( .C1(n3177), .C2(n4348), .A(n3183), .B(n3017), .ZN(n3018)
         );
  AOI21_X1 U3832 ( .B1(n3175), .B2(n4582), .A(n3018), .ZN(n3023) );
  INV_X1 U3833 ( .A(n4406), .ZN(n4574) );
  AND2_X1 U3834 ( .A1(n3118), .A2(n3108), .ZN(n3019) );
  NOR2_X1 U3835 ( .A1(n3085), .A2(n3019), .ZN(n3186) );
  AOI22_X1 U3836 ( .A1(n4574), .A2(n3186), .B1(REG0_REG_5__SCAN_IN), .B2(n4587), .ZN(n3020) );
  OAI21_X1 U3837 ( .B1(n3023), .B2(n4587), .A(n3020), .ZN(U3477) );
  NAND2_X1 U3838 ( .A1(n4596), .A2(REG1_REG_5__SCAN_IN), .ZN(n3022) );
  INV_X1 U3839 ( .A(n4338), .ZN(n4592) );
  NAND2_X1 U3840 ( .A1(n4592), .A2(n3186), .ZN(n3021) );
  OAI211_X1 U3841 ( .C1(n3023), .C2(n4596), .A(n3022), .B(n3021), .ZN(U3523)
         );
  OR2_X1 U3842 ( .A1(n3054), .A2(n3062), .ZN(n3024) );
  XNOR2_X1 U3843 ( .A(n3025), .B(n2145), .ZN(n3037) );
  XNOR2_X1 U3844 ( .A(n3026), .B(n2145), .ZN(n3031) );
  AOI22_X1 U3845 ( .A1(n3027), .A2(n4303), .B1(n4342), .B2(n3077), .ZN(n3028)
         );
  OAI21_X1 U3846 ( .B1(n3177), .B2(n4307), .A(n3028), .ZN(n3030) );
  NOR2_X1 U3847 ( .A1(n3037), .A2(n4210), .ZN(n3029) );
  AOI211_X1 U3848 ( .C1(n3031), .C2(n4254), .A(n3030), .B(n3029), .ZN(n3043)
         );
  OAI21_X1 U3849 ( .B1(n3037), .B2(n4565), .A(n3043), .ZN(n3034) );
  NAND2_X1 U3850 ( .A1(n3034), .A2(n4589), .ZN(n3033) );
  NAND2_X1 U3851 ( .A1(n4587), .A2(REG0_REG_3__SCAN_IN), .ZN(n3032) );
  OAI211_X1 U3852 ( .C1(n3039), .C2(n4406), .A(n3033), .B(n3032), .ZN(U3473)
         );
  NAND2_X1 U3853 ( .A1(n3034), .A2(n4599), .ZN(n3036) );
  NAND2_X1 U3854 ( .A1(n4596), .A2(REG1_REG_3__SCAN_IN), .ZN(n3035) );
  OAI211_X1 U3855 ( .C1(n4338), .C2(n3039), .A(n3036), .B(n3035), .ZN(U3521)
         );
  INV_X2 U3856 ( .A(n4421), .ZN(n4222) );
  INV_X1 U3857 ( .A(n3037), .ZN(n3041) );
  AOI22_X1 U3858 ( .A1(n4222), .A2(REG2_REG_3__SCAN_IN), .B1(n4539), .B2(n3074), .ZN(n3038) );
  OAI21_X1 U3859 ( .B1(n4238), .B2(n3039), .A(n3038), .ZN(n3040) );
  AOI21_X1 U3860 ( .B1(n3041), .B2(n4544), .A(n3040), .ZN(n3042) );
  OAI21_X1 U3861 ( .B1(n3043), .B2(n4222), .A(n3042), .ZN(U3287) );
  XNOR2_X1 U3862 ( .A(n3045), .B(n3044), .ZN(n4570) );
  OAI21_X1 U3863 ( .B1(n2683), .B2(n3047), .A(n3046), .ZN(n3052) );
  AOI22_X1 U3864 ( .A1(n3150), .A2(n4344), .B1(n3056), .B2(n4342), .ZN(n3048)
         );
  OAI21_X1 U3865 ( .B1(n3049), .B2(n4348), .A(n3048), .ZN(n3051) );
  NOR2_X1 U3866 ( .A1(n4570), .A2(n4210), .ZN(n3050) );
  AOI211_X1 U3867 ( .C1(n4254), .C2(n3052), .A(n3051), .B(n3050), .ZN(n4571)
         );
  MUX2_X1 U3868 ( .A(n3053), .B(n4571), .S(n4421), .Z(n3058) );
  AOI21_X1 U3869 ( .B1(n3056), .B2(n3055), .A(n3054), .ZN(n4591) );
  AOI22_X1 U3870 ( .A1(n4543), .A2(n4591), .B1(REG3_REG_2__SCAN_IN), .B2(n4539), .ZN(n3057) );
  OAI211_X1 U3871 ( .C1(n4570), .C2(n4219), .A(n3058), .B(n3057), .ZN(U3288)
         );
  NAND2_X1 U3872 ( .A1(n3150), .A2(n3604), .ZN(n3060) );
  NAND2_X1 U3873 ( .A1(n3594), .A2(n3077), .ZN(n3059) );
  NAND2_X1 U3874 ( .A1(n3060), .A2(n3059), .ZN(n3061) );
  XNOR2_X1 U3875 ( .A(n3061), .B(n2132), .ZN(n3095) );
  OAI22_X1 U3876 ( .A1(n3063), .A2(n3631), .B1(n3630), .B2(n3062), .ZN(n3094)
         );
  XNOR2_X1 U3877 ( .A(n3095), .B(n3094), .ZN(n3096) );
  NOR2_X2 U3878 ( .A1(n3067), .A2(n3066), .ZN(n3097) );
  XOR2_X1 U3879 ( .A(n3096), .B(n3097), .Z(n3079) );
  OAI22_X1 U3880 ( .A1(n3068), .A2(n3807), .B1(n3795), .B2(n3177), .ZN(n3076)
         );
  INV_X1 U3881 ( .A(n3069), .ZN(n3070) );
  NOR3_X1 U3882 ( .A1(n3071), .A2(n2775), .A3(n3070), .ZN(n3073) );
  MUX2_X1 U3883 ( .A(U3149), .B(n3746), .S(n3074), .Z(n3075) );
  AOI211_X1 U3884 ( .C1(n3077), .C2(n3729), .A(n3076), .B(n3075), .ZN(n3078)
         );
  OAI21_X1 U3885 ( .B1(n3079), .B2(n3800), .A(n3078), .ZN(U3215) );
  AND2_X1 U3886 ( .A1(n2208), .A2(n3903), .ZN(n3870) );
  XOR2_X1 U3887 ( .A(n3870), .B(n3080), .Z(n3203) );
  INV_X1 U3888 ( .A(n4582), .ZN(n4358) );
  XOR2_X1 U3889 ( .A(n3870), .B(n3081), .Z(n3201) );
  AOI22_X1 U3890 ( .A1(n3307), .A2(n4344), .B1(n3167), .B2(n4342), .ZN(n3082)
         );
  OAI21_X1 U3891 ( .B1(n3194), .B2(n4348), .A(n3082), .ZN(n3083) );
  AOI21_X1 U3892 ( .B1(n3201), .B2(n4254), .A(n3083), .ZN(n3084) );
  OAI21_X1 U3893 ( .B1(n3203), .B2(n4358), .A(n3084), .ZN(n3092) );
  OR2_X1 U3894 ( .A1(n3085), .A2(n3193), .ZN(n3086) );
  NAND2_X1 U3895 ( .A1(n3140), .A2(n3086), .ZN(n3198) );
  INV_X1 U3896 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3087) );
  OAI22_X1 U3897 ( .A1(n3198), .A2(n4406), .B1(n4589), .B2(n3087), .ZN(n3088)
         );
  AOI21_X1 U3898 ( .B1(n3092), .B2(n4589), .A(n3088), .ZN(n3089) );
  INV_X1 U3899 ( .A(n3089), .ZN(U3479) );
  OAI22_X1 U3900 ( .A1(n3198), .A2(n4338), .B1(n4599), .B2(n3090), .ZN(n3091)
         );
  AOI21_X1 U3901 ( .B1(n3092), .B2(n4599), .A(n3091), .ZN(n3093) );
  INV_X1 U3902 ( .A(n3093), .ZN(U3524) );
  INV_X1 U3903 ( .A(n3798), .ZN(n3815) );
  NOR2_X1 U3904 ( .A1(n3630), .A2(n3123), .ZN(n3098) );
  AOI21_X1 U3905 ( .B1(n3099), .B2(n2945), .A(n3098), .ZN(n3105) );
  NAND2_X1 U3906 ( .A1(n3099), .A2(n3604), .ZN(n3101) );
  NAND2_X1 U3907 ( .A1(n3594), .A2(n3151), .ZN(n3100) );
  NAND2_X1 U3908 ( .A1(n3101), .A2(n3100), .ZN(n3102) );
  XNOR2_X1 U3909 ( .A(n3102), .B(n2133), .ZN(n3104) );
  XOR2_X1 U3910 ( .A(n3105), .B(n3104), .Z(n3157) );
  INV_X1 U3911 ( .A(n3157), .ZN(n3103) );
  OR2_X1 U3912 ( .A1(n3194), .A2(n3631), .ZN(n3110) );
  NAND2_X1 U3913 ( .A1(n3604), .A2(n3108), .ZN(n3109) );
  NAND2_X1 U3914 ( .A1(n3110), .A2(n3109), .ZN(n3162) );
  OAI22_X1 U3915 ( .A1(n3194), .A2(n3630), .B1(n3627), .B2(n3176), .ZN(n3111)
         );
  XNOR2_X1 U3916 ( .A(n3111), .B(n2133), .ZN(n3163) );
  XOR2_X1 U3917 ( .A(n3162), .B(n3163), .Z(n3112) );
  OAI211_X1 U3918 ( .C1(n3113), .C2(n3112), .A(n3164), .B(n3805), .ZN(n3117)
         );
  INV_X1 U3919 ( .A(n3239), .ZN(n3178) );
  OAI22_X1 U3920 ( .A1(n2934), .A2(n3176), .B1(n3178), .B2(n3795), .ZN(n3114)
         );
  AOI211_X1 U3921 ( .C1(n3744), .C2(n3099), .A(n3115), .B(n3114), .ZN(n3116)
         );
  OAI211_X1 U3922 ( .C1(n3815), .C2(n3179), .A(n3117), .B(n3116), .ZN(U3224)
         );
  OAI211_X1 U3923 ( .C1(n3119), .C2(n3123), .A(n4354), .B(n3118), .ZN(n4576)
         );
  NOR2_X1 U3924 ( .A1(n4576), .A2(n4412), .ZN(n3131) );
  XNOR2_X1 U3925 ( .A(n3121), .B(n3120), .ZN(n3130) );
  NAND2_X1 U3926 ( .A1(n3150), .A2(n4303), .ZN(n3122) );
  OAI21_X1 U3927 ( .B1(n4273), .B2(n3123), .A(n3122), .ZN(n3128) );
  NAND2_X1 U3928 ( .A1(n3124), .A2(n3863), .ZN(n3125) );
  NAND2_X1 U3929 ( .A1(n3126), .A2(n3125), .ZN(n3132) );
  NOR2_X1 U3930 ( .A1(n3132), .A2(n4210), .ZN(n3127) );
  AOI211_X1 U3931 ( .C1(n4344), .C2(n3984), .A(n3128), .B(n3127), .ZN(n3129)
         );
  OAI21_X1 U3932 ( .B1(n4233), .B2(n3130), .A(n3129), .ZN(n4577) );
  AOI211_X1 U3933 ( .C1(n4539), .C2(n3160), .A(n3131), .B(n4577), .ZN(n3134)
         );
  INV_X1 U3934 ( .A(n3132), .ZN(n4580) );
  AOI22_X1 U3935 ( .A1(n4580), .A2(n4544), .B1(REG2_REG_4__SCAN_IN), .B2(n4222), .ZN(n3133) );
  OAI21_X1 U3936 ( .B1(n3134), .B2(n4222), .A(n3133), .ZN(U3286) );
  XNOR2_X1 U3937 ( .A(n3135), .B(n2363), .ZN(n3138) );
  AOI22_X1 U3938 ( .A1(n3983), .A2(n4344), .B1(n4342), .B2(n3231), .ZN(n3136)
         );
  OAI21_X1 U3939 ( .B1(n3178), .B2(n4348), .A(n3136), .ZN(n3137) );
  AOI21_X1 U3940 ( .B1(n3138), .B2(n4254), .A(n3137), .ZN(n4586) );
  NOR2_X1 U3941 ( .A1(n4421), .A2(n3987), .ZN(n3143) );
  AOI21_X1 U3942 ( .B1(n3140), .B2(n3231), .A(n3139), .ZN(n3141) );
  NAND2_X1 U3943 ( .A1(n3141), .A2(n3299), .ZN(n4585) );
  NOR2_X1 U3944 ( .A1(n4585), .A2(n4261), .ZN(n3142) );
  AOI211_X1 U3945 ( .C1(n4539), .C2(n3240), .A(n3143), .B(n3142), .ZN(n3149)
         );
  NAND2_X1 U3946 ( .A1(n3145), .A2(n2363), .ZN(n4583) );
  NAND2_X1 U3947 ( .A1(n4210), .A2(n3146), .ZN(n3147) );
  NAND3_X1 U3948 ( .A1(n3144), .A2(n4583), .A3(n4188), .ZN(n3148) );
  OAI211_X1 U3949 ( .C1(n4586), .C2(n4222), .A(n3149), .B(n3148), .ZN(U3283)
         );
  AOI22_X1 U3950 ( .A1(n3729), .A2(n3151), .B1(n3744), .B2(n3150), .ZN(n3153)
         );
  OAI211_X1 U3951 ( .C1(n3194), .C2(n3795), .A(n3153), .B(n3152), .ZN(n3159)
         );
  INV_X1 U3952 ( .A(n3155), .ZN(n3156) );
  AOI211_X1 U3953 ( .C1(n3157), .C2(n3154), .A(n3800), .B(n3156), .ZN(n3158)
         );
  AOI211_X1 U3954 ( .C1(n3160), .C2(n3798), .A(n3159), .B(n3158), .ZN(n3161)
         );
  INV_X1 U3955 ( .A(n3161), .ZN(U3227) );
  INV_X1 U3956 ( .A(n3162), .ZN(n3166) );
  INV_X1 U3957 ( .A(n3163), .ZN(n3165) );
  AOI22_X1 U3958 ( .A1(n3239), .A2(n3604), .B1(n3594), .B2(n3167), .ZN(n3168)
         );
  XOR2_X1 U3959 ( .A(n2133), .B(n3168), .Z(n3227) );
  OAI22_X1 U3960 ( .A1(n3178), .A2(n3631), .B1(n3630), .B2(n3193), .ZN(n3228)
         );
  INV_X1 U3961 ( .A(n3228), .ZN(n3230) );
  XNOR2_X1 U3962 ( .A(n3227), .B(n3230), .ZN(n3169) );
  XNOR2_X1 U3963 ( .A(n3229), .B(n3169), .ZN(n3174) );
  INV_X1 U3964 ( .A(n3307), .ZN(n3270) );
  OAI22_X1 U3965 ( .A1(n2934), .A2(n3193), .B1(n3270), .B2(n3795), .ZN(n3170)
         );
  AOI211_X1 U3966 ( .C1(n3744), .C2(n3984), .A(n3171), .B(n3170), .ZN(n3173)
         );
  NAND2_X1 U3967 ( .A1(n3746), .A2(n3189), .ZN(n3172) );
  OAI211_X1 U3968 ( .C1(n3174), .C2(n3800), .A(n3173), .B(n3172), .ZN(U3236)
         );
  INV_X1 U3969 ( .A(n3175), .ZN(n3188) );
  NAND2_X1 U3970 ( .A1(n4421), .A2(n4303), .ZN(n4197) );
  NAND2_X1 U3971 ( .A1(n4421), .A2(n4342), .ZN(n4196) );
  OAI22_X1 U3972 ( .A1(n3177), .A2(n4197), .B1(n4196), .B2(n3176), .ZN(n3182)
         );
  NAND2_X1 U3973 ( .A1(n4421), .A2(n4344), .ZN(n4193) );
  NOR2_X1 U3974 ( .A1(n4193), .A2(n3178), .ZN(n3181) );
  OAI22_X1 U3975 ( .A1(n4421), .A2(n2850), .B1(n3179), .B2(n4239), .ZN(n3180)
         );
  OR3_X1 U3976 ( .A1(n3182), .A2(n3181), .A3(n3180), .ZN(n3185) );
  NOR2_X1 U3977 ( .A1(n3183), .A2(n4222), .ZN(n3184) );
  AOI211_X1 U3978 ( .C1(n3186), .C2(n4543), .A(n3185), .B(n3184), .ZN(n3187)
         );
  OAI21_X1 U3979 ( .B1(n4265), .B2(n3188), .A(n3187), .ZN(U3285) );
  NAND2_X1 U3980 ( .A1(n4421), .A2(n4254), .ZN(n3298) );
  INV_X1 U3981 ( .A(n3298), .ZN(n3200) );
  INV_X1 U3982 ( .A(n4193), .ZN(n3292) );
  INV_X1 U3983 ( .A(n3189), .ZN(n3190) );
  OAI22_X1 U3984 ( .A1(n4421), .A2(n3191), .B1(n3190), .B2(n4239), .ZN(n3192)
         );
  AOI21_X1 U3985 ( .B1(n3292), .B2(n3307), .A(n3192), .ZN(n3197) );
  OAI22_X1 U3986 ( .A1(n3194), .A2(n4197), .B1(n4196), .B2(n3193), .ZN(n3195)
         );
  INV_X1 U3987 ( .A(n3195), .ZN(n3196) );
  OAI211_X1 U3988 ( .C1(n4238), .C2(n3198), .A(n3197), .B(n3196), .ZN(n3199)
         );
  AOI21_X1 U3989 ( .B1(n3201), .B2(n3200), .A(n3199), .ZN(n3202) );
  OAI21_X1 U3990 ( .B1(n4265), .B2(n3203), .A(n3202), .ZN(U3284) );
  AND2_X1 U3991 ( .A1(n2225), .A2(n3909), .ZN(n3864) );
  XNOR2_X1 U3992 ( .A(n3204), .B(n3864), .ZN(n3244) );
  INV_X1 U3993 ( .A(n3217), .ZN(n3205) );
  OAI21_X1 U3994 ( .B1(n3300), .B2(n3328), .A(n3205), .ZN(n3255) );
  INV_X1 U3995 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3206) );
  OAI22_X1 U3996 ( .A1(n3332), .A2(n4239), .B1(n3206), .B2(n4421), .ZN(n3208)
         );
  OAI22_X1 U3997 ( .A1(n3327), .A2(n4197), .B1(n4196), .B2(n3328), .ZN(n3207)
         );
  AOI211_X1 U3998 ( .C1(n3292), .C2(n3399), .A(n3208), .B(n3207), .ZN(n3209)
         );
  OAI21_X1 U3999 ( .B1(n3255), .B2(n4238), .A(n3209), .ZN(n3214) );
  INV_X1 U4000 ( .A(n3864), .ZN(n3210) );
  XNOR2_X1 U4001 ( .A(n3211), .B(n3210), .ZN(n3212) );
  NAND2_X1 U4002 ( .A1(n3212), .A2(n4254), .ZN(n3247) );
  NOR2_X1 U4003 ( .A1(n3247), .A2(n4222), .ZN(n3213) );
  AOI211_X1 U4004 ( .C1(n3244), .C2(n4188), .A(n3214), .B(n3213), .ZN(n3215)
         );
  INV_X1 U4005 ( .A(n3215), .ZN(U3281) );
  NAND2_X1 U4006 ( .A1(n3918), .A2(n3923), .ZN(n3223) );
  INV_X1 U4007 ( .A(n3223), .ZN(n3859) );
  XNOR2_X1 U4008 ( .A(n3216), .B(n3859), .ZN(n3277) );
  INV_X1 U4009 ( .A(n3277), .ZN(n3226) );
  OAI21_X1 U4010 ( .B1(n3217), .B2(n3397), .A(n3289), .ZN(n3284) );
  INV_X1 U4011 ( .A(n3284), .ZN(n3221) );
  AOI22_X1 U4012 ( .A1(n4222), .A2(REG2_REG_10__SCAN_IN), .B1(n3680), .B2(
        n4539), .ZN(n3218) );
  OAI21_X1 U4013 ( .B1(n3708), .B2(n4193), .A(n3218), .ZN(n3220) );
  OAI22_X1 U4014 ( .A1(n3673), .A2(n4197), .B1(n4196), .B2(n3397), .ZN(n3219)
         );
  AOI211_X1 U4015 ( .C1(n3221), .C2(n4543), .A(n3220), .B(n3219), .ZN(n3225)
         );
  XNOR2_X1 U4016 ( .A(n3222), .B(n3223), .ZN(n3278) );
  NAND2_X1 U4017 ( .A1(n3278), .A2(n4188), .ZN(n3224) );
  OAI211_X1 U4018 ( .C1(n3226), .C2(n3298), .A(n3225), .B(n3224), .ZN(U3280)
         );
  NAND2_X1 U4019 ( .A1(n3307), .A2(n3604), .ZN(n3233) );
  NAND2_X1 U4020 ( .A1(n3594), .A2(n3231), .ZN(n3232) );
  NAND2_X1 U4021 ( .A1(n3233), .A2(n3232), .ZN(n3234) );
  XNOR2_X1 U4022 ( .A(n3234), .B(n2133), .ZN(n3256) );
  NOR2_X1 U4023 ( .A1(n3630), .A2(n3236), .ZN(n3235) );
  AOI21_X1 U4024 ( .B1(n3307), .B2(n2945), .A(n3235), .ZN(n3257) );
  XNOR2_X1 U4025 ( .A(n3256), .B(n3257), .ZN(n3259) );
  XNOR2_X1 U4026 ( .A(n3260), .B(n3259), .ZN(n3243) );
  OAI22_X1 U4027 ( .A1(n2934), .A2(n3236), .B1(n3327), .B2(n3795), .ZN(n3237)
         );
  AOI211_X1 U4028 ( .C1(n3744), .C2(n3239), .A(n3238), .B(n3237), .ZN(n3242)
         );
  NAND2_X1 U4029 ( .A1(n3746), .A2(n3240), .ZN(n3241) );
  OAI211_X1 U4030 ( .C1(n3243), .C2(n3800), .A(n3242), .B(n3241), .ZN(U3210)
         );
  INV_X1 U4031 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3250) );
  NAND2_X1 U4032 ( .A1(n3244), .A2(n4582), .ZN(n3249) );
  OR2_X1 U4033 ( .A1(n3327), .A2(n4348), .ZN(n3246) );
  AOI22_X1 U4034 ( .A1(n3399), .A2(n4344), .B1(n4342), .B2(n3322), .ZN(n3245)
         );
  AND2_X1 U4035 ( .A1(n3246), .A2(n3245), .ZN(n3248) );
  AND3_X1 U4036 ( .A1(n3249), .A2(n3248), .A3(n3247), .ZN(n3252) );
  MUX2_X1 U4037 ( .A(n3250), .B(n3252), .S(n4599), .Z(n3251) );
  OAI21_X1 U4038 ( .B1(n4338), .B2(n3255), .A(n3251), .ZN(U3527) );
  INV_X1 U4039 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3253) );
  MUX2_X1 U4040 ( .A(n3253), .B(n3252), .S(n4589), .Z(n3254) );
  OAI21_X1 U4041 ( .B1(n3255), .B2(n4406), .A(n3254), .ZN(U3485) );
  INV_X1 U4042 ( .A(n3256), .ZN(n3258) );
  OR2_X1 U40430 ( .A1(n3327), .A2(n3631), .ZN(n3262) );
  NAND2_X1 U4044 ( .A1(n3553), .A2(n3306), .ZN(n3261) );
  NAND2_X1 U4045 ( .A1(n3262), .A2(n3261), .ZN(n3265) );
  OAI22_X1 U4046 ( .A1(n3327), .A2(n3630), .B1(n3627), .B2(n3302), .ZN(n3263)
         );
  XNOR2_X1 U4047 ( .A(n3263), .B(n2133), .ZN(n3264) );
  NAND2_X1 U4048 ( .A1(n3265), .A2(n3264), .ZN(n3318) );
  INV_X1 U4049 ( .A(n3264), .ZN(n3267) );
  INV_X1 U4050 ( .A(n3265), .ZN(n3266) );
  NAND2_X1 U4051 ( .A1(n3267), .A2(n3266), .ZN(n3320) );
  NAND2_X1 U4052 ( .A1(n3318), .A2(n3320), .ZN(n3268) );
  XNOR2_X1 U4053 ( .A(n3319), .B(n3268), .ZN(n3273) );
  AOI22_X1 U4054 ( .A1(n3729), .A2(n3306), .B1(n3811), .B2(n3982), .ZN(n3269)
         );
  NAND2_X1 U4055 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n4432) );
  OAI211_X1 U4056 ( .C1(n3270), .C2(n3807), .A(n3269), .B(n4432), .ZN(n3271)
         );
  AOI21_X1 U4057 ( .B1(n4540), .B2(n3746), .A(n3271), .ZN(n3272) );
  OAI21_X1 U4058 ( .B1(n3273), .B2(n3800), .A(n3272), .ZN(U3218) );
  INV_X1 U4059 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4727) );
  NAND2_X1 U4060 ( .A1(n3982), .A2(n4303), .ZN(n3275) );
  NAND2_X1 U4061 ( .A1(n3670), .A2(n4344), .ZN(n3274) );
  OAI211_X1 U4062 ( .C1(n4273), .C2(n3397), .A(n3275), .B(n3274), .ZN(n3276)
         );
  AOI21_X1 U4063 ( .B1(n3277), .B2(n4254), .A(n3276), .ZN(n3280) );
  NAND2_X1 U4064 ( .A1(n3278), .A2(n4582), .ZN(n3279) );
  AND2_X1 U4065 ( .A1(n3280), .A2(n3279), .ZN(n3282) );
  MUX2_X1 U4066 ( .A(n4727), .B(n3282), .S(n4599), .Z(n3281) );
  OAI21_X1 U4067 ( .B1(n3284), .B2(n4338), .A(n3281), .ZN(U3528) );
  INV_X1 U4068 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4699) );
  MUX2_X1 U4069 ( .A(n4699), .B(n3282), .S(n4589), .Z(n3283) );
  OAI21_X1 U4070 ( .B1(n3284), .B2(n4406), .A(n3283), .ZN(U3487) );
  XNOR2_X1 U4071 ( .A(n3285), .B(n3854), .ZN(n3355) );
  OAI21_X1 U4072 ( .B1(n3287), .B2(n3854), .A(n3286), .ZN(n3349) );
  NAND2_X1 U4073 ( .A1(n3289), .A2(n3288), .ZN(n3290) );
  NAND2_X1 U4074 ( .A1(n3338), .A2(n3290), .ZN(n3376) );
  INV_X1 U4075 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4747) );
  OAI22_X1 U4076 ( .A1(n3413), .A2(n4239), .B1(n4747), .B2(n4421), .ZN(n3291)
         );
  AOI21_X1 U4077 ( .B1(n3292), .B2(n3981), .A(n3291), .ZN(n3295) );
  INV_X1 U4078 ( .A(n3399), .ZN(n3408) );
  OAI22_X1 U4079 ( .A1(n3408), .A2(n4197), .B1(n4196), .B2(n3409), .ZN(n3293)
         );
  INV_X1 U4080 ( .A(n3293), .ZN(n3294) );
  OAI211_X1 U4081 ( .C1(n3376), .C2(n4238), .A(n3295), .B(n3294), .ZN(n3296)
         );
  AOI21_X1 U4082 ( .B1(n3349), .B2(n4188), .A(n3296), .ZN(n3297) );
  OAI21_X1 U4083 ( .B1(n3355), .B2(n3298), .A(n3297), .ZN(U3279) );
  INV_X1 U4084 ( .A(n3299), .ZN(n3303) );
  INV_X1 U4085 ( .A(n3300), .ZN(n3301) );
  OAI21_X1 U4086 ( .B1(n3303), .B2(n3302), .A(n3301), .ZN(n4541) );
  INV_X1 U4087 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4867) );
  NAND2_X1 U4088 ( .A1(n3908), .A2(n3906), .ZN(n3856) );
  XNOR2_X1 U4089 ( .A(n3304), .B(n3856), .ZN(n3309) );
  INV_X1 U4090 ( .A(n3309), .ZN(n4545) );
  XNOR2_X1 U4091 ( .A(n3305), .B(n3856), .ZN(n3312) );
  AOI22_X1 U4092 ( .A1(n3307), .A2(n4303), .B1(n3306), .B2(n4342), .ZN(n3308)
         );
  OAI21_X1 U4093 ( .B1(n3673), .B2(n4307), .A(n3308), .ZN(n3311) );
  NOR2_X1 U4094 ( .A1(n3309), .A2(n4210), .ZN(n3310) );
  AOI211_X1 U4095 ( .C1(n4254), .C2(n3312), .A(n3311), .B(n3310), .ZN(n4548)
         );
  INV_X1 U4096 ( .A(n4548), .ZN(n3313) );
  AOI21_X1 U4097 ( .B1(n4579), .B2(n4545), .A(n3313), .ZN(n3315) );
  MUX2_X1 U4098 ( .A(n4867), .B(n3315), .S(n4599), .Z(n3314) );
  OAI21_X1 U4099 ( .B1(n4541), .B2(n4338), .A(n3314), .ZN(U3526) );
  INV_X1 U4100 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3316) );
  MUX2_X1 U4101 ( .A(n3316), .B(n3315), .S(n4589), .Z(n3317) );
  OAI21_X1 U4102 ( .B1(n4541), .B2(n4406), .A(n3317), .ZN(U3483) );
  NAND2_X1 U4103 ( .A1(n3321), .A2(n3320), .ZN(n3387) );
  NAND2_X1 U4104 ( .A1(n3982), .A2(n3553), .ZN(n3324) );
  NAND2_X1 U4105 ( .A1(n3594), .A2(n3322), .ZN(n3323) );
  NAND2_X1 U4106 ( .A1(n3324), .A2(n3323), .ZN(n3325) );
  XNOR2_X1 U4107 ( .A(n3325), .B(n2132), .ZN(n3389) );
  OAI22_X1 U4108 ( .A1(n3673), .A2(n3631), .B1(n3630), .B2(n3328), .ZN(n3388)
         );
  XOR2_X1 U4109 ( .A(n3389), .B(n3388), .Z(n3386) );
  XNOR2_X1 U4110 ( .A(n3387), .B(n3386), .ZN(n3326) );
  NAND2_X1 U4111 ( .A1(n3326), .A2(n3805), .ZN(n3331) );
  AND2_X1 U4112 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4451) );
  OAI22_X1 U4113 ( .A1(n2934), .A2(n3328), .B1(n3327), .B2(n3807), .ZN(n3329)
         );
  AOI211_X1 U4114 ( .C1(n3811), .C2(n3399), .A(n4451), .B(n3329), .ZN(n3330)
         );
  OAI211_X1 U4115 ( .C1(n3815), .C2(n3332), .A(n3331), .B(n3330), .ZN(U3228)
         );
  NAND2_X1 U4116 ( .A1(n3334), .A2(n3333), .ZN(n3361) );
  NAND2_X1 U4117 ( .A1(n3358), .A2(n3359), .ZN(n3852) );
  INV_X1 U4118 ( .A(n3852), .ZN(n3335) );
  XNOR2_X1 U4119 ( .A(n3361), .B(n3335), .ZN(n3336) );
  NAND2_X1 U4120 ( .A1(n3336), .A2(n4254), .ZN(n3378) );
  XNOR2_X1 U4121 ( .A(n3337), .B(n3852), .ZN(n3380) );
  NAND2_X1 U4122 ( .A1(n3380), .A2(n4188), .ZN(n3348) );
  AND2_X1 U4123 ( .A1(n3338), .A2(n3706), .ZN(n3339) );
  OR2_X1 U4124 ( .A1(n3339), .A2(n3367), .ZN(n3385) );
  INV_X1 U4125 ( .A(n3385), .ZN(n3346) );
  OAI22_X1 U4126 ( .A1(n3708), .A2(n4197), .B1(n4196), .B2(n3505), .ZN(n3344)
         );
  INV_X1 U4127 ( .A(n3980), .ZN(n3656) );
  NOR2_X1 U4128 ( .A1(n4193), .A2(n3656), .ZN(n3343) );
  INV_X1 U4129 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3341) );
  INV_X1 U4130 ( .A(n3710), .ZN(n3340) );
  OAI22_X1 U4131 ( .A1(n4421), .A2(n3341), .B1(n3340), .B2(n4239), .ZN(n3342)
         );
  OR3_X1 U4132 ( .A1(n3344), .A2(n3343), .A3(n3342), .ZN(n3345) );
  AOI21_X1 U4133 ( .B1(n3346), .B2(n4543), .A(n3345), .ZN(n3347) );
  OAI211_X1 U4134 ( .C1(n4222), .C2(n3378), .A(n3348), .B(n3347), .ZN(U3278)
         );
  NAND2_X1 U4135 ( .A1(n3349), .A2(n4582), .ZN(n3354) );
  NAND2_X1 U4136 ( .A1(n3399), .A2(n4303), .ZN(n3351) );
  NAND2_X1 U4137 ( .A1(n3981), .A2(n4344), .ZN(n3350) );
  OAI211_X1 U4138 ( .C1(n4273), .C2(n3409), .A(n3351), .B(n3350), .ZN(n3352)
         );
  INV_X1 U4139 ( .A(n3352), .ZN(n3353) );
  OAI211_X1 U4140 ( .C1(n4233), .C2(n3355), .A(n3354), .B(n3353), .ZN(n3373)
         );
  MUX2_X1 U4141 ( .A(n3373), .B(REG1_REG_11__SCAN_IN), .S(n4596), .Z(n3356) );
  INV_X1 U4142 ( .A(n3356), .ZN(n3357) );
  OAI21_X1 U4143 ( .B1(n4338), .B2(n3376), .A(n3357), .ZN(U3529) );
  INV_X1 U4144 ( .A(n3358), .ZN(n3360) );
  OAI21_X1 U4145 ( .B1(n3361), .B2(n3360), .A(n3359), .ZN(n3362) );
  XNOR2_X1 U4146 ( .A(n3980), .B(n3494), .ZN(n3875) );
  XNOR2_X1 U4147 ( .A(n3362), .B(n3875), .ZN(n3365) );
  OAI22_X1 U4148 ( .A1(n3808), .A2(n4307), .B1(n4273), .B2(n3617), .ZN(n3363)
         );
  AOI21_X1 U4149 ( .B1(n4303), .B2(n3981), .A(n3363), .ZN(n3364) );
  OAI21_X1 U4150 ( .B1(n3365), .B2(n4233), .A(n3364), .ZN(n3414) );
  INV_X1 U4151 ( .A(n3414), .ZN(n3372) );
  XOR2_X1 U4152 ( .A(n3875), .B(n3366), .Z(n3415) );
  NOR2_X1 U4153 ( .A1(n3367), .A2(n3617), .ZN(n3368) );
  OR2_X1 U4154 ( .A1(n3441), .A2(n3368), .ZN(n3421) );
  AOI22_X1 U4155 ( .A1(n4222), .A2(REG2_REG_13__SCAN_IN), .B1(n3619), .B2(
        n4539), .ZN(n3369) );
  OAI21_X1 U4156 ( .B1(n3421), .B2(n4238), .A(n3369), .ZN(n3370) );
  AOI21_X1 U4157 ( .B1(n3415), .B2(n4188), .A(n3370), .ZN(n3371) );
  OAI21_X1 U4158 ( .B1(n4222), .B2(n3372), .A(n3371), .ZN(U3277) );
  MUX2_X1 U4159 ( .A(REG0_REG_11__SCAN_IN), .B(n3373), .S(n4589), .Z(n3374) );
  INV_X1 U4160 ( .A(n3374), .ZN(n3375) );
  OAI21_X1 U4161 ( .B1(n3376), .B2(n4406), .A(n3375), .ZN(U3489) );
  INV_X1 U4162 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4700) );
  AOI22_X1 U4163 ( .A1(n3980), .A2(n4344), .B1(n4342), .B2(n3706), .ZN(n3377)
         );
  OAI211_X1 U4164 ( .C1(n3708), .C2(n4348), .A(n3378), .B(n3377), .ZN(n3379)
         );
  AOI21_X1 U4165 ( .B1(n4582), .B2(n3380), .A(n3379), .ZN(n3382) );
  MUX2_X1 U4166 ( .A(n4700), .B(n3382), .S(n4589), .Z(n3381) );
  OAI21_X1 U4167 ( .B1(n3385), .B2(n4406), .A(n3381), .ZN(U3491) );
  INV_X1 U4168 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3383) );
  MUX2_X1 U4169 ( .A(n3383), .B(n3382), .S(n4599), .Z(n3384) );
  OAI21_X1 U4170 ( .B1(n3385), .B2(n4338), .A(n3384), .ZN(U3530) );
  NAND2_X1 U4171 ( .A1(n3387), .A2(n3386), .ZN(n3393) );
  NAND2_X1 U4172 ( .A1(n3399), .A2(n3604), .ZN(n3395) );
  NAND2_X1 U4173 ( .A1(n3594), .A2(n3671), .ZN(n3394) );
  NAND2_X1 U4174 ( .A1(n3395), .A2(n3394), .ZN(n3396) );
  XNOR2_X1 U4175 ( .A(n3396), .B(n2132), .ZN(n3403) );
  NOR2_X1 U4176 ( .A1(n3397), .A2(n3630), .ZN(n3398) );
  AOI21_X1 U4177 ( .B1(n3399), .B2(n2945), .A(n3398), .ZN(n3401) );
  XOR2_X1 U4178 ( .A(n3403), .B(n3401), .Z(n3677) );
  INV_X1 U4179 ( .A(n3401), .ZN(n3402) );
  NAND2_X1 U4180 ( .A1(n3403), .A2(n3402), .ZN(n3404) );
  OAI22_X1 U4181 ( .A1(n3708), .A2(n3630), .B1(n3627), .B2(n3409), .ZN(n3405)
         );
  XNOR2_X1 U4182 ( .A(n3405), .B(n2132), .ZN(n3496) );
  OAI22_X1 U4183 ( .A1(n3708), .A2(n3631), .B1(n3630), .B2(n3409), .ZN(n3497)
         );
  XNOR2_X1 U4184 ( .A(n3496), .B(n3497), .ZN(n3406) );
  XNOR2_X1 U4185 ( .A(n3498), .B(n3406), .ZN(n3407) );
  NAND2_X1 U4186 ( .A1(n3407), .A2(n3805), .ZN(n3412) );
  INV_X1 U4187 ( .A(REG3_REG_11__SCAN_IN), .ZN(n4804) );
  NOR2_X1 U4188 ( .A1(STATE_REG_SCAN_IN), .A2(n4804), .ZN(n4472) );
  OAI22_X1 U4189 ( .A1(n2934), .A2(n3409), .B1(n3408), .B2(n3807), .ZN(n3410)
         );
  AOI211_X1 U4190 ( .C1(n3811), .C2(n3981), .A(n4472), .B(n3410), .ZN(n3411)
         );
  OAI211_X1 U4191 ( .C1(n3815), .C2(n3413), .A(n3412), .B(n3411), .ZN(U3233)
         );
  INV_X1 U4192 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3416) );
  AOI21_X1 U4193 ( .B1(n3415), .B2(n4582), .A(n3414), .ZN(n3418) );
  MUX2_X1 U4194 ( .A(n3416), .B(n3418), .S(n4599), .Z(n3417) );
  OAI21_X1 U4195 ( .B1(n4338), .B2(n3421), .A(n3417), .ZN(U3531) );
  INV_X1 U4196 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3419) );
  MUX2_X1 U4197 ( .A(n3419), .B(n3418), .S(n4589), .Z(n3420) );
  OAI21_X1 U4198 ( .B1(n3421), .B2(n4406), .A(n3420), .ZN(U3493) );
  XNOR2_X1 U4199 ( .A(n3422), .B(n3866), .ZN(n3465) );
  INV_X1 U4200 ( .A(n3465), .ZN(n3432) );
  NAND2_X1 U4201 ( .A1(n3435), .A2(n3817), .ZN(n3423) );
  XNOR2_X1 U4202 ( .A(n3423), .B(n3866), .ZN(n3426) );
  INV_X1 U4203 ( .A(n3977), .ZN(n4349) );
  OAI22_X1 U4204 ( .A1(n4349), .A2(n4307), .B1(n4273), .B2(n3809), .ZN(n3424)
         );
  AOI21_X1 U4205 ( .B1(n4303), .B2(n3979), .A(n3424), .ZN(n3425) );
  OAI21_X1 U4206 ( .B1(n3426), .B2(n4233), .A(n3425), .ZN(n3464) );
  NAND2_X1 U4207 ( .A1(n3440), .A2(n3520), .ZN(n3427) );
  NAND2_X1 U4208 ( .A1(n3457), .A2(n3427), .ZN(n3471) );
  AOI22_X1 U4209 ( .A1(n4222), .A2(REG2_REG_15__SCAN_IN), .B1(n3428), .B2(
        n4539), .ZN(n3429) );
  OAI21_X1 U4210 ( .B1(n3471), .B2(n4238), .A(n3429), .ZN(n3430) );
  AOI21_X1 U4211 ( .B1(n3464), .B2(n4421), .A(n3430), .ZN(n3431) );
  OAI21_X1 U4212 ( .B1(n3432), .B2(n4265), .A(n3431), .ZN(U3275) );
  OAI21_X1 U4213 ( .B1(n3434), .B2(n3437), .A(n3433), .ZN(n3475) );
  INV_X1 U4214 ( .A(n3475), .ZN(n3448) );
  INV_X1 U4215 ( .A(n3821), .ZN(n3438) );
  INV_X1 U4216 ( .A(n3435), .ZN(n3436) );
  AOI21_X1 U4217 ( .B1(n3438), .B2(n3437), .A(n3436), .ZN(n3439) );
  OAI22_X1 U4218 ( .A1(n3448), .A2(n4210), .B1(n4233), .B2(n3439), .ZN(n3473)
         );
  NAND2_X1 U4219 ( .A1(n3473), .A2(n4421), .ZN(n3447) );
  OAI21_X1 U4220 ( .B1(n3441), .B2(n3515), .A(n3440), .ZN(n3481) );
  INV_X1 U4221 ( .A(n3481), .ZN(n3445) );
  INV_X1 U4222 ( .A(n3978), .ZN(n3731) );
  AOI22_X1 U4223 ( .A1(n4222), .A2(REG2_REG_14__SCAN_IN), .B1(n3658), .B2(
        n4539), .ZN(n3442) );
  OAI21_X1 U4224 ( .B1(n3731), .B2(n4193), .A(n3442), .ZN(n3444) );
  OAI22_X1 U4225 ( .A1(n3656), .A2(n4197), .B1(n4196), .B2(n3515), .ZN(n3443)
         );
  AOI211_X1 U4226 ( .C1(n3445), .C2(n4543), .A(n3444), .B(n3443), .ZN(n3446)
         );
  OAI211_X1 U4227 ( .C1(n3448), .C2(n4219), .A(n3447), .B(n3446), .ZN(U3276)
         );
  OAI21_X1 U4228 ( .B1(n3450), .B2(n3451), .A(n3449), .ZN(n4359) );
  XNOR2_X1 U4229 ( .A(n3452), .B(n3451), .ZN(n3456) );
  NAND2_X1 U4230 ( .A1(n3728), .A2(n4342), .ZN(n3454) );
  NAND2_X1 U4231 ( .A1(n3978), .A2(n4303), .ZN(n3453) );
  OAI211_X1 U4232 ( .C1(n4250), .C2(n4307), .A(n3454), .B(n3453), .ZN(n3455)
         );
  AOI21_X1 U4233 ( .B1(n3456), .B2(n4254), .A(n3455), .ZN(n4357) );
  INV_X1 U4234 ( .A(n4357), .ZN(n3462) );
  INV_X1 U4235 ( .A(REG2_REG_16__SCAN_IN), .ZN(n3460) );
  NAND2_X1 U4236 ( .A1(n3457), .A2(n3728), .ZN(n4353) );
  NAND3_X1 U4237 ( .A1(n4355), .A2(n4543), .A3(n4353), .ZN(n3459) );
  NAND2_X1 U4238 ( .A1(n4539), .A2(n3733), .ZN(n3458) );
  OAI211_X1 U4239 ( .C1(n4421), .C2(n3460), .A(n3459), .B(n3458), .ZN(n3461)
         );
  AOI21_X1 U4240 ( .B1(n3462), .B2(n4421), .A(n3461), .ZN(n3463) );
  OAI21_X1 U4241 ( .B1(n4359), .B2(n4265), .A(n3463), .ZN(U3274) );
  AOI21_X1 U4242 ( .B1(n3465), .B2(n4582), .A(n3464), .ZN(n3469) );
  INV_X1 U4243 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3466) );
  MUX2_X1 U4244 ( .A(n3469), .B(n3466), .S(n4596), .Z(n3467) );
  OAI21_X1 U4245 ( .B1(n4338), .B2(n3471), .A(n3467), .ZN(U3533) );
  INV_X1 U4246 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3468) );
  MUX2_X1 U4247 ( .A(n3469), .B(n3468), .S(n4587), .Z(n3470) );
  OAI21_X1 U4248 ( .B1(n3471), .B2(n4406), .A(n3470), .ZN(U3497) );
  INV_X1 U4249 ( .A(REG1_REG_14__SCAN_IN), .ZN(n3476) );
  INV_X1 U4250 ( .A(n3515), .ZN(n3654) );
  AOI22_X1 U4251 ( .A1(n3978), .A2(n4344), .B1(n4342), .B2(n3654), .ZN(n3472)
         );
  OAI21_X1 U4252 ( .B1(n3656), .B2(n4348), .A(n3472), .ZN(n3474) );
  AOI211_X1 U4253 ( .C1(n4579), .C2(n3475), .A(n3474), .B(n3473), .ZN(n3478)
         );
  MUX2_X1 U4254 ( .A(n3476), .B(n3478), .S(n4599), .Z(n3477) );
  OAI21_X1 U4255 ( .B1(n4338), .B2(n3481), .A(n3477), .ZN(U3532) );
  INV_X1 U4256 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3479) );
  MUX2_X1 U4257 ( .A(n3479), .B(n3478), .S(n4589), .Z(n3480) );
  OAI21_X1 U4258 ( .B1(n3481), .B2(n4406), .A(n3480), .ZN(U3495) );
  AND2_X1 U4259 ( .A1(n2166), .A2(n4224), .ZN(n3865) );
  INV_X1 U4260 ( .A(n3865), .ZN(n3482) );
  XNOR2_X1 U4261 ( .A(n3483), .B(n3482), .ZN(n3484) );
  NAND2_X1 U4262 ( .A1(n3484), .A2(n4254), .ZN(n4347) );
  XNOR2_X1 U4263 ( .A(n3485), .B(n3865), .ZN(n4351) );
  NAND2_X1 U4264 ( .A1(n4351), .A2(n4188), .ZN(n3493) );
  INV_X1 U4265 ( .A(n4355), .ZN(n3487) );
  INV_X1 U4266 ( .A(n4258), .ZN(n3486) );
  OAI21_X1 U4267 ( .B1(n3487), .B2(n3742), .A(n3486), .ZN(n4407) );
  INV_X1 U4268 ( .A(n4407), .ZN(n3491) );
  AOI22_X1 U4269 ( .A1(n4222), .A2(REG2_REG_17__SCAN_IN), .B1(n3745), .B2(
        n4539), .ZN(n3488) );
  OAI21_X1 U4270 ( .B1(n3741), .B2(n4193), .A(n3488), .ZN(n3490) );
  OAI22_X1 U4271 ( .A1(n4349), .A2(n4197), .B1(n4196), .B2(n3742), .ZN(n3489)
         );
  AOI211_X1 U4272 ( .C1(n3491), .C2(n4543), .A(n3490), .B(n3489), .ZN(n3492)
         );
  OAI211_X1 U4273 ( .C1(n4222), .C2(n4347), .A(n3493), .B(n3492), .ZN(U3273)
         );
  AOI22_X1 U4274 ( .A1(n3980), .A2(n3553), .B1(n3594), .B2(n3494), .ZN(n3495)
         );
  XOR2_X1 U4275 ( .A(n2133), .B(n3495), .Z(n3511) );
  INV_X1 U4276 ( .A(n3498), .ZN(n3501) );
  INV_X1 U4277 ( .A(n3497), .ZN(n3500) );
  OAI21_X1 U4278 ( .B1(n3501), .B2(n3500), .A(n3499), .ZN(n3705) );
  INV_X1 U4279 ( .A(n3705), .ZN(n3510) );
  NAND2_X1 U4280 ( .A1(n3981), .A2(n3553), .ZN(n3503) );
  NAND2_X1 U4281 ( .A1(n3594), .A2(n3706), .ZN(n3502) );
  NAND2_X1 U4282 ( .A1(n3503), .A2(n3502), .ZN(n3504) );
  XNOR2_X1 U4283 ( .A(n3504), .B(n2952), .ZN(n3508) );
  NOR2_X1 U4284 ( .A1(n3505), .A2(n3630), .ZN(n3506) );
  AOI21_X1 U4285 ( .B1(n3981), .B2(n2945), .A(n3506), .ZN(n3507) );
  NOR2_X1 U4286 ( .A1(n3508), .A2(n3507), .ZN(n3703) );
  OAI22_X1 U4287 ( .A1(n3656), .A2(n3631), .B1(n3630), .B2(n3617), .ZN(n3613)
         );
  NAND2_X1 U4288 ( .A1(n3979), .A2(n3553), .ZN(n3513) );
  NAND2_X1 U4289 ( .A1(n3594), .A2(n3654), .ZN(n3512) );
  NAND2_X1 U4290 ( .A1(n3513), .A2(n3512), .ZN(n3514) );
  XNOR2_X1 U4291 ( .A(n3514), .B(n2952), .ZN(n3518) );
  NOR2_X1 U4292 ( .A1(n3630), .A2(n3515), .ZN(n3516) );
  AOI21_X1 U4293 ( .B1(n3979), .B2(n2945), .A(n3516), .ZN(n3517) );
  NOR2_X1 U4294 ( .A1(n3518), .A2(n3517), .ZN(n3651) );
  AOI22_X1 U4295 ( .A1(n3978), .A2(n3553), .B1(n3594), .B2(n3520), .ZN(n3519)
         );
  XNOR2_X1 U4296 ( .A(n3519), .B(n2132), .ZN(n3530) );
  NAND2_X1 U4297 ( .A1(n3531), .A2(n3530), .ZN(n3724) );
  NAND2_X1 U4298 ( .A1(n3978), .A2(n2945), .ZN(n3522) );
  NAND2_X1 U4299 ( .A1(n3553), .A2(n3520), .ZN(n3521) );
  NAND2_X1 U4300 ( .A1(n3522), .A2(n3521), .ZN(n3803) );
  NAND2_X1 U4301 ( .A1(n3724), .A2(n3803), .ZN(n3532) );
  NAND2_X1 U4302 ( .A1(n3977), .A2(n3553), .ZN(n3524) );
  NAND2_X1 U4303 ( .A1(n3594), .A2(n3728), .ZN(n3523) );
  NAND2_X1 U4304 ( .A1(n3524), .A2(n3523), .ZN(n3525) );
  XNOR2_X1 U4305 ( .A(n3525), .B(n2133), .ZN(n3529) );
  NAND2_X1 U4306 ( .A1(n3977), .A2(n2945), .ZN(n3527) );
  NAND2_X1 U4307 ( .A1(n3553), .A2(n3728), .ZN(n3526) );
  NAND2_X1 U4308 ( .A1(n3527), .A2(n3526), .ZN(n3528) );
  NOR2_X1 U4309 ( .A1(n3529), .A2(n3528), .ZN(n3533) );
  OR2_X2 U4310 ( .A1(n3531), .A2(n3530), .ZN(n3802) );
  NAND3_X1 U4311 ( .A1(n3532), .A2(n3727), .A3(n3802), .ZN(n3535) );
  INV_X1 U4312 ( .A(n3533), .ZN(n3534) );
  NAND2_X1 U4313 ( .A1(n3535), .A2(n3534), .ZN(n3740) );
  OAI22_X1 U4314 ( .A1(n4250), .A2(n3630), .B1(n3627), .B2(n3742), .ZN(n3536)
         );
  XNOR2_X1 U4315 ( .A(n3536), .B(n2133), .ZN(n3540) );
  OR2_X1 U4316 ( .A1(n4250), .A2(n3631), .ZN(n3538) );
  NAND2_X1 U4317 ( .A1(n3553), .A2(n4343), .ZN(n3537) );
  NAND2_X1 U4318 ( .A1(n3538), .A2(n3537), .ZN(n3539) );
  NAND2_X1 U4319 ( .A1(n3540), .A2(n3539), .ZN(n3737) );
  NOR2_X1 U4320 ( .A1(n3540), .A2(n3539), .ZN(n3736) );
  OAI22_X1 U4321 ( .A1(n3741), .A2(n3631), .B1(n3630), .B2(n4257), .ZN(n3781)
         );
  OAI22_X1 U4322 ( .A1(n3741), .A2(n3630), .B1(n3627), .B2(n4257), .ZN(n3541)
         );
  XNOR2_X1 U4323 ( .A(n3541), .B(n2132), .ZN(n3780) );
  NAND2_X1 U4324 ( .A1(n3975), .A2(n3553), .ZN(n3543) );
  NAND2_X1 U4325 ( .A1(n3594), .A2(n3686), .ZN(n3542) );
  NAND2_X1 U4326 ( .A1(n3543), .A2(n3542), .ZN(n3544) );
  XNOR2_X1 U4327 ( .A(n3544), .B(n2952), .ZN(n3547) );
  NOR2_X1 U4328 ( .A1(n4236), .A2(n3630), .ZN(n3545) );
  AOI21_X1 U4329 ( .B1(n3975), .B2(n2945), .A(n3545), .ZN(n3546) );
  NAND2_X1 U4330 ( .A1(n3547), .A2(n3546), .ZN(n3549) );
  OAI21_X1 U4331 ( .B1(n3547), .B2(n3546), .A(n3549), .ZN(n3685) );
  NAND2_X1 U4332 ( .A1(n3683), .A2(n3549), .ZN(n3693) );
  NAND2_X1 U4333 ( .A1(n3974), .A2(n3553), .ZN(n3551) );
  NAND2_X1 U4334 ( .A1(n3594), .A2(n4216), .ZN(n3550) );
  NAND2_X1 U4335 ( .A1(n3551), .A2(n3550), .ZN(n3552) );
  XNOR2_X1 U4336 ( .A(n3552), .B(n2133), .ZN(n3556) );
  NAND2_X1 U4337 ( .A1(n3974), .A2(n2945), .ZN(n3555) );
  NAND2_X1 U4338 ( .A1(n3553), .A2(n4216), .ZN(n3554) );
  NAND2_X1 U4339 ( .A1(n3555), .A2(n3554), .ZN(n3557) );
  NAND2_X1 U4340 ( .A1(n3556), .A2(n3557), .ZN(n3761) );
  NAND2_X1 U4341 ( .A1(n3693), .A2(n3761), .ZN(n3760) );
  INV_X1 U4342 ( .A(n3556), .ZN(n3559) );
  INV_X1 U4343 ( .A(n3557), .ZN(n3558) );
  NAND2_X1 U4344 ( .A1(n3559), .A2(n3558), .ZN(n3763) );
  NAND2_X1 U4345 ( .A1(n3760), .A2(n3763), .ZN(n3697) );
  NAND2_X1 U4346 ( .A1(n4206), .A2(n3553), .ZN(n3561) );
  NAND2_X1 U4347 ( .A1(n3594), .A2(n4321), .ZN(n3560) );
  NAND2_X1 U4348 ( .A1(n3561), .A2(n3560), .ZN(n3562) );
  XNOR2_X1 U4349 ( .A(n3562), .B(n2952), .ZN(n3564) );
  NOR2_X1 U4350 ( .A1(n3630), .A2(n4195), .ZN(n3563) );
  AOI21_X1 U4351 ( .B1(n4206), .B2(n2945), .A(n3563), .ZN(n3565) );
  INV_X1 U4352 ( .A(n3564), .ZN(n3567) );
  INV_X1 U4353 ( .A(n3565), .ZN(n3566) );
  NAND2_X1 U4354 ( .A1(n3567), .A2(n3566), .ZN(n3692) );
  OAI22_X1 U4355 ( .A1(n4194), .A2(n3630), .B1(n3627), .B2(n4177), .ZN(n3568)
         );
  XNOR2_X1 U4356 ( .A(n3568), .B(n2132), .ZN(n3570) );
  OAI22_X1 U4357 ( .A1(n4194), .A2(n3631), .B1(n3630), .B2(n4177), .ZN(n3569)
         );
  XNOR2_X1 U4358 ( .A(n3570), .B(n3569), .ZN(n3773) );
  NOR2_X1 U4359 ( .A1(n3570), .A2(n3569), .ZN(n3663) );
  NAND2_X1 U4360 ( .A1(n4304), .A2(n3553), .ZN(n3572) );
  NAND2_X1 U4361 ( .A1(n3594), .A2(n4155), .ZN(n3571) );
  NAND2_X1 U4362 ( .A1(n3572), .A2(n3571), .ZN(n3573) );
  XNOR2_X1 U4363 ( .A(n3573), .B(n2952), .ZN(n3576) );
  NOR2_X1 U4364 ( .A1(n3630), .A2(n4160), .ZN(n3574) );
  AOI21_X1 U4365 ( .B1(n4304), .B2(n2945), .A(n3574), .ZN(n3577) );
  XNOR2_X1 U4366 ( .A(n3576), .B(n3577), .ZN(n3662) );
  NOR2_X1 U4367 ( .A1(n3663), .A2(n3662), .ZN(n3575) );
  INV_X1 U4368 ( .A(n3576), .ZN(n3579) );
  INV_X1 U4369 ( .A(n3577), .ZN(n3578) );
  NAND2_X1 U4370 ( .A1(n3579), .A2(n3578), .ZN(n3583) );
  NOR2_X1 U4371 ( .A1(n3630), .A2(n4140), .ZN(n3580) );
  AOI21_X1 U4372 ( .B1(n4116), .B2(n2945), .A(n3580), .ZN(n3584) );
  OAI22_X1 U4373 ( .A1(n4158), .A2(n3630), .B1(n3627), .B2(n4140), .ZN(n3582)
         );
  XNOR2_X1 U4374 ( .A(n3582), .B(n2133), .ZN(n3753) );
  NAND2_X1 U4375 ( .A1(n3750), .A2(n3753), .ZN(n3587) );
  INV_X1 U4376 ( .A(n3584), .ZN(n3585) );
  NAND2_X1 U4377 ( .A1(n3586), .A2(n3585), .ZN(n3751) );
  NAND2_X1 U4378 ( .A1(n3587), .A2(n3751), .ZN(n3717) );
  NAND2_X1 U4379 ( .A1(n4101), .A2(n3553), .ZN(n3589) );
  NAND2_X1 U4380 ( .A1(n3594), .A2(n4115), .ZN(n3588) );
  NAND2_X1 U4381 ( .A1(n3589), .A2(n3588), .ZN(n3590) );
  XNOR2_X1 U4382 ( .A(n3590), .B(n2952), .ZN(n3593) );
  NOR2_X1 U4383 ( .A1(n3630), .A2(n4122), .ZN(n3591) );
  AOI21_X1 U4384 ( .B1(n4101), .B2(n2945), .A(n3591), .ZN(n3592) );
  NAND2_X1 U4385 ( .A1(n3593), .A2(n3592), .ZN(n3713) );
  NOR2_X1 U4386 ( .A1(n3593), .A2(n3592), .ZN(n3715) );
  NAND2_X1 U4387 ( .A1(n4287), .A2(n3553), .ZN(n3596) );
  NAND2_X1 U4388 ( .A1(n3594), .A2(n4100), .ZN(n3595) );
  NAND2_X1 U4389 ( .A1(n3596), .A2(n3595), .ZN(n3597) );
  XNOR2_X1 U4390 ( .A(n3597), .B(n2952), .ZN(n3602) );
  INV_X1 U4391 ( .A(n3602), .ZN(n3600) );
  NOR2_X1 U4392 ( .A1(n3630), .A2(n4105), .ZN(n3598) );
  AOI21_X1 U4393 ( .B1(n4287), .B2(n2945), .A(n3598), .ZN(n3601) );
  INV_X1 U4394 ( .A(n3601), .ZN(n3599) );
  NAND2_X1 U4395 ( .A1(n3600), .A2(n3599), .ZN(n3790) );
  AND2_X1 U4396 ( .A1(n3602), .A2(n3601), .ZN(n3789) );
  OAI22_X1 U4397 ( .A1(n4281), .A2(n3630), .B1(n3627), .B2(n2643), .ZN(n3603)
         );
  XNOR2_X1 U4398 ( .A(n3603), .B(n2952), .ZN(n3636) );
  OR2_X1 U4399 ( .A1(n4281), .A2(n3631), .ZN(n3606) );
  NAND2_X1 U4400 ( .A1(n3553), .A2(n4286), .ZN(n3605) );
  NAND2_X1 U4401 ( .A1(n3606), .A2(n3605), .ZN(n3634) );
  XNOR2_X1 U4402 ( .A(n3636), .B(n3634), .ZN(n3625) );
  XNOR2_X1 U4403 ( .A(n3626), .B(n3625), .ZN(n3611) );
  OAI22_X1 U4404 ( .A1(n2934), .A2(n2643), .B1(n4119), .B2(n3807), .ZN(n3609)
         );
  OAI22_X1 U4405 ( .A1(n4290), .A2(n3795), .B1(STATE_REG_SCAN_IN), .B2(n3607), 
        .ZN(n3608) );
  AOI211_X1 U4406 ( .C1(n4088), .C2(n3798), .A(n3609), .B(n3608), .ZN(n3610)
         );
  OAI21_X1 U4407 ( .B1(n3611), .B2(n3800), .A(n3610), .ZN(U3211) );
  XNOR2_X1 U4408 ( .A(n2300), .B(n3613), .ZN(n3614) );
  XNOR2_X1 U4409 ( .A(n3612), .B(n3614), .ZN(n3622) );
  NOR2_X1 U4410 ( .A1(STATE_REG_SCAN_IN), .A2(n3615), .ZN(n4487) );
  INV_X1 U4411 ( .A(n3981), .ZN(n3616) );
  OAI22_X1 U4412 ( .A1(n2934), .A2(n3617), .B1(n3616), .B2(n3807), .ZN(n3618)
         );
  AOI211_X1 U4413 ( .C1(n3811), .C2(n3979), .A(n4487), .B(n3618), .ZN(n3621)
         );
  NAND2_X1 U4414 ( .A1(n3746), .A2(n3619), .ZN(n3620) );
  OAI211_X1 U4415 ( .C1(n3622), .C2(n3800), .A(n3621), .B(n3620), .ZN(U3231)
         );
  NAND2_X1 U4416 ( .A1(U3149), .A2(DATAI_25_), .ZN(n3623) );
  OAI21_X1 U4417 ( .B1(n3624), .B2(U3149), .A(n3623), .ZN(U3327) );
  NAND2_X1 U4418 ( .A1(n3626), .A2(n3625), .ZN(n3650) );
  OAI22_X1 U4419 ( .A1(n4290), .A2(n3630), .B1(n3627), .B2(n4077), .ZN(n3629)
         );
  XNOR2_X1 U4420 ( .A(n3629), .B(n2132), .ZN(n3633) );
  OAI22_X1 U4421 ( .A1(n4290), .A2(n3631), .B1(n3630), .B2(n4077), .ZN(n3632)
         );
  XNOR2_X1 U4422 ( .A(n3633), .B(n3632), .ZN(n3638) );
  NAND2_X1 U4423 ( .A1(n3638), .A2(n3805), .ZN(n3649) );
  INV_X1 U4424 ( .A(n3634), .ZN(n3635) );
  NOR2_X1 U4425 ( .A1(n3636), .A2(n3635), .ZN(n3639) );
  NOR3_X1 U4426 ( .A1(n3638), .A2(n3639), .A3(n3800), .ZN(n3637) );
  NAND2_X1 U4427 ( .A1(n3650), .A2(n3637), .ZN(n3648) );
  INV_X1 U4428 ( .A(n3638), .ZN(n3641) );
  INV_X1 U4429 ( .A(n3639), .ZN(n3640) );
  NOR3_X1 U4430 ( .A1(n3641), .A2(n3640), .A3(n3800), .ZN(n3646) );
  AOI22_X1 U4431 ( .A1(n4278), .A2(n3811), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3644) );
  AOI22_X1 U4432 ( .A1(n3642), .A2(n3744), .B1(n3729), .B2(n4277), .ZN(n3643)
         );
  OAI211_X1 U4433 ( .C1(n3815), .C2(n4073), .A(n3644), .B(n3643), .ZN(n3645)
         );
  NOR2_X1 U4434 ( .A1(n3646), .A2(n3645), .ZN(n3647) );
  OAI211_X1 U4435 ( .C1(n3650), .C2(n3649), .A(n3648), .B(n3647), .ZN(U3217)
         );
  NOR2_X1 U4436 ( .A1(n3651), .A2(n2169), .ZN(n3652) );
  XNOR2_X1 U4437 ( .A(n3653), .B(n3652), .ZN(n3660) );
  AOI22_X1 U4438 ( .A1(n3729), .A2(n3654), .B1(n3811), .B2(n3978), .ZN(n3655)
         );
  NAND2_X1 U4439 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4494) );
  OAI211_X1 U4440 ( .C1(n3656), .C2(n3807), .A(n3655), .B(n4494), .ZN(n3657)
         );
  AOI21_X1 U4441 ( .B1(n3658), .B2(n3746), .A(n3657), .ZN(n3659) );
  OAI21_X1 U4442 ( .B1(n3660), .B2(n3800), .A(n3659), .ZN(U3212) );
  INV_X1 U4443 ( .A(n3661), .ZN(n3771) );
  OAI21_X1 U4444 ( .B1(n3771), .B2(n3663), .A(n3662), .ZN(n3665) );
  NAND3_X1 U4445 ( .A1(n3665), .A2(n3805), .A3(n3664), .ZN(n3669) );
  NOR2_X1 U4446 ( .A1(n4158), .A2(n3795), .ZN(n3667) );
  OAI22_X1 U4447 ( .A1(n2934), .A2(n4160), .B1(n4194), .B2(n3807), .ZN(n3666)
         );
  AOI211_X1 U4448 ( .C1(REG3_REG_23__SCAN_IN), .C2(U3149), .A(n3667), .B(n3666), .ZN(n3668) );
  OAI211_X1 U4449 ( .C1(n3815), .C2(n4162), .A(n3669), .B(n3668), .ZN(U3213)
         );
  AOI22_X1 U4450 ( .A1(n3729), .A2(n3671), .B1(n3811), .B2(n3670), .ZN(n3672)
         );
  NAND2_X1 U4451 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4455) );
  OAI211_X1 U4452 ( .C1(n3673), .C2(n3807), .A(n3672), .B(n4455), .ZN(n3679)
         );
  INV_X1 U4453 ( .A(n3675), .ZN(n3676) );
  AOI211_X1 U4454 ( .C1(n3677), .C2(n3674), .A(n3800), .B(n3676), .ZN(n3678)
         );
  AOI211_X1 U4455 ( .C1(n3680), .C2(n3746), .A(n3679), .B(n3678), .ZN(n3681)
         );
  INV_X1 U4456 ( .A(n3681), .ZN(U3214) );
  INV_X1 U4457 ( .A(n3683), .ZN(n3684) );
  AOI21_X1 U4458 ( .B1(n3685), .B2(n3682), .A(n3684), .ZN(n3691) );
  AOI22_X1 U4459 ( .A1(n3729), .A2(n3686), .B1(n3744), .B2(n4345), .ZN(n3687)
         );
  NAND2_X1 U4460 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4049) );
  OAI211_X1 U4461 ( .C1(n4325), .C2(n3795), .A(n3687), .B(n4049), .ZN(n3688)
         );
  AOI21_X1 U4462 ( .B1(n3689), .B2(n3746), .A(n3688), .ZN(n3690) );
  OAI21_X1 U4463 ( .B1(n3691), .B2(n3800), .A(n3690), .ZN(U3216) );
  NAND2_X1 U4464 ( .A1(n2167), .A2(n3692), .ZN(n3696) );
  INV_X1 U4465 ( .A(n3763), .ZN(n3694) );
  OAI211_X1 U4466 ( .C1(n3693), .C2(n3694), .A(n3761), .B(n3696), .ZN(n3695)
         );
  OAI211_X1 U4467 ( .C1(n3697), .C2(n3696), .A(n3805), .B(n3695), .ZN(n3702)
         );
  OAI22_X1 U4468 ( .A1(n3795), .A2(n4194), .B1(STATE_REG_SCAN_IN), .B2(n3698), 
        .ZN(n3700) );
  OAI22_X1 U4469 ( .A1(n2934), .A2(n4195), .B1(n4325), .B2(n3807), .ZN(n3699)
         );
  AOI211_X1 U4470 ( .C1(n4191), .C2(n3798), .A(n3700), .B(n3699), .ZN(n3701)
         );
  NAND2_X1 U4471 ( .A1(n3702), .A2(n3701), .ZN(U3220) );
  NOR2_X1 U4472 ( .A1(n3703), .A2(n2362), .ZN(n3704) );
  XNOR2_X1 U4473 ( .A(n3705), .B(n3704), .ZN(n3712) );
  AOI22_X1 U4474 ( .A1(n3729), .A2(n3706), .B1(n3811), .B2(n3980), .ZN(n3707)
         );
  NAND2_X1 U4475 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4476) );
  OAI211_X1 U4476 ( .C1(n3708), .C2(n3807), .A(n3707), .B(n4476), .ZN(n3709)
         );
  AOI21_X1 U4477 ( .B1(n3710), .B2(n3746), .A(n3709), .ZN(n3711) );
  OAI21_X1 U4478 ( .B1(n3712), .B2(n3800), .A(n3711), .ZN(U3221) );
  INV_X1 U4479 ( .A(n3713), .ZN(n3714) );
  NOR2_X1 U4480 ( .A1(n3715), .A2(n3714), .ZN(n3716) );
  XNOR2_X1 U4481 ( .A(n3717), .B(n3716), .ZN(n3723) );
  INV_X1 U4482 ( .A(n3718), .ZN(n4123) );
  OAI22_X1 U4483 ( .A1(n4119), .A2(n3795), .B1(STATE_REG_SCAN_IN), .B2(n3719), 
        .ZN(n3721) );
  OAI22_X1 U4484 ( .A1(n2934), .A2(n4122), .B1(n4158), .B2(n3807), .ZN(n3720)
         );
  AOI211_X1 U4485 ( .C1(n4123), .C2(n3798), .A(n3721), .B(n3720), .ZN(n3722)
         );
  OAI21_X1 U4486 ( .B1(n3723), .B2(n3800), .A(n3722), .ZN(U3222) );
  INV_X1 U4487 ( .A(n3802), .ZN(n3725) );
  OAI21_X1 U4488 ( .B1(n3725), .B2(n3803), .A(n3724), .ZN(n3726) );
  XOR2_X1 U4489 ( .A(n3727), .B(n3726), .Z(n3735) );
  AOI22_X1 U4490 ( .A1(n3729), .A2(n3728), .B1(n3811), .B2(n3976), .ZN(n3730)
         );
  NAND2_X1 U4491 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4523) );
  OAI211_X1 U4492 ( .C1(n3731), .C2(n3807), .A(n3730), .B(n4523), .ZN(n3732)
         );
  AOI21_X1 U4493 ( .B1(n3733), .B2(n3746), .A(n3732), .ZN(n3734) );
  OAI21_X1 U4494 ( .B1(n3735), .B2(n3800), .A(n3734), .ZN(U3223) );
  INV_X1 U4495 ( .A(n3736), .ZN(n3738) );
  NAND2_X1 U4496 ( .A1(n3738), .A2(n3737), .ZN(n3739) );
  XNOR2_X1 U4497 ( .A(n3740), .B(n3739), .ZN(n3749) );
  AND2_X1 U4498 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4031) );
  OAI22_X1 U4499 ( .A1(n2934), .A2(n3742), .B1(n3741), .B2(n3795), .ZN(n3743)
         );
  AOI211_X1 U4500 ( .C1(n3744), .C2(n3977), .A(n4031), .B(n3743), .ZN(n3748)
         );
  NAND2_X1 U4501 ( .A1(n3746), .A2(n3745), .ZN(n3747) );
  OAI211_X1 U4502 ( .C1(n3749), .C2(n3800), .A(n3748), .B(n3747), .ZN(U3225)
         );
  NAND2_X1 U4503 ( .A1(n3751), .A2(n3750), .ZN(n3752) );
  XOR2_X1 U4504 ( .A(n3753), .B(n3752), .Z(n3759) );
  INV_X1 U4505 ( .A(n3754), .ZN(n4138) );
  OAI22_X1 U4506 ( .A1(n4308), .A2(n3795), .B1(STATE_REG_SCAN_IN), .B2(n3755), 
        .ZN(n3757) );
  OAI22_X1 U4507 ( .A1(n2934), .A2(n4140), .B1(n4172), .B2(n3807), .ZN(n3756)
         );
  AOI211_X1 U4508 ( .C1(n4138), .C2(n3798), .A(n3757), .B(n3756), .ZN(n3758)
         );
  OAI21_X1 U4509 ( .B1(n3759), .B2(n3800), .A(n3758), .ZN(U3226) );
  INV_X1 U4510 ( .A(n3760), .ZN(n3764) );
  AOI21_X1 U4511 ( .B1(n3761), .B2(n3763), .A(n3693), .ZN(n3762) );
  AOI21_X1 U4512 ( .B1(n3764), .B2(n3763), .A(n3762), .ZN(n3770) );
  INV_X1 U4513 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3765) );
  OAI22_X1 U4514 ( .A1(n3795), .A2(n3774), .B1(STATE_REG_SCAN_IN), .B2(n3765), 
        .ZN(n3768) );
  INV_X1 U4515 ( .A(n3975), .ZN(n4251) );
  OAI22_X1 U4516 ( .A1(n2934), .A2(n3766), .B1(n4251), .B2(n3807), .ZN(n3767)
         );
  AOI211_X1 U4517 ( .C1(n4214), .C2(n3798), .A(n3768), .B(n3767), .ZN(n3769)
         );
  OAI21_X1 U4518 ( .B1(n3770), .B2(n3800), .A(n3769), .ZN(U3230) );
  AOI21_X1 U4519 ( .B1(n3773), .B2(n3772), .A(n3771), .ZN(n3779) );
  INV_X1 U4520 ( .A(n4178), .ZN(n3777) );
  OAI22_X1 U4521 ( .A1(n3795), .A2(n4172), .B1(STATE_REG_SCAN_IN), .B2(n4805), 
        .ZN(n3776) );
  OAI22_X1 U4522 ( .A1(n2934), .A2(n4177), .B1(n3774), .B2(n3807), .ZN(n3775)
         );
  AOI211_X1 U4523 ( .C1(n3777), .C2(n3798), .A(n3776), .B(n3775), .ZN(n3778)
         );
  OAI21_X1 U4524 ( .B1(n3779), .B2(n3800), .A(n3778), .ZN(U3232) );
  XOR2_X1 U4525 ( .A(n3781), .B(n3780), .Z(n3782) );
  XNOR2_X1 U4526 ( .A(n3783), .B(n3782), .ZN(n3787) );
  NAND2_X1 U4527 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4526) );
  OAI21_X1 U4528 ( .B1(n3795), .B2(n4251), .A(n4526), .ZN(n3785) );
  OAI22_X1 U4529 ( .A1(n2934), .A2(n4257), .B1(n4250), .B2(n3807), .ZN(n3784)
         );
  AOI211_X1 U4530 ( .C1(n4259), .C2(n3798), .A(n3785), .B(n3784), .ZN(n3786)
         );
  OAI21_X1 U4531 ( .B1(n3787), .B2(n3800), .A(n3786), .ZN(U3235) );
  INV_X1 U4532 ( .A(n3789), .ZN(n3791) );
  NAND2_X1 U4533 ( .A1(n3791), .A2(n3790), .ZN(n3792) );
  XNOR2_X1 U4534 ( .A(n3788), .B(n3792), .ZN(n3801) );
  INV_X1 U4535 ( .A(n3793), .ZN(n4106) );
  OAI22_X1 U4536 ( .A1(n2934), .A2(n4105), .B1(n4308), .B2(n3807), .ZN(n3797)
         );
  INV_X1 U4537 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3794) );
  OAI22_X1 U4538 ( .A1(n4281), .A2(n3795), .B1(STATE_REG_SCAN_IN), .B2(n3794), 
        .ZN(n3796) );
  AOI211_X1 U4539 ( .C1(n4106), .C2(n3798), .A(n3797), .B(n3796), .ZN(n3799)
         );
  OAI21_X1 U4540 ( .B1(n3801), .B2(n3800), .A(n3799), .ZN(U3237) );
  NAND2_X1 U4541 ( .A1(n3802), .A2(n3724), .ZN(n3804) );
  XNOR2_X1 U4542 ( .A(n3804), .B(n3803), .ZN(n3806) );
  NAND2_X1 U4543 ( .A1(n3806), .A2(n3805), .ZN(n3813) );
  AND2_X1 U4544 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4508) );
  OAI22_X1 U4545 ( .A1(n2934), .A2(n3809), .B1(n3808), .B2(n3807), .ZN(n3810)
         );
  AOI211_X1 U4546 ( .C1(n3811), .C2(n3977), .A(n4508), .B(n3810), .ZN(n3812)
         );
  OAI211_X1 U4547 ( .C1(n3815), .C2(n3814), .A(n3813), .B(n3812), .ZN(U3238)
         );
  INV_X1 U4548 ( .A(n3816), .ZN(n3884) );
  NOR2_X1 U4549 ( .A1(n3846), .A2(n3884), .ZN(n3948) );
  INV_X1 U4550 ( .A(n3948), .ZN(n3829) );
  NAND2_X1 U4551 ( .A1(n3817), .A2(n3820), .ZN(n3929) );
  NAND2_X1 U4552 ( .A1(n3819), .A2(n3818), .ZN(n3911) );
  NAND2_X1 U4553 ( .A1(n3911), .A2(n3820), .ZN(n3928) );
  OAI21_X1 U4554 ( .B1(n3821), .B2(n3929), .A(n3928), .ZN(n3822) );
  NAND2_X1 U4555 ( .A1(n3822), .A2(n3935), .ZN(n3823) );
  NAND4_X1 U4556 ( .A1(n3823), .A2(n3936), .A3(n3931), .A4(n2166), .ZN(n3825)
         );
  INV_X1 U4557 ( .A(n3824), .ZN(n3939) );
  AOI21_X1 U4558 ( .B1(n3825), .B2(n3940), .A(n3939), .ZN(n3827) );
  OAI21_X1 U4559 ( .B1(n3827), .B2(n3942), .A(n3826), .ZN(n3828) );
  OAI221_X1 U4560 ( .B1(n3829), .B2(n3944), .C1(n3829), .C2(n3828), .A(n3953), 
        .ZN(n3831) );
  INV_X1 U4561 ( .A(n4278), .ZN(n4076) );
  NAND2_X1 U4562 ( .A1(n2138), .A2(DATAI_30_), .ZN(n4274) );
  NAND2_X1 U4563 ( .A1(n2137), .A2(DATAI_31_), .ZN(n4057) );
  NAND2_X1 U4564 ( .A1(n4056), .A2(n4057), .ZN(n3956) );
  OAI21_X1 U4565 ( .B1(n3843), .B2(n4274), .A(n3956), .ZN(n3850) );
  AOI21_X1 U4566 ( .B1(n4076), .B2(n3833), .A(n3850), .ZN(n3837) );
  INV_X1 U4567 ( .A(n3837), .ZN(n3830) );
  NOR4_X1 U4568 ( .A1(n3831), .A2(n3836), .A3(n3835), .A4(n3830), .ZN(n3842)
         );
  INV_X1 U4569 ( .A(n4086), .ZN(n3840) );
  OAI21_X1 U4570 ( .B1(n4076), .B2(n3833), .A(n3832), .ZN(n3838) );
  NOR2_X1 U4571 ( .A1(n3834), .A2(n3838), .ZN(n3949) );
  NOR2_X1 U4572 ( .A1(n3836), .A2(n3835), .ZN(n3839) );
  OAI21_X1 U4573 ( .B1(n3839), .B2(n3838), .A(n3837), .ZN(n3954) );
  AOI21_X1 U4574 ( .B1(n3840), .B2(n3949), .A(n3954), .ZN(n3841) );
  OAI22_X1 U4575 ( .A1(n3842), .A2(n3841), .B1(n4274), .B2(n4056), .ZN(n3964)
         );
  NAND2_X1 U4576 ( .A1(n3843), .A2(n4274), .ZN(n3849) );
  AOI21_X1 U4577 ( .B1(n3849), .B2(n4056), .A(n4057), .ZN(n3845) );
  NOR2_X1 U4578 ( .A1(n3845), .A2(n3844), .ZN(n3963) );
  INV_X1 U4579 ( .A(n3846), .ZN(n3848) );
  NAND2_X1 U4580 ( .A1(n3848), .A2(n3847), .ZN(n4112) );
  OAI21_X1 U4581 ( .B1(n4056), .B2(n4057), .A(n3849), .ZN(n3957) );
  NOR2_X1 U4582 ( .A1(n3850), .A2(n4410), .ZN(n3851) );
  NAND2_X1 U4583 ( .A1(n4566), .A2(n3851), .ZN(n3853) );
  NOR4_X1 U4584 ( .A1(n4112), .A2(n3957), .A3(n3853), .A4(n3852), .ZN(n3876)
         );
  INV_X1 U4585 ( .A(n3854), .ZN(n3855) );
  NAND4_X1 U4586 ( .A1(n4248), .A2(n3855), .A3(n2683), .A4(n2145), .ZN(n3862)
         );
  INV_X1 U4587 ( .A(n3856), .ZN(n3858) );
  NAND4_X1 U4588 ( .A1(n3860), .A2(n3859), .A3(n3858), .A4(n3857), .ZN(n3861)
         );
  NOR2_X1 U4589 ( .A1(n3862), .A2(n3861), .ZN(n3874) );
  NAND4_X1 U4590 ( .A1(n3865), .A2(n3864), .A3(n2363), .A4(n3863), .ZN(n3872)
         );
  INV_X1 U4591 ( .A(n3866), .ZN(n3867) );
  NAND4_X1 U4592 ( .A1(n3870), .A2(n3869), .A3(n3868), .A4(n3867), .ZN(n3871)
         );
  NOR2_X1 U4593 ( .A1(n3872), .A2(n3871), .ZN(n3873) );
  NAND4_X1 U4594 ( .A1(n3876), .A2(n3875), .A3(n3874), .A4(n3873), .ZN(n3877)
         );
  XNOR2_X1 U4595 ( .A(n4287), .B(n4105), .ZN(n4097) );
  OR4_X1 U4596 ( .A1(n4068), .A2(n3878), .A3(n3877), .A4(n4097), .ZN(n3887) );
  INV_X1 U4597 ( .A(n4148), .ZN(n3879) );
  AND2_X1 U4598 ( .A1(n3879), .A2(n4147), .ZN(n4187) );
  INV_X1 U4599 ( .A(n3880), .ZN(n3882) );
  AND2_X1 U4600 ( .A1(n3882), .A2(n3881), .ZN(n4208) );
  XNOR2_X1 U4601 ( .A(n4304), .B(n4160), .ZN(n4152) );
  OR2_X1 U4602 ( .A1(n3884), .A2(n3883), .ZN(n4133) );
  XNOR2_X1 U4603 ( .A(n3975), .B(n4236), .ZN(n4230) );
  NOR4_X1 U4604 ( .A1(n4208), .A2(n4152), .A3(n4133), .A4(n4230), .ZN(n3885)
         );
  NAND3_X1 U4605 ( .A1(n4151), .A2(n4187), .A3(n3885), .ZN(n3886) );
  NOR3_X1 U4606 ( .A1(n3887), .A2(n3886), .A3(n4086), .ZN(n3961) );
  OAI211_X1 U4607 ( .C1(n2321), .C2(n4410), .A(n3890), .B(n3889), .ZN(n3893)
         );
  NAND3_X1 U4608 ( .A1(n3893), .A2(n3892), .A3(n3891), .ZN(n3896) );
  NAND3_X1 U4609 ( .A1(n3896), .A2(n3895), .A3(n3894), .ZN(n3899) );
  NAND3_X1 U4610 ( .A1(n3899), .A2(n3898), .A3(n3897), .ZN(n3902) );
  NAND4_X1 U4611 ( .A1(n3902), .A2(n3901), .A3(n2208), .A4(n3900), .ZN(n3905)
         );
  AND3_X1 U4612 ( .A1(n3905), .A2(n3904), .A3(n3903), .ZN(n3910) );
  NAND2_X1 U4613 ( .A1(n3907), .A2(n3906), .ZN(n3916) );
  OAI211_X1 U4614 ( .C1(n3910), .C2(n3916), .A(n3909), .B(n3908), .ZN(n3913)
         );
  INV_X1 U4615 ( .A(n3911), .ZN(n3912) );
  NAND3_X1 U4616 ( .A1(n3913), .A2(n3912), .A3(n2225), .ZN(n3922) );
  NOR4_X1 U4617 ( .A1(n3917), .A2(n3916), .A3(n3915), .A4(n3914), .ZN(n3920)
         );
  INV_X1 U4618 ( .A(n3918), .ZN(n3919) );
  OAI21_X1 U4619 ( .B1(n3920), .B2(n3919), .A(n3928), .ZN(n3921) );
  NAND2_X1 U4620 ( .A1(n3922), .A2(n3921), .ZN(n3926) );
  NAND4_X1 U4621 ( .A1(n3926), .A2(n3925), .A3(n3924), .A4(n3923), .ZN(n3934)
         );
  INV_X1 U4622 ( .A(n3927), .ZN(n3930) );
  OAI21_X1 U4623 ( .B1(n3930), .B2(n3929), .A(n3928), .ZN(n3933) );
  INV_X1 U4624 ( .A(n3931), .ZN(n3932) );
  AOI21_X1 U4625 ( .B1(n3934), .B2(n3933), .A(n3932), .ZN(n3938) );
  INV_X1 U4626 ( .A(n3935), .ZN(n3937) );
  OAI211_X1 U4627 ( .C1(n3938), .C2(n3937), .A(n3936), .B(n2166), .ZN(n3941)
         );
  AOI211_X1 U4628 ( .C1(n3941), .C2(n3940), .A(n3939), .B(n4148), .ZN(n3943)
         );
  NOR2_X1 U4629 ( .A1(n3943), .A2(n3942), .ZN(n3946) );
  OAI21_X1 U4630 ( .B1(n3946), .B2(n3945), .A(n3944), .ZN(n3947) );
  NAND2_X1 U4631 ( .A1(n3948), .A2(n3947), .ZN(n3952) );
  INV_X1 U4632 ( .A(n3949), .ZN(n3950) );
  AOI211_X1 U4633 ( .C1(n3953), .C2(n3952), .A(n3951), .B(n3950), .ZN(n3955)
         );
  OR2_X1 U4634 ( .A1(n3955), .A2(n3954), .ZN(n3959) );
  NAND2_X1 U4635 ( .A1(n3957), .A2(n3956), .ZN(n3958) );
  AND2_X1 U4636 ( .A1(n3959), .A2(n3958), .ZN(n3960) );
  MUX2_X1 U4637 ( .A(n3961), .B(n3960), .S(n2676), .Z(n3962) );
  AOI21_X1 U4638 ( .B1(n3964), .B2(n3963), .A(n3962), .ZN(n3965) );
  XNOR2_X1 U4639 ( .A(n3965), .B(n4050), .ZN(n3972) );
  NAND2_X1 U4640 ( .A1(n3967), .A2(n3966), .ZN(n3968) );
  OAI211_X1 U4641 ( .C1(n3969), .C2(n3971), .A(n3968), .B(B_REG_SCAN_IN), .ZN(
        n3970) );
  OAI21_X1 U4642 ( .B1(n3972), .B2(n3971), .A(n3970), .ZN(U3239) );
  MUX2_X1 U4643 ( .A(DATAO_REG_28__SCAN_IN), .B(n3973), .S(n3985), .Z(U3578)
         );
  MUX2_X1 U4644 ( .A(DATAO_REG_24__SCAN_IN), .B(n4116), .S(n3985), .Z(U3574)
         );
  MUX2_X1 U4645 ( .A(DATAO_REG_21__SCAN_IN), .B(n4206), .S(n3985), .Z(U3571)
         );
  MUX2_X1 U4646 ( .A(DATAO_REG_20__SCAN_IN), .B(n3974), .S(n3985), .Z(U3570)
         );
  MUX2_X1 U4647 ( .A(DATAO_REG_19__SCAN_IN), .B(n3975), .S(n3985), .Z(U3569)
         );
  MUX2_X1 U4648 ( .A(DATAO_REG_17__SCAN_IN), .B(n3976), .S(n3985), .Z(U3567)
         );
  MUX2_X1 U4649 ( .A(DATAO_REG_16__SCAN_IN), .B(n3977), .S(n3985), .Z(U3566)
         );
  MUX2_X1 U4650 ( .A(DATAO_REG_15__SCAN_IN), .B(n3978), .S(n3985), .Z(U3565)
         );
  MUX2_X1 U4651 ( .A(DATAO_REG_14__SCAN_IN), .B(n3979), .S(n3985), .Z(U3564)
         );
  MUX2_X1 U4652 ( .A(DATAO_REG_13__SCAN_IN), .B(n3980), .S(n3985), .Z(U3563)
         );
  MUX2_X1 U4653 ( .A(DATAO_REG_12__SCAN_IN), .B(n3981), .S(n3985), .Z(U3562)
         );
  MUX2_X1 U4654 ( .A(DATAO_REG_9__SCAN_IN), .B(n3982), .S(n3985), .Z(U3559) );
  MUX2_X1 U4655 ( .A(DATAO_REG_8__SCAN_IN), .B(n3983), .S(n3985), .Z(U3558) );
  MUX2_X1 U4656 ( .A(DATAO_REG_5__SCAN_IN), .B(n3984), .S(n3985), .Z(U3555) );
  MUX2_X1 U4657 ( .A(DATAO_REG_4__SCAN_IN), .B(n3099), .S(n3985), .Z(U3554) );
  MUX2_X1 U4658 ( .A(DATAO_REG_1__SCAN_IN), .B(n2948), .S(n3985), .Z(U3551) );
  XNOR2_X1 U4659 ( .A(n4037), .B(REG2_REG_17__SCAN_IN), .ZN(n4002) );
  INV_X1 U4660 ( .A(n4470), .ZN(n4004) );
  NAND2_X1 U4661 ( .A1(n4004), .A2(REG2_REG_11__SCAN_IN), .ZN(n3993) );
  MUX2_X1 U4662 ( .A(n4747), .B(REG2_REG_11__SCAN_IN), .S(n4470), .Z(n4466) );
  NAND2_X1 U4663 ( .A1(n4440), .A2(REG2_REG_9__SCAN_IN), .ZN(n3990) );
  MUX2_X1 U4664 ( .A(REG2_REG_9__SCAN_IN), .B(n3206), .S(n4440), .Z(n4445) );
  OAI21_X1 U4665 ( .B1(n4414), .B2(n3987), .A(n3986), .ZN(n3988) );
  NAND2_X1 U4666 ( .A1(n4600), .A2(n3988), .ZN(n3989) );
  XNOR2_X1 U4667 ( .A(n3988), .B(n4439), .ZN(n4431) );
  NAND2_X1 U4668 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4431), .ZN(n4430) );
  NAND2_X1 U4669 ( .A1(n3989), .A2(n4430), .ZN(n4446) );
  NAND2_X1 U4670 ( .A1(n4445), .A2(n4446), .ZN(n4444) );
  NAND2_X1 U4671 ( .A1(n3990), .A2(n4444), .ZN(n3991) );
  NAND2_X1 U4672 ( .A1(n4013), .A2(n3991), .ZN(n3992) );
  INV_X1 U4673 ( .A(n4013), .ZN(n4561) );
  XNOR2_X1 U4674 ( .A(n3991), .B(n4561), .ZN(n4454) );
  NAND2_X1 U4675 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4454), .ZN(n4453) );
  NAND2_X1 U4676 ( .A1(n3992), .A2(n4453), .ZN(n4467) );
  NAND2_X1 U4677 ( .A1(n4466), .A2(n4467), .ZN(n4465) );
  NAND2_X1 U4678 ( .A1(n3993), .A2(n4465), .ZN(n3994) );
  NAND2_X1 U4679 ( .A1(n4016), .A2(n3994), .ZN(n3995) );
  INV_X1 U4680 ( .A(n4016), .ZN(n4560) );
  XNOR2_X1 U4681 ( .A(n3994), .B(n4560), .ZN(n4475) );
  NAND2_X1 U4682 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4475), .ZN(n4474) );
  NAND2_X1 U4683 ( .A1(n3995), .A2(n4474), .ZN(n4485) );
  NOR2_X1 U4684 ( .A1(n4558), .A2(n3996), .ZN(n3997) );
  INV_X1 U4685 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4497) );
  NAND2_X1 U4686 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4003), .ZN(n3998) );
  OAI21_X1 U4687 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4003), .A(n3998), .ZN(n4505) );
  NOR2_X1 U4688 ( .A1(n4506), .A2(n4505), .ZN(n4504) );
  NAND2_X1 U4689 ( .A1(n3999), .A2(n4555), .ZN(n4000) );
  NAND2_X1 U4690 ( .A1(n4001), .A2(n4002), .ZN(n4038) );
  AOI221_X1 U4691 ( .B1(n4002), .B2(n4038), .C1(n4001), .C2(n4038), .A(n4527), 
        .ZN(n4035) );
  NAND2_X1 U4692 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4003), .ZN(n4023) );
  INV_X1 U4693 ( .A(n4003), .ZN(n4557) );
  AOI22_X1 U4694 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4003), .B1(n4557), .B2(
        n3466), .ZN(n4511) );
  NAND2_X1 U4695 ( .A1(n4004), .A2(REG1_REG_11__SCAN_IN), .ZN(n4015) );
  INV_X1 U4696 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4005) );
  MUX2_X1 U4697 ( .A(REG1_REG_11__SCAN_IN), .B(n4005), .S(n4470), .Z(n4006) );
  INV_X1 U4698 ( .A(n4006), .ZN(n4463) );
  NAND2_X1 U4699 ( .A1(n4440), .A2(REG1_REG_9__SCAN_IN), .ZN(n4011) );
  MUX2_X1 U4700 ( .A(n3250), .B(REG1_REG_9__SCAN_IN), .S(n4440), .Z(n4007) );
  INV_X1 U4701 ( .A(n4007), .ZN(n4442) );
  NAND2_X1 U4702 ( .A1(n4009), .A2(n4600), .ZN(n4010) );
  NAND2_X1 U4703 ( .A1(n4442), .A2(n4443), .ZN(n4441) );
  NAND2_X1 U4704 ( .A1(n4013), .A2(n4012), .ZN(n4014) );
  NAND2_X1 U4705 ( .A1(n4463), .A2(n4464), .ZN(n4462) );
  NAND2_X1 U4706 ( .A1(n4016), .A2(n4017), .ZN(n4018) );
  INV_X1 U4707 ( .A(n4483), .ZN(n4559) );
  AOI22_X1 U4708 ( .A1(n4483), .A2(REG1_REG_13__SCAN_IN), .B1(n3416), .B2(
        n4559), .ZN(n4491) );
  NAND2_X1 U4709 ( .A1(n4483), .A2(REG1_REG_13__SCAN_IN), .ZN(n4019) );
  NAND2_X1 U4710 ( .A1(n4020), .A2(n4021), .ZN(n4022) );
  XNOR2_X1 U4711 ( .A(n4021), .B(n4558), .ZN(n4501) );
  NAND2_X1 U4712 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4501), .ZN(n4500) );
  NOR2_X1 U4713 ( .A1(n4024), .A2(n4025), .ZN(n4026) );
  INV_X1 U4714 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4027) );
  NAND2_X1 U4715 ( .A1(n4037), .A2(n4027), .ZN(n4041) );
  OAI21_X1 U4716 ( .B1(n4037), .B2(n4027), .A(n4041), .ZN(n4028) );
  AOI21_X1 U4717 ( .B1(n4029), .B2(n4028), .A(n4042), .ZN(n4030) );
  NOR2_X1 U4718 ( .A1(n4030), .A2(n4518), .ZN(n4034) );
  AOI21_X1 U4719 ( .B1(n4531), .B2(ADDR_REG_17__SCAN_IN), .A(n4031), .ZN(n4032) );
  OAI21_X1 U4720 ( .B1(n4538), .B2(n4037), .A(n4032), .ZN(n4033) );
  OR3_X1 U4721 ( .A1(n4035), .A2(n4034), .A3(n4033), .ZN(U3257) );
  INV_X1 U4722 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4862) );
  MUX2_X1 U4723 ( .A(REG2_REG_19__SCAN_IN), .B(n4862), .S(n4412), .Z(n4040) );
  INV_X1 U4724 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4036) );
  AOI22_X1 U4725 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4537), .B1(n4553), .B2(
        n4036), .ZN(n4529) );
  INV_X1 U4726 ( .A(n4037), .ZN(n4413) );
  AOI21_X1 U4727 ( .B1(n4553), .B2(REG2_REG_18__SCAN_IN), .A(n4528), .ZN(n4039) );
  XOR2_X1 U4728 ( .A(n4040), .B(n4039), .Z(n4054) );
  INV_X1 U4729 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U4730 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4553), .B1(n4537), .B2(
        n4044), .ZN(n4534) );
  INV_X1 U4731 ( .A(n4041), .ZN(n4043) );
  OAI21_X1 U4732 ( .B1(n4044), .B2(n4537), .A(n4532), .ZN(n4047) );
  INV_X1 U4733 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4045) );
  MUX2_X1 U4734 ( .A(n4045), .B(REG1_REG_19__SCAN_IN), .S(n4412), .Z(n4046) );
  XNOR2_X1 U4735 ( .A(n4047), .B(n4046), .ZN(n4052) );
  NAND2_X1 U4736 ( .A1(n4531), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4048) );
  OAI211_X1 U4737 ( .C1(n4538), .C2(n4050), .A(n4049), .B(n4048), .ZN(n4051)
         );
  AOI21_X1 U4738 ( .B1(n4052), .B2(n4533), .A(n4051), .ZN(n4053) );
  OAI21_X1 U4739 ( .B1(n4054), .B2(n4527), .A(n4053), .ZN(U3259) );
  INV_X1 U4740 ( .A(n4274), .ZN(n4271) );
  XNOR2_X1 U4741 ( .A(n4269), .B(n4057), .ZN(n4363) );
  NAND2_X1 U4742 ( .A1(n4056), .A2(n4055), .ZN(n4272) );
  OAI21_X1 U4743 ( .B1(n4057), .B2(n4273), .A(n4272), .ZN(n4360) );
  NAND2_X1 U4744 ( .A1(n4421), .A2(n4360), .ZN(n4059) );
  NAND2_X1 U4745 ( .A1(n4222), .A2(REG2_REG_31__SCAN_IN), .ZN(n4058) );
  OAI211_X1 U4746 ( .C1(n4363), .C2(n4238), .A(n4059), .B(n4058), .ZN(U3260)
         );
  INV_X1 U4747 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4065) );
  NAND2_X1 U4748 ( .A1(n4060), .A2(n4188), .ZN(n4064) );
  XOR2_X1 U4749 ( .A(n4068), .B(n4066), .Z(n4067) );
  NAND2_X1 U4750 ( .A1(n4067), .A2(n4254), .ZN(n4280) );
  INV_X1 U4751 ( .A(n4068), .ZN(n4069) );
  XNOR2_X1 U4752 ( .A(n4070), .B(n4069), .ZN(n4283) );
  NAND2_X1 U4753 ( .A1(n4283), .A2(n4188), .ZN(n4082) );
  AND2_X1 U4754 ( .A1(n2144), .A2(n4277), .ZN(n4071) );
  OR2_X1 U4755 ( .A1(n4072), .A2(n4071), .ZN(n4369) );
  INV_X1 U4756 ( .A(n4369), .ZN(n4080) );
  INV_X1 U4757 ( .A(n4073), .ZN(n4074) );
  AOI22_X1 U4758 ( .A1(n4074), .A2(n4539), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4222), .ZN(n4075) );
  OAI21_X1 U4759 ( .B1(n4076), .B2(n4193), .A(n4075), .ZN(n4079) );
  OAI22_X1 U4760 ( .A1(n4281), .A2(n4197), .B1(n4196), .B2(n4077), .ZN(n4078)
         );
  AOI211_X1 U4761 ( .C1(n4080), .C2(n4543), .A(n4079), .B(n4078), .ZN(n4081)
         );
  OAI211_X1 U4762 ( .C1(n4222), .C2(n4280), .A(n4082), .B(n4081), .ZN(U3262)
         );
  XNOR2_X1 U4763 ( .A(n4083), .B(n4086), .ZN(n4084) );
  NAND2_X1 U4764 ( .A1(n4084), .A2(n4254), .ZN(n4289) );
  XOR2_X1 U4765 ( .A(n4086), .B(n4085), .Z(n4292) );
  NAND2_X1 U4766 ( .A1(n4292), .A2(n4188), .ZN(n4094) );
  NAND2_X1 U4767 ( .A1(n4104), .A2(n4286), .ZN(n4087) );
  NAND2_X1 U4768 ( .A1(n2144), .A2(n4087), .ZN(n4373) );
  INV_X1 U4769 ( .A(n4373), .ZN(n4092) );
  AOI22_X1 U4770 ( .A1(n4088), .A2(n4539), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4222), .ZN(n4089) );
  OAI21_X1 U4771 ( .B1(n4290), .B2(n4193), .A(n4089), .ZN(n4091) );
  OAI22_X1 U4772 ( .A1(n4119), .A2(n4197), .B1(n2643), .B2(n4196), .ZN(n4090)
         );
  AOI211_X1 U4773 ( .C1(n4092), .C2(n4543), .A(n4091), .B(n4090), .ZN(n4093)
         );
  OAI211_X1 U4774 ( .C1(n4222), .C2(n4289), .A(n4094), .B(n4093), .ZN(U3263)
         );
  XNOR2_X1 U4775 ( .A(n2153), .B(n4097), .ZN(n4296) );
  INV_X1 U4776 ( .A(n4296), .ZN(n4110) );
  NOR2_X1 U4777 ( .A1(n4096), .A2(n4095), .ZN(n4098) );
  XNOR2_X1 U4778 ( .A(n4098), .B(n4097), .ZN(n4099) );
  NAND2_X1 U4779 ( .A1(n4099), .A2(n4254), .ZN(n4103) );
  AOI22_X1 U4780 ( .A1(n4101), .A2(n4303), .B1(n4100), .B2(n4342), .ZN(n4102)
         );
  OAI211_X1 U4781 ( .C1(n4281), .C2(n4307), .A(n4103), .B(n4102), .ZN(n4295)
         );
  OAI21_X1 U4782 ( .B1(n4120), .B2(n4105), .A(n4104), .ZN(n4377) );
  AOI22_X1 U4783 ( .A1(n4106), .A2(n4539), .B1(n4222), .B2(
        REG2_REG_26__SCAN_IN), .ZN(n4107) );
  OAI21_X1 U4784 ( .B1(n4377), .B2(n4238), .A(n4107), .ZN(n4108) );
  AOI21_X1 U4785 ( .B1(n4295), .B2(n4421), .A(n4108), .ZN(n4109) );
  OAI21_X1 U4786 ( .B1(n4110), .B2(n4265), .A(n4109), .ZN(U3264) );
  XOR2_X1 U4787 ( .A(n4112), .B(n4111), .Z(n4299) );
  INV_X1 U4788 ( .A(n4299), .ZN(n4127) );
  XNOR2_X1 U4789 ( .A(n4113), .B(n4112), .ZN(n4114) );
  NAND2_X1 U4790 ( .A1(n4114), .A2(n4254), .ZN(n4118) );
  AOI22_X1 U4791 ( .A1(n4116), .A2(n4303), .B1(n4115), .B2(n4342), .ZN(n4117)
         );
  OAI211_X1 U4792 ( .C1(n4119), .C2(n4307), .A(n4118), .B(n4117), .ZN(n4298)
         );
  INV_X1 U4793 ( .A(n4120), .ZN(n4121) );
  OAI21_X1 U4794 ( .B1(n4135), .B2(n4122), .A(n4121), .ZN(n4381) );
  AOI22_X1 U4795 ( .A1(n4222), .A2(REG2_REG_25__SCAN_IN), .B1(n4123), .B2(
        n4539), .ZN(n4124) );
  OAI21_X1 U4796 ( .B1(n4381), .B2(n4238), .A(n4124), .ZN(n4125) );
  AOI21_X1 U4797 ( .B1(n4298), .B2(n4421), .A(n4125), .ZN(n4126) );
  OAI21_X1 U4798 ( .B1(n4127), .B2(n4265), .A(n4126), .ZN(U3265) );
  OR2_X1 U4799 ( .A1(n4129), .A2(n4128), .ZN(n4131) );
  INV_X1 U4800 ( .A(n4133), .ZN(n4130) );
  XNOR2_X1 U4801 ( .A(n4131), .B(n4130), .ZN(n4132) );
  NAND2_X1 U4802 ( .A1(n4132), .A2(n4254), .ZN(n4306) );
  XNOR2_X1 U4803 ( .A(n4134), .B(n4133), .ZN(n4310) );
  NAND2_X1 U4804 ( .A1(n4310), .A2(n4188), .ZN(n4145) );
  INV_X1 U4805 ( .A(n4159), .ZN(n4137) );
  INV_X1 U4806 ( .A(n4135), .ZN(n4136) );
  OAI21_X1 U4807 ( .B1(n4137), .B2(n4140), .A(n4136), .ZN(n4385) );
  INV_X1 U4808 ( .A(n4385), .ZN(n4143) );
  AOI22_X1 U4809 ( .A1(n4222), .A2(REG2_REG_24__SCAN_IN), .B1(n4138), .B2(
        n4539), .ZN(n4139) );
  OAI21_X1 U4810 ( .B1(n4308), .B2(n4193), .A(n4139), .ZN(n4142) );
  OAI22_X1 U4811 ( .A1(n4172), .A2(n4197), .B1(n4196), .B2(n4140), .ZN(n4141)
         );
  AOI211_X1 U4812 ( .C1(n4143), .C2(n4543), .A(n4142), .B(n4141), .ZN(n4144)
         );
  OAI211_X1 U4813 ( .C1(n4222), .C2(n4306), .A(n4145), .B(n4144), .ZN(U3266)
         );
  XOR2_X1 U4814 ( .A(n4152), .B(n4146), .Z(n4313) );
  INV_X1 U4815 ( .A(n4313), .ZN(n4167) );
  OAI21_X1 U4816 ( .B1(n4184), .B2(n4148), .A(n4147), .ZN(n4171) );
  INV_X1 U4817 ( .A(n4149), .ZN(n4150) );
  AOI21_X1 U4818 ( .B1(n4171), .B2(n4151), .A(n4150), .ZN(n4153) );
  XNOR2_X1 U4819 ( .A(n4153), .B(n4152), .ZN(n4154) );
  NAND2_X1 U4820 ( .A1(n4154), .A2(n4254), .ZN(n4157) );
  AOI22_X1 U4821 ( .A1(n4322), .A2(n4303), .B1(n4342), .B2(n4155), .ZN(n4156)
         );
  OAI211_X1 U4822 ( .C1(n4158), .C2(n4307), .A(n4157), .B(n4156), .ZN(n4312)
         );
  INV_X1 U4823 ( .A(n4176), .ZN(n4161) );
  OAI21_X1 U4824 ( .B1(n4161), .B2(n4160), .A(n4159), .ZN(n4388) );
  NOR2_X1 U4825 ( .A1(n4388), .A2(n4238), .ZN(n4165) );
  INV_X1 U4826 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4163) );
  OAI22_X1 U4827 ( .A1(n4421), .A2(n4163), .B1(n4162), .B2(n4239), .ZN(n4164)
         );
  AOI211_X1 U4828 ( .C1(n4312), .C2(n4421), .A(n4165), .B(n4164), .ZN(n4166)
         );
  OAI21_X1 U4829 ( .B1(n4167), .B2(n4265), .A(n4166), .ZN(U3267) );
  OAI21_X1 U4830 ( .B1(n4169), .B2(n4170), .A(n4168), .ZN(n4316) );
  XNOR2_X1 U4831 ( .A(n4171), .B(n4170), .ZN(n4175) );
  OAI22_X1 U4832 ( .A1(n4172), .A2(n4307), .B1(n4177), .B2(n4273), .ZN(n4173)
         );
  AOI21_X1 U4833 ( .B1(n4303), .B2(n4206), .A(n4173), .ZN(n4174) );
  OAI21_X1 U4834 ( .B1(n4175), .B2(n4233), .A(n4174), .ZN(n4317) );
  OAI21_X1 U4835 ( .B1(n4189), .B2(n4177), .A(n4176), .ZN(n4392) );
  NOR2_X1 U4836 ( .A1(n4392), .A2(n4238), .ZN(n4181) );
  INV_X1 U4837 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4179) );
  OAI22_X1 U4838 ( .A1(n4421), .A2(n4179), .B1(n4178), .B2(n4239), .ZN(n4180)
         );
  AOI211_X1 U4839 ( .C1(n4317), .C2(n4421), .A(n4181), .B(n4180), .ZN(n4182)
         );
  OAI21_X1 U4840 ( .B1(n4316), .B2(n4265), .A(n4182), .ZN(U3268) );
  INV_X1 U4841 ( .A(n4187), .ZN(n4183) );
  XNOR2_X1 U4842 ( .A(n4184), .B(n4183), .ZN(n4185) );
  NAND2_X1 U4843 ( .A1(n4185), .A2(n4254), .ZN(n4324) );
  XOR2_X1 U4844 ( .A(n4187), .B(n4186), .Z(n4327) );
  NAND2_X1 U4845 ( .A1(n4327), .A2(n4188), .ZN(n4202) );
  INV_X1 U4846 ( .A(n4189), .ZN(n4190) );
  OAI21_X1 U4847 ( .B1(n4215), .B2(n4195), .A(n4190), .ZN(n4396) );
  INV_X1 U4848 ( .A(n4396), .ZN(n4200) );
  AOI22_X1 U4849 ( .A1(n4222), .A2(REG2_REG_21__SCAN_IN), .B1(n4191), .B2(
        n4539), .ZN(n4192) );
  OAI21_X1 U4850 ( .B1(n4194), .B2(n4193), .A(n4192), .ZN(n4199) );
  OAI22_X1 U4851 ( .A1(n4325), .A2(n4197), .B1(n4196), .B2(n4195), .ZN(n4198)
         );
  AOI211_X1 U4852 ( .C1(n4200), .C2(n4543), .A(n4199), .B(n4198), .ZN(n4201)
         );
  OAI211_X1 U4853 ( .C1(n4222), .C2(n4324), .A(n4202), .B(n4201), .ZN(U3269)
         );
  NAND2_X1 U4854 ( .A1(n4204), .A2(n4203), .ZN(n4205) );
  XOR2_X1 U4855 ( .A(n4205), .B(n4208), .Z(n4213) );
  AOI22_X1 U4856 ( .A1(n4206), .A2(n4344), .B1(n4342), .B2(n4216), .ZN(n4207)
         );
  OAI21_X1 U4857 ( .B1(n4251), .B2(n4348), .A(n4207), .ZN(n4212) );
  XNOR2_X1 U4858 ( .A(n4209), .B(n4208), .ZN(n4334) );
  NOR2_X1 U4859 ( .A1(n4334), .A2(n4210), .ZN(n4211) );
  AOI211_X1 U4860 ( .C1(n4254), .C2(n4213), .A(n4212), .B(n4211), .ZN(n4333)
         );
  AOI22_X1 U4861 ( .A1(n4222), .A2(REG2_REG_20__SCAN_IN), .B1(n4214), .B2(
        n4539), .ZN(n4218) );
  INV_X1 U4862 ( .A(n4215), .ZN(n4331) );
  NAND2_X1 U4863 ( .A1(n4235), .A2(n4216), .ZN(n4330) );
  NAND3_X1 U4864 ( .A1(n4331), .A2(n4543), .A3(n4330), .ZN(n4217) );
  OAI211_X1 U4865 ( .C1(n4334), .C2(n4219), .A(n4218), .B(n4217), .ZN(n4220)
         );
  INV_X1 U4866 ( .A(n4220), .ZN(n4221) );
  OAI21_X1 U4867 ( .B1(n4333), .B2(n4222), .A(n4221), .ZN(U3270) );
  XNOR2_X1 U4868 ( .A(n4223), .B(n4230), .ZN(n4336) );
  INV_X1 U4869 ( .A(n4336), .ZN(n4244) );
  NAND2_X1 U4870 ( .A1(n4225), .A2(n4224), .ZN(n4249) );
  INV_X1 U4871 ( .A(n4226), .ZN(n4228) );
  OAI21_X1 U4872 ( .B1(n4249), .B2(n4228), .A(n4227), .ZN(n4229) );
  XOR2_X1 U4873 ( .A(n4230), .B(n4229), .Z(n4234) );
  OAI22_X1 U4874 ( .A1(n4325), .A2(n4307), .B1(n4273), .B2(n4236), .ZN(n4231)
         );
  AOI21_X1 U4875 ( .B1(n4303), .B2(n4345), .A(n4231), .ZN(n4232) );
  OAI21_X1 U4876 ( .B1(n4234), .B2(n4233), .A(n4232), .ZN(n4335) );
  INV_X1 U4877 ( .A(n4256), .ZN(n4237) );
  OAI21_X1 U4878 ( .B1(n4237), .B2(n4236), .A(n4235), .ZN(n4401) );
  NOR2_X1 U4879 ( .A1(n4401), .A2(n4238), .ZN(n4242) );
  OAI22_X1 U4880 ( .A1(n4421), .A2(n4862), .B1(n4240), .B2(n4239), .ZN(n4241)
         );
  AOI211_X1 U4881 ( .C1(n4335), .C2(n4421), .A(n4242), .B(n4241), .ZN(n4243)
         );
  OAI21_X1 U4882 ( .B1(n4244), .B2(n4265), .A(n4243), .ZN(U3271) );
  INV_X1 U4883 ( .A(n4245), .ZN(n4246) );
  AOI21_X1 U4884 ( .B1(n4248), .B2(n4247), .A(n4246), .ZN(n4341) );
  XNOR2_X1 U4885 ( .A(n4249), .B(n4248), .ZN(n4255) );
  NOR2_X1 U4886 ( .A1(n4250), .A2(n4348), .ZN(n4253) );
  OAI22_X1 U4887 ( .A1(n4251), .A2(n4307), .B1(n4273), .B2(n4257), .ZN(n4252)
         );
  AOI211_X1 U4888 ( .C1(n4255), .C2(n4254), .A(n4253), .B(n4252), .ZN(n4340)
         );
  INV_X1 U4889 ( .A(n4340), .ZN(n4263) );
  OAI211_X1 U4890 ( .C1(n4258), .C2(n4257), .A(n4256), .B(n4354), .ZN(n4339)
         );
  AOI22_X1 U4891 ( .A1(n4222), .A2(REG2_REG_18__SCAN_IN), .B1(n4259), .B2(
        n4539), .ZN(n4260) );
  OAI21_X1 U4892 ( .B1(n4339), .B2(n4261), .A(n4260), .ZN(n4262) );
  AOI21_X1 U4893 ( .B1(n4263), .B2(n4421), .A(n4262), .ZN(n4264) );
  OAI21_X1 U4894 ( .B1(n4341), .B2(n4265), .A(n4264), .ZN(U3272) );
  NOR2_X1 U4895 ( .A1(n4599), .A2(n4266), .ZN(n4267) );
  AOI21_X1 U4896 ( .B1(n4599), .B2(n4360), .A(n4267), .ZN(n4268) );
  OAI21_X1 U4897 ( .B1(n4363), .B2(n4338), .A(n4268), .ZN(U3549) );
  AOI21_X1 U4898 ( .B1(n4271), .B2(n4270), .A(n4269), .ZN(n4419) );
  NAND2_X1 U4899 ( .A1(n4419), .A2(n4592), .ZN(n4276) );
  OAI21_X1 U4900 ( .B1(n4274), .B2(n4273), .A(n4272), .ZN(n4418) );
  NAND2_X1 U4901 ( .A1(n4599), .A2(n4418), .ZN(n4275) );
  OAI211_X1 U4902 ( .C1(n4599), .C2(n2717), .A(n4276), .B(n4275), .ZN(U3548)
         );
  AOI22_X1 U4903 ( .A1(n4278), .A2(n4344), .B1(n4342), .B2(n4277), .ZN(n4279)
         );
  OAI211_X1 U4904 ( .C1(n4281), .C2(n4348), .A(n4280), .B(n4279), .ZN(n4282)
         );
  AOI21_X1 U4905 ( .B1(n4283), .B2(n4582), .A(n4282), .ZN(n4366) );
  MUX2_X1 U4906 ( .A(n4284), .B(n4366), .S(n4599), .Z(n4285) );
  OAI21_X1 U4907 ( .B1(n4338), .B2(n4369), .A(n4285), .ZN(U3546) );
  AOI22_X1 U4908 ( .A1(n4287), .A2(n4303), .B1(n4286), .B2(n4342), .ZN(n4288)
         );
  OAI211_X1 U4909 ( .C1(n4290), .C2(n4307), .A(n4289), .B(n4288), .ZN(n4291)
         );
  AOI21_X1 U4910 ( .B1(n4292), .B2(n4582), .A(n4291), .ZN(n4370) );
  MUX2_X1 U4911 ( .A(n4293), .B(n4370), .S(n4599), .Z(n4294) );
  OAI21_X1 U4912 ( .B1(n4338), .B2(n4373), .A(n4294), .ZN(U3545) );
  AOI21_X1 U4913 ( .B1(n4296), .B2(n4582), .A(n4295), .ZN(n4374) );
  MUX2_X1 U4914 ( .A(n4732), .B(n4374), .S(n4599), .Z(n4297) );
  OAI21_X1 U4915 ( .B1(n4338), .B2(n4377), .A(n4297), .ZN(U3544) );
  AOI21_X1 U4916 ( .B1(n4299), .B2(n4582), .A(n4298), .ZN(n4378) );
  MUX2_X1 U4917 ( .A(n4300), .B(n4378), .S(n4599), .Z(n4301) );
  OAI21_X1 U4918 ( .B1(n4338), .B2(n4381), .A(n4301), .ZN(U3543) );
  AOI22_X1 U4919 ( .A1(n4304), .A2(n4303), .B1(n4342), .B2(n4302), .ZN(n4305)
         );
  OAI211_X1 U4920 ( .C1(n4308), .C2(n4307), .A(n4306), .B(n4305), .ZN(n4309)
         );
  AOI21_X1 U4921 ( .B1(n4310), .B2(n4582), .A(n4309), .ZN(n4382) );
  MUX2_X1 U4922 ( .A(n4730), .B(n4382), .S(n4599), .Z(n4311) );
  OAI21_X1 U4923 ( .B1(n4338), .B2(n4385), .A(n4311), .ZN(U3542) );
  AOI21_X1 U4924 ( .B1(n4313), .B2(n4582), .A(n4312), .ZN(n4386) );
  MUX2_X1 U4925 ( .A(n4314), .B(n4386), .S(n4599), .Z(n4315) );
  OAI21_X1 U4926 ( .B1(n4338), .B2(n4388), .A(n4315), .ZN(U3541) );
  INV_X1 U4927 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4319) );
  INV_X1 U4928 ( .A(n4316), .ZN(n4318) );
  AOI21_X1 U4929 ( .B1(n4318), .B2(n4582), .A(n4317), .ZN(n4389) );
  MUX2_X1 U4930 ( .A(n4319), .B(n4389), .S(n4599), .Z(n4320) );
  OAI21_X1 U4931 ( .B1(n4338), .B2(n4392), .A(n4320), .ZN(U3540) );
  INV_X1 U4932 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4328) );
  AOI22_X1 U4933 ( .A1(n4322), .A2(n4344), .B1(n4342), .B2(n4321), .ZN(n4323)
         );
  OAI211_X1 U4934 ( .C1(n4325), .C2(n4348), .A(n4324), .B(n4323), .ZN(n4326)
         );
  AOI21_X1 U4935 ( .B1(n4327), .B2(n4582), .A(n4326), .ZN(n4393) );
  MUX2_X1 U4936 ( .A(n4328), .B(n4393), .S(n4599), .Z(n4329) );
  OAI21_X1 U4937 ( .B1(n4338), .B2(n4396), .A(n4329), .ZN(U3539) );
  NAND3_X1 U4938 ( .A1(n4331), .A2(n4330), .A3(n4354), .ZN(n4332) );
  OAI211_X1 U4939 ( .C1(n4334), .C2(n4565), .A(n4333), .B(n4332), .ZN(n4397)
         );
  MUX2_X1 U4940 ( .A(REG1_REG_20__SCAN_IN), .B(n4397), .S(n4599), .Z(U3538) );
  AOI21_X1 U4941 ( .B1(n4336), .B2(n4582), .A(n4335), .ZN(n4398) );
  MUX2_X1 U4942 ( .A(n4045), .B(n4398), .S(n4599), .Z(n4337) );
  OAI21_X1 U4943 ( .B1(n4338), .B2(n4401), .A(n4337), .ZN(U3537) );
  OAI211_X1 U4944 ( .C1(n4341), .C2(n4358), .A(n4340), .B(n4339), .ZN(n4402)
         );
  MUX2_X1 U4945 ( .A(REG1_REG_18__SCAN_IN), .B(n4402), .S(n4599), .Z(U3536) );
  AOI22_X1 U4946 ( .A1(n4345), .A2(n4344), .B1(n4343), .B2(n4342), .ZN(n4346)
         );
  OAI211_X1 U4947 ( .C1(n4349), .C2(n4348), .A(n4347), .B(n4346), .ZN(n4350)
         );
  AOI21_X1 U4948 ( .B1(n4351), .B2(n4582), .A(n4350), .ZN(n4403) );
  MUX2_X1 U4949 ( .A(n4027), .B(n4403), .S(n4599), .Z(n4352) );
  OAI21_X1 U4950 ( .B1(n4338), .B2(n4407), .A(n4352), .ZN(U3535) );
  NAND3_X1 U4951 ( .A1(n4355), .A2(n4354), .A3(n4353), .ZN(n4356) );
  OAI211_X1 U4952 ( .C1(n4359), .C2(n4358), .A(n4357), .B(n4356), .ZN(n4408)
         );
  MUX2_X1 U4953 ( .A(REG1_REG_16__SCAN_IN), .B(n4408), .S(n4599), .Z(U3534) );
  NAND2_X1 U4954 ( .A1(n4589), .A2(n4360), .ZN(n4362) );
  NAND2_X1 U4955 ( .A1(n4587), .A2(REG0_REG_31__SCAN_IN), .ZN(n4361) );
  OAI211_X1 U4956 ( .C1(n4363), .C2(n4406), .A(n4362), .B(n4361), .ZN(U3517)
         );
  INV_X1 U4957 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4717) );
  NAND2_X1 U4958 ( .A1(n4419), .A2(n4574), .ZN(n4365) );
  NAND2_X1 U4959 ( .A1(n4589), .A2(n4418), .ZN(n4364) );
  OAI211_X1 U4960 ( .C1(n4589), .C2(n4717), .A(n4365), .B(n4364), .ZN(U3516)
         );
  INV_X1 U4961 ( .A(REG0_REG_28__SCAN_IN), .ZN(n4367) );
  MUX2_X1 U4962 ( .A(n4367), .B(n4366), .S(n4589), .Z(n4368) );
  OAI21_X1 U4963 ( .B1(n4369), .B2(n4406), .A(n4368), .ZN(U3514) );
  INV_X1 U4964 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4371) );
  MUX2_X1 U4965 ( .A(n4371), .B(n4370), .S(n4589), .Z(n4372) );
  OAI21_X1 U4966 ( .B1(n4373), .B2(n4406), .A(n4372), .ZN(U3513) );
  INV_X1 U4967 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4375) );
  MUX2_X1 U4968 ( .A(n4375), .B(n4374), .S(n4589), .Z(n4376) );
  OAI21_X1 U4969 ( .B1(n4377), .B2(n4406), .A(n4376), .ZN(U3512) );
  INV_X1 U4970 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4379) );
  MUX2_X1 U4971 ( .A(n4379), .B(n4378), .S(n4589), .Z(n4380) );
  OAI21_X1 U4972 ( .B1(n4381), .B2(n4406), .A(n4380), .ZN(U3511) );
  INV_X1 U4973 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4383) );
  MUX2_X1 U4974 ( .A(n4383), .B(n4382), .S(n4589), .Z(n4384) );
  OAI21_X1 U4975 ( .B1(n4385), .B2(n4406), .A(n4384), .ZN(U3510) );
  MUX2_X1 U4976 ( .A(n4703), .B(n4386), .S(n4589), .Z(n4387) );
  OAI21_X1 U4977 ( .B1(n4388), .B2(n4406), .A(n4387), .ZN(U3509) );
  INV_X1 U4978 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4390) );
  MUX2_X1 U4979 ( .A(n4390), .B(n4389), .S(n4589), .Z(n4391) );
  OAI21_X1 U4980 ( .B1(n4392), .B2(n4406), .A(n4391), .ZN(U3508) );
  INV_X1 U4981 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4394) );
  MUX2_X1 U4982 ( .A(n4394), .B(n4393), .S(n4589), .Z(n4395) );
  OAI21_X1 U4983 ( .B1(n4396), .B2(n4406), .A(n4395), .ZN(U3507) );
  MUX2_X1 U4984 ( .A(REG0_REG_20__SCAN_IN), .B(n4397), .S(n4589), .Z(U3506) );
  INV_X1 U4985 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4399) );
  MUX2_X1 U4986 ( .A(n4399), .B(n4398), .S(n4589), .Z(n4400) );
  OAI21_X1 U4987 ( .B1(n4401), .B2(n4406), .A(n4400), .ZN(U3505) );
  MUX2_X1 U4988 ( .A(REG0_REG_18__SCAN_IN), .B(n4402), .S(n4589), .Z(U3503) );
  INV_X1 U4989 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4404) );
  MUX2_X1 U4990 ( .A(n4404), .B(n4403), .S(n4589), .Z(n4405) );
  OAI21_X1 U4991 ( .B1(n4407), .B2(n4406), .A(n4405), .ZN(U3501) );
  MUX2_X1 U4992 ( .A(REG0_REG_16__SCAN_IN), .B(n4408), .S(n4589), .Z(U3499) );
  MUX2_X1 U4993 ( .A(n2381), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U4994 ( .A(n4409), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U4995 ( .A(n4410), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U4996 ( .A(DATAI_20_), .B(n4411), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4997 ( .A(n4412), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4998 ( .A(n4413), .B(DATAI_17_), .S(U3149), .Z(U3335) );
  MUX2_X1 U4999 ( .A(n4440), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U5000 ( .A(DATAI_7_), .B(n2265), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U5001 ( .A(n4415), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5002 ( .A(n4416), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5003 ( .A(n4417), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  INV_X1 U5004 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4762) );
  AOI22_X1 U5005 ( .A1(n4419), .A2(n4543), .B1(n4421), .B2(n4418), .ZN(n4420)
         );
  OAI21_X1 U5006 ( .B1(n4762), .B2(n4421), .A(n4420), .ZN(U3261) );
  INV_X1 U5007 ( .A(n4424), .ZN(n4422) );
  OAI211_X1 U5008 ( .C1(n4423), .C2(REG1_REG_0__SCAN_IN), .A(n4425), .B(n4422), 
        .ZN(n4429) );
  AOI22_X1 U5009 ( .A1(n4425), .A2(n4424), .B1(n4533), .B2(n2774), .ZN(n4427)
         );
  AOI22_X1 U5010 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4531), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4426) );
  OAI221_X1 U5011 ( .B1(IR_REG_0__SCAN_IN), .B2(n4429), .C1(n4428), .C2(n4427), 
        .A(n4426), .ZN(U3240) );
  OAI211_X1 U5012 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4431), .A(n4522), .B(n4430), 
        .ZN(n4433) );
  NAND2_X1 U5013 ( .A1(n4433), .A2(n4432), .ZN(n4434) );
  AOI21_X1 U5014 ( .B1(n4531), .B2(ADDR_REG_8__SCAN_IN), .A(n4434), .ZN(n4438)
         );
  OAI211_X1 U5015 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4436), .A(n4533), .B(n4435), 
        .ZN(n4437) );
  OAI211_X1 U5016 ( .C1(n4538), .C2(n4439), .A(n4438), .B(n4437), .ZN(U3248)
         );
  INV_X1 U5017 ( .A(n4440), .ZN(n4449) );
  OAI211_X1 U5018 ( .C1(n4443), .C2(n4442), .A(n4533), .B(n4441), .ZN(n4448)
         );
  OAI211_X1 U5019 ( .C1(n4446), .C2(n4445), .A(n4522), .B(n4444), .ZN(n4447)
         );
  OAI211_X1 U5020 ( .C1(n4538), .C2(n4449), .A(n4448), .B(n4447), .ZN(n4450)
         );
  AOI211_X1 U5021 ( .C1(n4531), .C2(ADDR_REG_9__SCAN_IN), .A(n4451), .B(n4450), 
        .ZN(n4452) );
  INV_X1 U5022 ( .A(n4452), .ZN(U3249) );
  OAI211_X1 U5023 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4454), .A(n4522), .B(n4453), .ZN(n4456) );
  NAND2_X1 U5024 ( .A1(n4456), .A2(n4455), .ZN(n4457) );
  AOI21_X1 U5025 ( .B1(n4531), .B2(ADDR_REG_10__SCAN_IN), .A(n4457), .ZN(n4461) );
  OAI211_X1 U5026 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4459), .A(n4533), .B(n4458), .ZN(n4460) );
  OAI211_X1 U5027 ( .C1(n4538), .C2(n4561), .A(n4461), .B(n4460), .ZN(U3250)
         );
  OAI211_X1 U5028 ( .C1(n4464), .C2(n4463), .A(n4533), .B(n4462), .ZN(n4469)
         );
  OAI211_X1 U5029 ( .C1(n4467), .C2(n4466), .A(n4522), .B(n4465), .ZN(n4468)
         );
  OAI211_X1 U5030 ( .C1(n4538), .C2(n4470), .A(n4469), .B(n4468), .ZN(n4471)
         );
  AOI211_X1 U5031 ( .C1(n4531), .C2(ADDR_REG_11__SCAN_IN), .A(n4472), .B(n4471), .ZN(n4473) );
  INV_X1 U5032 ( .A(n4473), .ZN(U3251) );
  OAI211_X1 U5033 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4475), .A(n4522), .B(n4474), .ZN(n4477) );
  NAND2_X1 U5034 ( .A1(n4477), .A2(n4476), .ZN(n4478) );
  AOI21_X1 U5035 ( .B1(n4531), .B2(ADDR_REG_12__SCAN_IN), .A(n4478), .ZN(n4482) );
  OAI211_X1 U5036 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4480), .A(n4533), .B(n4479), .ZN(n4481) );
  OAI211_X1 U5037 ( .C1(n4538), .C2(n4560), .A(n4482), .B(n4481), .ZN(U3252)
         );
  INV_X1 U5038 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4748) );
  AOI22_X1 U5039 ( .A1(n4483), .A2(REG2_REG_13__SCAN_IN), .B1(n4748), .B2(
        n4559), .ZN(n4486) );
  OAI21_X1 U5040 ( .B1(n4486), .B2(n4485), .A(n4522), .ZN(n4484) );
  AOI21_X1 U5041 ( .B1(n4486), .B2(n4485), .A(n4484), .ZN(n4488) );
  AOI211_X1 U5042 ( .C1(n4531), .C2(ADDR_REG_13__SCAN_IN), .A(n4488), .B(n4487), .ZN(n4493) );
  OAI211_X1 U5043 ( .C1(n4491), .C2(n4490), .A(n4533), .B(n4489), .ZN(n4492)
         );
  OAI211_X1 U5044 ( .C1(n4538), .C2(n4559), .A(n4493), .B(n4492), .ZN(U3253)
         );
  INV_X1 U5045 ( .A(n4494), .ZN(n4499) );
  AOI211_X1 U5046 ( .C1(n4497), .C2(n4496), .A(n4495), .B(n4527), .ZN(n4498)
         );
  AOI211_X1 U5047 ( .C1(n4531), .C2(ADDR_REG_14__SCAN_IN), .A(n4499), .B(n4498), .ZN(n4503) );
  OAI211_X1 U5048 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4501), .A(n4533), .B(n4500), .ZN(n4502) );
  OAI211_X1 U5049 ( .C1(n4538), .C2(n4558), .A(n4503), .B(n4502), .ZN(U3254)
         );
  AOI211_X1 U5050 ( .C1(n4506), .C2(n4505), .A(n4504), .B(n4527), .ZN(n4507)
         );
  AOI211_X1 U5051 ( .C1(n4531), .C2(ADDR_REG_15__SCAN_IN), .A(n4508), .B(n4507), .ZN(n4513) );
  OAI211_X1 U5052 ( .C1(n4511), .C2(n4510), .A(n4533), .B(n4509), .ZN(n4512)
         );
  OAI211_X1 U5053 ( .C1(n4538), .C2(n4557), .A(n4513), .B(n4512), .ZN(U3255)
         );
  INV_X1 U5054 ( .A(n4531), .ZN(n4525) );
  INV_X1 U5055 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n4766) );
  OAI21_X1 U5056 ( .B1(n4515), .B2(n3460), .A(n4514), .ZN(n4521) );
  AOI21_X1 U5057 ( .B1(REG1_REG_16__SCAN_IN), .B2(n4517), .A(n4516), .ZN(n4519) );
  OAI22_X1 U5058 ( .A1(n4519), .A2(n4518), .B1(n4555), .B2(n4538), .ZN(n4520)
         );
  AOI21_X1 U5059 ( .B1(n4522), .B2(n4521), .A(n4520), .ZN(n4524) );
  OAI211_X1 U5060 ( .C1(n4525), .C2(n4766), .A(n4524), .B(n4523), .ZN(U3256)
         );
  INV_X1 U5061 ( .A(n4526), .ZN(n4530) );
  OAI211_X1 U5062 ( .C1(n4534), .C2(n2151), .A(n4533), .B(n4532), .ZN(n4535)
         );
  OAI211_X1 U5063 ( .C1(n4538), .C2(n4537), .A(n4536), .B(n4535), .ZN(U3258)
         );
  AOI22_X1 U5064 ( .A1(n4222), .A2(REG2_REG_8__SCAN_IN), .B1(n4540), .B2(n4539), .ZN(n4547) );
  INV_X1 U5065 ( .A(n4541), .ZN(n4542) );
  AOI22_X1 U5066 ( .A1(n4545), .A2(n4544), .B1(n4543), .B2(n4542), .ZN(n4546)
         );
  OAI211_X1 U5067 ( .C1(n4222), .C2(n4548), .A(n4547), .B(n4546), .ZN(U3282)
         );
  INV_X1 U5068 ( .A(D_REG_31__SCAN_IN), .ZN(n4868) );
  NOR2_X1 U5069 ( .A1(n4550), .A2(n4868), .ZN(U3291) );
  INV_X1 U5070 ( .A(D_REG_30__SCAN_IN), .ZN(n4688) );
  NOR2_X1 U5071 ( .A1(n4550), .A2(n4688), .ZN(U3292) );
  INV_X1 U5072 ( .A(D_REG_29__SCAN_IN), .ZN(n4686) );
  NOR2_X1 U5073 ( .A1(n4550), .A2(n4686), .ZN(U3293) );
  AND2_X1 U5074 ( .A1(D_REG_28__SCAN_IN), .A2(n4549), .ZN(U3294) );
  INV_X1 U5075 ( .A(D_REG_27__SCAN_IN), .ZN(n4685) );
  NOR2_X1 U5076 ( .A1(n4550), .A2(n4685), .ZN(U3295) );
  INV_X1 U5077 ( .A(D_REG_26__SCAN_IN), .ZN(n4683) );
  NOR2_X1 U5078 ( .A1(n4550), .A2(n4683), .ZN(U3296) );
  AND2_X1 U5079 ( .A1(D_REG_25__SCAN_IN), .A2(n4549), .ZN(U3297) );
  AND2_X1 U5080 ( .A1(D_REG_24__SCAN_IN), .A2(n4549), .ZN(U3298) );
  AND2_X1 U5081 ( .A1(D_REG_23__SCAN_IN), .A2(n4549), .ZN(U3299) );
  INV_X1 U5082 ( .A(D_REG_22__SCAN_IN), .ZN(n4682) );
  NOR2_X1 U5083 ( .A1(n4550), .A2(n4682), .ZN(U3300) );
  AND2_X1 U5084 ( .A1(D_REG_21__SCAN_IN), .A2(n4549), .ZN(U3301) );
  AND2_X1 U5085 ( .A1(D_REG_20__SCAN_IN), .A2(n4549), .ZN(U3302) );
  AND2_X1 U5086 ( .A1(D_REG_19__SCAN_IN), .A2(n4549), .ZN(U3303) );
  AND2_X1 U5087 ( .A1(D_REG_18__SCAN_IN), .A2(n4549), .ZN(U3304) );
  INV_X1 U5088 ( .A(D_REG_17__SCAN_IN), .ZN(n4676) );
  NOR2_X1 U5089 ( .A1(n4550), .A2(n4676), .ZN(U3305) );
  AND2_X1 U5090 ( .A1(D_REG_16__SCAN_IN), .A2(n4549), .ZN(U3306) );
  INV_X1 U5091 ( .A(D_REG_15__SCAN_IN), .ZN(n4675) );
  NOR2_X1 U5092 ( .A1(n4550), .A2(n4675), .ZN(U3307) );
  AND2_X1 U5093 ( .A1(D_REG_14__SCAN_IN), .A2(n4549), .ZN(U3308) );
  INV_X1 U5094 ( .A(D_REG_13__SCAN_IN), .ZN(n4673) );
  NOR2_X1 U5095 ( .A1(n4550), .A2(n4673), .ZN(U3309) );
  INV_X1 U5096 ( .A(D_REG_12__SCAN_IN), .ZN(n4672) );
  NOR2_X1 U5097 ( .A1(n4550), .A2(n4672), .ZN(U3310) );
  AND2_X1 U5098 ( .A1(D_REG_11__SCAN_IN), .A2(n4549), .ZN(U3311) );
  INV_X1 U5099 ( .A(D_REG_10__SCAN_IN), .ZN(n4670) );
  NOR2_X1 U5100 ( .A1(n4550), .A2(n4670), .ZN(U3312) );
  AND2_X1 U5101 ( .A1(D_REG_9__SCAN_IN), .A2(n4549), .ZN(U3313) );
  AND2_X1 U5102 ( .A1(D_REG_8__SCAN_IN), .A2(n4549), .ZN(U3314) );
  INV_X1 U5103 ( .A(D_REG_7__SCAN_IN), .ZN(n4669) );
  NOR2_X1 U5104 ( .A1(n4550), .A2(n4669), .ZN(U3315) );
  AND2_X1 U5105 ( .A1(D_REG_6__SCAN_IN), .A2(n4549), .ZN(U3316) );
  AND2_X1 U5106 ( .A1(D_REG_5__SCAN_IN), .A2(n4549), .ZN(U3317) );
  AND2_X1 U5107 ( .A1(D_REG_4__SCAN_IN), .A2(n4549), .ZN(U3318) );
  AND2_X1 U5108 ( .A1(D_REG_3__SCAN_IN), .A2(n4549), .ZN(U3319) );
  INV_X1 U5109 ( .A(D_REG_2__SCAN_IN), .ZN(n4667) );
  NOR2_X1 U5110 ( .A1(n4550), .A2(n4667), .ZN(U3320) );
  OAI21_X1 U5111 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4551), .ZN(
        n4552) );
  INV_X1 U5112 ( .A(n4552), .ZN(U3329) );
  OAI22_X1 U5113 ( .A1(U3149), .A2(n4553), .B1(DATAI_18_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4554) );
  INV_X1 U5114 ( .A(n4554), .ZN(U3334) );
  AOI22_X1 U5115 ( .A1(STATE_REG_SCAN_IN), .A2(n4555), .B1(n2566), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5116 ( .A(DATAI_15_), .ZN(n4556) );
  AOI22_X1 U5117 ( .A1(STATE_REG_SCAN_IN), .A2(n4557), .B1(n4556), .B2(U3149), 
        .ZN(U3337) );
  AOI22_X1 U5118 ( .A1(STATE_REG_SCAN_IN), .A2(n4558), .B1(n2542), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5119 ( .A(DATAI_13_), .ZN(n4619) );
  AOI22_X1 U5120 ( .A1(STATE_REG_SCAN_IN), .A2(n4559), .B1(n4619), .B2(U3149), 
        .ZN(U3339) );
  INV_X1 U5121 ( .A(DATAI_12_), .ZN(n4622) );
  AOI22_X1 U5122 ( .A1(STATE_REG_SCAN_IN), .A2(n4560), .B1(n4622), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5123 ( .A(DATAI_10_), .ZN(n4621) );
  AOI22_X1 U5124 ( .A1(STATE_REG_SCAN_IN), .A2(n4561), .B1(n4621), .B2(U3149), 
        .ZN(U3342) );
  OAI22_X1 U5125 ( .A1(U3149), .A2(IR_REG_0__SCAN_IN), .B1(DATAI_0_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4562) );
  INV_X1 U5126 ( .A(n4562), .ZN(U3352) );
  OAI211_X1 U5127 ( .C1(n4566), .C2(n4565), .A(n4564), .B(n4563), .ZN(n4567)
         );
  INV_X1 U5128 ( .A(n4567), .ZN(n4590) );
  INV_X1 U5129 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4691) );
  AOI22_X1 U5130 ( .A1(n4589), .A2(n4590), .B1(n4691), .B2(n4587), .ZN(U3467)
         );
  INV_X1 U5131 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4568) );
  AOI22_X1 U5132 ( .A1(n4589), .A2(n4569), .B1(n4568), .B2(n4587), .ZN(U3469)
         );
  INV_X1 U5133 ( .A(n4570), .ZN(n4573) );
  INV_X1 U5134 ( .A(n4571), .ZN(n4572) );
  AOI21_X1 U5135 ( .B1(n4579), .B2(n4573), .A(n4572), .ZN(n4594) );
  AOI22_X1 U5136 ( .A1(n4574), .A2(n4591), .B1(REG0_REG_2__SCAN_IN), .B2(n4587), .ZN(n4575) );
  OAI21_X1 U5137 ( .B1(n4594), .B2(n4587), .A(n4575), .ZN(U3471) );
  INV_X1 U5138 ( .A(n4576), .ZN(n4578) );
  AOI211_X1 U5139 ( .C1(n4580), .C2(n4579), .A(n4578), .B(n4577), .ZN(n4595)
         );
  INV_X1 U5140 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4581) );
  AOI22_X1 U5141 ( .A1(n4589), .A2(n4595), .B1(n4581), .B2(n4587), .ZN(U3475)
         );
  NAND3_X1 U5142 ( .A1(n3144), .A2(n4583), .A3(n4582), .ZN(n4584) );
  INV_X1 U5143 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4588) );
  AOI22_X1 U5144 ( .A1(n4589), .A2(n4598), .B1(n4588), .B2(n4587), .ZN(U3481)
         );
  AOI22_X1 U5145 ( .A1(n4599), .A2(n4590), .B1(n2774), .B2(n4596), .ZN(U3518)
         );
  AOI22_X1 U5146 ( .A1(n4592), .A2(n4591), .B1(REG1_REG_2__SCAN_IN), .B2(n4596), .ZN(n4593) );
  OAI21_X1 U5147 ( .B1(n4594), .B2(n4596), .A(n4593), .ZN(U3520) );
  AOI22_X1 U5148 ( .A1(n4599), .A2(n4595), .B1(n4718), .B2(n4596), .ZN(U3522)
         );
  AOI22_X1 U5149 ( .A1(n4599), .A2(n4598), .B1(n4597), .B2(n4596), .ZN(U3525)
         );
  AOI22_X1 U5150 ( .A1(STATE_REG_SCAN_IN), .A2(n4600), .B1(DATAI_8_), .B2(
        U3149), .ZN(n4824) );
  INV_X1 U5151 ( .A(DATAI_29_), .ZN(n4603) );
  AOI22_X1 U5152 ( .A1(n4603), .A2(keyinput30), .B1(keyinput58), .B2(n4602), 
        .ZN(n4601) );
  OAI221_X1 U5153 ( .B1(n4603), .B2(keyinput30), .C1(n4602), .C2(keyinput58), 
        .A(n4601), .ZN(n4615) );
  AOI22_X1 U5154 ( .A1(n4606), .A2(keyinput53), .B1(keyinput95), .B2(n4605), 
        .ZN(n4604) );
  OAI221_X1 U5155 ( .B1(n4606), .B2(keyinput53), .C1(n4605), .C2(keyinput95), 
        .A(n4604), .ZN(n4614) );
  AOI22_X1 U5156 ( .A1(n4861), .A2(keyinput49), .B1(n4608), .B2(keyinput67), 
        .ZN(n4607) );
  OAI221_X1 U5157 ( .B1(n4861), .B2(keyinput49), .C1(n4608), .C2(keyinput67), 
        .A(n4607), .ZN(n4613) );
  INV_X1 U5158 ( .A(DATAI_19_), .ZN(n4610) );
  AOI22_X1 U5159 ( .A1(n4611), .A2(keyinput47), .B1(keyinput64), .B2(n4610), 
        .ZN(n4609) );
  OAI221_X1 U5160 ( .B1(n4611), .B2(keyinput47), .C1(n4610), .C2(keyinput64), 
        .A(n4609), .ZN(n4612) );
  NOR4_X1 U5161 ( .A1(n4615), .A2(n4614), .A3(n4613), .A4(n4612), .ZN(n4654)
         );
  AOI22_X1 U5162 ( .A1(n4617), .A2(keyinput43), .B1(keyinput114), .B2(n2566), 
        .ZN(n4616) );
  OAI221_X1 U5163 ( .B1(n4617), .B2(keyinput43), .C1(n2566), .C2(keyinput114), 
        .A(n4616), .ZN(n4629) );
  AOI22_X1 U5164 ( .A1(n2542), .A2(keyinput125), .B1(keyinput89), .B2(n4619), 
        .ZN(n4618) );
  OAI221_X1 U5165 ( .B1(n2542), .B2(keyinput125), .C1(n4619), .C2(keyinput89), 
        .A(n4618), .ZN(n4628) );
  AOI22_X1 U5166 ( .A1(n4622), .A2(keyinput92), .B1(keyinput121), .B2(n4621), 
        .ZN(n4620) );
  OAI221_X1 U5167 ( .B1(n4622), .B2(keyinput92), .C1(n4621), .C2(keyinput121), 
        .A(n4620), .ZN(n4627) );
  AOI22_X1 U5168 ( .A1(n4625), .A2(keyinput27), .B1(keyinput87), .B2(n4624), 
        .ZN(n4623) );
  OAI221_X1 U5169 ( .B1(n4625), .B2(keyinput27), .C1(n4624), .C2(keyinput87), 
        .A(n4623), .ZN(n4626) );
  NOR4_X1 U5170 ( .A1(n4629), .A2(n4628), .A3(n4627), .A4(n4626), .ZN(n4653)
         );
  AOI22_X1 U5171 ( .A1(n3698), .A2(keyinput75), .B1(keyinput32), .B2(n4631), 
        .ZN(n4630) );
  OAI221_X1 U5172 ( .B1(n3698), .B2(keyinput75), .C1(n4631), .C2(keyinput32), 
        .A(n4630), .ZN(n4640) );
  AOI22_X1 U5173 ( .A1(n2645), .A2(keyinput54), .B1(keyinput13), .B2(n4633), 
        .ZN(n4632) );
  OAI221_X1 U5174 ( .B1(n2645), .B2(keyinput54), .C1(n4633), .C2(keyinput13), 
        .A(n4632), .ZN(n4639) );
  XNOR2_X1 U5175 ( .A(DATAI_3_), .B(keyinput105), .ZN(n4637) );
  XNOR2_X1 U5176 ( .A(STATE_REG_SCAN_IN), .B(keyinput102), .ZN(n4636) );
  XNOR2_X1 U5177 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput127), .ZN(n4635) );
  XNOR2_X1 U5178 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput68), .ZN(n4634) );
  NAND4_X1 U5179 ( .A1(n4637), .A2(n4636), .A3(n4635), .A4(n4634), .ZN(n4638)
         );
  NOR3_X1 U5180 ( .A1(n4640), .A2(n4639), .A3(n4638), .ZN(n4652) );
  XNOR2_X1 U5181 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput112), .ZN(n4644) );
  XNOR2_X1 U5182 ( .A(REG3_REG_16__SCAN_IN), .B(keyinput72), .ZN(n4643) );
  XNOR2_X1 U5183 ( .A(REG3_REG_20__SCAN_IN), .B(keyinput45), .ZN(n4642) );
  XNOR2_X1 U5184 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput60), .ZN(n4641) );
  NAND4_X1 U5185 ( .A1(n4644), .A2(n4643), .A3(n4642), .A4(n4641), .ZN(n4650)
         );
  XNOR2_X1 U5186 ( .A(IR_REG_4__SCAN_IN), .B(keyinput108), .ZN(n4648) );
  XNOR2_X1 U5187 ( .A(IR_REG_3__SCAN_IN), .B(keyinput46), .ZN(n4647) );
  XNOR2_X1 U5188 ( .A(IR_REG_9__SCAN_IN), .B(keyinput17), .ZN(n4646) );
  XNOR2_X1 U5189 ( .A(IR_REG_8__SCAN_IN), .B(keyinput10), .ZN(n4645) );
  NAND4_X1 U5190 ( .A1(n4648), .A2(n4647), .A3(n4646), .A4(n4645), .ZN(n4649)
         );
  NOR2_X1 U5191 ( .A1(n4650), .A2(n4649), .ZN(n4651) );
  NAND4_X1 U5192 ( .A1(n4654), .A2(n4653), .A3(n4652), .A4(n4651), .ZN(n4822)
         );
  XNOR2_X1 U5193 ( .A(IR_REG_15__SCAN_IN), .B(keyinput41), .ZN(n4658) );
  XNOR2_X1 U5194 ( .A(IR_REG_11__SCAN_IN), .B(keyinput55), .ZN(n4657) );
  XNOR2_X1 U5195 ( .A(IR_REG_19__SCAN_IN), .B(keyinput86), .ZN(n4656) );
  XNOR2_X1 U5196 ( .A(IR_REG_17__SCAN_IN), .B(keyinput96), .ZN(n4655) );
  NAND4_X1 U5197 ( .A1(n4658), .A2(n4657), .A3(n4656), .A4(n4655), .ZN(n4664)
         );
  XNOR2_X1 U5198 ( .A(IR_REG_24__SCAN_IN), .B(keyinput37), .ZN(n4662) );
  XNOR2_X1 U5199 ( .A(IR_REG_22__SCAN_IN), .B(keyinput19), .ZN(n4661) );
  XNOR2_X1 U5200 ( .A(IR_REG_28__SCAN_IN), .B(keyinput85), .ZN(n4660) );
  XNOR2_X1 U5201 ( .A(IR_REG_25__SCAN_IN), .B(keyinput80), .ZN(n4659) );
  NAND4_X1 U5202 ( .A1(n4662), .A2(n4661), .A3(n4660), .A4(n4659), .ZN(n4663)
         );
  NOR2_X1 U5203 ( .A1(n4664), .A2(n4663), .ZN(n4712) );
  AOI22_X1 U5204 ( .A1(n4667), .A2(keyinput56), .B1(keyinput126), .B2(n4666), 
        .ZN(n4665) );
  OAI221_X1 U5205 ( .B1(n4667), .B2(keyinput56), .C1(n4666), .C2(keyinput126), 
        .A(n4665), .ZN(n4680) );
  AOI22_X1 U5206 ( .A1(n4670), .A2(keyinput57), .B1(n4669), .B2(keyinput98), 
        .ZN(n4668) );
  OAI221_X1 U5207 ( .B1(n4670), .B2(keyinput57), .C1(n4669), .C2(keyinput98), 
        .A(n4668), .ZN(n4679) );
  AOI22_X1 U5208 ( .A1(n4673), .A2(keyinput88), .B1(keyinput71), .B2(n4672), 
        .ZN(n4671) );
  OAI221_X1 U5209 ( .B1(n4673), .B2(keyinput88), .C1(n4672), .C2(keyinput71), 
        .A(n4671), .ZN(n4678) );
  AOI22_X1 U5210 ( .A1(n4676), .A2(keyinput40), .B1(n4675), .B2(keyinput61), 
        .ZN(n4674) );
  OAI221_X1 U5211 ( .B1(n4676), .B2(keyinput40), .C1(n4675), .C2(keyinput61), 
        .A(n4674), .ZN(n4677) );
  NOR4_X1 U5212 ( .A1(n4680), .A2(n4679), .A3(n4678), .A4(n4677), .ZN(n4711)
         );
  AOI22_X1 U5213 ( .A1(n4683), .A2(keyinput103), .B1(keyinput113), .B2(n4682), 
        .ZN(n4681) );
  OAI221_X1 U5214 ( .B1(n4683), .B2(keyinput103), .C1(n4682), .C2(keyinput113), 
        .A(n4681), .ZN(n4695) );
  AOI22_X1 U5215 ( .A1(n4686), .A2(keyinput42), .B1(n4685), .B2(keyinput20), 
        .ZN(n4684) );
  OAI221_X1 U5216 ( .B1(n4686), .B2(keyinput42), .C1(n4685), .C2(keyinput20), 
        .A(n4684), .ZN(n4694) );
  AOI22_X1 U5217 ( .A1(n4868), .A2(keyinput52), .B1(n4688), .B2(keyinput44), 
        .ZN(n4687) );
  OAI221_X1 U5218 ( .B1(n4868), .B2(keyinput52), .C1(n4688), .C2(keyinput44), 
        .A(n4687), .ZN(n4693) );
  INV_X1 U5219 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4690) );
  AOI22_X1 U5220 ( .A1(n4691), .A2(keyinput35), .B1(n4690), .B2(keyinput1), 
        .ZN(n4689) );
  OAI221_X1 U5221 ( .B1(n4691), .B2(keyinput35), .C1(n4690), .C2(keyinput1), 
        .A(n4689), .ZN(n4692) );
  NOR4_X1 U5222 ( .A1(n4695), .A2(n4694), .A3(n4693), .A4(n4692), .ZN(n4710)
         );
  INV_X1 U5223 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4697) );
  AOI22_X1 U5224 ( .A1(n4697), .A2(keyinput117), .B1(n3253), .B2(keyinput97), 
        .ZN(n4696) );
  OAI221_X1 U5225 ( .B1(n4697), .B2(keyinput117), .C1(n3253), .C2(keyinput97), 
        .A(n4696), .ZN(n4708) );
  AOI22_X1 U5226 ( .A1(n4700), .A2(keyinput39), .B1(keyinput83), .B2(n4699), 
        .ZN(n4698) );
  OAI221_X1 U5227 ( .B1(n4700), .B2(keyinput39), .C1(n4699), .C2(keyinput83), 
        .A(n4698), .ZN(n4707) );
  AOI22_X1 U5228 ( .A1(n3468), .A2(keyinput94), .B1(n4399), .B2(keyinput15), 
        .ZN(n4701) );
  OAI221_X1 U5229 ( .B1(n3468), .B2(keyinput94), .C1(n4399), .C2(keyinput15), 
        .A(n4701), .ZN(n4706) );
  INV_X1 U5230 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4704) );
  INV_X1 U5231 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4703) );
  AOI22_X1 U5232 ( .A1(n4704), .A2(keyinput82), .B1(n4703), .B2(keyinput50), 
        .ZN(n4702) );
  OAI221_X1 U5233 ( .B1(n4704), .B2(keyinput82), .C1(n4703), .C2(keyinput50), 
        .A(n4702), .ZN(n4705) );
  NOR4_X1 U5234 ( .A1(n4708), .A2(n4707), .A3(n4706), .A4(n4705), .ZN(n4709)
         );
  NAND4_X1 U5235 ( .A1(n4712), .A2(n4711), .A3(n4710), .A4(n4709), .ZN(n4821)
         );
  INV_X1 U5236 ( .A(REG1_REG_5__SCAN_IN), .ZN(n4714) );
  AOI22_X1 U5237 ( .A1(n4714), .A2(keyinput65), .B1(n4867), .B2(keyinput6), 
        .ZN(n4713) );
  OAI221_X1 U5238 ( .B1(n4714), .B2(keyinput65), .C1(n4867), .C2(keyinput6), 
        .A(n4713), .ZN(n4725) );
  INV_X1 U5239 ( .A(REG0_REG_29__SCAN_IN), .ZN(n4716) );
  AOI22_X1 U5240 ( .A1(n4371), .A2(keyinput18), .B1(n4716), .B2(keyinput116), 
        .ZN(n4715) );
  OAI221_X1 U5241 ( .B1(n4371), .B2(keyinput18), .C1(n4716), .C2(keyinput116), 
        .A(n4715), .ZN(n4724) );
  XOR2_X1 U5242 ( .A(n4717), .B(keyinput99), .Z(n4722) );
  XOR2_X1 U5243 ( .A(n4718), .B(keyinput70), .Z(n4721) );
  XNOR2_X1 U5244 ( .A(REG1_REG_1__SCAN_IN), .B(keyinput90), .ZN(n4720) );
  XNOR2_X1 U5245 ( .A(REG1_REG_2__SCAN_IN), .B(keyinput100), .ZN(n4719) );
  NAND4_X1 U5246 ( .A1(n4722), .A2(n4721), .A3(n4720), .A4(n4719), .ZN(n4723)
         );
  NOR3_X1 U5247 ( .A1(n4725), .A2(n4724), .A3(n4723), .ZN(n4760) );
  AOI22_X1 U5248 ( .A1(n3416), .A2(keyinput77), .B1(keyinput124), .B2(n4727), 
        .ZN(n4726) );
  OAI221_X1 U5249 ( .B1(n3416), .B2(keyinput77), .C1(n4727), .C2(keyinput124), 
        .A(n4726), .ZN(n4736) );
  AOI22_X1 U5250 ( .A1(n3466), .A2(keyinput84), .B1(n4328), .B2(keyinput118), 
        .ZN(n4728) );
  OAI221_X1 U5251 ( .B1(n3466), .B2(keyinput84), .C1(n4328), .C2(keyinput118), 
        .A(n4728), .ZN(n4735) );
  AOI22_X1 U5252 ( .A1(n4314), .A2(keyinput109), .B1(keyinput91), .B2(n4730), 
        .ZN(n4729) );
  OAI221_X1 U5253 ( .B1(n4314), .B2(keyinput109), .C1(n4730), .C2(keyinput91), 
        .A(n4729), .ZN(n4734) );
  AOI22_X1 U5254 ( .A1(n4300), .A2(keyinput14), .B1(n4732), .B2(keyinput38), 
        .ZN(n4731) );
  OAI221_X1 U5255 ( .B1(n4300), .B2(keyinput14), .C1(n4732), .C2(keyinput38), 
        .A(n4731), .ZN(n4733) );
  NOR4_X1 U5256 ( .A1(n4736), .A2(n4735), .A3(n4734), .A4(n4733), .ZN(n4759)
         );
  AOI22_X1 U5257 ( .A1(n2761), .A2(keyinput93), .B1(keyinput23), .B2(n2717), 
        .ZN(n4737) );
  OAI221_X1 U5258 ( .B1(n2761), .B2(keyinput93), .C1(n2717), .C2(keyinput23), 
        .A(n4737), .ZN(n4745) );
  AOI22_X1 U5259 ( .A1(n2784), .A2(keyinput123), .B1(keyinput115), .B2(n4266), 
        .ZN(n4738) );
  OAI221_X1 U5260 ( .B1(n2784), .B2(keyinput123), .C1(n4266), .C2(keyinput115), 
        .A(n4738), .ZN(n4744) );
  AOI22_X1 U5261 ( .A1(n2252), .A2(keyinput21), .B1(keyinput120), .B2(n3053), 
        .ZN(n4739) );
  OAI221_X1 U5262 ( .B1(n2252), .B2(keyinput21), .C1(n3053), .C2(keyinput120), 
        .A(n4739), .ZN(n4743) );
  INV_X1 U5263 ( .A(REG2_REG_10__SCAN_IN), .ZN(n4741) );
  AOI22_X1 U5264 ( .A1(n3191), .A2(keyinput16), .B1(n4741), .B2(keyinput101), 
        .ZN(n4740) );
  OAI221_X1 U5265 ( .B1(n3191), .B2(keyinput16), .C1(n4741), .C2(keyinput101), 
        .A(n4740), .ZN(n4742) );
  NOR4_X1 U5266 ( .A1(n4745), .A2(n4744), .A3(n4743), .A4(n4742), .ZN(n4758)
         );
  AOI22_X1 U5267 ( .A1(n4748), .A2(keyinput62), .B1(keyinput119), .B2(n4747), 
        .ZN(n4746) );
  OAI221_X1 U5268 ( .B1(n4748), .B2(keyinput62), .C1(n4747), .C2(keyinput119), 
        .A(n4746), .ZN(n4756) );
  AOI22_X1 U5269 ( .A1(n4862), .A2(keyinput73), .B1(keyinput106), .B2(n3460), 
        .ZN(n4749) );
  OAI221_X1 U5270 ( .B1(n4862), .B2(keyinput73), .C1(n3460), .C2(keyinput106), 
        .A(n4749), .ZN(n4755) );
  INV_X1 U5271 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4751) );
  AOI22_X1 U5272 ( .A1(n4163), .A2(keyinput4), .B1(keyinput36), .B2(n4751), 
        .ZN(n4750) );
  OAI221_X1 U5273 ( .B1(n4163), .B2(keyinput4), .C1(n4751), .C2(keyinput36), 
        .A(n4750), .ZN(n4754) );
  INV_X1 U5274 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4863) );
  AOI22_X1 U5275 ( .A1(n4863), .A2(keyinput2), .B1(n4065), .B2(keyinput76), 
        .ZN(n4752) );
  OAI221_X1 U5276 ( .B1(n4863), .B2(keyinput2), .C1(n4065), .C2(keyinput76), 
        .A(n4752), .ZN(n4753) );
  NOR4_X1 U5277 ( .A1(n4756), .A2(n4755), .A3(n4754), .A4(n4753), .ZN(n4757)
         );
  NAND4_X1 U5278 ( .A1(n4760), .A2(n4759), .A3(n4758), .A4(n4757), .ZN(n4820)
         );
  INV_X1 U5279 ( .A(ADDR_REG_19__SCAN_IN), .ZN(n4763) );
  AOI22_X1 U5280 ( .A1(n4763), .A2(keyinput12), .B1(n4762), .B2(keyinput25), 
        .ZN(n4761) );
  OAI221_X1 U5281 ( .B1(n4763), .B2(keyinput12), .C1(n4762), .C2(keyinput25), 
        .A(n4761), .ZN(n4774) );
  INV_X1 U5282 ( .A(ADDR_REG_18__SCAN_IN), .ZN(n4765) );
  AOI22_X1 U5283 ( .A1(n4766), .A2(keyinput81), .B1(n4765), .B2(keyinput26), 
        .ZN(n4764) );
  OAI221_X1 U5284 ( .B1(n4766), .B2(keyinput81), .C1(n4765), .C2(keyinput26), 
        .A(n4764), .ZN(n4773) );
  INV_X1 U5285 ( .A(ADDR_REG_15__SCAN_IN), .ZN(n4835) );
  INV_X1 U5286 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n4768) );
  AOI22_X1 U5287 ( .A1(n4835), .A2(keyinput28), .B1(keyinput3), .B2(n4768), 
        .ZN(n4767) );
  OAI221_X1 U5288 ( .B1(n4835), .B2(keyinput28), .C1(n4768), .C2(keyinput3), 
        .A(n4767), .ZN(n4772) );
  INV_X1 U5289 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n4860) );
  INV_X1 U5290 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n4770) );
  AOI22_X1 U5291 ( .A1(n4860), .A2(keyinput59), .B1(keyinput104), .B2(n4770), 
        .ZN(n4769) );
  OAI221_X1 U5292 ( .B1(n4860), .B2(keyinput59), .C1(n4770), .C2(keyinput104), 
        .A(n4769), .ZN(n4771) );
  NOR4_X1 U5293 ( .A1(n4774), .A2(n4773), .A3(n4772), .A4(n4771), .ZN(n4818)
         );
  INV_X1 U5294 ( .A(ADDR_REG_1__SCAN_IN), .ZN(n4777) );
  INV_X1 U5295 ( .A(ADDR_REG_2__SCAN_IN), .ZN(n4776) );
  AOI22_X1 U5296 ( .A1(n4777), .A2(keyinput48), .B1(n4776), .B2(keyinput8), 
        .ZN(n4775) );
  OAI221_X1 U5297 ( .B1(n4777), .B2(keyinput48), .C1(n4776), .C2(keyinput8), 
        .A(n4775), .ZN(n4785) );
  INV_X1 U5298 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n4779) );
  AOI22_X1 U5299 ( .A1(n4779), .A2(keyinput5), .B1(n4834), .B2(keyinput29), 
        .ZN(n4778) );
  OAI221_X1 U5300 ( .B1(n4779), .B2(keyinput5), .C1(n4834), .C2(keyinput29), 
        .A(n4778), .ZN(n4784) );
  AOI22_X1 U5301 ( .A1(n4832), .A2(keyinput110), .B1(n4833), .B2(keyinput31), 
        .ZN(n4780) );
  OAI221_X1 U5302 ( .B1(n4832), .B2(keyinput110), .C1(n4833), .C2(keyinput31), 
        .A(n4780), .ZN(n4783) );
  AOI22_X1 U5303 ( .A1(n4831), .A2(keyinput22), .B1(keyinput122), .B2(n4829), 
        .ZN(n4781) );
  OAI221_X1 U5304 ( .B1(n4831), .B2(keyinput22), .C1(n4829), .C2(keyinput122), 
        .A(n4781), .ZN(n4782) );
  NOR4_X1 U5305 ( .A1(n4785), .A2(n4784), .A3(n4783), .A4(n4782), .ZN(n4817)
         );
  AOI22_X1 U5306 ( .A1(n4787), .A2(keyinput69), .B1(keyinput11), .B2(n4830), 
        .ZN(n4786) );
  OAI221_X1 U5307 ( .B1(n4787), .B2(keyinput69), .C1(n4830), .C2(keyinput11), 
        .A(n4786), .ZN(n4799) );
  AOI22_X1 U5308 ( .A1(n4789), .A2(keyinput107), .B1(keyinput111), .B2(n4828), 
        .ZN(n4788) );
  OAI221_X1 U5309 ( .B1(n4789), .B2(keyinput107), .C1(n4828), .C2(keyinput111), 
        .A(n4788), .ZN(n4798) );
  AOI22_X1 U5310 ( .A1(n4792), .A2(keyinput51), .B1(keyinput0), .B2(n4791), 
        .ZN(n4790) );
  OAI221_X1 U5311 ( .B1(n4792), .B2(keyinput51), .C1(n4791), .C2(keyinput0), 
        .A(n4790), .ZN(n4797) );
  AOI22_X1 U5312 ( .A1(n4795), .A2(keyinput78), .B1(n4794), .B2(keyinput63), 
        .ZN(n4793) );
  OAI221_X1 U5313 ( .B1(n4795), .B2(keyinput78), .C1(n4794), .C2(keyinput63), 
        .A(n4793), .ZN(n4796) );
  NOR4_X1 U5314 ( .A1(n4799), .A2(n4798), .A3(n4797), .A4(n4796), .ZN(n4816)
         );
  INV_X1 U5315 ( .A(REG3_REG_2__SCAN_IN), .ZN(n4802) );
  AOI22_X1 U5316 ( .A1(n4802), .A2(keyinput9), .B1(keyinput79), .B2(n4801), 
        .ZN(n4800) );
  OAI221_X1 U5317 ( .B1(n4802), .B2(keyinput9), .C1(n4801), .C2(keyinput79), 
        .A(n4800), .ZN(n4814) );
  AOI22_X1 U5318 ( .A1(n4805), .A2(keyinput66), .B1(keyinput34), .B2(n4804), 
        .ZN(n4803) );
  OAI221_X1 U5319 ( .B1(n4805), .B2(keyinput66), .C1(n4804), .C2(keyinput34), 
        .A(n4803), .ZN(n4813) );
  AOI22_X1 U5320 ( .A1(n4808), .A2(keyinput24), .B1(keyinput7), .B2(n4807), 
        .ZN(n4806) );
  OAI221_X1 U5321 ( .B1(n4808), .B2(keyinput24), .C1(n4807), .C2(keyinput7), 
        .A(n4806), .ZN(n4812) );
  XNOR2_X1 U5322 ( .A(IR_REG_2__SCAN_IN), .B(keyinput33), .ZN(n4810) );
  XNOR2_X1 U5323 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput74), .ZN(n4809) );
  NAND2_X1 U5324 ( .A1(n4810), .A2(n4809), .ZN(n4811) );
  NOR4_X1 U5325 ( .A1(n4814), .A2(n4813), .A3(n4812), .A4(n4811), .ZN(n4815)
         );
  NAND4_X1 U5326 ( .A1(n4818), .A2(n4817), .A3(n4816), .A4(n4815), .ZN(n4819)
         );
  NOR4_X1 U5327 ( .A1(n4822), .A2(n4821), .A3(n4820), .A4(n4819), .ZN(n4823)
         );
  XNOR2_X1 U5328 ( .A(n4824), .B(n4823), .ZN(n4884) );
  AND4_X1 U5329 ( .A1(n4602), .A2(n4825), .A3(STATE_REG_SCAN_IN), .A4(
        IR_REG_3__SCAN_IN), .ZN(n4827) );
  NAND4_X1 U5330 ( .A1(n4827), .A2(IR_REG_8__SCAN_IN), .A3(
        ADDR_REG_19__SCAN_IN), .A4(n4826), .ZN(n4843) );
  NAND4_X1 U5331 ( .A1(n4831), .A2(n4830), .A3(n4829), .A4(n4828), .ZN(n4842)
         );
  NAND4_X1 U5332 ( .A1(n4835), .A2(n4834), .A3(n4833), .A4(n4832), .ZN(n4841)
         );
  NOR4_X1 U5333 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_0__SCAN_IN), .A3(
        REG0_REG_30__SCAN_IN), .A4(REG1_REG_31__SCAN_IN), .ZN(n4839) );
  NOR4_X1 U5334 ( .A1(REG3_REG_10__SCAN_IN), .A2(ADDR_REG_18__SCAN_IN), .A3(
        DATAO_REG_23__SCAN_IN), .A4(DATAO_REG_25__SCAN_IN), .ZN(n4838) );
  NOR4_X1 U5335 ( .A1(IR_REG_22__SCAN_IN), .A2(REG3_REG_19__SCAN_IN), .A3(
        REG1_REG_21__SCAN_IN), .A4(REG0_REG_19__SCAN_IN), .ZN(n4837) );
  NOR4_X1 U5336 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG0_REG_27__SCAN_IN), .A3(
        REG1_REG_25__SCAN_IN), .A4(REG1_REG_24__SCAN_IN), .ZN(n4836) );
  NAND4_X1 U5337 ( .A1(n4839), .A2(n4838), .A3(n4837), .A4(n4836), .ZN(n4840)
         );
  NOR4_X1 U5338 ( .A1(n4843), .A2(n4842), .A3(n4841), .A4(n4840), .ZN(n4882)
         );
  NAND4_X1 U5339 ( .A1(D_REG_7__SCAN_IN), .A2(REG1_REG_26__SCAN_IN), .A3(
        REG1_REG_23__SCAN_IN), .A4(REG0_REG_20__SCAN_IN), .ZN(n4847) );
  NAND4_X1 U5340 ( .A1(REG1_REG_29__SCAN_IN), .A2(REG0_REG_29__SCAN_IN), .A3(
        REG0_REG_23__SCAN_IN), .A4(DATAO_REG_26__SCAN_IN), .ZN(n4846) );
  NAND4_X1 U5341 ( .A1(IR_REG_19__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_30__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n4845) );
  NAND4_X1 U5342 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n4844) );
  NOR4_X1 U5343 ( .A1(n4847), .A2(n4846), .A3(n4845), .A4(n4844), .ZN(n4881)
         );
  NAND4_X1 U5344 ( .A1(IR_REG_24__SCAN_IN), .A2(REG3_REG_16__SCAN_IN), .A3(
        REG3_REG_12__SCAN_IN), .A4(DATAO_REG_18__SCAN_IN), .ZN(n4851) );
  NAND4_X1 U5345 ( .A1(IR_REG_25__SCAN_IN), .A2(REG3_REG_8__SCAN_IN), .A3(
        DATAI_16_), .A4(DATAI_13_), .ZN(n4850) );
  NAND4_X1 U5346 ( .A1(REG1_REG_30__SCAN_IN), .A2(DATAO_REG_27__SCAN_IN), .A3(
        DATAO_REG_29__SCAN_IN), .A4(DATAO_REG_30__SCAN_IN), .ZN(n4849) );
  NAND4_X1 U5347 ( .A1(DATAI_29_), .A2(ADDR_REG_13__SCAN_IN), .A3(
        DATAO_REG_10__SCAN_IN), .A4(DATAO_REG_31__SCAN_IN), .ZN(n4848) );
  NOR4_X1 U5348 ( .A1(n4851), .A2(n4850), .A3(n4849), .A4(n4848), .ZN(n4880)
         );
  NOR4_X1 U5349 ( .A1(REG3_REG_11__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        DATAI_17_), .A4(ADDR_REG_1__SCAN_IN), .ZN(n4855) );
  NOR4_X1 U5350 ( .A1(REG1_REG_4__SCAN_IN), .A2(REG2_REG_4__SCAN_IN), .A3(
        ADDR_REG_2__SCAN_IN), .A4(ADDR_REG_5__SCAN_IN), .ZN(n4854) );
  NOR4_X1 U5351 ( .A1(REG3_REG_28__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .A3(
        REG3_REG_20__SCAN_IN), .A4(REG2_REG_30__SCAN_IN), .ZN(n4853) );
  NOR4_X1 U5352 ( .A1(REG2_REG_23__SCAN_IN), .A2(DATAI_22_), .A3(
        REG2_REG_21__SCAN_IN), .A4(REG2_REG_16__SCAN_IN), .ZN(n4852) );
  NAND4_X1 U5353 ( .A1(n4855), .A2(n4854), .A3(n4853), .A4(n4852), .ZN(n4878)
         );
  NOR4_X1 U5354 ( .A1(DATAI_14_), .A2(DATAI_12_), .A3(REG0_REG_12__SCAN_IN), 
        .A4(DATAI_10_), .ZN(n4859) );
  NOR4_X1 U5355 ( .A1(IR_REG_9__SCAN_IN), .A2(DATAI_5_), .A3(
        REG0_REG_5__SCAN_IN), .A4(DATAI_3_), .ZN(n4858) );
  NOR4_X1 U5356 ( .A1(REG1_REG_13__SCAN_IN), .A2(REG2_REG_11__SCAN_IN), .A3(
        REG2_REG_10__SCAN_IN), .A4(REG2_REG_6__SCAN_IN), .ZN(n4857) );
  NOR4_X1 U5357 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .A3(
        REG0_REG_15__SCAN_IN), .A4(REG1_REG_2__SCAN_IN), .ZN(n4856) );
  NAND4_X1 U5358 ( .A1(n4859), .A2(n4858), .A3(n4857), .A4(n4856), .ZN(n4877)
         );
  NOR4_X1 U5359 ( .A1(n4863), .A2(n4862), .A3(n4861), .A4(n4860), .ZN(n4864)
         );
  NAND4_X1 U5360 ( .A1(n4865), .A2(REG2_REG_29__SCAN_IN), .A3(
        REG3_REG_0__SCAN_IN), .A4(n4864), .ZN(n4876) );
  NAND4_X1 U5361 ( .A1(REG1_REG_10__SCAN_IN), .A2(DATAI_7_), .A3(
        REG0_REG_2__SCAN_IN), .A4(REG0_REG_0__SCAN_IN), .ZN(n4866) );
  NOR3_X1 U5362 ( .A1(n4868), .A2(n4867), .A3(n4866), .ZN(n4874) );
  NAND4_X1 U5363 ( .A1(REG1_REG_15__SCAN_IN), .A2(REG2_REG_2__SCAN_IN), .A3(
        REG1_REG_1__SCAN_IN), .A4(REG2_REG_1__SCAN_IN), .ZN(n4872) );
  NAND4_X1 U5364 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_28__SCAN_IN), .A3(
        REG0_REG_10__SCAN_IN), .A4(REG1_REG_5__SCAN_IN), .ZN(n4871) );
  NAND4_X1 U5365 ( .A1(DATAI_28_), .A2(DATAI_27_), .A3(DATAI_26_), .A4(
        DATAI_19_), .ZN(n4870) );
  NAND4_X1 U5366 ( .A1(REG2_REG_13__SCAN_IN), .A2(REG3_REG_2__SCAN_IN), .A3(
        ADDR_REG_16__SCAN_IN), .A4(ADDR_REG_0__SCAN_IN), .ZN(n4869) );
  NOR4_X1 U5367 ( .A1(n4872), .A2(n4871), .A3(n4870), .A4(n4869), .ZN(n4873)
         );
  NAND4_X1 U5368 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG0_REG_9__SCAN_IN), .A3(
        n4874), .A4(n4873), .ZN(n4875) );
  NOR4_X1 U5369 ( .A1(n4878), .A2(n4877), .A3(n4876), .A4(n4875), .ZN(n4879)
         );
  NAND4_X1 U5370 ( .A1(n4882), .A2(n4881), .A3(n4880), .A4(n4879), .ZN(n4883)
         );
  XNOR2_X1 U5371 ( .A(n4884), .B(n4883), .ZN(U3344) );
  CLKBUF_X2 U2382 ( .A(n3628), .Z(n2132) );
  CLKBUF_X1 U2379 ( .A(n3628), .Z(n2133) );
endmodule

