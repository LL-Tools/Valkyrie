

module b20_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7824, n7825, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10858;

  INV_X2 U5006 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5007 ( .A(n8890), .ZN(n9041) );
  NAND2_X1 U5008 ( .A1(n8034), .A2(n8033), .ZN(n9788) );
  NAND2_X1 U5009 ( .A1(n8851), .A2(n8850), .ZN(n8849) );
  OR2_X1 U5010 ( .A1(n5545), .A2(n7610), .ZN(n5544) );
  INV_X1 U5011 ( .A(n9962), .ZN(n10720) );
  CLKBUF_X2 U5013 ( .A(n8218), .Z(n9705) );
  INV_X1 U5014 ( .A(n6306), .ZN(n6016) );
  INV_X2 U5015 ( .A(n6046), .ZN(n8473) );
  CLKBUF_X2 U5016 ( .A(n6835), .Z(n8324) );
  AND2_X1 U5017 ( .A1(n8690), .A2(n6431), .ZN(n6813) );
  CLKBUF_X1 U5019 ( .A(n10842), .Z(n4942) );
  NOR2_X1 U5020 ( .A1(n10731), .A2(n9882), .ZN(n10842) );
  INV_X1 U5021 ( .A(n6751), .ZN(n8739) );
  INV_X2 U5022 ( .A(n8655), .ZN(n8610) );
  INV_X1 U5023 ( .A(n7750), .ZN(n5323) );
  NAND2_X1 U5024 ( .A1(n10720), .A2(n8204), .ZN(n10716) );
  OR2_X1 U5025 ( .A1(n8750), .A2(n8654), .ZN(n6274) );
  NAND2_X1 U5026 ( .A1(n6268), .A2(n8651), .ZN(n8650) );
  NAND2_X1 U5027 ( .A1(n8675), .A2(n9011), .ZN(n6747) );
  INV_X1 U5028 ( .A(n10297), .ZN(n9638) );
  NAND2_X1 U5029 ( .A1(n8369), .A2(n8368), .ZN(n9647) );
  CLKBUF_X3 U5030 ( .A(n7274), .Z(n9700) );
  INV_X1 U5031 ( .A(n7502), .ZN(n10660) );
  INV_X2 U5032 ( .A(n5674), .ZN(n5575) );
  AOI22_X1 U5033 ( .A1(P2_REG1_REG_1__SCAN_IN), .A2(n5459), .B1(n5460), .B2(
        n5699), .ZN(n5461) );
  CLKBUF_X2 U5034 ( .A(n5575), .Z(n4945) );
  NAND4_X1 U5035 ( .A1(n7524), .A2(n7523), .A3(n7522), .A4(n7521), .ZN(n10746)
         );
  INV_X2 U5036 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  OR2_X1 U5037 ( .A1(n6316), .A2(n6315), .ZN(n4943) );
  INV_X1 U5038 ( .A(n7012), .ZN(n4946) );
  NAND2_X1 U5039 ( .A1(n8447), .A2(n6828), .ZN(n7012) );
  AOI21_X2 U5040 ( .B1(n8209), .B2(n9686), .A(n8208), .ZN(n10247) );
  OAI21_X2 U5041 ( .B1(n5398), .B2(n5397), .A(n8124), .ZN(n8209) );
  OAI21_X2 U5042 ( .B1(n10233), .B2(n8315), .A(n9721), .ZN(n10224) );
  OAI21_X2 U5043 ( .B1(n10250), .B2(n8314), .A(n9922), .ZN(n10233) );
  XNOR2_X2 U5044 ( .A(n6388), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6607) );
  OAI22_X2 U5045 ( .A1(n7892), .A2(n7891), .B1(n7890), .B2(n7889), .ZN(n7947)
         );
  AOI21_X2 U5046 ( .B1(n7829), .B2(n7828), .A(n7827), .ZN(n7892) );
  AOI21_X2 U5047 ( .B1(n10169), .B2(n10168), .A(n8318), .ZN(n10151) );
  NAND2_X2 U5048 ( .A1(n5450), .A2(n9855), .ZN(n10169) );
  INV_X1 U5049 ( .A(n10746), .ZN(n8201) );
  OAI21_X1 U5050 ( .B1(n8432), .B2(n8433), .A(n5316), .ZN(n9636) );
  OAI21_X1 U5051 ( .B1(n9023), .B2(n7539), .A(n5052), .ZN(n9015) );
  NAND2_X1 U5052 ( .A1(n8734), .A2(n8733), .ZN(n8786) );
  OR2_X1 U5053 ( .A1(n9042), .A2(n6259), .ZN(n6262) );
  AND2_X1 U5054 ( .A1(n10278), .A2(n5259), .ZN(n5258) );
  NAND2_X1 U5055 ( .A1(n9647), .A2(n5340), .ZN(n5338) );
  NAND2_X1 U5056 ( .A1(n8770), .A2(n8715), .ZN(n8824) );
  INV_X1 U5057 ( .A(n10276), .ZN(n5257) );
  NAND2_X1 U5058 ( .A1(n8710), .A2(n4951), .ZN(n8770) );
  AND2_X1 U5059 ( .A1(n7990), .A2(n7983), .ZN(n7988) );
  NAND2_X1 U5060 ( .A1(n5355), .A2(n7841), .ZN(n7977) );
  OAI21_X1 U5061 ( .B1(n10809), .B2(n10826), .A(n8031), .ZN(n10815) );
  NAND2_X1 U5062 ( .A1(n5714), .A2(n5713), .ZN(n9052) );
  NAND2_X1 U5063 ( .A1(n7195), .A2(n7194), .ZN(n5353) );
  NAND2_X1 U5064 ( .A1(n7633), .A2(n7632), .ZN(n10790) );
  NAND2_X1 U5065 ( .A1(n7510), .A2(n7509), .ZN(n8204) );
  NAND2_X1 U5066 ( .A1(n7546), .A2(n7545), .ZN(n10748) );
  NAND2_X1 U5067 ( .A1(n5866), .A2(n5865), .ZN(n7626) );
  NAND2_X1 U5068 ( .A1(n5835), .A2(n5834), .ZN(n7405) );
  NAND2_X2 U5069 ( .A1(n10684), .A2(n9739), .ZN(n10674) );
  XNOR2_X1 U5070 ( .A(n5216), .B(n5846), .ZN(n7555) );
  INV_X1 U5071 ( .A(n10698), .ZN(n10680) );
  OR2_X1 U5072 ( .A1(n9964), .A2(n7343), .ZN(n9899) );
  NAND2_X2 U5073 ( .A1(n7017), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9654) );
  NAND2_X1 U5074 ( .A1(n9729), .A2(n9894), .ZN(n7130) );
  INV_X1 U5075 ( .A(n7061), .ZN(n10636) );
  NAND2_X1 U5076 ( .A1(n5791), .A2(n5790), .ZN(n7061) );
  OR2_X1 U5077 ( .A1(n9965), .A2(n7412), .ZN(n9729) );
  NAND2_X1 U5078 ( .A1(n5824), .A2(n5823), .ZN(n5822) );
  INV_X2 U5079 ( .A(n8448), .ZN(n8438) );
  INV_X2 U5080 ( .A(n6829), .ZN(n8460) );
  OR2_X1 U5081 ( .A1(n6746), .A2(n6745), .ZN(n6750) );
  INV_X1 U5082 ( .A(n6806), .ZN(n8448) );
  CLKBUF_X2 U5083 ( .A(n6968), .Z(n10591) );
  NAND4_X1 U5084 ( .A1(n7210), .A2(n7209), .A3(n7208), .A4(n7207), .ZN(n9963)
         );
  AND2_X1 U5085 ( .A1(n6727), .A2(n6611), .ZN(n6806) );
  BUF_X2 U5086 ( .A(n6813), .Z(n7274) );
  INV_X1 U5087 ( .A(n10592), .ZN(n9890) );
  NAND2_X1 U5088 ( .A1(n6410), .A2(n6337), .ZN(n6727) );
  XNOR2_X1 U5089 ( .A(n6107), .B(n6106), .ZN(n6746) );
  NAND2_X1 U5090 ( .A1(n6192), .A2(n6191), .ZN(n7866) );
  XNOR2_X1 U5091 ( .A(n6189), .B(n6188), .ZN(n7868) );
  AND2_X1 U5092 ( .A1(n6327), .A2(n6334), .ZN(n6410) );
  NAND2_X1 U5093 ( .A1(n5529), .A2(n5528), .ZN(n6107) );
  NAND2_X1 U5094 ( .A1(n6332), .A2(n6331), .ZN(n7882) );
  INV_X2 U5095 ( .A(n5760), .ZN(n6252) );
  INV_X1 U5096 ( .A(n6431), .ZN(n10402) );
  MUX2_X1 U5097 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6330), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n6332) );
  MUX2_X1 U5098 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6321), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n6327) );
  XNOR2_X1 U5099 ( .A(n6105), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9011) );
  AND2_X1 U5100 ( .A1(n6391), .A2(n6390), .ZN(n9881) );
  INV_X4 U5101 ( .A(n6797), .ZN(n7007) );
  NAND2_X1 U5102 ( .A1(n8471), .A2(n9262), .ZN(n5760) );
  NAND2_X1 U5103 ( .A1(n5699), .A2(n5698), .ZN(n5930) );
  NAND2_X2 U5104 ( .A1(n5700), .A2(n9262), .ZN(n8182) );
  MUX2_X1 U5105 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6604), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n6606) );
  NAND2_X1 U5106 ( .A1(n6186), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6195) );
  NOR2_X1 U5107 ( .A1(n6605), .A2(n6319), .ZN(n6328) );
  NAND2_X1 U5108 ( .A1(n6605), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6602) );
  AND2_X1 U5109 ( .A1(n6394), .A2(n6426), .ZN(n6429) );
  NOR2_X1 U5110 ( .A1(n6334), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U5111 ( .A1(n6326), .A2(n6318), .ZN(n6605) );
  INV_X2 U5112 ( .A(n7819), .ZN(n4944) );
  AND2_X1 U5113 ( .A1(n5534), .A2(n5533), .ZN(n6003) );
  NOR2_X1 U5114 ( .A1(n5860), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n6183) );
  NOR2_X1 U5115 ( .A1(n4949), .A2(n5940), .ZN(n5671) );
  NAND2_X1 U5116 ( .A1(n5154), .A2(n5152), .ZN(n5674) );
  NOR2_X1 U5117 ( .A1(n6361), .A2(n5453), .ZN(n6379) );
  NAND2_X1 U5118 ( .A1(n6173), .A2(n5537), .ZN(n5536) );
  OAI21_X1 U5119 ( .B1(P1_ADDR_REG_19__SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        n5153), .ZN(n5152) );
  AND4_X1 U5120 ( .A1(n5518), .A2(n5662), .A3(n6174), .A4(n5282), .ZN(n5278)
         );
  AND3_X1 U5121 ( .A1(n5832), .A2(n5281), .A3(n5280), .ZN(n5279) );
  INV_X1 U5122 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6309) );
  NOR2_X1 U5123 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n6308) );
  INV_X1 U5124 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n6472) );
  NOR2_X1 U5125 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n6312) );
  INV_X1 U5126 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5456) );
  INV_X1 U5127 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6376) );
  INV_X1 U5128 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5153) );
  INV_X1 U5129 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n7048) );
  INV_X1 U5130 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6473) );
  INV_X1 U5131 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5662) );
  INV_X1 U5132 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5282) );
  INV_X1 U5133 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5285) );
  INV_X1 U5134 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5517) );
  INV_X1 U5135 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5518) );
  NOR2_X2 U5136 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n6175) );
  NOR2_X2 U5137 ( .A1(n10151), .A2(n10153), .ZN(n10150) );
  NOR2_X2 U5138 ( .A1(n7339), .A2(n10641), .ZN(n7490) );
  AOI22_X2 U5139 ( .A1(n7575), .A2(n7574), .B1(n10720), .B2(n5271), .ZN(n10712) );
  NAND2_X2 U5140 ( .A1(n7506), .A2(n7505), .ZN(n7575) );
  INV_X4 U5141 ( .A(n8739), .ZN(n8744) );
  INV_X4 U5142 ( .A(n4946), .ZN(n4947) );
  OR2_X1 U5143 ( .A1(n8578), .A2(n8897), .ZN(n6148) );
  AND2_X1 U5144 ( .A1(n10778), .A2(n7896), .ZN(n8569) );
  INV_X1 U5145 ( .A(n8269), .ZN(n5379) );
  AOI21_X1 U5146 ( .B1(n5403), .B2(n5405), .A(n4997), .ZN(n5402) );
  INV_X1 U5147 ( .A(n5951), .ZN(n5403) );
  XNOR2_X1 U5148 ( .A(n8766), .B(n8892), .ZN(n8709) );
  AOI211_X1 U5149 ( .C1(n8655), .C2(n9206), .A(n8602), .B(n9154), .ZN(n8606)
         );
  AND2_X1 U5150 ( .A1(n5295), .A2(n8478), .ZN(n5293) );
  NAND2_X1 U5151 ( .A1(n6727), .A2(n6615), .ZN(n6828) );
  NAND2_X1 U5152 ( .A1(n5510), .A2(n4965), .ZN(n5120) );
  INV_X1 U5153 ( .A(n5481), .ZN(n5480) );
  NOR2_X1 U5154 ( .A1(n9236), .A2(n9085), .ZN(n8622) );
  OR2_X1 U5155 ( .A1(n8708), .A2(n9137), .ZN(n6155) );
  AND2_X1 U5156 ( .A1(n5489), .A2(n8903), .ZN(n5073) );
  AND2_X1 U5157 ( .A1(n5078), .A2(n5798), .ZN(n5490) );
  NAND2_X1 U5158 ( .A1(n6885), .A2(n5079), .ZN(n5078) );
  INV_X1 U5159 ( .A(n5536), .ZN(n5535) );
  INV_X1 U5160 ( .A(n9587), .ZN(n5336) );
  OR2_X1 U5161 ( .A1(n10272), .A2(n10280), .ZN(n9853) );
  OR2_X1 U5162 ( .A1(n10291), .A2(n10281), .ZN(n9847) );
  NAND2_X1 U5163 ( .A1(n10291), .A2(n10281), .ZN(n10086) );
  AND2_X1 U5164 ( .A1(n10308), .A2(n9638), .ZN(n9813) );
  OR2_X1 U5165 ( .A1(n10204), .A2(n10339), .ZN(n10170) );
  INV_X1 U5166 ( .A(n5366), .ZN(n5365) );
  OAI21_X1 U5167 ( .B1(n5367), .B2(n5369), .A(n5555), .ZN(n5366) );
  OR2_X1 U5168 ( .A1(n10222), .A2(n10237), .ZN(n5555) );
  NAND2_X1 U5169 ( .A1(n5365), .A2(n5367), .ZN(n5363) );
  NOR2_X1 U5170 ( .A1(n10360), .A2(n10355), .ZN(n5268) );
  NAND2_X1 U5171 ( .A1(n8267), .A2(n9695), .ZN(n5436) );
  NAND2_X1 U5172 ( .A1(n6797), .A2(n5575), .ZN(n7185) );
  AND2_X1 U5173 ( .A1(n5603), .A2(n4973), .ZN(n5163) );
  XNOR2_X1 U5174 ( .A(n5597), .B(SI_8_), .ZN(n5846) );
  NAND2_X1 U5175 ( .A1(n5594), .A2(SI_7_), .ZN(n5844) );
  NAND2_X1 U5176 ( .A1(n5581), .A2(SI_4_), .ZN(n5584) );
  NAND2_X1 U5177 ( .A1(n5576), .A2(SI_3_), .ZN(n5580) );
  XNOR2_X1 U5178 ( .A(n6751), .B(n7116), .ZN(n6762) );
  NAND2_X1 U5179 ( .A1(n8508), .A2(n6746), .ZN(n8509) );
  INV_X1 U5180 ( .A(n5930), .ZN(n6250) );
  NOR2_X1 U5182 ( .A1(n10532), .A2(n6675), .ZN(n6676) );
  NAND2_X1 U5183 ( .A1(n5131), .A2(n5133), .ZN(n7711) );
  AND2_X1 U5184 ( .A1(n5132), .A2(n5032), .ZN(n5131) );
  NAND2_X1 U5185 ( .A1(n7918), .A2(n7919), .ZN(n8908) );
  NAND2_X1 U5186 ( .A1(n8929), .A2(n5512), .ZN(n5510) );
  OR2_X1 U5187 ( .A1(n8907), .A2(n5511), .ZN(n5124) );
  OAI22_X1 U5188 ( .A1(n9050), .A2(n6102), .B1(n9171), .B2(n8891), .ZN(n9039)
         );
  NAND2_X1 U5189 ( .A1(n9078), .A2(n9077), .ZN(n5290) );
  NOR2_X1 U5190 ( .A1(n9114), .A2(n5302), .ZN(n5301) );
  INV_X1 U5191 ( .A(n6156), .ZN(n5302) );
  NOR2_X1 U5192 ( .A1(n5305), .A2(n8099), .ZN(n5304) );
  INV_X1 U5193 ( .A(n6151), .ZN(n5305) );
  NAND2_X1 U5194 ( .A1(n5069), .A2(n6148), .ZN(n5068) );
  NAND2_X1 U5195 ( .A1(n8577), .A2(n5935), .ZN(n5069) );
  INV_X1 U5196 ( .A(n5067), .ZN(n5066) );
  OAI21_X1 U5197 ( .B1(n5068), .B2(n5935), .A(n8584), .ZN(n5067) );
  NAND2_X1 U5198 ( .A1(n5274), .A2(n5277), .ZN(n5273) );
  NAND2_X1 U5199 ( .A1(n7667), .A2(n6144), .ZN(n7741) );
  AOI21_X1 U5200 ( .B1(n10339), .B2(n8438), .A(n8397), .ZN(n8403) );
  NOR2_X1 U5201 ( .A1(n8416), .A2(n8415), .ZN(n8417) );
  INV_X1 U5202 ( .A(n5317), .ZN(n5316) );
  OAI21_X1 U5203 ( .B1(n8431), .B2(n8433), .A(n9569), .ZN(n5317) );
  AND2_X1 U5204 ( .A1(n10267), .A2(n10076), .ZN(n9939) );
  NOR2_X1 U5205 ( .A1(n10125), .A2(n10291), .ZN(n10070) );
  OAI21_X1 U5206 ( .B1(n10124), .B2(n10123), .A(n9816), .ZN(n8320) );
  NAND2_X1 U5207 ( .A1(n5262), .A2(n10305), .ZN(n8299) );
  INV_X1 U5208 ( .A(n5376), .ZN(n5375) );
  OAI21_X1 U5209 ( .B1(n8275), .B2(n5377), .A(n8274), .ZN(n5376) );
  OR2_X1 U5210 ( .A1(n5380), .A2(n5379), .ZN(n5377) );
  OR2_X1 U5211 ( .A1(n10314), .A2(n10318), .ZN(n9841) );
  AND2_X1 U5212 ( .A1(n10365), .A2(n10368), .ZN(n8208) );
  NOR2_X1 U5213 ( .A1(n9788), .A2(n9957), .ZN(n5397) );
  OR2_X1 U5214 ( .A1(n10371), .A2(n10824), .ZN(n8124) );
  AOI21_X1 U5215 ( .B1(n10786), .B2(n10801), .A(n7811), .ZN(n8030) );
  XNOR2_X1 U5217 ( .A(n6247), .B(n6246), .ZN(n8687) );
  NOR2_X1 U5218 ( .A1(n6043), .A2(n5415), .ZN(n5414) );
  INV_X1 U5219 ( .A(n5634), .ZN(n5415) );
  NOR2_X1 U5220 ( .A1(n5400), .A2(n5175), .ZN(n5174) );
  INV_X1 U5221 ( .A(n5556), .ZN(n5175) );
  NAND2_X1 U5222 ( .A1(n5164), .A2(n5163), .ZN(n5876) );
  NAND2_X1 U5223 ( .A1(n5803), .A2(n5589), .ZN(n5824) );
  CLKBUF_X1 U5224 ( .A(n6361), .Z(n6362) );
  CLKBUF_X1 U5225 ( .A(n5674), .Z(n8169) );
  INV_X1 U5226 ( .A(n9051), .ZN(n9076) );
  INV_X1 U5227 ( .A(n8891), .ZN(n9064) );
  AND2_X1 U5228 ( .A1(n6284), .A2(n6283), .ZN(n5052) );
  NAND2_X1 U5229 ( .A1(n5250), .A2(n8655), .ZN(n5249) );
  NAND2_X1 U5230 ( .A1(n8549), .A2(n8610), .ZN(n5248) );
  NAND2_X1 U5231 ( .A1(n8547), .A2(n8548), .ZN(n5250) );
  OAI211_X1 U5232 ( .C1(n5245), .C2(n4983), .A(n5242), .B(n4961), .ZN(n5241)
         );
  OAI21_X1 U5233 ( .B1(n8572), .B2(n5244), .A(n5243), .ZN(n5242) );
  AOI211_X1 U5234 ( .C1(n8572), .C2(n8571), .A(n8569), .B(n8570), .ZN(n5245)
         );
  NOR2_X1 U5235 ( .A1(n5240), .A2(n5277), .ZN(n5239) );
  INV_X1 U5236 ( .A(n8576), .ZN(n5240) );
  NAND2_X1 U5237 ( .A1(n9854), .A2(n9831), .ZN(n5432) );
  NAND2_X1 U5238 ( .A1(n4970), .A2(n5232), .ZN(n5231) );
  NAND2_X1 U5239 ( .A1(n5004), .A2(n5233), .ZN(n5232) );
  NOR2_X1 U5240 ( .A1(n9043), .A2(n8645), .ZN(n5233) );
  INV_X1 U5241 ( .A(n6246), .ZN(n5193) );
  INV_X1 U5242 ( .A(n8888), .ZN(n6296) );
  OR2_X1 U5243 ( .A1(n9171), .A2(n9064), .ZN(n8642) );
  NAND2_X1 U5244 ( .A1(n9179), .A2(n9076), .ZN(n5497) );
  INV_X1 U5245 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6173) );
  INV_X1 U5246 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5281) );
  INV_X1 U5247 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5280) );
  NOR2_X1 U5248 ( .A1(n5846), .A2(n5196), .ZN(n5409) );
  NAND2_X1 U5249 ( .A1(n5410), .A2(n5844), .ZN(n5196) );
  NAND2_X1 U5250 ( .A1(n5829), .A2(n5411), .ZN(n5410) );
  INV_X1 U5251 ( .A(n5593), .ZN(n5411) );
  OAI21_X1 U5252 ( .B1(n5674), .B2(n5047), .A(n5046), .ZN(n5563) );
  INV_X1 U5253 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5047) );
  NAND2_X1 U5254 ( .A1(n5674), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5046) );
  INV_X1 U5255 ( .A(n5551), .ZN(n5548) );
  NOR2_X1 U5256 ( .A1(n9222), .A2(n8887), .ZN(n8665) );
  AOI21_X1 U5257 ( .B1(n8662), .B2(n8661), .A(n8660), .ZN(n8671) );
  OAI21_X1 U5258 ( .B1(n8640), .B2(n5229), .A(n5225), .ZN(n8662) );
  NAND2_X1 U5259 ( .A1(n5230), .A2(n5222), .ZN(n5229) );
  NOR2_X1 U5260 ( .A1(n8507), .A2(n5182), .ZN(n5181) );
  NAND2_X1 U5261 ( .A1(n5292), .A2(n5183), .ZN(n5182) );
  NAND2_X1 U5262 ( .A1(n10493), .A2(n6669), .ZN(n6671) );
  AND2_X1 U5263 ( .A1(n6671), .A2(n6670), .ZN(n6673) );
  NAND2_X1 U5264 ( .A1(n10535), .A2(n6642), .ZN(n6643) );
  NAND2_X1 U5265 ( .A1(n6939), .A2(n5200), .ZN(n7160) );
  OR2_X1 U5266 ( .A1(n6940), .A2(n6647), .ZN(n5200) );
  AND2_X1 U5267 ( .A1(n8651), .A2(n8646), .ZN(n6263) );
  AND2_X1 U5268 ( .A1(n6241), .A2(n4950), .ZN(n5080) );
  OR2_X1 U5269 ( .A1(n8750), .A2(n8889), .ZN(n6241) );
  NOR2_X1 U5270 ( .A1(n6296), .A2(n9150), .ZN(n6298) );
  NOR2_X1 U5271 ( .A1(n9041), .A2(n9148), .ZN(n6297) );
  OR2_X1 U5272 ( .A1(n6264), .A2(n6263), .ZN(n6267) );
  AND2_X1 U5273 ( .A1(n8868), .A2(n9052), .ZN(n5481) );
  INV_X1 U5274 ( .A(n5061), .ZN(n5060) );
  NAND2_X1 U5275 ( .A1(n5057), .A2(n5060), .ZN(n5055) );
  AND2_X1 U5276 ( .A1(n5058), .A2(n5482), .ZN(n5057) );
  NAND2_X1 U5277 ( .A1(n4955), .A2(n5483), .ZN(n5482) );
  NAND2_X1 U5278 ( .A1(n5061), .A2(n5059), .ZN(n5058) );
  NAND2_X1 U5279 ( .A1(n6028), .A2(n5485), .ZN(n5483) );
  AOI21_X1 U5280 ( .B1(n8493), .B2(n5466), .A(n4991), .ZN(n5465) );
  INV_X1 U5281 ( .A(n7417), .ZN(n5466) );
  INV_X1 U5282 ( .A(n5490), .ZN(n5488) );
  AND2_X1 U5283 ( .A1(n7358), .A2(n8556), .ZN(n8551) );
  OAI21_X1 U5284 ( .B1(n7099), .B2(n8532), .A(n8550), .ZN(n7292) );
  NOR2_X1 U5285 ( .A1(n6344), .A2(n4945), .ZN(n5070) );
  XNOR2_X1 U5286 ( .A(n6803), .B(n6828), .ZN(n6808) );
  XNOR2_X1 U5287 ( .A(n8412), .B(n8460), .ZN(n9295) );
  NOR2_X1 U5288 ( .A1(n10107), .A2(n5420), .ZN(n5419) );
  INV_X1 U5289 ( .A(n9824), .ZN(n5420) );
  OR2_X1 U5290 ( .A1(n10131), .A2(n10305), .ZN(n9846) );
  AND2_X1 U5291 ( .A1(n9844), .A2(n9815), .ZN(n9818) );
  NAND2_X1 U5292 ( .A1(n5436), .A2(n5434), .ZN(n9809) );
  NOR2_X1 U5293 ( .A1(n10176), .A2(n5435), .ZN(n5434) );
  INV_X1 U5294 ( .A(n8268), .ZN(n5435) );
  NAND2_X1 U5295 ( .A1(n10321), .A2(n10176), .ZN(n9838) );
  NOR2_X1 U5296 ( .A1(n10170), .A2(n10178), .ZN(n10154) );
  INV_X1 U5297 ( .A(n9772), .ZN(n5443) );
  AOI21_X1 U5298 ( .B1(n9772), .B2(n5442), .A(n5441), .ZN(n5440) );
  INV_X1 U5299 ( .A(n9761), .ZN(n5441) );
  NAND2_X1 U5300 ( .A1(n4979), .A2(n5393), .ZN(n5386) );
  INV_X1 U5301 ( .A(n5388), .ZN(n5383) );
  NAND2_X1 U5302 ( .A1(n7849), .A2(n10757), .ZN(n5395) );
  AND2_X1 U5303 ( .A1(n5396), .A2(n5395), .ZN(n5388) );
  OR2_X1 U5304 ( .A1(n8200), .A2(n10680), .ZN(n9746) );
  XNOR2_X1 U5305 ( .A(n7347), .B(n6968), .ZN(n9670) );
  INV_X1 U5306 ( .A(n5187), .ZN(n5186) );
  AOI21_X1 U5307 ( .B1(n5187), .B2(n5185), .A(n5034), .ZN(n5184) );
  AOI21_X1 U5308 ( .B1(n6058), .B2(n5643), .A(n5001), .ZN(n5187) );
  OAI21_X1 U5309 ( .B1(n6012), .B2(n6011), .A(n5631), .ZN(n6030) );
  INV_X1 U5310 ( .A(n5859), .ZN(n5157) );
  NOR2_X1 U5311 ( .A1(n5161), .A2(n5424), .ZN(n5160) );
  INV_X1 U5312 ( .A(n5163), .ZN(n5161) );
  INV_X1 U5313 ( .A(n5425), .ZN(n5424) );
  INV_X1 U5314 ( .A(n5429), .ZN(n5423) );
  INV_X1 U5315 ( .A(n5607), .ZN(n5422) );
  NOR2_X1 U5316 ( .A1(n5888), .A2(n5430), .ZN(n5429) );
  INV_X1 U5317 ( .A(n5604), .ZN(n5430) );
  XNOR2_X1 U5318 ( .A(n5605), .B(SI_11_), .ZN(n5888) );
  XNOR2_X1 U5319 ( .A(n5599), .B(n9472), .ZN(n5859) );
  NAND2_X1 U5320 ( .A1(n5408), .A2(n5407), .ZN(n5858) );
  AOI21_X1 U5321 ( .B1(n5409), .B2(n5412), .A(n4999), .ZN(n5407) );
  NAND2_X1 U5322 ( .A1(n5822), .A2(n5409), .ZN(n5408) );
  INV_X1 U5323 ( .A(n5829), .ZN(n5412) );
  NAND2_X1 U5324 ( .A1(n5590), .A2(SI_6_), .ZN(n5593) );
  NAND2_X1 U5325 ( .A1(n5585), .A2(SI_5_), .ZN(n5589) );
  NAND2_X1 U5326 ( .A1(n5563), .A2(SI_1_), .ZN(n5569) );
  XNOR2_X1 U5327 ( .A(n5082), .B(P2_IR_REG_27__SCAN_IN), .ZN(n6127) );
  NOR2_X1 U5328 ( .A1(n5671), .A2(n5672), .ZN(n5082) );
  XNOR2_X1 U5329 ( .A(n5670), .B(n5669), .ZN(n6125) );
  INV_X1 U5330 ( .A(n8903), .ZN(n7088) );
  NOR2_X1 U5331 ( .A1(n5171), .A2(n7614), .ZN(n5170) );
  INV_X1 U5332 ( .A(n5544), .ZN(n5171) );
  AND2_X1 U5333 ( .A1(n5148), .A2(n5147), .ZN(n8851) );
  AND2_X1 U5334 ( .A1(n5149), .A2(n5017), .ZN(n5147) );
  NAND2_X1 U5335 ( .A1(n8147), .A2(n5165), .ZN(n8697) );
  NOR2_X1 U5336 ( .A1(n8150), .A2(n5166), .ZN(n5165) );
  INV_X1 U5337 ( .A(n8146), .ZN(n5166) );
  XNOR2_X1 U5338 ( .A(n10503), .B(n6666), .ZN(n10495) );
  NAND2_X1 U5339 ( .A1(n10495), .A2(n10494), .ZN(n10493) );
  NOR2_X1 U5340 ( .A1(n5768), .A2(n10515), .ZN(n10514) );
  NOR2_X1 U5341 ( .A1(n10545), .A2(n10546), .ZN(n10544) );
  OR2_X1 U5342 ( .A1(n10544), .A2(n5088), .ZN(n5087) );
  NOR2_X1 U5343 ( .A1(n5089), .A2(n10543), .ZN(n5088) );
  INV_X1 U5344 ( .A(n6657), .ZN(n5089) );
  XNOR2_X1 U5345 ( .A(n6643), .B(n10566), .ZN(n10556) );
  NAND2_X1 U5346 ( .A1(n10556), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10555) );
  OR2_X1 U5347 ( .A1(n5804), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5825) );
  XNOR2_X1 U5348 ( .A(n7160), .B(n7143), .ZN(n6941) );
  NAND2_X1 U5349 ( .A1(n6941), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7162) );
  OR2_X1 U5350 ( .A1(n6926), .A2(n7143), .ZN(n5126) );
  NAND2_X1 U5351 ( .A1(n6926), .A2(n5023), .ZN(n5125) );
  OR2_X1 U5352 ( .A1(n6925), .A2(n7143), .ZN(n5127) );
  NAND2_X1 U5353 ( .A1(n5505), .A2(n5504), .ZN(n7443) );
  AND2_X1 U5354 ( .A1(n7710), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5116) );
  OR2_X1 U5355 ( .A1(n7711), .A2(n7720), .ZN(n5513) );
  NAND2_X1 U5356 ( .A1(n10573), .A2(n7717), .ZN(n7718) );
  NAND2_X1 U5357 ( .A1(n7718), .A2(n7719), .ZN(n7777) );
  NAND2_X1 U5358 ( .A1(n5114), .A2(n5116), .ZN(n5112) );
  AND2_X1 U5359 ( .A1(n5513), .A2(n5115), .ZN(n5114) );
  NAND2_X1 U5360 ( .A1(n5111), .A2(n5115), .ZN(n5110) );
  NAND2_X1 U5361 ( .A1(n7777), .A2(n5199), .ZN(n7915) );
  NAND2_X1 U5362 ( .A1(n7780), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5199) );
  NAND2_X1 U5363 ( .A1(n8908), .A2(n8909), .ZN(n8931) );
  NAND2_X1 U5364 ( .A1(n5120), .A2(n8974), .ZN(n5119) );
  OR2_X1 U5365 ( .A1(n5511), .A2(n8984), .ZN(n5121) );
  OR2_X1 U5366 ( .A1(n8977), .A2(n8978), .ZN(n8979) );
  INV_X1 U5367 ( .A(n5120), .ZN(n5123) );
  NAND2_X1 U5368 ( .A1(n8979), .A2(n8980), .ZN(n8994) );
  AOI21_X1 U5369 ( .B1(n5297), .B2(n6273), .A(n5296), .ZN(n5295) );
  INV_X1 U5370 ( .A(n6274), .ZN(n5296) );
  INV_X1 U5371 ( .A(n6271), .ZN(n5297) );
  NOR2_X1 U5372 ( .A1(n6129), .A2(n6785), .ZN(n6131) );
  OR2_X1 U5373 ( .A1(n8868), .A2(n8790), .ZN(n8485) );
  NAND2_X1 U5374 ( .A1(n6266), .A2(n8641), .ZN(n9042) );
  NAND2_X1 U5375 ( .A1(n8634), .A2(n5495), .ZN(n5494) );
  NAND2_X1 U5376 ( .A1(n5496), .A2(n6161), .ZN(n5495) );
  NAND2_X1 U5377 ( .A1(n6070), .A2(n8631), .ZN(n5496) );
  NAND2_X1 U5378 ( .A1(n9084), .A2(n4959), .ZN(n5493) );
  OR2_X1 U5379 ( .A1(n9184), .A2(n9104), .ZN(n8631) );
  OAI22_X1 U5380 ( .A1(n9088), .A2(n6160), .B1(n6159), .B2(n9104), .ZN(n9078)
         );
  NOR2_X1 U5381 ( .A1(n9102), .A2(n8622), .ZN(n9084) );
  NOR2_X1 U5382 ( .A1(n9095), .A2(n8616), .ZN(n5299) );
  OR2_X1 U5383 ( .A1(n9194), .A2(n9103), .ZN(n9099) );
  NAND2_X1 U5384 ( .A1(n9139), .A2(n8709), .ZN(n6157) );
  NAND2_X1 U5385 ( .A1(n6150), .A2(n5059), .ZN(n7965) );
  AOI21_X1 U5386 ( .B1(n7857), .B2(n5066), .A(n5064), .ZN(n5063) );
  NAND2_X1 U5387 ( .A1(n5065), .A2(n8582), .ZN(n5064) );
  NAND2_X1 U5388 ( .A1(n5066), .A2(n5068), .ZN(n5065) );
  AOI21_X1 U5389 ( .B1(n8577), .B2(n5276), .A(n5275), .ZN(n5274) );
  INV_X1 U5390 ( .A(n8575), .ZN(n5276) );
  NAND2_X1 U5391 ( .A1(n7741), .A2(n6146), .ZN(n6147) );
  NAND2_X1 U5392 ( .A1(n7619), .A2(n6143), .ZN(n7667) );
  OR2_X1 U5393 ( .A1(n7626), .A2(n7700), .ZN(n8548) );
  NAND2_X1 U5394 ( .A1(n7360), .A2(n7417), .ZN(n5464) );
  AOI21_X1 U5395 ( .B1(n5799), .B2(n5490), .A(n4994), .ZN(n5489) );
  OR2_X1 U5396 ( .A1(n8610), .A2(n6786), .ZN(n9148) );
  INV_X1 U5397 ( .A(n9150), .ZN(n10608) );
  NAND2_X1 U5398 ( .A1(n8175), .A2(n8174), .ZN(n8481) );
  NAND2_X1 U5399 ( .A1(n6019), .A2(n6018), .ZN(n8766) );
  NAND2_X1 U5400 ( .A1(n6006), .A2(n6005), .ZN(n8708) );
  INV_X1 U5401 ( .A(n7116), .ZN(n10628) );
  NAND2_X1 U5402 ( .A1(n9255), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5696) );
  INV_X1 U5403 ( .A(n5532), .ZN(n5531) );
  OAI21_X1 U5404 ( .B1(n6104), .B2(n5672), .A(n6112), .ZN(n5532) );
  NAND2_X1 U5405 ( .A1(n5530), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6108) );
  AND2_X1 U5406 ( .A1(n5775), .A2(n5804), .ZN(n10520) );
  AND2_X1 U5407 ( .A1(n5672), .A2(n5662), .ZN(n5508) );
  AND2_X1 U5408 ( .A1(n5518), .A2(n5517), .ZN(n6556) );
  NAND2_X1 U5409 ( .A1(n5319), .A2(n4982), .ZN(n7762) );
  NAND2_X1 U5410 ( .A1(n5323), .A2(n5320), .ZN(n5319) );
  NAND2_X1 U5411 ( .A1(n7763), .A2(n7764), .ZN(n5355) );
  AOI21_X1 U5412 ( .B1(n5325), .B2(n5322), .A(n5324), .ZN(n5321) );
  NAND2_X1 U5413 ( .A1(n5332), .A2(n5330), .ZN(n5329) );
  INV_X1 U5414 ( .A(n8390), .ZN(n5330) );
  AND2_X1 U5415 ( .A1(n9607), .A2(n5022), .ZN(n5332) );
  NOR2_X1 U5416 ( .A1(n8374), .A2(n9648), .ZN(n5340) );
  NAND2_X1 U5417 ( .A1(n8432), .A2(n8431), .ZN(n9596) );
  XNOR2_X1 U5418 ( .A(n7192), .B(n6829), .ZN(n7217) );
  NAND2_X1 U5419 ( .A1(n5309), .A2(n5308), .ZN(n8366) );
  AOI21_X1 U5420 ( .B1(n5310), .B2(n5313), .A(n5000), .ZN(n5308) );
  INV_X1 U5421 ( .A(n8116), .ZN(n5313) );
  NAND2_X1 U5422 ( .A1(n10078), .A2(n9663), .ZN(n9942) );
  XNOR2_X1 U5423 ( .A(n9973), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n9970) );
  OR2_X1 U5424 ( .A1(n9970), .A2(n9971), .ZN(n5142) );
  OR2_X1 U5425 ( .A1(n6590), .A2(n6589), .ZN(n5138) );
  NOR2_X1 U5426 ( .A1(n6536), .A2(n5020), .ZN(n6497) );
  NOR2_X1 U5427 ( .A1(n6497), .A2(n5040), .ZN(n6575) );
  NOR2_X1 U5428 ( .A1(n6533), .A2(n5021), .ZN(n6483) );
  AOI21_X1 U5429 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n8063), .A(n8059), .ZN(
        n10004) );
  NAND2_X1 U5430 ( .A1(n9666), .A2(n9665), .ZN(n10272) );
  NAND2_X1 U5431 ( .A1(n10154), .A2(n5261), .ZN(n10125) );
  AND2_X1 U5432 ( .A1(n4957), .A2(n5262), .ZN(n5261) );
  AOI21_X1 U5433 ( .B1(n5446), .B2(n9691), .A(n9813), .ZN(n5444) );
  INV_X1 U5434 ( .A(n5446), .ZN(n5445) );
  AOI21_X1 U5435 ( .B1(n4958), .B2(n5378), .A(n5005), .ZN(n5371) );
  OR2_X1 U5436 ( .A1(n8275), .A2(n5379), .ZN(n5378) );
  INV_X1 U5437 ( .A(n9818), .ZN(n10137) );
  NOR2_X1 U5438 ( .A1(n10137), .A2(n5447), .ZN(n5446) );
  INV_X1 U5439 ( .A(n9841), .ZN(n5447) );
  NAND2_X1 U5440 ( .A1(n8342), .A2(n9811), .ZN(n8341) );
  NOR2_X1 U5441 ( .A1(n8270), .A2(n5381), .ZN(n5380) );
  INV_X1 U5442 ( .A(n8265), .ZN(n5381) );
  NOR2_X1 U5443 ( .A1(n4969), .A2(n5370), .ZN(n5369) );
  INV_X1 U5444 ( .A(n8213), .ZN(n5370) );
  INV_X1 U5445 ( .A(n9688), .ZN(n10225) );
  AOI21_X1 U5446 ( .B1(n8229), .B2(n5368), .A(n4969), .ZN(n5367) );
  INV_X1 U5447 ( .A(n5557), .ZN(n5368) );
  NOR2_X1 U5448 ( .A1(n10817), .A2(n9788), .ZN(n8128) );
  NAND2_X1 U5449 ( .A1(n9921), .A2(n9919), .ZN(n9686) );
  NAND2_X1 U5450 ( .A1(n10846), .A2(n8046), .ZN(n5399) );
  NAND2_X1 U5451 ( .A1(n5394), .A2(n10787), .ZN(n5393) );
  NAND2_X1 U5452 ( .A1(n5390), .A2(n5395), .ZN(n5389) );
  INV_X1 U5453 ( .A(n5391), .ZN(n5390) );
  AOI21_X1 U5454 ( .B1(n10718), .B2(n5396), .A(n5392), .ZN(n5391) );
  INV_X1 U5455 ( .A(n7595), .ZN(n5392) );
  NAND2_X1 U5456 ( .A1(n7504), .A2(n5562), .ZN(n7505) );
  NOR2_X1 U5457 ( .A1(n7204), .A2(n6446), .ZN(n7276) );
  NAND2_X1 U5458 ( .A1(n8200), .A2(n10680), .ZN(n10687) );
  BUF_X1 U5459 ( .A(n9670), .Z(n5042) );
  AOI21_X1 U5460 ( .B1(n9662), .B2(n9695), .A(n5561), .ZN(n10267) );
  INV_X1 U5461 ( .A(n10084), .ZN(n10270) );
  INV_X1 U5462 ( .A(n10296), .ZN(n10281) );
  NAND2_X1 U5463 ( .A1(n8127), .A2(n8126), .ZN(n10365) );
  NAND2_X1 U5464 ( .A1(n6977), .A2(n6976), .ZN(n10828) );
  AND2_X1 U5465 ( .A1(n6710), .A2(n10395), .ZN(n7300) );
  NAND2_X1 U5466 ( .A1(n10397), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6428) );
  XNOR2_X1 U5467 ( .A(n8470), .B(n8469), .ZN(n9696) );
  XNOR2_X1 U5468 ( .A(n6430), .B(P1_IR_REG_29__SCAN_IN), .ZN(n6431) );
  OR2_X1 U5469 ( .A1(n6429), .A2(n10396), .ZN(n6430) );
  XNOR2_X1 U5470 ( .A(n6392), .B(n6426), .ZN(n6417) );
  OR2_X1 U5471 ( .A1(n6394), .A2(n10396), .ZN(n6392) );
  OAI21_X1 U5472 ( .B1(n6335), .B2(n5253), .A(n5251), .ZN(n6418) );
  NAND2_X1 U5473 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n5253) );
  NOR2_X1 U5474 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5252) );
  XNOR2_X1 U5475 ( .A(n5718), .B(n5717), .ZN(n8288) );
  NAND2_X1 U5476 ( .A1(n6086), .A2(n5643), .ZN(n5716) );
  XNOR2_X1 U5477 ( .A(n6090), .B(n6089), .ZN(n8276) );
  AND2_X1 U5478 ( .A1(n6088), .A2(n6087), .ZN(n6090) );
  OR2_X1 U5479 ( .A1(n6059), .A2(n6058), .ZN(n6086) );
  AND2_X2 U5480 ( .A1(n7067), .A2(n6317), .ZN(n6326) );
  INV_X1 U5481 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6317) );
  INV_X1 U5482 ( .A(n5984), .ZN(n5401) );
  NAND2_X1 U5483 ( .A1(n5939), .A2(n5177), .ZN(n5176) );
  AND2_X1 U5484 ( .A1(n4960), .A2(n5615), .ZN(n5177) );
  OAI21_X1 U5485 ( .B1(n5952), .B2(n5404), .A(n5402), .ZN(n5985) );
  NAND2_X1 U5486 ( .A1(n5952), .A2(n5951), .ZN(n5954) );
  OAI21_X1 U5487 ( .B1(n5606), .B2(SI_12_), .A(n5607), .ZN(n5904) );
  NOR2_X1 U5488 ( .A1(n5904), .A2(n5428), .ZN(n5425) );
  NAND2_X1 U5489 ( .A1(n5876), .A2(n5429), .ZN(n5426) );
  NAND2_X1 U5490 ( .A1(n5604), .A2(n5602), .ZN(n5874) );
  NAND2_X1 U5491 ( .A1(n5858), .A2(n5859), .ZN(n5164) );
  NAND2_X1 U5492 ( .A1(n5845), .A2(n5844), .ZN(n5216) );
  NAND2_X1 U5493 ( .A1(n5822), .A2(n5593), .ZN(n5830) );
  OAI21_X1 U5494 ( .B1(n5360), .B2(n5580), .A(n5584), .ZN(n5211) );
  INV_X1 U5495 ( .A(n6362), .ZN(n5455) );
  NAND2_X1 U5496 ( .A1(n5776), .A2(n5777), .ZN(n5779) );
  AND2_X1 U5497 ( .A1(n6356), .A2(n6355), .ZN(n6821) );
  OR2_X1 U5498 ( .A1(n7087), .A2(n7088), .ZN(n5551) );
  INV_X1 U5499 ( .A(n5550), .ZN(n7316) );
  AOI21_X1 U5500 ( .B1(n8862), .B2(n5024), .A(n5144), .ZN(n5146) );
  NAND2_X1 U5501 ( .A1(n5145), .A2(n8848), .ZN(n5144) );
  NAND2_X1 U5502 ( .A1(n8753), .A2(n5030), .ZN(n5145) );
  NAND2_X1 U5503 ( .A1(n6075), .A2(n6074), .ZN(n8763) );
  AOI21_X1 U5504 ( .B1(n5541), .B2(n5540), .A(n5539), .ZN(n5538) );
  INV_X1 U5505 ( .A(n8742), .ZN(n5539) );
  INV_X1 U5506 ( .A(n8863), .ZN(n5540) );
  AND2_X1 U5507 ( .A1(n6758), .A2(n6756), .ZN(n6954) );
  NAND2_X1 U5508 ( .A1(n5911), .A2(n5910), .ZN(n7903) );
  NAND2_X1 U5509 ( .A1(n5974), .A2(n5973), .ZN(n8801) );
  NAND2_X1 U5510 ( .A1(n5728), .A2(n5727), .ZN(n8819) );
  NAND2_X1 U5511 ( .A1(n6864), .A2(n5526), .ZN(n5524) );
  AND3_X1 U5512 ( .A1(n5996), .A2(n5995), .A3(n5994), .ZN(n9147) );
  NOR2_X1 U5513 ( .A1(n8676), .A2(n5178), .ZN(n8678) );
  AOI21_X1 U5514 ( .B1(n5217), .B2(n8673), .A(n6745), .ZN(n8676) );
  AOI21_X1 U5515 ( .B1(n8509), .B2(n5179), .A(n8675), .ZN(n5178) );
  NAND2_X1 U5516 ( .A1(n6101), .A2(n6100), .ZN(n8891) );
  NAND2_X1 U5517 ( .A1(n5734), .A2(n5733), .ZN(n9051) );
  AND2_X1 U5518 ( .A1(n6084), .A2(n6083), .ZN(n9063) );
  OR2_X1 U5519 ( .A1(n6680), .A2(n6679), .ZN(n6926) );
  XNOR2_X1 U5520 ( .A(n5849), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7391) );
  NAND2_X1 U5521 ( .A1(n5112), .A2(n5110), .ZN(n7774) );
  XNOR2_X1 U5522 ( .A(n8926), .B(n8927), .ZN(n8907) );
  NAND2_X1 U5523 ( .A1(n5104), .A2(n8997), .ZN(n5103) );
  OAI21_X1 U5524 ( .B1(n8988), .B2(n8989), .A(n10504), .ZN(n5104) );
  AOI21_X1 U5525 ( .B1(n8988), .B2(n5102), .A(n5100), .ZN(n5099) );
  NOR2_X1 U5526 ( .A1(n10562), .A2(n8997), .ZN(n5102) );
  INV_X1 U5527 ( .A(n5101), .ZN(n5100) );
  AOI21_X1 U5528 ( .B1(n10572), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8990), .ZN(
        n5101) );
  NAND2_X1 U5529 ( .A1(n5879), .A2(n5878), .ZN(n10771) );
  AND2_X1 U5530 ( .A1(n6285), .A2(n10655), .ZN(n6286) );
  OR2_X1 U5531 ( .A1(n8302), .A2(n6046), .ZN(n5677) );
  NAND2_X1 U5532 ( .A1(n6048), .A2(n6047), .ZN(n9236) );
  OR2_X1 U5533 ( .A1(n8244), .A2(n6046), .ZN(n6048) );
  NAND2_X1 U5534 ( .A1(n8304), .A2(n8303), .ZN(n10291) );
  OR2_X1 U5535 ( .A1(n8302), .A2(n8301), .ZN(n8304) );
  INV_X1 U5536 ( .A(n10161), .ZN(n10336) );
  NOR2_X1 U5537 ( .A1(n5346), .A2(n9632), .ZN(n5344) );
  NOR2_X1 U5538 ( .A1(n5347), .A2(n5349), .ZN(n5346) );
  INV_X1 U5539 ( .A(n5350), .ZN(n5347) );
  NAND2_X1 U5540 ( .A1(n5350), .A2(n5351), .ZN(n5348) );
  NAND2_X1 U5541 ( .A1(n8458), .A2(n8457), .ZN(n10284) );
  NAND2_X1 U5542 ( .A1(n8687), .A2(n9695), .ZN(n8458) );
  NAND2_X1 U5543 ( .A1(n8246), .A2(n8245), .ZN(n10339) );
  OR2_X1 U5544 ( .A1(n8244), .A2(n8301), .ZN(n8246) );
  INV_X1 U5545 ( .A(n10144), .ZN(n10318) );
  INV_X1 U5546 ( .A(n10226), .ZN(n10253) );
  NAND2_X1 U5547 ( .A1(n8273), .A2(n8272), .ZN(n10314) );
  NAND2_X1 U5548 ( .A1(n8271), .A2(n9695), .ZN(n8273) );
  NAND2_X1 U5549 ( .A1(n8414), .A2(n8413), .ZN(n9617) );
  NAND2_X1 U5550 ( .A1(n8216), .A2(n8215), .ZN(n10355) );
  OR2_X1 U5551 ( .A1(n8214), .A2(n8301), .ZN(n8216) );
  AOI21_X1 U5552 ( .B1(n5316), .B2(n8433), .A(n5003), .ZN(n5314) );
  NOR2_X1 U5553 ( .A1(n6483), .A2(n6484), .ZN(n6570) );
  INV_X1 U5554 ( .A(n10058), .ZN(n5045) );
  NAND2_X1 U5555 ( .A1(n7679), .A2(n7678), .ZN(n8078) );
  OR2_X1 U5556 ( .A1(n7676), .A2(n8301), .ZN(n7679) );
  NAND2_X1 U5557 ( .A1(n7566), .A2(n7565), .ZN(n10759) );
  OAI21_X1 U5558 ( .B1(n7263), .B2(n8301), .A(n7267), .ZN(n10698) );
  AND2_X1 U5559 ( .A1(n7266), .A2(n4987), .ZN(n7267) );
  NAND2_X1 U5560 ( .A1(n6730), .A2(n6982), .ZN(n10847) );
  INV_X1 U5561 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10396) );
  INV_X1 U5562 ( .A(n6136), .ZN(n8513) );
  NOR2_X1 U5563 ( .A1(n8565), .A2(n5246), .ZN(n8559) );
  NOR2_X1 U5564 ( .A1(n8549), .A2(n5247), .ZN(n5246) );
  INV_X1 U5565 ( .A(n8556), .ZN(n5247) );
  NAND2_X1 U5566 ( .A1(n5901), .A2(n8564), .ZN(n5244) );
  NAND2_X1 U5567 ( .A1(n5241), .A2(n5239), .ZN(n8586) );
  NAND2_X1 U5568 ( .A1(n5237), .A2(n5492), .ZN(n5236) );
  NAND2_X1 U5569 ( .A1(n4970), .A2(n5235), .ZN(n5234) );
  NOR2_X1 U5570 ( .A1(n8639), .A2(n8638), .ZN(n5235) );
  NAND2_X1 U5571 ( .A1(n9839), .A2(n9820), .ZN(n5433) );
  AND2_X1 U5572 ( .A1(n9756), .A2(n7592), .ZN(n9744) );
  INV_X1 U5573 ( .A(n5234), .ZN(n5230) );
  INV_X1 U5574 ( .A(n5226), .ZN(n5225) );
  OAI211_X1 U5575 ( .C1(n8658), .C2(n5231), .A(n5227), .B(n5238), .ZN(n5226)
         );
  NAND2_X1 U5576 ( .A1(n8653), .A2(n5222), .ZN(n5227) );
  AND2_X1 U5577 ( .A1(n8982), .A2(n5098), .ZN(n8986) );
  NAND2_X1 U5578 ( .A1(n8983), .A2(n8984), .ZN(n5098) );
  OR2_X1 U5579 ( .A1(n8099), .A2(n5486), .ZN(n5485) );
  NOR2_X1 U5580 ( .A1(n5484), .A2(n5062), .ZN(n5061) );
  INV_X1 U5581 ( .A(n5983), .ZN(n5062) );
  NAND2_X1 U5582 ( .A1(n4955), .A2(n5997), .ZN(n5484) );
  INV_X1 U5583 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5284) );
  INV_X1 U5584 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5283) );
  AOI21_X1 U5585 ( .B1(n9817), .B2(n9857), .A(n9812), .ZN(n9814) );
  INV_X1 U5586 ( .A(n9813), .ZN(n9815) );
  NOR2_X1 U5587 ( .A1(n10759), .A2(n10787), .ZN(n9904) );
  NAND2_X1 U5588 ( .A1(n5192), .A2(n6245), .ZN(n8162) );
  INV_X1 U5589 ( .A(n5643), .ZN(n5185) );
  NOR2_X2 U5590 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n6349) );
  NAND2_X1 U5591 ( .A1(n5209), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5155) );
  INV_X1 U5592 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5209) );
  NOR2_X1 U5593 ( .A1(n8665), .A2(n5298), .ZN(n5197) );
  NAND2_X1 U5594 ( .A1(n5293), .A2(n8743), .ZN(n5291) );
  INV_X1 U5595 ( .A(n8667), .ZN(n5298) );
  INV_X1 U5596 ( .A(n8673), .ZN(n8507) );
  INV_X1 U5597 ( .A(n8665), .ZN(n8668) );
  INV_X1 U5598 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5533) );
  OAI21_X1 U5599 ( .B1(n8679), .B2(P2_REG2_REG_1__SCAN_IN), .A(n5084), .ZN(
        n5083) );
  XNOR2_X1 U5600 ( .A(n6640), .B(n10520), .ZN(n10517) );
  NAND2_X1 U5601 ( .A1(n10501), .A2(n5198), .ZN(n6640) );
  OR2_X1 U5602 ( .A1(n6654), .A2(n6639), .ZN(n5198) );
  NAND2_X1 U5603 ( .A1(n4974), .A2(n10533), .ZN(n5130) );
  INV_X1 U5604 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5832) );
  NOR2_X1 U5605 ( .A1(n5097), .A2(n7447), .ZN(n5096) );
  INV_X1 U5606 ( .A(n7455), .ZN(n5097) );
  INV_X1 U5607 ( .A(n7446), .ZN(n5134) );
  INV_X1 U5608 ( .A(n7384), .ZN(n5092) );
  NAND2_X1 U5609 ( .A1(n5094), .A2(n7722), .ZN(n5093) );
  INV_X1 U5610 ( .A(n5096), .ZN(n5094) );
  INV_X1 U5611 ( .A(n8930), .ZN(n5512) );
  NAND2_X1 U5612 ( .A1(n5512), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5511) );
  NOR2_X1 U5613 ( .A1(n8986), .A2(n8985), .ZN(n8998) );
  INV_X1 U5614 ( .A(n8660), .ZN(n8505) );
  OR2_X1 U5615 ( .A1(n6095), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5708) );
  NOR2_X1 U5616 ( .A1(n6076), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5050) );
  INV_X1 U5617 ( .A(n5050), .ZN(n6078) );
  OR2_X1 U5618 ( .A1(n6062), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6076) );
  OR2_X1 U5619 ( .A1(n6034), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6049) );
  INV_X1 U5620 ( .A(n5051), .ZN(n5992) );
  NOR2_X1 U5621 ( .A1(n5895), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5049) );
  NAND2_X1 U5622 ( .A1(n7061), .A2(n8904), .ZN(n5798) );
  OR2_X1 U5623 ( .A1(n10609), .A2(n10628), .ZN(n8528) );
  AND2_X1 U5624 ( .A1(n6203), .A2(n5190), .ZN(n5189) );
  NAND2_X1 U5625 ( .A1(n5053), .A2(n4992), .ZN(n9050) );
  NAND2_X1 U5626 ( .A1(n9084), .A2(n4986), .ZN(n5053) );
  INV_X1 U5627 ( .A(n5497), .ZN(n5491) );
  INV_X1 U5628 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5537) );
  INV_X1 U5629 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9523) );
  NOR2_X1 U5630 ( .A1(n5324), .A2(n5322), .ZN(n5320) );
  NAND2_X1 U5631 ( .A1(n8195), .A2(n8196), .ZN(n5326) );
  NOR2_X1 U5632 ( .A1(n8195), .A2(n8196), .ZN(n5324) );
  INV_X1 U5633 ( .A(n5039), .ZN(n5322) );
  INV_X1 U5634 ( .A(n8374), .ZN(n5342) );
  AND2_X1 U5635 ( .A1(n8421), .A2(n8420), .ZN(n9292) );
  OR2_X1 U5636 ( .A1(n7981), .A2(n7984), .ZN(n7989) );
  AND2_X1 U5637 ( .A1(n8355), .A2(n5311), .ZN(n5310) );
  NAND2_X1 U5638 ( .A1(n8116), .A2(n5312), .ZN(n5311) );
  INV_X1 U5639 ( .A(n8113), .ZN(n5312) );
  NAND2_X1 U5640 ( .A1(n10284), .A2(n10288), .ZN(n9862) );
  OR2_X1 U5641 ( .A1(n10284), .A2(n10288), .ZN(n9850) );
  NOR2_X1 U5642 ( .A1(n10321), .A2(n10314), .ZN(n5263) );
  NOR2_X1 U5643 ( .A1(n8316), .A2(n5452), .ZN(n5451) );
  INV_X1 U5644 ( .A(n9929), .ZN(n5452) );
  OR2_X1 U5645 ( .A1(n10339), .A2(n10214), .ZN(n9930) );
  AND2_X1 U5646 ( .A1(n8219), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8234) );
  OR2_X1 U5647 ( .A1(n10365), .A2(n10252), .ZN(n9921) );
  OR2_X1 U5648 ( .A1(n7638), .A2(n10790), .ZN(n7686) );
  OR2_X1 U5649 ( .A1(n10748), .A2(n10757), .ZN(n9756) );
  AND2_X1 U5650 ( .A1(n10674), .A2(n7504), .ZN(n7500) );
  NAND2_X1 U5651 ( .A1(n7499), .A2(n7503), .ZN(n7504) );
  CLKBUF_X1 U5652 ( .A(n10682), .Z(n5043) );
  NAND2_X1 U5653 ( .A1(n7128), .A2(n9723), .ZN(n9731) );
  NAND2_X1 U5654 ( .A1(n9966), .A2(n6972), .ZN(n9893) );
  NAND2_X1 U5655 ( .A1(n10254), .A2(n10262), .ZN(n10255) );
  NOR2_X1 U5656 ( .A1(n7686), .A2(n8078), .ZN(n7814) );
  NOR2_X1 U5657 ( .A1(n10714), .A2(n10748), .ZN(n7587) );
  NAND3_X1 U5658 ( .A1(n4956), .A2(n5270), .A3(n7490), .ZN(n10714) );
  XNOR2_X1 U5659 ( .A(n8162), .B(n8161), .ZN(n8159) );
  AND2_X1 U5660 ( .A1(n6325), .A2(n5458), .ZN(n5457) );
  NOR2_X1 U5661 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n5458) );
  OR2_X1 U5662 ( .A1(n5654), .A2(n5653), .ZN(n5715) );
  OR2_X1 U5663 ( .A1(n6389), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n6391) );
  NAND2_X1 U5664 ( .A1(n6000), .A2(n5628), .ZN(n6012) );
  INV_X1 U5665 ( .A(n5620), .ZN(n5406) );
  INV_X1 U5666 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6310) );
  INV_X1 U5667 ( .A(n5563), .ZN(n5565) );
  NAND2_X1 U5668 ( .A1(n7317), .A2(n7318), .ZN(n5549) );
  NAND2_X1 U5669 ( .A1(n8849), .A2(n5547), .ZN(n5550) );
  NAND2_X1 U5670 ( .A1(n5150), .A2(n6766), .ZN(n5148) );
  AND2_X1 U5671 ( .A1(n6765), .A2(n5151), .ZN(n5150) );
  NAND2_X1 U5672 ( .A1(n6763), .A2(n10609), .ZN(n5526) );
  NAND2_X1 U5673 ( .A1(n8849), .A2(n4952), .ZN(n5172) );
  INV_X1 U5674 ( .A(n8772), .ZN(n8713) );
  NOR2_X1 U5675 ( .A1(n8849), .A2(n5169), .ZN(n5167) );
  OAI21_X1 U5676 ( .B1(n4952), .B2(n5169), .A(n4995), .ZN(n5168) );
  NAND2_X1 U5677 ( .A1(n5051), .A2(n9418), .ZN(n6007) );
  OR2_X1 U5678 ( .A1(n6007), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6020) );
  NAND2_X1 U5679 ( .A1(n5687), .A2(n5686), .ZN(n5975) );
  INV_X1 U5680 ( .A(n5960), .ZN(n5687) );
  NAND2_X1 U5681 ( .A1(n8484), .A2(n8886), .ZN(n8673) );
  OR2_X1 U5682 ( .A1(n8666), .A2(n5221), .ZN(n5220) );
  INV_X1 U5683 ( .A(n8674), .ZN(n5218) );
  NAND2_X1 U5684 ( .A1(n5105), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6668) );
  INV_X1 U5685 ( .A(n6559), .ZN(n5105) );
  XNOR2_X1 U5686 ( .A(n5083), .B(n6652), .ZN(n6653) );
  NAND2_X1 U5687 ( .A1(n10496), .A2(n10497), .ZN(n10501) );
  NAND2_X1 U5688 ( .A1(n6668), .A2(n6667), .ZN(n10494) );
  OAI22_X1 U5689 ( .A1(n10489), .A2(n6653), .B1(n6652), .B2(n5083), .ZN(n10508) );
  OR2_X1 U5690 ( .A1(n6673), .A2(n6672), .ZN(n10515) );
  OR2_X1 U5691 ( .A1(n5774), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5804) );
  INV_X1 U5692 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U5693 ( .A1(n5085), .A2(n6658), .ZN(n6659) );
  NAND2_X1 U5694 ( .A1(n5087), .A2(n5086), .ZN(n5085) );
  INV_X1 U5695 ( .A(n10551), .ZN(n5086) );
  NAND2_X1 U5696 ( .A1(n10555), .A2(n6644), .ZN(n6646) );
  NAND2_X1 U5697 ( .A1(n7162), .A2(n7163), .ZN(n7164) );
  NOR2_X1 U5698 ( .A1(n7385), .A2(n7384), .ZN(n7454) );
  AND2_X1 U5699 ( .A1(n7443), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5501) );
  NAND2_X1 U5700 ( .A1(n5503), .A2(n5029), .ZN(n5502) );
  INV_X1 U5701 ( .A(n7376), .ZN(n5503) );
  NOR2_X1 U5702 ( .A1(n7454), .A2(n5096), .ZN(n7723) );
  NAND2_X1 U5703 ( .A1(n7445), .A2(n5134), .ZN(n5132) );
  OAI21_X1 U5704 ( .B1(n7385), .B2(n5091), .A(n5090), .ZN(n10576) );
  NAND2_X1 U5705 ( .A1(n5093), .A2(n5095), .ZN(n5090) );
  NAND2_X1 U5706 ( .A1(n5092), .A2(n5095), .ZN(n5091) );
  INV_X1 U5707 ( .A(n7721), .ZN(n5095) );
  NAND2_X1 U5708 ( .A1(n10576), .A2(n10577), .ZN(n10575) );
  AND3_X1 U5709 ( .A1(n5112), .A2(n5110), .A3(n5036), .ZN(n7909) );
  NAND2_X1 U5710 ( .A1(n7916), .A2(n7917), .ZN(n7918) );
  AOI21_X1 U5711 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8911), .A(n8906), .ZN(
        n8926) );
  NAND2_X1 U5712 ( .A1(n8932), .A2(n8933), .ZN(n8934) );
  NAND2_X1 U5713 ( .A1(n8934), .A2(n8935), .ZN(n8953) );
  NAND2_X1 U5714 ( .A1(n8962), .A2(n8963), .ZN(n8982) );
  XNOR2_X1 U5715 ( .A(n8973), .B(n8984), .ZN(n8955) );
  NAND2_X1 U5716 ( .A1(n8953), .A2(n5201), .ZN(n8973) );
  OR2_X1 U5717 ( .A1(n8954), .A2(n9211), .ZN(n5201) );
  NAND2_X1 U5718 ( .A1(n8478), .A2(n8667), .ZN(n8660) );
  OR2_X1 U5719 ( .A1(n6117), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8191) );
  OAI21_X1 U5720 ( .B1(n5471), .B2(n5473), .A(n6299), .ZN(n5470) );
  NOR2_X1 U5721 ( .A1(n6298), .A2(n6297), .ZN(n6299) );
  NAND2_X1 U5722 ( .A1(n5475), .A2(n5479), .ZN(n5471) );
  INV_X1 U5723 ( .A(n5476), .ZN(n5475) );
  OAI21_X1 U5724 ( .B1(n8743), .B2(n4950), .A(n10611), .ZN(n5476) );
  OR2_X1 U5725 ( .A1(n6270), .A2(n6269), .ZN(n6271) );
  NAND2_X1 U5726 ( .A1(n5050), .A2(n9524), .ZN(n6093) );
  NAND2_X1 U5727 ( .A1(n5691), .A2(n9517), .ZN(n6095) );
  INV_X1 U5728 ( .A(n6093), .ZN(n5691) );
  OR2_X1 U5729 ( .A1(n5288), .A2(n8637), .ZN(n5286) );
  NOR2_X1 U5730 ( .A1(n5492), .A2(n5289), .ZN(n5288) );
  INV_X1 U5731 ( .A(n6162), .ZN(n5289) );
  NAND2_X1 U5732 ( .A1(n5054), .A2(n5057), .ZN(n9117) );
  OR2_X1 U5733 ( .A1(n7962), .A2(n5060), .ZN(n5054) );
  NAND2_X1 U5734 ( .A1(n5056), .A2(n4989), .ZN(n9118) );
  AND2_X1 U5735 ( .A1(n9116), .A2(n9114), .ZN(n6042) );
  NAND2_X1 U5736 ( .A1(n7961), .A2(n5983), .ZN(n8100) );
  NAND2_X1 U5737 ( .A1(n8100), .A2(n8099), .ZN(n8098) );
  NAND2_X1 U5738 ( .A1(n7962), .A2(n8594), .ZN(n7961) );
  OR2_X1 U5739 ( .A1(n5944), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5960) );
  NAND2_X1 U5740 ( .A1(n5685), .A2(n5684), .ZN(n5944) );
  INV_X1 U5741 ( .A(n5928), .ZN(n5685) );
  NAND2_X1 U5742 ( .A1(n5049), .A2(n9515), .ZN(n5928) );
  INV_X1 U5743 ( .A(n5049), .ZN(n5913) );
  AND2_X1 U5744 ( .A1(n5901), .A2(n6145), .ZN(n8497) );
  AOI21_X1 U5745 ( .B1(n5465), .B2(n5467), .A(n4988), .ZN(n5463) );
  OR2_X1 U5746 ( .A1(n5880), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5895) );
  OAI21_X1 U5747 ( .B1(n7360), .B2(n5467), .A(n5465), .ZN(n7535) );
  NAND2_X1 U5748 ( .A1(n5683), .A2(n5682), .ZN(n5880) );
  INV_X1 U5749 ( .A(n5867), .ZN(n5683) );
  NAND2_X1 U5750 ( .A1(n6142), .A2(n8557), .ZN(n7422) );
  NAND2_X1 U5751 ( .A1(n5681), .A2(n5680), .ZN(n5851) );
  INV_X1 U5752 ( .A(n5837), .ZN(n5681) );
  OR2_X1 U5753 ( .A1(n5851), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5867) );
  AND2_X1 U5754 ( .A1(n5075), .A2(n5074), .ZN(n7290) );
  OR2_X1 U5755 ( .A1(n5489), .A2(n8903), .ZN(n5076) );
  NAND2_X1 U5756 ( .A1(n5679), .A2(n5678), .ZN(n5816) );
  INV_X1 U5757 ( .A(n5809), .ZN(n5679) );
  OR2_X1 U5758 ( .A1(n5816), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5837) );
  NAND2_X1 U5759 ( .A1(n9500), .A2(n9523), .ZN(n5809) );
  AND2_X1 U5760 ( .A1(n8528), .A2(n8535), .ZN(n8486) );
  INV_X1 U5761 ( .A(n6991), .ZN(n8512) );
  OR2_X1 U5762 ( .A1(n6134), .A2(n6923), .ZN(n6989) );
  NAND2_X1 U5763 ( .A1(n8477), .A2(n8476), .ZN(n8480) );
  NAND2_X1 U5764 ( .A1(n5959), .A2(n5958), .ZN(n8698) );
  OR2_X1 U5765 ( .A1(n8032), .A2(n6046), .ZN(n5959) );
  INV_X1 U5766 ( .A(n6885), .ZN(n10651) );
  NAND2_X1 U5767 ( .A1(n5072), .A2(n5071), .ZN(n5307) );
  NOR2_X1 U5768 ( .A1(n8475), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5306) );
  CLKBUF_X1 U5769 ( .A(n6125), .Z(n6126) );
  XNOR2_X1 U5770 ( .A(n5826), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6940) );
  NAND2_X1 U5771 ( .A1(n8029), .A2(n8028), .ZN(n8351) );
  OR2_X1 U5772 ( .A1(n8027), .A2(n8301), .ZN(n8029) );
  AND2_X1 U5773 ( .A1(n8113), .A2(n8083), .ZN(n8088) );
  NAND2_X1 U5774 ( .A1(n5342), .A2(n9576), .ZN(n5341) );
  INV_X1 U5775 ( .A(n9293), .ZN(n8416) );
  NAND2_X1 U5776 ( .A1(n5353), .A2(n5352), .ZN(n7222) );
  AND2_X1 U5777 ( .A1(n7200), .A2(n7199), .ZN(n5352) );
  NOR2_X1 U5778 ( .A1(n7548), .A2(n7547), .ZN(n7568) );
  NAND2_X1 U5779 ( .A1(n5334), .A2(n8390), .ZN(n5333) );
  NAND2_X1 U5780 ( .A1(n8114), .A2(n8113), .ZN(n8115) );
  AND2_X1 U5781 ( .A1(n7568), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7577) );
  AND2_X1 U5782 ( .A1(n8086), .A2(n7999), .ZN(n8003) );
  INV_X1 U5783 ( .A(n6808), .ZN(n6811) );
  NOR2_X1 U5784 ( .A1(n7803), .A2(n7802), .ZN(n8036) );
  INV_X1 U5785 ( .A(n8367), .ZN(n8368) );
  NAND2_X1 U5786 ( .A1(n9827), .A2(n5416), .ZN(n9829) );
  NAND2_X1 U5787 ( .A1(n5418), .A2(n5417), .ZN(n5416) );
  AOI21_X1 U5788 ( .B1(n9825), .B2(n5419), .A(n9826), .ZN(n5418) );
  NOR4_X1 U5789 ( .A1(n9939), .A2(n9832), .A3(n9708), .A4(n9707), .ZN(n9837)
         );
  OR2_X1 U5790 ( .A1(n6524), .A2(n6523), .ZN(n5136) );
  NOR2_X1 U5791 ( .A1(n6575), .A2(n6574), .ZN(n6576) );
  NOR2_X1 U5792 ( .A1(n5140), .A2(n7250), .ZN(n7251) );
  AND2_X1 U5793 ( .A1(n7631), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5140) );
  NAND2_X1 U5794 ( .A1(n7251), .A2(n7252), .ZN(n7432) );
  XNOR2_X1 U5795 ( .A(n9995), .B(n10003), .ZN(n8065) );
  NOR2_X1 U5796 ( .A1(n8062), .A2(n5143), .ZN(n9995) );
  AND2_X1 U5797 ( .A1(n8063), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5143) );
  NOR2_X1 U5798 ( .A1(n8065), .A2(n8035), .ZN(n9996) );
  NOR2_X1 U5799 ( .A1(n10006), .A2(n10005), .ZN(n10009) );
  AOI21_X1 U5800 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n10020), .A(n10015), .ZN(
        n10016) );
  AND2_X1 U5801 ( .A1(n10092), .A2(n5028), .ZN(n5356) );
  NOR2_X1 U5802 ( .A1(n10111), .A2(n10272), .ZN(n10096) );
  INV_X1 U5803 ( .A(n10107), .ZN(n10109) );
  INV_X1 U5804 ( .A(n10089), .ZN(n10090) );
  NAND2_X1 U5805 ( .A1(n9850), .A2(n9862), .ZN(n10107) );
  INV_X1 U5806 ( .A(n8218), .ZN(n8305) );
  AND2_X1 U5807 ( .A1(n9847), .A2(n10086), .ZN(n10089) );
  INV_X1 U5808 ( .A(n6702), .ZN(n6703) );
  INV_X1 U5809 ( .A(n10314), .ZN(n8337) );
  NAND2_X1 U5810 ( .A1(n10154), .A2(n10163), .ZN(n10155) );
  AND2_X1 U5811 ( .A1(n9714), .A2(n9713), .ZN(n10168) );
  AND2_X1 U5812 ( .A1(n9930), .A2(n9805), .ZN(n10188) );
  OR2_X1 U5813 ( .A1(n10345), .A2(n10335), .ZN(n9929) );
  NAND2_X1 U5814 ( .A1(n8234), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8233) );
  NOR2_X1 U5815 ( .A1(n10345), .A2(n5267), .ZN(n5265) );
  AOI21_X1 U5816 ( .B1(n10247), .B2(n5365), .A(n5362), .ZN(n5361) );
  NAND2_X1 U5817 ( .A1(n5363), .A2(n8240), .ZN(n5362) );
  OR2_X1 U5818 ( .A1(n10349), .A2(n9955), .ZN(n8240) );
  NAND2_X1 U5819 ( .A1(n10254), .A2(n5268), .ZN(n10238) );
  AND3_X1 U5820 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .A3(n8132), .ZN(n8219) );
  INV_X1 U5821 ( .A(n8037), .ZN(n8132) );
  AND2_X1 U5822 ( .A1(n8128), .A2(n9790), .ZN(n10254) );
  OR2_X1 U5823 ( .A1(n8032), .A2(n8301), .ZN(n8034) );
  INV_X1 U5824 ( .A(n9702), .ZN(n8258) );
  OR2_X1 U5825 ( .A1(n10816), .A2(n8351), .ZN(n10817) );
  AND2_X1 U5826 ( .A1(n9911), .A2(n9912), .ZN(n10821) );
  OR2_X1 U5827 ( .A1(n7643), .A2(n7436), .ZN(n7803) );
  OR2_X1 U5828 ( .A1(n7641), .A2(n7640), .ZN(n7643) );
  NAND2_X1 U5829 ( .A1(n5440), .A2(n5443), .ZN(n5438) );
  NAND2_X1 U5830 ( .A1(n7675), .A2(n9772), .ZN(n7681) );
  OAI211_X1 U5831 ( .C1(n4954), .C2(n5386), .A(n4990), .B(n5385), .ZN(n7810)
         );
  NOR2_X1 U5832 ( .A1(n5386), .A2(n5383), .ZN(n5382) );
  AND2_X1 U5833 ( .A1(n9773), .A2(n9767), .ZN(n9680) );
  NAND2_X1 U5834 ( .A1(n7635), .A2(n9757), .ZN(n7675) );
  OR2_X1 U5835 ( .A1(n7518), .A2(n7517), .ZN(n7548) );
  AND2_X1 U5836 ( .A1(n7592), .A2(n9751), .ZN(n10718) );
  NAND2_X1 U5837 ( .A1(n7490), .A2(n4953), .ZN(n10678) );
  NAND2_X1 U5838 ( .A1(n4956), .A2(n7490), .ZN(n10713) );
  INV_X1 U5839 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6446) );
  INV_X1 U5840 ( .A(n10683), .ZN(n7499) );
  OR2_X1 U5841 ( .A1(n9963), .A2(n10660), .ZN(n10684) );
  NAND2_X1 U5842 ( .A1(n9746), .A2(n10687), .ZN(n10683) );
  AND2_X1 U5843 ( .A1(n7490), .A2(n10660), .ZN(n10679) );
  AND2_X1 U5844 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n7205) );
  NAND2_X1 U5845 ( .A1(n5254), .A2(n7412), .ZN(n7339) );
  INV_X1 U5846 ( .A(n7135), .ZN(n5254) );
  OAI211_X1 U5847 ( .C1(n7228), .C2(n6825), .A(n6824), .B(n6823), .ZN(n7472)
         );
  NAND2_X1 U5848 ( .A1(n6972), .A2(n6971), .ZN(n7135) );
  NOR2_X1 U5849 ( .A1(n9968), .A2(n9890), .ZN(n7175) );
  NAND2_X1 U5850 ( .A1(n6737), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6738) );
  INV_X1 U5851 ( .A(n10275), .ZN(n5259) );
  INV_X1 U5852 ( .A(n10093), .ZN(n10288) );
  NAND2_X1 U5853 ( .A1(n8278), .A2(n8277), .ZN(n10308) );
  NAND2_X1 U5854 ( .A1(n8276), .A2(n9695), .ZN(n8278) );
  OR2_X1 U5855 ( .A1(n8688), .A2(n9868), .ZN(n10825) );
  INV_X1 U5856 ( .A(n7472), .ZN(n6972) );
  OR2_X1 U5857 ( .A1(n9945), .A2(n6965), .ZN(n10820) );
  NAND2_X1 U5858 ( .A1(n10831), .A2(n10673), .ZN(n10811) );
  NAND2_X1 U5859 ( .A1(n7264), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6799) );
  AND2_X1 U5860 ( .A1(n6413), .A2(n6412), .ZN(n6723) );
  XNOR2_X1 U5861 ( .A(n8173), .B(n8172), .ZN(n9662) );
  OAI21_X1 U5862 ( .B1(n8470), .B2(n8469), .A(n8168), .ZN(n8173) );
  XNOR2_X1 U5863 ( .A(n5725), .B(n5724), .ZN(n8271) );
  AND2_X1 U5864 ( .A1(n5723), .A2(n5722), .ZN(n5725) );
  NAND2_X1 U5865 ( .A1(n6387), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6388) );
  NAND2_X1 U5866 ( .A1(n5954), .A2(n5620), .ZN(n5969) );
  NAND2_X1 U5867 ( .A1(n5939), .A2(n5615), .ZN(n5952) );
  AND2_X1 U5868 ( .A1(n5620), .A2(n5619), .ZN(n5951) );
  AND2_X1 U5869 ( .A1(n5615), .A2(n5614), .ZN(n5936) );
  AOI21_X1 U5870 ( .B1(n5423), .B2(n5425), .A(n5422), .ZN(n5421) );
  NAND2_X1 U5871 ( .A1(n5159), .A2(n5160), .ZN(n5158) );
  NAND2_X1 U5872 ( .A1(n5160), .A2(n5157), .ZN(n5156) );
  AND2_X1 U5873 ( .A1(n5611), .A2(n5610), .ZN(n5920) );
  CLKBUF_X1 U5874 ( .A(n6397), .Z(n6398) );
  AND2_X1 U5875 ( .A1(n5844), .A2(n5596), .ZN(n5829) );
  NAND2_X1 U5876 ( .A1(n5830), .A2(n5829), .ZN(n5845) );
  AND2_X1 U5877 ( .A1(n5593), .A2(n5592), .ZN(n5823) );
  AND2_X1 U5878 ( .A1(n5589), .A2(n5588), .ZN(n5800) );
  NAND2_X1 U5879 ( .A1(n5787), .A2(n5786), .ZN(n5789) );
  NAND2_X1 U5880 ( .A1(n5779), .A2(n5580), .ZN(n5787) );
  NAND2_X1 U5881 ( .A1(n5756), .A2(n5574), .ZN(n5777) );
  AND2_X1 U5882 ( .A1(n5580), .A2(n5579), .ZN(n5776) );
  NAND2_X1 U5883 ( .A1(n5543), .A2(n5541), .ZN(n8754) );
  NAND2_X1 U5884 ( .A1(n5943), .A2(n5942), .ZN(n8578) );
  OR2_X1 U5885 ( .A1(n8027), .A2(n6046), .ZN(n5943) );
  INV_X1 U5886 ( .A(n6864), .ZN(n5520) );
  AND2_X1 U5887 ( .A1(n6946), .A2(n6761), .ZN(n5521) );
  NAND2_X1 U5888 ( .A1(n6946), .A2(n6761), .ZN(n6863) );
  INV_X1 U5889 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9500) );
  NAND2_X1 U5890 ( .A1(n6240), .A2(n6239), .ZN(n8750) );
  AND2_X1 U5891 ( .A1(n5550), .A2(n5549), .ZN(n7612) );
  AOI21_X1 U5892 ( .B1(n6923), .B2(n6751), .A(n6757), .ZN(n6955) );
  NAND2_X1 U5893 ( .A1(n6092), .A2(n6091), .ZN(n9171) );
  NAND2_X1 U5894 ( .A1(n5148), .A2(n5149), .ZN(n7085) );
  OR2_X1 U5895 ( .A1(n8703), .A2(n8810), .ZN(n8704) );
  AND2_X1 U5896 ( .A1(n5172), .A2(n5170), .ZN(n7699) );
  NAND2_X1 U5897 ( .A1(n5172), .A2(n5544), .ZN(n7613) );
  NAND2_X1 U5898 ( .A1(n5926), .A2(n5925), .ZN(n7948) );
  OR2_X1 U5899 ( .A1(n7794), .A2(n6046), .ZN(n5926) );
  AND2_X1 U5900 ( .A1(n6787), .A2(n6786), .ZN(n8876) );
  NAND2_X1 U5901 ( .A1(n5720), .A2(n5719), .ZN(n8868) );
  NAND2_X1 U5902 ( .A1(n8697), .A2(n8696), .ZN(n8873) );
  NAND2_X1 U5903 ( .A1(n5706), .A2(n5705), .ZN(n8890) );
  NAND4_X1 U5904 ( .A1(n5765), .A2(n5764), .A3(n5763), .A4(n5762), .ZN(n8905)
         );
  OR2_X1 U5905 ( .A1(n5760), .A2(n5761), .ZN(n5763) );
  AND2_X1 U5906 ( .A1(n5698), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5460) );
  OR2_X1 U5907 ( .A1(n6775), .A2(n6343), .ZN(n8989) );
  INV_X1 U5908 ( .A(n5087), .ZN(n10552) );
  AND2_X1 U5909 ( .A1(n5128), .A2(n4972), .ZN(n7146) );
  AND2_X1 U5910 ( .A1(n6926), .A2(n6925), .ZN(n7142) );
  NAND2_X1 U5911 ( .A1(n7443), .A2(n5502), .ZN(n7377) );
  AND2_X1 U5912 ( .A1(n5501), .A2(n5502), .ZN(n7444) );
  NAND2_X1 U5913 ( .A1(n5133), .A2(n5132), .ZN(n7709) );
  NAND2_X1 U5914 ( .A1(n5513), .A2(n7710), .ZN(n10582) );
  XNOR2_X1 U5915 ( .A(n7915), .B(n7910), .ZN(n7779) );
  XNOR2_X1 U5916 ( .A(n7909), .B(n7910), .ZN(n7775) );
  NOR2_X1 U5917 ( .A1(n7775), .A2(n7776), .ZN(n7911) );
  OAI21_X1 U5918 ( .B1(n7775), .B2(n5515), .A(n5514), .ZN(n8906) );
  NAND2_X1 U5919 ( .A1(n5516), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5515) );
  NAND2_X1 U5920 ( .A1(n7912), .A2(n5516), .ZN(n5514) );
  INV_X1 U5921 ( .A(n7914), .ZN(n5516) );
  XNOR2_X1 U5922 ( .A(n8931), .B(n8927), .ZN(n8910) );
  NOR2_X1 U5923 ( .A1(n8907), .A2(n5962), .ZN(n8928) );
  NAND2_X1 U5924 ( .A1(n5124), .A2(n5510), .ZN(n8951) );
  NAND2_X1 U5925 ( .A1(n5118), .A2(n5117), .ZN(n8952) );
  NAND2_X1 U5926 ( .A1(n4962), .A2(n5124), .ZN(n5117) );
  AND2_X1 U5927 ( .A1(n5119), .A2(n5122), .ZN(n5118) );
  NAND2_X1 U5928 ( .A1(n8994), .A2(n5109), .ZN(n5108) );
  NAND2_X1 U5929 ( .A1(n9006), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5109) );
  XNOR2_X1 U5930 ( .A(n5206), .B(n9009), .ZN(n5205) );
  NAND2_X1 U5931 ( .A1(n5208), .A2(n5207), .ZN(n5206) );
  NAND2_X1 U5932 ( .A1(n9006), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5207) );
  NAND2_X1 U5933 ( .A1(n9008), .A2(n9007), .ZN(n5208) );
  NAND2_X1 U5934 ( .A1(n5204), .A2(n5203), .ZN(n5202) );
  NAND2_X1 U5935 ( .A1(n10571), .A2(n9011), .ZN(n5203) );
  INV_X1 U5936 ( .A(n9010), .ZN(n5204) );
  OAI211_X1 U5937 ( .C1(n5477), .C2(n5472), .A(n5469), .B(n5468), .ZN(n9024)
         );
  NAND2_X1 U5938 ( .A1(n5474), .A2(n5475), .ZN(n5472) );
  NAND2_X1 U5939 ( .A1(n5477), .A2(n4985), .ZN(n5468) );
  INV_X1 U5940 ( .A(n5470), .ZN(n5469) );
  OAI21_X1 U5941 ( .B1(n6133), .B2(n9145), .A(n6132), .ZN(n9032) );
  NOR2_X1 U5942 ( .A1(n6131), .A2(n6130), .ZN(n6132) );
  NOR2_X1 U5943 ( .A1(n9148), .A2(n8790), .ZN(n6130) );
  INV_X1 U5944 ( .A(n8819), .ZN(n9179) );
  NAND2_X1 U5945 ( .A1(n5290), .A2(n5288), .ZN(n9068) );
  NAND2_X1 U5946 ( .A1(n5290), .A2(n6162), .ZN(n9069) );
  NAND2_X1 U5947 ( .A1(n5493), .A2(n5494), .ZN(n9061) );
  OAI21_X1 U5948 ( .B1(n9084), .B2(n6070), .A(n8631), .ZN(n9073) );
  NAND2_X1 U5949 ( .A1(n6061), .A2(n6060), .ZN(n9184) );
  NAND2_X1 U5950 ( .A1(n5300), .A2(n8615), .ZN(n9096) );
  NAND2_X1 U5951 ( .A1(n6033), .A2(n6032), .ZN(n9194) );
  NAND2_X1 U5952 ( .A1(n6157), .A2(n6156), .ZN(n9115) );
  NAND2_X1 U5953 ( .A1(n5303), .A2(n6152), .ZN(n9153) );
  NAND2_X1 U5954 ( .A1(n5991), .A2(n5990), .ZN(n9206) );
  NAND2_X1 U5955 ( .A1(n7965), .A2(n6151), .ZN(n8097) );
  OAI21_X1 U5956 ( .B1(n7857), .B2(n5068), .A(n5066), .ZN(n7870) );
  OAI21_X1 U5957 ( .B1(n6147), .B2(n5277), .A(n5274), .ZN(n7942) );
  NAND2_X1 U5958 ( .A1(n7863), .A2(n8577), .ZN(n7862) );
  NAND2_X1 U5959 ( .A1(n6147), .A2(n8575), .ZN(n7863) );
  NAND2_X1 U5960 ( .A1(n5892), .A2(n5891), .ZN(n10778) );
  NAND2_X1 U5961 ( .A1(n5464), .A2(n8493), .ZN(n7419) );
  AND2_X1 U5962 ( .A1(n10626), .A2(n10625), .ZN(n9161) );
  NAND2_X1 U5963 ( .A1(n7555), .A2(n8473), .ZN(n5215) );
  NAND2_X1 U5964 ( .A1(n5487), .A2(n5489), .ZN(n7100) );
  OR2_X1 U5965 ( .A1(n7008), .A2(n6046), .ZN(n5781) );
  INV_X1 U5966 ( .A(n8481), .ZN(n8484) );
  INV_X1 U5967 ( .A(n8480), .ZN(n9222) );
  INV_X1 U5968 ( .A(n8750), .ZN(n9027) );
  AOI21_X1 U5969 ( .B1(n10632), .B2(n9029), .A(n9024), .ZN(n6302) );
  AOI21_X1 U5970 ( .B1(n9036), .B2(n10632), .A(n9032), .ZN(n6232) );
  INV_X1 U5971 ( .A(n8868), .ZN(n9226) );
  AOI21_X1 U5972 ( .B1(n5531), .B2(n5672), .A(n5672), .ZN(n5528) );
  NAND2_X1 U5973 ( .A1(n5527), .A2(n5531), .ZN(n6110) );
  INV_X1 U5974 ( .A(n10520), .ZN(n6670) );
  INV_X1 U5975 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U5976 ( .A1(n5507), .A2(n5509), .ZN(n10503) );
  NAND2_X1 U5977 ( .A1(n5752), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n5509) );
  NAND2_X1 U5978 ( .A1(n5327), .A2(n7749), .ZN(n8194) );
  NAND2_X1 U5979 ( .A1(n5323), .A2(n5039), .ZN(n5327) );
  NAND2_X1 U5980 ( .A1(n5354), .A2(n7841), .ZN(n7842) );
  INV_X1 U5981 ( .A(n5355), .ZN(n5354) );
  NAND2_X1 U5982 ( .A1(n5333), .A2(n5332), .ZN(n9606) );
  NAND2_X1 U5983 ( .A1(n5331), .A2(n5328), .ZN(n9559) );
  AND2_X1 U5984 ( .A1(n8401), .A2(n5329), .ZN(n5328) );
  AND2_X1 U5985 ( .A1(n9560), .A2(n9561), .ZN(n8401) );
  NAND2_X1 U5986 ( .A1(n9596), .A2(n8434), .ZN(n9568) );
  INV_X1 U5987 ( .A(n9957), .ZN(n10824) );
  AND2_X1 U5988 ( .A1(n5339), .A2(n9575), .ZN(n9579) );
  NOR2_X1 U5989 ( .A1(n9652), .A2(n9576), .ZN(n5339) );
  NAND2_X1 U5990 ( .A1(n5353), .A2(n7199), .ZN(n7202) );
  INV_X1 U5991 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U5992 ( .A1(n6797), .A2(n10407), .ZN(n5255) );
  INV_X1 U5993 ( .A(n9958), .ZN(n10786) );
  NAND4_X1 U5994 ( .A1(n6452), .A2(n6451), .A3(n6450), .A4(n6449), .ZN(n8200)
         );
  INV_X1 U5995 ( .A(n5142), .ZN(n9969) );
  NAND2_X1 U5996 ( .A1(n9973), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5141) );
  OR2_X1 U5997 ( .A1(n6689), .A2(n6490), .ZN(n9990) );
  INV_X1 U5998 ( .A(n5138), .ZN(n6588) );
  AND2_X1 U5999 ( .A1(n5138), .A2(n5137), .ZN(n6524) );
  NAND2_X1 U6000 ( .A1(n7186), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5137) );
  INV_X1 U6001 ( .A(n5136), .ZN(n6522) );
  AOI21_X1 U6002 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n7186), .A(n6493), .ZN(
        n6527) );
  AND2_X1 U6003 ( .A1(n5136), .A2(n5135), .ZN(n6512) );
  NAND2_X1 U6004 ( .A1(n7223), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5135) );
  AOI21_X1 U6005 ( .B1(n7223), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6525), .ZN(
        n6515) );
  NOR2_X1 U6006 ( .A1(n6570), .A2(n5031), .ZN(n6572) );
  NAND2_X1 U6007 ( .A1(n6572), .A2(n6571), .ZN(n6868) );
  NOR2_X1 U6008 ( .A1(n7071), .A2(n5139), .ZN(n7073) );
  AND2_X1 U6009 ( .A1(n7564), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5139) );
  NOR2_X1 U6010 ( .A1(n7072), .A2(n7073), .ZN(n7250) );
  AOI21_X1 U6011 ( .B1(n7564), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7074), .ZN(
        n7077) );
  AOI21_X1 U6012 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n7795), .A(n7658), .ZN(
        n7659) );
  INV_X1 U6013 ( .A(n10267), .ZN(n10078) );
  NAND2_X1 U6014 ( .A1(n9699), .A2(n9698), .ZN(n10084) );
  AOI211_X1 U6015 ( .C1(n10111), .C2(n10272), .A(n10096), .B(n10257), .ZN(
        n10276) );
  AOI211_X1 U6016 ( .C1(n10284), .C2(n10113), .A(n10257), .B(n10112), .ZN(
        n10282) );
  NAND2_X1 U6017 ( .A1(n8288), .A2(n9695), .ZN(n8290) );
  NAND2_X1 U6018 ( .A1(n5373), .A2(n5375), .ZN(n10138) );
  OR2_X1 U6019 ( .A1(n8266), .A2(n5378), .ZN(n5373) );
  NAND2_X1 U6020 ( .A1(n8341), .A2(n9841), .ZN(n10136) );
  AND2_X1 U6021 ( .A1(n8341), .A2(n5446), .ZN(n10135) );
  NAND2_X1 U6022 ( .A1(n5374), .A2(n8269), .ZN(n8336) );
  NAND2_X1 U6023 ( .A1(n8266), .A2(n5380), .ZN(n5374) );
  NAND2_X1 U6024 ( .A1(n8266), .A2(n8265), .ZN(n10152) );
  NAND2_X1 U6025 ( .A1(n8255), .A2(n8254), .ZN(n10178) );
  INV_X1 U6026 ( .A(n10227), .ZN(n10335) );
  INV_X1 U6027 ( .A(n5364), .ZN(n10217) );
  AOI21_X1 U6028 ( .B1(n10247), .B2(n5369), .A(n5367), .ZN(n5364) );
  INV_X1 U6029 ( .A(n10355), .ZN(n10244) );
  AOI21_X1 U6030 ( .B1(n10247), .B2(n8213), .A(n5557), .ZN(n10232) );
  INV_X1 U6031 ( .A(n9788), .ZN(n10371) );
  INV_X1 U6032 ( .A(n5398), .ZN(n8123) );
  NAND2_X1 U6033 ( .A1(n7797), .A2(n7796), .ZN(n8112) );
  OR2_X1 U6034 ( .A1(n7794), .A2(n8301), .ZN(n7797) );
  NAND2_X1 U6035 ( .A1(n5384), .A2(n5393), .ZN(n7684) );
  NAND2_X1 U6036 ( .A1(n5387), .A2(n4954), .ZN(n5384) );
  NAND2_X1 U6037 ( .A1(n5387), .A2(n5389), .ZN(n7637) );
  INV_X1 U6038 ( .A(n10732), .ZN(n10845) );
  CLKBUF_X1 U6039 ( .A(n6417), .Z(n8688) );
  NAND2_X1 U6040 ( .A1(n5558), .A2(n5661), .ZN(n8302) );
  CLKBUF_X1 U6041 ( .A(n6418), .Z(n10074) );
  XNOR2_X1 U6042 ( .A(n6073), .B(n6072), .ZN(n8267) );
  NAND2_X1 U6043 ( .A1(n5635), .A2(n5634), .ZN(n6044) );
  INV_X1 U6044 ( .A(n6326), .ZN(n6603) );
  OR2_X1 U6045 ( .A1(n5998), .A2(n5556), .ZN(n5999) );
  NOR2_X1 U6046 ( .A1(n5173), .A2(n5400), .ZN(n5998) );
  INV_X1 U6047 ( .A(n5176), .ZN(n5173) );
  NAND2_X1 U6048 ( .A1(n5426), .A2(n5425), .ZN(n5906) );
  NAND2_X1 U6049 ( .A1(n5426), .A2(n5427), .ZN(n5905) );
  NAND2_X1 U6050 ( .A1(n5164), .A2(n4973), .ZN(n5162) );
  OAI21_X1 U6051 ( .B1(n5824), .B2(n5823), .A(n5822), .ZN(n7263) );
  NOR2_X1 U6052 ( .A1(n6362), .A2(n5454), .ZN(n6375) );
  NAND2_X1 U6053 ( .A1(n6309), .A2(n5456), .ZN(n5454) );
  XNOR2_X1 U6054 ( .A(n6352), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9988) );
  NAND2_X1 U6055 ( .A1(n8849), .A2(n5551), .ZN(n7089) );
  AND2_X1 U6056 ( .A1(n7710), .A2(n5113), .ZN(n7713) );
  AND2_X1 U6057 ( .A1(n5103), .A2(n5099), .ZN(n8991) );
  NAND2_X1 U6058 ( .A1(n9012), .A2(n5106), .ZN(P2_U3201) );
  NAND2_X1 U6059 ( .A1(n5107), .A2(n10583), .ZN(n5106) );
  AOI21_X1 U6060 ( .B1(n5205), .B2(n10580), .A(n5202), .ZN(n9012) );
  XNOR2_X1 U6061 ( .A(n5108), .B(n9000), .ZN(n5107) );
  AOI21_X1 U6062 ( .B1(n9019), .B2(n9237), .A(n6288), .ZN(n6289) );
  NOR2_X1 U6063 ( .A1(n10785), .A2(n6287), .ZN(n6288) );
  NAND2_X1 U6064 ( .A1(n5348), .A2(n9651), .ZN(n5345) );
  AND2_X1 U6065 ( .A1(n10154), .A2(n4957), .ZN(n4948) );
  INV_X1 U6066 ( .A(n5774), .ZN(n5195) );
  OR2_X1 U6067 ( .A1(n5668), .A2(n5667), .ZN(n4949) );
  OAI21_X1 U6068 ( .B1(n5402), .B2(n5401), .A(n4998), .ZN(n5400) );
  NOR2_X1 U6069 ( .A1(n8429), .A2(n8428), .ZN(n8433) );
  INV_X1 U6070 ( .A(n9960), .ZN(n10787) );
  AND2_X1 U6071 ( .A1(n6797), .A2(n8169), .ZN(n7264) );
  INV_X1 U6072 ( .A(n7264), .ZN(n7228) );
  NAND2_X1 U6073 ( .A1(n5048), .A2(n9041), .ZN(n4950) );
  INV_X2 U6074 ( .A(n5745), .ZN(n5459) );
  NOR2_X1 U6075 ( .A1(n8841), .A2(n8713), .ZN(n4951) );
  AND2_X1 U6076 ( .A1(n5547), .A2(n5546), .ZN(n4952) );
  XNOR2_X1 U6077 ( .A(n8801), .B(n8810), .ZN(n8594) );
  INV_X1 U6078 ( .A(n8594), .ZN(n5059) );
  AND2_X1 U6079 ( .A1(n10660), .A2(n10680), .ZN(n4953) );
  AND2_X1 U6080 ( .A1(n5389), .A2(n9677), .ZN(n4954) );
  OR2_X1 U6081 ( .A1(n8709), .A2(n9132), .ZN(n4955) );
  INV_X1 U6082 ( .A(n8740), .ZN(n5048) );
  AND2_X1 U6083 ( .A1(n4953), .A2(n5271), .ZN(n4956) );
  AND2_X1 U6084 ( .A1(n5263), .A2(n10146), .ZN(n4957) );
  AND2_X1 U6085 ( .A1(n5375), .A2(n4976), .ZN(n4958) );
  AND2_X1 U6086 ( .A1(n8634), .A2(n8631), .ZN(n4959) );
  INV_X1 U6087 ( .A(n8658), .ZN(n5222) );
  AND2_X1 U6088 ( .A1(n5405), .A2(n5984), .ZN(n4960) );
  NAND2_X1 U6089 ( .A1(n8890), .A2(n5048), .ZN(n6268) );
  NAND2_X1 U6090 ( .A1(n5659), .A2(SI_27_), .ZN(n5194) );
  NAND2_X1 U6091 ( .A1(n7738), .A2(n7737), .ZN(n4961) );
  INV_X1 U6092 ( .A(n9100), .ZN(n9095) );
  NAND2_X1 U6093 ( .A1(n6057), .A2(n6056), .ZN(n9100) );
  INV_X1 U6094 ( .A(n5267), .ZN(n5266) );
  NAND2_X1 U6095 ( .A1(n5268), .A2(n10222), .ZN(n5267) );
  AND2_X1 U6096 ( .A1(n5510), .A2(n5037), .ZN(n4962) );
  OR2_X1 U6097 ( .A1(n10533), .A2(n10566), .ZN(n4963) );
  AND2_X1 U6098 ( .A1(n5333), .A2(n5022), .ZN(n4964) );
  INV_X1 U6099 ( .A(n6127), .ZN(n8999) );
  INV_X1 U6100 ( .A(n8493), .ZN(n5467) );
  OAI21_X1 U6101 ( .B1(n7056), .B2(n5799), .A(n5798), .ZN(n7035) );
  OR2_X1 U6102 ( .A1(n8954), .A2(n5978), .ZN(n4965) );
  NAND2_X2 U6103 ( .A1(n6750), .A2(n6749), .ZN(n6751) );
  XNOR2_X1 U6104 ( .A(n6347), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9973) );
  OR2_X1 U6105 ( .A1(n5658), .A2(n5657), .ZN(n4966) );
  NAND2_X1 U6106 ( .A1(n6326), .A2(n6325), .ZN(n6334) );
  NAND2_X1 U6107 ( .A1(n7711), .A2(n7720), .ZN(n7710) );
  AND4_X1 U6108 ( .A1(n5517), .A2(n5285), .A3(n5283), .A4(n5284), .ZN(n4967)
         );
  AND2_X1 U6109 ( .A1(n5494), .A2(n5492), .ZN(n4968) );
  AND2_X1 U6110 ( .A1(n10355), .A2(n10226), .ZN(n4969) );
  NOR2_X1 U6111 ( .A1(n8650), .A2(n8649), .ZN(n4970) );
  OR2_X1 U6112 ( .A1(n8763), .A2(n9086), .ZN(n8634) );
  NAND2_X1 U6113 ( .A1(n5455), .A2(n6309), .ZN(n6360) );
  AND3_X1 U6114 ( .A1(n7024), .A2(n7023), .A3(n7022), .ZN(n4971) );
  XNOR2_X1 U6115 ( .A(n8819), .B(n9051), .ZN(n9060) );
  INV_X1 U6116 ( .A(n9060), .ZN(n5492) );
  OR2_X1 U6117 ( .A1(n7143), .A2(n7142), .ZN(n4972) );
  INV_X1 U6118 ( .A(n9757), .ZN(n5442) );
  OR2_X1 U6119 ( .A1(n5599), .A2(SI_9_), .ZN(n4973) );
  INV_X1 U6120 ( .A(n5786), .ZN(n5360) );
  NOR2_X1 U6121 ( .A1(n6675), .A2(n6650), .ZN(n4974) );
  NOR4_X1 U6122 ( .A1(n9154), .A2(n8499), .A3(n8582), .A4(n8498), .ZN(n4975)
         );
  AND2_X1 U6123 ( .A1(n8579), .A2(n8580), .ZN(n8577) );
  INV_X1 U6124 ( .A(n8577), .ZN(n5277) );
  NAND2_X1 U6125 ( .A1(n6274), .A2(n6260), .ZN(n8743) );
  NAND2_X1 U6126 ( .A1(n8098), .A2(n5997), .ZN(n9130) );
  INV_X1 U6127 ( .A(n8204), .ZN(n5271) );
  INV_X1 U6128 ( .A(n10759), .ZN(n5394) );
  OR2_X1 U6129 ( .A1(n10308), .A2(n10297), .ZN(n4976) );
  INV_X1 U6130 ( .A(n8653), .ZN(n5228) );
  AND2_X1 U6131 ( .A1(n5142), .A2(n5141), .ZN(n4977) );
  AND2_X1 U6132 ( .A1(n5294), .A2(n5295), .ZN(n4978) );
  NAND2_X1 U6133 ( .A1(n9934), .A2(n9853), .ZN(n10095) );
  INV_X1 U6134 ( .A(n10095), .ZN(n5417) );
  OR2_X1 U6135 ( .A1(n10790), .A2(n9959), .ZN(n4979) );
  NAND2_X1 U6136 ( .A1(n5436), .A2(n8268), .ZN(n10321) );
  AND3_X1 U6137 ( .A1(n6837), .A2(n6838), .A3(n6839), .ZN(n4980) );
  AND2_X1 U6138 ( .A1(n8743), .A2(n5478), .ZN(n4981) );
  AND2_X1 U6139 ( .A1(n9841), .A2(n9857), .ZN(n9811) );
  OR2_X1 U6140 ( .A1(n5325), .A2(n5324), .ZN(n4982) );
  INV_X1 U6141 ( .A(n5213), .ZN(n5741) );
  OR2_X1 U6142 ( .A1(n8573), .A2(n8655), .ZN(n4983) );
  INV_X1 U6143 ( .A(n10360), .ZN(n10262) );
  NAND2_X1 U6144 ( .A1(n8212), .A2(n8211), .ZN(n10360) );
  INV_X1 U6145 ( .A(n5997), .ZN(n5486) );
  NOR2_X1 U6146 ( .A1(n7986), .A2(n7985), .ZN(n4984) );
  AND2_X1 U6147 ( .A1(n5475), .A2(n4981), .ZN(n4985) );
  AND2_X1 U6148 ( .A1(n4959), .A2(n5497), .ZN(n4986) );
  OR2_X1 U6149 ( .A1(n6797), .A2(n7265), .ZN(n4987) );
  AND2_X1 U6150 ( .A1(n10771), .A2(n8899), .ZN(n4988) );
  AND2_X1 U6151 ( .A1(n5055), .A2(n6042), .ZN(n4989) );
  OR2_X1 U6152 ( .A1(n8011), .A2(n10756), .ZN(n4990) );
  NOR2_X1 U6153 ( .A1(n7626), .A2(n8900), .ZN(n4991) );
  OR2_X1 U6154 ( .A1(n4968), .A2(n5491), .ZN(n4992) );
  NAND2_X1 U6155 ( .A1(n6675), .A2(n6650), .ZN(n4993) );
  INV_X1 U6156 ( .A(n5428), .ZN(n5427) );
  NOR2_X1 U6157 ( .A1(n5605), .A2(SI_11_), .ZN(n5428) );
  AND2_X1 U6158 ( .A1(n10651), .A2(n8854), .ZN(n4994) );
  NAND2_X1 U6159 ( .A1(n7698), .A2(n8900), .ZN(n4995) );
  NAND2_X1 U6160 ( .A1(n5673), .A2(n5669), .ZN(n4996) );
  AND2_X1 U6161 ( .A1(n5622), .A2(n9427), .ZN(n4997) );
  OR2_X1 U6162 ( .A1(n5624), .A2(SI_17_), .ZN(n4998) );
  AND2_X1 U6163 ( .A1(n5598), .A2(n9475), .ZN(n4999) );
  INV_X1 U6164 ( .A(n5405), .ZN(n5404) );
  NOR2_X1 U6165 ( .A1(n5968), .A2(n5406), .ZN(n5405) );
  NAND2_X1 U6166 ( .A1(n5635), .A2(n5414), .ZN(n5413) );
  AND2_X1 U6167 ( .A1(n8358), .A2(n8357), .ZN(n5000) );
  NAND2_X1 U6168 ( .A1(n5717), .A2(n5715), .ZN(n5001) );
  AND4_X1 U6169 ( .A1(n5285), .A2(n5283), .A3(n5282), .A4(n5284), .ZN(n5002)
         );
  NAND2_X1 U6170 ( .A1(n9634), .A2(n9635), .ZN(n5003) );
  OR2_X1 U6171 ( .A1(n5236), .A2(n8639), .ZN(n5004) );
  NOR2_X1 U6172 ( .A1(n10146), .A2(n9638), .ZN(n5005) );
  NAND2_X1 U6173 ( .A1(n5315), .A2(n5314), .ZN(n9269) );
  INV_X1 U6174 ( .A(n8580), .ZN(n5275) );
  INV_X1 U6175 ( .A(n5474), .ZN(n5473) );
  NAND2_X1 U6176 ( .A1(n8743), .A2(n4950), .ZN(n5474) );
  AND2_X1 U6177 ( .A1(n6163), .A2(n9077), .ZN(n5006) );
  AND2_X1 U6178 ( .A1(n8483), .A2(n8516), .ZN(n5007) );
  INV_X1 U6179 ( .A(n9677), .ZN(n7636) );
  NOR2_X1 U6180 ( .A1(n5488), .A2(n8903), .ZN(n5008) );
  AND2_X1 U6181 ( .A1(n5273), .A2(n8589), .ZN(n5009) );
  AND2_X1 U6182 ( .A1(n9680), .A2(n5438), .ZN(n5010) );
  AND2_X1 U6183 ( .A1(n6154), .A2(n6152), .ZN(n5011) );
  AND2_X1 U6184 ( .A1(n8699), .A2(n8696), .ZN(n5012) );
  AND2_X1 U6185 ( .A1(n5197), .A2(n5291), .ZN(n5013) );
  OR2_X1 U6186 ( .A1(n9019), .A2(n6296), .ZN(n8478) );
  AND2_X1 U6187 ( .A1(n5341), .A2(n5336), .ZN(n5014) );
  AND2_X1 U6188 ( .A1(n5493), .A2(n4968), .ZN(n5015) );
  NAND2_X1 U6189 ( .A1(n10168), .A2(n9808), .ZN(n5016) );
  NAND2_X1 U6190 ( .A1(n7086), .A2(n8854), .ZN(n5017) );
  AND2_X1 U6191 ( .A1(n5130), .A2(n4993), .ZN(n5018) );
  AND2_X1 U6192 ( .A1(n5123), .A2(n5124), .ZN(n5019) );
  AND2_X1 U6193 ( .A1(n5326), .A2(n7749), .ZN(n5325) );
  AND2_X2 U6194 ( .A1(n6326), .A2(n5457), .ZN(n6394) );
  INV_X1 U6195 ( .A(n5479), .ZN(n5478) );
  NAND2_X1 U6196 ( .A1(n8115), .A2(n8116), .ZN(n8356) );
  NAND2_X1 U6197 ( .A1(n5677), .A2(n5676), .ZN(n8740) );
  AND2_X1 U6198 ( .A1(n7508), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5020) );
  AND2_X1 U6199 ( .A1(n7508), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5021) );
  NAND2_X1 U6200 ( .A1(n8389), .A2(n8388), .ZN(n5022) );
  OAI21_X1 U6201 ( .B1(n7857), .B2(n8577), .A(n5935), .ZN(n7938) );
  INV_X1 U6202 ( .A(n10543), .ZN(n6665) );
  AND2_X1 U6203 ( .A1(n6925), .A2(n7143), .ZN(n5023) );
  AND2_X1 U6204 ( .A1(n8753), .A2(n8863), .ZN(n5024) );
  NAND2_X1 U6205 ( .A1(n8232), .A2(n8231), .ZN(n10349) );
  NAND2_X1 U6206 ( .A1(n8147), .A2(n8146), .ZN(n8148) );
  NOR2_X1 U6207 ( .A1(n7911), .A2(n7912), .ZN(n5025) );
  NOR2_X1 U6208 ( .A1(n8928), .A2(n8929), .ZN(n5026) );
  AND2_X1 U6209 ( .A1(n8351), .A2(n10369), .ZN(n5027) );
  INV_X1 U6210 ( .A(n10345), .ZN(n10206) );
  NAND2_X1 U6211 ( .A1(n8243), .A2(n8242), .ZN(n10345) );
  NAND2_X1 U6212 ( .A1(n10154), .A2(n5263), .ZN(n5264) );
  NAND2_X1 U6213 ( .A1(n10254), .A2(n5266), .ZN(n5269) );
  OR2_X1 U6214 ( .A1(n10291), .A2(n10296), .ZN(n5028) );
  NOR2_X1 U6215 ( .A1(n7375), .A2(n7447), .ZN(n5029) );
  NAND2_X1 U6216 ( .A1(n9647), .A2(n8371), .ZN(n9575) );
  AND2_X1 U6217 ( .A1(n8738), .A2(n8790), .ZN(n5030) );
  NAND2_X1 U6218 ( .A1(n8290), .A2(n8289), .ZN(n10131) );
  INV_X1 U6219 ( .A(n10131), .ZN(n5262) );
  NAND2_X1 U6220 ( .A1(n6249), .A2(n6248), .ZN(n9019) );
  INV_X1 U6221 ( .A(n5542), .ZN(n5541) );
  OR2_X1 U6222 ( .A1(n8753), .A2(n5030), .ZN(n5542) );
  NAND2_X1 U6223 ( .A1(n7558), .A2(n7557), .ZN(n10733) );
  INV_X1 U6224 ( .A(n10733), .ZN(n5270) );
  AND2_X1 U6225 ( .A1(n7556), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5031) );
  NAND2_X1 U6226 ( .A1(n5784), .A2(n5783), .ZN(n7056) );
  OR2_X1 U6227 ( .A1(n7715), .A2(n7708), .ZN(n5032) );
  NOR2_X1 U6228 ( .A1(n7444), .A2(n7445), .ZN(n5033) );
  AND2_X1 U6229 ( .A1(n5656), .A2(n9444), .ZN(n5034) );
  AND2_X1 U6230 ( .A1(n7841), .A2(n7763), .ZN(n5035) );
  OR2_X1 U6231 ( .A1(n7778), .A2(n7743), .ZN(n5036) );
  INV_X1 U6232 ( .A(n10609), .ZN(n5525) );
  AND4_X1 U6233 ( .A1(n5815), .A2(n5814), .A3(n5813), .A4(n5812), .ZN(n8854)
         );
  INV_X1 U6234 ( .A(n8854), .ZN(n5079) );
  NOR2_X1 U6235 ( .A1(n7347), .A2(n10592), .ZN(n6971) );
  NAND2_X1 U6236 ( .A1(n6947), .A2(n6948), .ZN(n6946) );
  INV_X1 U6237 ( .A(n7610), .ZN(n5546) );
  AND2_X1 U6238 ( .A1(n4965), .A2(n8984), .ZN(n5037) );
  AND2_X1 U6239 ( .A1(n5521), .A2(n5520), .ZN(n5038) );
  NAND2_X1 U6240 ( .A1(n7272), .A2(n7271), .ZN(n5039) );
  XOR2_X1 U6241 ( .A(n7556), .B(n7516), .Z(n5040) );
  NAND2_X1 U6242 ( .A1(n6110), .A2(n6109), .ZN(n8675) );
  NAND2_X1 U6243 ( .A1(n8672), .A2(n8610), .ZN(n5219) );
  OR2_X1 U6244 ( .A1(n8665), .A2(n8610), .ZN(n5221) );
  OR2_X1 U6245 ( .A1(n8610), .A2(n6785), .ZN(n9150) );
  NOR2_X1 U6246 ( .A1(n8569), .A2(n8610), .ZN(n5243) );
  MUX2_X1 U6247 ( .A(n8521), .B(n8520), .S(n8610), .Z(n8527) );
  NAND2_X2 U6248 ( .A1(n6415), .A2(n6730), .ZN(n10408) );
  NAND2_X1 U6249 ( .A1(n6308), .A2(n6349), .ZN(n6361) );
  INV_X1 U6250 ( .A(n5042), .ZN(n6974) );
  OAI21_X1 U6251 ( .B1(n10122), .B2(n8300), .A(n8299), .ZN(n10091) );
  OAI22_X1 U6252 ( .A1(n10189), .A2(n10188), .B1(n10339), .B2(n10325), .ZN(
        n10167) );
  XNOR2_X1 U6253 ( .A(n5358), .B(n5417), .ZN(n10271) );
  NAND2_X1 U6254 ( .A1(n7335), .A2(n9732), .ZN(n7485) );
  NAND2_X1 U6255 ( .A1(n7634), .A2(n7636), .ZN(n7635) );
  NAND2_X1 U6256 ( .A1(n10212), .A2(n5451), .ZN(n5450) );
  AOI21_X1 U6257 ( .B1(n10108), .B2(n10109), .A(n10088), .ZN(n5041) );
  NOR2_X1 U6258 ( .A1(n10150), .A2(n8319), .ZN(n8342) );
  OR2_X1 U6259 ( .A1(n8140), .A2(n9685), .ZN(n8141) );
  NAND2_X1 U6260 ( .A1(n7484), .A2(n9668), .ZN(n10685) );
  XNOR2_X1 U6261 ( .A(n5041), .B(n10095), .ZN(n10277) );
  NAND2_X1 U6262 ( .A1(n7562), .A2(n7561), .ZN(n7634) );
  NAND2_X1 U6263 ( .A1(n5439), .A2(n5010), .ZN(n7799) );
  NAND2_X1 U6264 ( .A1(n5801), .A2(n5800), .ZN(n5803) );
  OAI21_X1 U6265 ( .B1(n10822), .B2(n8045), .A(n9911), .ZN(n8140) );
  INV_X1 U6266 ( .A(n5211), .ZN(n5210) );
  NAND2_X2 U6267 ( .A1(n6840), .A2(n4980), .ZN(n9965) );
  NAND2_X1 U6268 ( .A1(n10223), .A2(n9925), .ZN(n10212) );
  NAND2_X1 U6269 ( .A1(n8044), .A2(n9768), .ZN(n10822) );
  OAI21_X1 U6270 ( .B1(n8342), .B2(n5445), .A(n5444), .ZN(n5448) );
  NAND2_X1 U6271 ( .A1(n7175), .A2(n9670), .ZN(n7174) );
  NOR2_X1 U6272 ( .A1(n6394), .A2(n5252), .ZN(n5251) );
  NAND2_X1 U6273 ( .A1(n5449), .A2(n9919), .ZN(n10250) );
  NAND2_X1 U6274 ( .A1(n10685), .A2(n7511), .ZN(n10682) );
  NAND2_X4 U6275 ( .A1(n6306), .A2(n4945), .ZN(n8475) );
  NAND2_X2 U6276 ( .A1(n6125), .A2(n6127), .ZN(n6306) );
  NAND4_X2 U6277 ( .A1(n5279), .A2(n5535), .A3(n5278), .A4(n4967), .ZN(n5940)
         );
  OR2_X2 U6278 ( .A1(n7422), .A2(n8493), .ZN(n7619) );
  NAND2_X1 U6279 ( .A1(n9057), .A2(n8642), .ZN(n6266) );
  NAND2_X1 U6280 ( .A1(n10277), .A2(n10828), .ZN(n5260) );
  INV_X1 U6281 ( .A(n5448), .ZN(n10124) );
  NAND2_X1 U6282 ( .A1(n8313), .A2(n9921), .ZN(n5449) );
  AOI21_X1 U6283 ( .B1(n5044), .B2(n10065), .A(n10064), .ZN(n10066) );
  XNOR2_X1 U6284 ( .A(n10057), .B(n5045), .ZN(n5044) );
  NAND2_X1 U6285 ( .A1(n5155), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5154) );
  NAND2_X1 U6286 ( .A1(n5372), .A2(n5371), .ZN(n10122) );
  NAND2_X1 U6287 ( .A1(n5212), .A2(n5210), .ZN(n5801) );
  NAND2_X1 U6288 ( .A1(n5359), .A2(n10094), .ZN(n5358) );
  OAI21_X2 U6289 ( .B1(n10815), .B2(n5027), .A(n5399), .ZN(n5398) );
  NAND2_X1 U6290 ( .A1(n5692), .A2(n9376), .ZN(n6117) );
  NAND2_X1 U6291 ( .A1(n5688), .A2(n9502), .ZN(n6034) );
  NAND2_X1 U6292 ( .A1(n5690), .A2(n5689), .ZN(n6062) );
  NOR2_X2 U6293 ( .A1(n5975), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5051) );
  NAND2_X1 U6294 ( .A1(n5287), .A2(n5286), .ZN(n9057) );
  NAND2_X1 U6295 ( .A1(n5303), .A2(n5011), .ZN(n9151) );
  NAND2_X1 U6296 ( .A1(n5300), .A2(n5299), .ZN(n9098) );
  NAND2_X1 U6297 ( .A1(n5671), .A2(n5673), .ZN(n5694) );
  NAND2_X1 U6298 ( .A1(n7962), .A2(n5057), .ZN(n5056) );
  INV_X1 U6299 ( .A(n5063), .ZN(n7869) );
  NAND2_X1 U6301 ( .A1(n6306), .A2(n5070), .ZN(n5072) );
  OR2_X1 U6302 ( .A1(n6306), .A2(n6652), .ZN(n5071) );
  NAND2_X1 U6303 ( .A1(n5487), .A2(n5073), .ZN(n5074) );
  NAND2_X1 U6304 ( .A1(n5008), .A2(n7056), .ZN(n5077) );
  NAND3_X1 U6305 ( .A1(n5077), .A2(n5076), .A3(n10670), .ZN(n5075) );
  INV_X1 U6306 ( .A(n6103), .ZN(n5477) );
  NAND2_X1 U6307 ( .A1(n5081), .A2(n5080), .ZN(n6242) );
  OR2_X1 U6308 ( .A1(n6103), .A2(n5479), .ZN(n5081) );
  NAND2_X1 U6309 ( .A1(n8679), .A2(n6552), .ZN(n5084) );
  INV_X1 U6310 ( .A(n7710), .ZN(n5111) );
  NAND2_X1 U6311 ( .A1(n5116), .A2(n5513), .ZN(n5113) );
  INV_X1 U6312 ( .A(n7712), .ZN(n5115) );
  NOR2_X1 U6313 ( .A1(n8952), .A2(n8957), .ZN(n8977) );
  OR2_X1 U6314 ( .A1(n8907), .A2(n5121), .ZN(n5122) );
  NAND3_X1 U6315 ( .A1(n5126), .A2(n5127), .A3(n5125), .ZN(n6927) );
  NAND4_X1 U6316 ( .A1(n5126), .A2(n5127), .A3(n5125), .A4(
        P2_REG2_REG_7__SCAN_IN), .ZN(n5128) );
  INV_X1 U6317 ( .A(n5128), .ZN(n7144) );
  OAI211_X1 U6318 ( .C1(n10534), .C2(n4963), .A(n5129), .B(n5018), .ZN(n10554)
         );
  NAND2_X1 U6319 ( .A1(n10534), .A2(n4974), .ZN(n5129) );
  NOR2_X1 U6320 ( .A1(n10534), .A2(n10533), .ZN(n10532) );
  NOR2_X1 U6321 ( .A1(n10554), .A2(n5811), .ZN(n10553) );
  NAND3_X1 U6322 ( .A1(n5501), .A2(n5134), .A3(n5502), .ZN(n5133) );
  NAND2_X1 U6323 ( .A1(n8862), .A2(n8863), .ZN(n5543) );
  NAND2_X1 U6324 ( .A1(n8754), .A2(n5146), .ZN(n8758) );
  INV_X1 U6325 ( .A(n6882), .ZN(n5151) );
  NAND2_X1 U6326 ( .A1(n6766), .A2(n6765), .ZN(n6883) );
  NAND2_X1 U6327 ( .A1(n5151), .A2(n6880), .ZN(n5149) );
  NAND3_X1 U6328 ( .A1(n5524), .A2(n5522), .A3(n5523), .ZN(n6766) );
  INV_X1 U6329 ( .A(n5858), .ZN(n5159) );
  NAND3_X1 U6330 ( .A1(n5158), .A2(n5421), .A3(n5156), .ZN(n5921) );
  NAND2_X1 U6331 ( .A1(n5921), .A2(n5920), .ZN(n5923) );
  NAND2_X1 U6332 ( .A1(n8697), .A2(n5012), .ZN(n8874) );
  NOR2_X2 U6333 ( .A1(n5167), .A2(n5168), .ZN(n7824) );
  INV_X1 U6334 ( .A(n5170), .ZN(n5169) );
  NAND2_X1 U6335 ( .A1(n5176), .A2(n5174), .ZN(n6000) );
  NAND2_X1 U6336 ( .A1(n5180), .A2(n5007), .ZN(n5179) );
  NAND2_X1 U6337 ( .A1(n5013), .A2(n5181), .ZN(n5180) );
  NAND2_X1 U6338 ( .A1(n8484), .A2(n8480), .ZN(n5183) );
  OAI21_X1 U6339 ( .B1(n6059), .B2(n5186), .A(n5184), .ZN(n5658) );
  AND2_X1 U6340 ( .A1(n5188), .A2(n6371), .ZN(n6748) );
  NAND4_X1 U6341 ( .A1(n5188), .A2(n6747), .A3(n6746), .A4(n6371), .ZN(n6749)
         );
  NAND2_X1 U6342 ( .A1(n7907), .A2(n7866), .ZN(n6371) );
  NAND2_X1 U6343 ( .A1(n5189), .A2(n6198), .ZN(n5188) );
  NAND2_X1 U6344 ( .A1(n6198), .A2(n6203), .ZN(n6370) );
  INV_X1 U6345 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5190) );
  INV_X1 U6346 ( .A(n5194), .ZN(n5191) );
  NAND2_X1 U6347 ( .A1(n4966), .A2(n5194), .ZN(n6247) );
  NAND2_X1 U6348 ( .A1(n5191), .A2(n4966), .ZN(n5558) );
  NAND2_X1 U6349 ( .A1(n4966), .A2(n5659), .ZN(n5660) );
  NAND3_X1 U6350 ( .A1(n4966), .A2(n5194), .A3(n5193), .ZN(n5192) );
  NAND3_X1 U6351 ( .A1(n5002), .A2(n5195), .A3(n5279), .ZN(n5860) );
  XNOR2_X1 U6352 ( .A(n6751), .B(n6759), .ZN(n6760) );
  MUX2_X1 U6353 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6639), .S(n10503), .Z(n10496) );
  NAND3_X1 U6354 ( .A1(n5518), .A2(n5662), .A3(n5517), .ZN(n5774) );
  NAND3_X1 U6355 ( .A1(n5786), .A2(n5776), .A3(n5777), .ZN(n5212) );
  OAI211_X1 U6356 ( .C1(n5674), .C2(P2_DATAO_REG_0__SCAN_IN), .A(SI_0_), .B(
        n5214), .ZN(n5213) );
  NAND2_X1 U6357 ( .A1(n5674), .A2(n5567), .ZN(n5214) );
  NAND2_X2 U6358 ( .A1(n5215), .A2(n5850), .ZN(n10743) );
  NAND3_X1 U6359 ( .A1(n5220), .A2(n5219), .A3(n5218), .ZN(n5217) );
  NOR2_X1 U6360 ( .A1(n5224), .A2(n5223), .ZN(n8659) );
  NOR2_X1 U6361 ( .A1(n8640), .A2(n5234), .ZN(n5223) );
  NAND2_X1 U6362 ( .A1(n5231), .A2(n5228), .ZN(n5224) );
  INV_X1 U6363 ( .A(n8638), .ZN(n5237) );
  OR2_X1 U6364 ( .A1(n8656), .A2(n8657), .ZN(n5238) );
  NAND3_X1 U6365 ( .A1(n5249), .A2(n5873), .A3(n5248), .ZN(n8565) );
  NAND2_X2 U6366 ( .A1(n6417), .A2(n6418), .ZN(n6797) );
  OAI21_X2 U6367 ( .B1(n6797), .B2(n5256), .A(n5255), .ZN(n10592) );
  NAND3_X1 U6368 ( .A1(n5260), .A2(n5258), .A3(n5257), .ZN(n10380) );
  INV_X1 U6369 ( .A(n5264), .ZN(n10139) );
  NAND2_X1 U6370 ( .A1(n10254), .A2(n5265), .ZN(n10204) );
  INV_X1 U6371 ( .A(n5269), .ZN(n10218) );
  NAND2_X1 U6372 ( .A1(n6147), .A2(n5274), .ZN(n5272) );
  NAND2_X1 U6373 ( .A1(n5272), .A2(n5009), .ZN(n7941) );
  INV_X1 U6374 ( .A(n5940), .ZN(n5534) );
  NAND2_X1 U6375 ( .A1(n9078), .A2(n5006), .ZN(n5287) );
  NOR2_X2 U6376 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n6113) );
  OR2_X1 U6377 ( .A1(n6272), .A2(n8743), .ZN(n5294) );
  NAND2_X1 U6378 ( .A1(n6272), .A2(n5293), .ZN(n5292) );
  NAND2_X1 U6379 ( .A1(n6272), .A2(n6271), .ZN(n6295) );
  NAND2_X1 U6380 ( .A1(n5498), .A2(n5499), .ZN(n5500) );
  NAND3_X1 U6381 ( .A1(n5498), .A2(n5695), .A3(n5499), .ZN(n9255) );
  NAND2_X1 U6382 ( .A1(n6157), .A2(n5301), .ZN(n5300) );
  NAND2_X1 U6383 ( .A1(n7965), .A2(n5304), .ZN(n5303) );
  OR2_X1 U6384 ( .A1(n6754), .A2(n10598), .ZN(n6136) );
  OR2_X2 U6385 ( .A1(n5307), .A2(n5306), .ZN(n10598) );
  OAI211_X2 U6386 ( .C1(n5735), .C2(n8182), .A(n5461), .B(n5737), .ZN(n6754)
         );
  NAND2_X1 U6387 ( .A1(n9151), .A2(n6155), .ZN(n9139) );
  NAND2_X1 U6388 ( .A1(n7112), .A2(n8486), .ZN(n7114) );
  NAND2_X1 U6389 ( .A1(n7941), .A2(n6149), .ZN(n7875) );
  MUX2_X2 U6390 ( .A(n6275), .B(n4978), .S(n8660), .Z(n9023) );
  NAND2_X1 U6391 ( .A1(n7875), .A2(n7874), .ZN(n7873) );
  NAND2_X1 U6392 ( .A1(n9098), .A2(n6158), .ZN(n9088) );
  NAND2_X1 U6393 ( .A1(n7034), .A2(n7036), .ZN(n7033) );
  INV_X1 U6394 ( .A(n5940), .ZN(n5498) );
  OAI21_X1 U6395 ( .B1(n7715), .B2(n7457), .A(n7714), .ZN(n7716) );
  OAI21_X1 U6396 ( .B1(n7391), .B2(n7149), .A(n7390), .ZN(n7448) );
  NOR2_X1 U6397 ( .A1(n5195), .A2(n5508), .ZN(n5507) );
  NAND2_X1 U6398 ( .A1(n6136), .A2(n8517), .ZN(n6991) );
  NAND2_X1 U6399 ( .A1(n8114), .A2(n5310), .ZN(n5309) );
  NAND2_X1 U6400 ( .A1(n8432), .A2(n5316), .ZN(n5315) );
  NAND2_X1 U6401 ( .A1(n5318), .A2(n5321), .ZN(n7760) );
  NAND2_X1 U6402 ( .A1(n7750), .A2(n5325), .ZN(n5318) );
  NAND2_X1 U6403 ( .A1(n9549), .A2(n5332), .ZN(n5331) );
  INV_X1 U6404 ( .A(n9549), .ZN(n5334) );
  NAND2_X1 U6405 ( .A1(n9652), .A2(n5342), .ZN(n5337) );
  NAND2_X1 U6406 ( .A1(n5335), .A2(n9585), .ZN(n8383) );
  NAND3_X1 U6407 ( .A1(n5338), .A2(n5337), .A3(n5014), .ZN(n5335) );
  NAND3_X1 U6408 ( .A1(n5338), .A2(n5337), .A3(n5341), .ZN(n9589) );
  NAND2_X1 U6409 ( .A1(n9268), .A2(n5344), .ZN(n5343) );
  OAI211_X1 U6410 ( .C1(n9268), .C2(n5345), .A(n8468), .B(n5343), .ZN(P1_U3220) );
  NOR2_X1 U6411 ( .A1(n8464), .A2(n8456), .ZN(n5349) );
  NAND2_X1 U6412 ( .A1(n8464), .A2(n8456), .ZN(n5350) );
  INV_X1 U6413 ( .A(n8464), .ZN(n5351) );
  NAND2_X1 U6414 ( .A1(n7977), .A2(n7976), .ZN(n7990) );
  AND2_X1 U6415 ( .A1(n5357), .A2(n5028), .ZN(n10110) );
  NAND2_X1 U6416 ( .A1(n5357), .A2(n5356), .ZN(n5359) );
  NAND2_X1 U6417 ( .A1(n10091), .A2(n10090), .ZN(n5357) );
  INV_X1 U6418 ( .A(n5361), .ZN(n10203) );
  NAND2_X1 U6419 ( .A1(n8266), .A2(n4958), .ZN(n5372) );
  NAND2_X2 U6420 ( .A1(n4945), .A2(P2_U3151), .ZN(n8472) );
  MUX2_X1 U6421 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5575), .Z(n5576) );
  MUX2_X1 U6422 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5575), .Z(n5585) );
  MUX2_X1 U6423 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5575), .Z(n5594) );
  MUX2_X1 U6424 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n4945), .Z(n5599) );
  MUX2_X1 U6425 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n4945), .Z(n5605) );
  MUX2_X1 U6426 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n4945), .Z(n5616) );
  MUX2_X1 U6427 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n4945), .Z(n5624) );
  MUX2_X1 U6428 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n4945), .Z(n5649) );
  MUX2_X1 U6429 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n4945), .Z(n5647) );
  MUX2_X1 U6430 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n4945), .Z(n5636) );
  MUX2_X1 U6431 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n4945), .Z(n5638) );
  MUX2_X1 U6432 ( .A(n5675), .B(n7960), .S(n4945), .Z(n5657) );
  NAND2_X1 U6433 ( .A1(n10712), .A2(n5382), .ZN(n5385) );
  NAND2_X1 U6434 ( .A1(n10712), .A2(n5388), .ZN(n5387) );
  OAI21_X1 U6435 ( .B1(n10712), .B2(n10718), .A(n5396), .ZN(n7596) );
  OR2_X1 U6436 ( .A1(n10733), .A2(n10746), .ZN(n5396) );
  NAND2_X1 U6437 ( .A1(n5413), .A2(n5637), .ZN(n6059) );
  NAND2_X1 U6438 ( .A1(n5876), .A2(n5604), .ZN(n5889) );
  NAND3_X1 U6439 ( .A1(n9811), .A2(n9810), .A3(n5431), .ZN(n9817) );
  NAND3_X1 U6440 ( .A1(n5016), .A2(n5433), .A3(n5432), .ZN(n5431) );
  NAND2_X1 U6441 ( .A1(n5575), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5437) );
  OAI21_X1 U6442 ( .B1(n5575), .B2(n5570), .A(n5437), .ZN(n5571) );
  NAND2_X2 U6443 ( .A1(n4945), .A2(P1_U3086), .ZN(n10404) );
  MUX2_X1 U6444 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5575), .Z(n5581) );
  MUX2_X1 U6445 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5575), .Z(n5590) );
  MUX2_X1 U6446 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n4945), .Z(n5597) );
  MUX2_X1 U6447 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n4945), .Z(n5600) );
  MUX2_X1 U6448 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n4945), .Z(n5606) );
  MUX2_X1 U6449 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n4945), .Z(n5608) );
  MUX2_X1 U6450 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4945), .Z(n5612) );
  MUX2_X1 U6451 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n4945), .Z(n5621) );
  MUX2_X1 U6452 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4945), .Z(n5625) );
  MUX2_X1 U6453 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n4945), .Z(n5629) );
  MUX2_X1 U6454 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n4945), .Z(n5632) );
  MUX2_X1 U6455 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n4945), .Z(n5645) );
  MUX2_X1 U6456 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .S(n4945), .Z(n5655) );
  MUX2_X1 U6457 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n4945), .Z(n6243) );
  NAND2_X1 U6458 ( .A1(n7635), .A2(n5440), .ZN(n5439) );
  NAND2_X1 U6459 ( .A1(n10212), .A2(n9929), .ZN(n10185) );
  INV_X1 U6460 ( .A(n5450), .ZN(n9863) );
  NAND3_X1 U6461 ( .A1(n6309), .A2(n5456), .A3(n6376), .ZN(n5453) );
  NAND2_X1 U6462 ( .A1(n7360), .A2(n5465), .ZN(n5462) );
  NAND2_X1 U6463 ( .A1(n5462), .A2(n5463), .ZN(n5887) );
  NOR2_X1 U6464 ( .A1(n6103), .A2(n5481), .ZN(n6237) );
  NAND2_X1 U6465 ( .A1(n6236), .A2(n5480), .ZN(n5479) );
  NAND2_X1 U6466 ( .A1(n7056), .A2(n5490), .ZN(n5487) );
  NAND2_X1 U6467 ( .A1(n5500), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5697) );
  NOR2_X2 U6468 ( .A1(n4949), .A2(n4996), .ZN(n5499) );
  NOR2_X1 U6469 ( .A1(n7146), .A2(n7145), .ZN(n7376) );
  AOI21_X1 U6470 ( .B1(n7145), .B2(n5506), .A(n7456), .ZN(n5504) );
  NAND2_X1 U6471 ( .A1(n7146), .A2(n5506), .ZN(n5505) );
  INV_X1 U6472 ( .A(n7375), .ZN(n5506) );
  NOR2_X1 U6473 ( .A1(n10553), .A2(n6677), .ZN(n6680) );
  NAND2_X1 U6474 ( .A1(n5519), .A2(n5526), .ZN(n5523) );
  INV_X1 U6475 ( .A(n6761), .ZN(n5519) );
  NAND3_X1 U6476 ( .A1(n6947), .A2(n5526), .A3(n6948), .ZN(n5522) );
  XNOR2_X1 U6477 ( .A(n6762), .B(n5525), .ZN(n6864) );
  OR2_X1 U6478 ( .A1(n6105), .A2(n5672), .ZN(n5527) );
  NAND2_X1 U6479 ( .A1(n6105), .A2(n6104), .ZN(n5530) );
  NAND2_X1 U6480 ( .A1(n6105), .A2(n5531), .ZN(n5529) );
  OAI21_X2 U6481 ( .B1(n8824), .B2(n8718), .A(n8723), .ZN(n8831) );
  NOR2_X1 U6482 ( .A1(n5860), .A2(n5536), .ZN(n5908) );
  OAI21_X1 U6483 ( .B1(n8862), .B2(n5542), .A(n5538), .ZN(n8746) );
  AND2_X1 U6484 ( .A1(n7611), .A2(n5549), .ZN(n5545) );
  NOR2_X1 U6485 ( .A1(n7090), .A2(n5548), .ZN(n5547) );
  NAND2_X1 U6486 ( .A1(n6607), .A2(n9879), .ZN(n6614) );
  CLKBUF_X1 U6487 ( .A(n7293), .Z(n7397) );
  INV_X1 U6488 ( .A(n6809), .ZN(n6810) );
  XNOR2_X1 U6489 ( .A(n8159), .B(SI_29_), .ZN(n9664) );
  OR2_X1 U6490 ( .A1(n6815), .A2(n6596), .ZN(n6597) );
  NAND2_X1 U6491 ( .A1(n9968), .A2(n10592), .ZN(n7170) );
  INV_X1 U6492 ( .A(n9262), .ZN(n5698) );
  AOI21_X1 U6493 ( .B1(n8527), .B2(n10612), .A(n8526), .ZN(n8540) );
  NAND2_X1 U6494 ( .A1(n6754), .A2(n10598), .ZN(n8517) );
  NAND2_X1 U6495 ( .A1(n5571), .A2(SI_2_), .ZN(n5574) );
  OR2_X1 U6496 ( .A1(n5571), .A2(SI_2_), .ZN(n5572) );
  INV_X1 U6497 ( .A(n6746), .ZN(n8516) );
  OR2_X1 U6498 ( .A1(n8729), .A2(n8728), .ZN(n8730) );
  INV_X2 U6499 ( .A(n6828), .ZN(n6829) );
  OR2_X1 U6500 ( .A1(n8654), .A2(n9027), .ZN(n5552) );
  AND2_X1 U6501 ( .A1(n6293), .A2(n6292), .ZN(n5553) );
  INV_X1 U6502 ( .A(n8569), .ZN(n6145) );
  OR2_X1 U6503 ( .A1(n8560), .A2(n8610), .ZN(n5554) );
  AND2_X1 U6504 ( .A1(n5628), .A2(n5627), .ZN(n5556) );
  AND2_X1 U6505 ( .A1(n10262), .A2(n10236), .ZN(n5557) );
  OR2_X1 U6506 ( .A1(n9027), .A2(n9252), .ZN(n5559) );
  INV_X1 U6507 ( .A(n9154), .ZN(n6154) );
  OR2_X1 U6508 ( .A1(n9027), .A2(n9213), .ZN(n5560) );
  AND2_X1 U6509 ( .A1(n9697), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n5561) );
  INV_X1 U6510 ( .A(n9954), .ZN(n10305) );
  NAND2_X1 U6511 ( .A1(n6974), .A2(n7170), .ZN(n7171) );
  NAND2_X1 U6512 ( .A1(n10675), .A2(n7503), .ZN(n5562) );
  INV_X1 U6513 ( .A(n10070), .ZN(n10113) );
  INV_X1 U6514 ( .A(n8517), .ZN(n8518) );
  INV_X1 U6515 ( .A(n8551), .ZN(n8552) );
  NAND2_X1 U6516 ( .A1(n8555), .A2(n8554), .ZN(n8561) );
  NAND2_X1 U6517 ( .A1(n8561), .A2(n5554), .ZN(n8562) );
  OAI21_X1 U6518 ( .B1(n8629), .B2(n8628), .A(n8627), .ZN(n8630) );
  INV_X1 U6519 ( .A(n10168), .ZN(n9689) );
  AND2_X1 U6520 ( .A1(n9236), .A2(n9085), .ZN(n8626) );
  NOR2_X1 U6521 ( .A1(n9295), .A2(n9617), .ZN(n8415) );
  INV_X1 U6522 ( .A(n8403), .ZN(n8404) );
  AND4_X1 U6523 ( .A1(n6338), .A2(n6324), .A3(n6323), .A4(n6322), .ZN(n6325)
         );
  OR2_X1 U6524 ( .A1(n8145), .A2(n8155), .ZN(n8146) );
  AOI21_X1 U6525 ( .B1(n8831), .B2(n8832), .A(n8726), .ZN(n8729) );
  INV_X1 U6526 ( .A(n8897), .ZN(n8695) );
  INV_X1 U6527 ( .A(n6049), .ZN(n5690) );
  NOR2_X1 U6528 ( .A1(n9049), .A2(n9064), .ZN(n6102) );
  OR2_X1 U6529 ( .A1(n8422), .A2(n8416), .ZN(n8430) );
  NAND2_X1 U6530 ( .A1(n9964), .A2(n6806), .ZN(n7191) );
  NAND2_X1 U6531 ( .A1(n8402), .A2(n8404), .ZN(n8405) );
  INV_X1 U6532 ( .A(n6614), .ZN(n6611) );
  INV_X1 U6533 ( .A(n10687), .ZN(n9747) );
  INV_X1 U6534 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6847) );
  NAND2_X1 U6535 ( .A1(n6760), .A2(n7111), .ZN(n6761) );
  AND2_X1 U6536 ( .A1(n6134), .A2(n6135), .ZN(n6757) );
  INV_X1 U6538 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5673) );
  INV_X1 U6539 ( .A(n9213), .ZN(n6290) );
  OR2_X1 U6540 ( .A1(n8610), .A2(n6169), .ZN(n6915) );
  AND2_X1 U6541 ( .A1(n9270), .A2(n9271), .ZN(n8455) );
  AOI21_X1 U6542 ( .B1(n10349), .B2(n8438), .A(n8387), .ZN(n9550) );
  NAND2_X1 U6543 ( .A1(n6811), .A2(n6810), .ZN(n6852) );
  INV_X1 U6544 ( .A(n9648), .ZN(n8371) );
  AND2_X1 U6545 ( .A1(n8430), .A2(n9595), .ZN(n8431) );
  NAND2_X1 U6546 ( .A1(n9551), .A2(n9550), .ZN(n8390) );
  AND2_X1 U6547 ( .A1(n7990), .A2(n7989), .ZN(n9305) );
  NOR2_X1 U6548 ( .A1(n8257), .A2(n9618), .ZN(n8256) );
  NAND2_X1 U6549 ( .A1(n7577), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7641) );
  INV_X1 U6550 ( .A(n10284), .ZN(n10069) );
  NAND2_X1 U6551 ( .A1(n9965), .A2(n7412), .ZN(n9894) );
  OR2_X1 U6552 ( .A1(n8162), .A2(n8161), .ZN(n8163) );
  OR2_X1 U6553 ( .A1(n5652), .A2(n5651), .ZN(n6087) );
  NAND2_X1 U6554 ( .A1(n5606), .A2(SI_12_), .ZN(n5607) );
  NAND2_X1 U6555 ( .A1(n5600), .A2(SI_10_), .ZN(n5604) );
  AND2_X1 U6556 ( .A1(n5584), .A2(n5583), .ZN(n5786) );
  INV_X1 U6557 ( .A(n9052), .ZN(n8790) );
  AND2_X1 U6558 ( .A1(n8769), .A2(n8714), .ZN(n8715) );
  INV_X1 U6559 ( .A(n8709), .ZN(n9138) );
  XNOR2_X1 U6560 ( .A(n6759), .B(n8905), .ZN(n10612) );
  OR2_X1 U6561 ( .A1(n10781), .A2(n6291), .ZN(n6292) );
  AND2_X1 U6562 ( .A1(n8373), .A2(n8372), .ZN(n8374) );
  NOR2_X1 U6563 ( .A1(n8233), .A2(n9609), .ZN(n8247) );
  NAND2_X1 U6564 ( .A1(n10070), .A2(n10069), .ZN(n10111) );
  INV_X1 U6565 ( .A(n10154), .ZN(n10171) );
  AOI22_X1 U6566 ( .A1(n10203), .A2(n10211), .B1(n10206), .B2(n10335), .ZN(
        n10189) );
  OR2_X1 U6567 ( .A1(n6965), .A2(n9946), .ZN(n10257) );
  OR2_X1 U6568 ( .A1(n6614), .A2(n10062), .ZN(n7350) );
  INV_X1 U6569 ( .A(n10820), .ZN(n10791) );
  INV_X1 U6570 ( .A(n5874), .ZN(n5603) );
  INV_X1 U6571 ( .A(n5753), .ZN(n5755) );
  OR2_X1 U6572 ( .A1(n8767), .A2(n8841), .ZN(n8842) );
  INV_X1 U6573 ( .A(n9011), .ZN(n8677) );
  AND2_X1 U6574 ( .A1(n6124), .A2(n6123), .ZN(n8654) );
  AND4_X1 U6575 ( .A1(n5885), .A2(n5884), .A3(n5883), .A4(n5882), .ZN(n7828)
         );
  OR2_X1 U6576 ( .A1(n5977), .A2(n5767), .ZN(n5770) );
  INV_X1 U6577 ( .A(n9063), .ZN(n9086) );
  INV_X1 U6578 ( .A(n8497), .ZN(n7668) );
  INV_X1 U6579 ( .A(n9148), .ZN(n10607) );
  OR2_X1 U6580 ( .A1(n8176), .A2(n6747), .ZN(n10620) );
  AND2_X1 U6581 ( .A1(n6729), .A2(n6724), .ZN(n9651) );
  NAND2_X1 U6582 ( .A1(n9846), .A2(n9816), .ZN(n10123) );
  NAND2_X1 U6583 ( .A1(n9929), .A2(n10184), .ZN(n10211) );
  INV_X1 U6584 ( .A(n10852), .ZN(n10731) );
  INV_X1 U6585 ( .A(n7828), .ZN(n8899) );
  INV_X1 U6586 ( .A(n9111), .ZN(n9159) );
  NAND2_X1 U6587 ( .A1(n8740), .A2(n6290), .ZN(n6222) );
  OR2_X1 U6588 ( .A1(n6220), .A2(n6219), .ZN(n10780) );
  AND2_X1 U6589 ( .A1(n6231), .A2(n6230), .ZN(n10782) );
  INV_X1 U6590 ( .A(n8351), .ZN(n10846) );
  INV_X1 U6591 ( .A(n10308), .ZN(n10146) );
  INV_X1 U6592 ( .A(n8112), .ZN(n10809) );
  INV_X1 U6593 ( .A(n9642), .ZN(n9661) );
  AND4_X1 U6594 ( .A1(n6903), .A2(n6902), .A3(n6901), .A4(n6900), .ZN(n10280)
         );
  INV_X1 U6595 ( .A(n10190), .ZN(n10265) );
  OR2_X1 U6596 ( .A1(n7121), .A2(n6986), .ZN(n10835) );
  INV_X1 U6597 ( .A(n10839), .ZN(n10836) );
  AND2_X1 U6598 ( .A1(n6616), .A2(n6414), .ZN(P1_U3973) );
  INV_X1 U6599 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6221) );
  INV_X1 U6600 ( .A(SI_1_), .ZN(n5564) );
  NAND2_X1 U6601 ( .A1(n5565), .A2(n5564), .ZN(n5566) );
  NAND2_X1 U6602 ( .A1(n5569), .A2(n5566), .ZN(n5742) );
  INV_X1 U6603 ( .A(n5742), .ZN(n5568) );
  INV_X1 U6604 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5567) );
  INV_X1 U6605 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6609) );
  INV_X1 U6606 ( .A(SI_0_), .ZN(n6608) );
  NAND2_X1 U6607 ( .A1(n5568), .A2(n5741), .ZN(n5744) );
  NAND2_X1 U6608 ( .A1(n5744), .A2(n5569), .ZN(n5753) );
  NAND2_X1 U6609 ( .A1(n5572), .A2(n5574), .ZN(n5754) );
  INV_X1 U6610 ( .A(n5754), .ZN(n5573) );
  NAND2_X1 U6611 ( .A1(n5753), .A2(n5573), .ZN(n5756) );
  INV_X1 U6612 ( .A(n5576), .ZN(n5578) );
  INV_X1 U6613 ( .A(SI_3_), .ZN(n5577) );
  NAND2_X1 U6614 ( .A1(n5578), .A2(n5577), .ZN(n5579) );
  INV_X1 U6615 ( .A(n5581), .ZN(n5582) );
  INV_X1 U6616 ( .A(SI_4_), .ZN(n9483) );
  NAND2_X1 U6617 ( .A1(n5582), .A2(n9483), .ZN(n5583) );
  INV_X1 U6618 ( .A(n5585), .ZN(n5587) );
  INV_X1 U6619 ( .A(SI_5_), .ZN(n5586) );
  NAND2_X1 U6620 ( .A1(n5587), .A2(n5586), .ZN(n5588) );
  INV_X1 U6621 ( .A(n5590), .ZN(n5591) );
  INV_X1 U6622 ( .A(SI_6_), .ZN(n9482) );
  NAND2_X1 U6623 ( .A1(n5591), .A2(n9482), .ZN(n5592) );
  INV_X1 U6624 ( .A(n5594), .ZN(n5595) );
  INV_X1 U6625 ( .A(SI_7_), .ZN(n9476) );
  NAND2_X1 U6626 ( .A1(n5595), .A2(n9476), .ZN(n5596) );
  INV_X1 U6627 ( .A(n5597), .ZN(n5598) );
  INV_X1 U6628 ( .A(SI_8_), .ZN(n9475) );
  INV_X1 U6629 ( .A(SI_9_), .ZN(n9472) );
  INV_X1 U6630 ( .A(n5600), .ZN(n5601) );
  INV_X1 U6631 ( .A(SI_10_), .ZN(n9356) );
  NAND2_X1 U6632 ( .A1(n5601), .A2(n9356), .ZN(n5602) );
  NAND2_X1 U6633 ( .A1(n5608), .A2(SI_13_), .ZN(n5611) );
  INV_X1 U6634 ( .A(n5608), .ZN(n5609) );
  INV_X1 U6635 ( .A(SI_13_), .ZN(n9467) );
  NAND2_X1 U6636 ( .A1(n5609), .A2(n9467), .ZN(n5610) );
  NAND2_X1 U6637 ( .A1(n5923), .A2(n5611), .ZN(n5937) );
  NAND2_X1 U6638 ( .A1(n5612), .A2(SI_14_), .ZN(n5615) );
  INV_X1 U6639 ( .A(n5612), .ZN(n5613) );
  INV_X1 U6640 ( .A(SI_14_), .ZN(n9425) );
  NAND2_X1 U6641 ( .A1(n5613), .A2(n9425), .ZN(n5614) );
  NAND2_X1 U6642 ( .A1(n5937), .A2(n5936), .ZN(n5939) );
  NAND2_X1 U6643 ( .A1(n5616), .A2(SI_15_), .ZN(n5620) );
  INV_X1 U6644 ( .A(n5616), .ZN(n5618) );
  INV_X1 U6645 ( .A(SI_15_), .ZN(n5617) );
  NAND2_X1 U6646 ( .A1(n5618), .A2(n5617), .ZN(n5619) );
  XNOR2_X1 U6647 ( .A(n5621), .B(SI_16_), .ZN(n5968) );
  INV_X1 U6648 ( .A(n5621), .ZN(n5622) );
  INV_X1 U6649 ( .A(SI_16_), .ZN(n9427) );
  INV_X1 U6650 ( .A(SI_17_), .ZN(n5623) );
  XNOR2_X1 U6651 ( .A(n5624), .B(n5623), .ZN(n5984) );
  NAND2_X1 U6652 ( .A1(n5625), .A2(SI_18_), .ZN(n5628) );
  INV_X1 U6653 ( .A(n5625), .ZN(n5626) );
  INV_X1 U6654 ( .A(SI_18_), .ZN(n9428) );
  NAND2_X1 U6655 ( .A1(n5626), .A2(n9428), .ZN(n5627) );
  XNOR2_X1 U6656 ( .A(n5629), .B(SI_19_), .ZN(n6011) );
  INV_X1 U6657 ( .A(n5629), .ZN(n5630) );
  INV_X1 U6658 ( .A(SI_19_), .ZN(n9430) );
  NAND2_X1 U6659 ( .A1(n5630), .A2(n9430), .ZN(n5631) );
  INV_X1 U6660 ( .A(SI_20_), .ZN(n9459) );
  XNOR2_X1 U6661 ( .A(n5632), .B(n9459), .ZN(n6029) );
  NAND2_X1 U6662 ( .A1(n6030), .A2(n6029), .ZN(n5635) );
  INV_X1 U6663 ( .A(n5632), .ZN(n5633) );
  NAND2_X1 U6664 ( .A1(n5633), .A2(n9459), .ZN(n5634) );
  NAND2_X1 U6665 ( .A1(n5636), .A2(SI_21_), .ZN(n5637) );
  OAI21_X1 U6666 ( .B1(n5636), .B2(SI_21_), .A(n5637), .ZN(n6043) );
  XNOR2_X1 U6667 ( .A(n5638), .B(SI_22_), .ZN(n6058) );
  INV_X1 U6668 ( .A(n5638), .ZN(n5639) );
  INV_X1 U6669 ( .A(SI_22_), .ZN(n9453) );
  NAND2_X1 U6670 ( .A1(n5639), .A2(n9453), .ZN(n6071) );
  INV_X1 U6671 ( .A(n5649), .ZN(n5640) );
  INV_X1 U6672 ( .A(SI_23_), .ZN(n9447) );
  NAND2_X1 U6673 ( .A1(n5640), .A2(n9447), .ZN(n5648) );
  AND2_X1 U6674 ( .A1(n6071), .A2(n5648), .ZN(n5721) );
  INV_X1 U6675 ( .A(n5647), .ZN(n5641) );
  INV_X1 U6676 ( .A(SI_24_), .ZN(n9446) );
  NAND2_X1 U6677 ( .A1(n5641), .A2(n9446), .ZN(n5646) );
  AND2_X1 U6678 ( .A1(n5721), .A2(n5646), .ZN(n6085) );
  INV_X1 U6679 ( .A(n5645), .ZN(n5642) );
  INV_X1 U6680 ( .A(SI_25_), .ZN(n9451) );
  NAND2_X1 U6681 ( .A1(n5642), .A2(n9451), .ZN(n5644) );
  AND2_X1 U6682 ( .A1(n6085), .A2(n5644), .ZN(n5643) );
  INV_X1 U6683 ( .A(SI_26_), .ZN(n9444) );
  XNOR2_X1 U6684 ( .A(n5655), .B(n9444), .ZN(n5717) );
  INV_X1 U6685 ( .A(n5644), .ZN(n5654) );
  XNOR2_X1 U6686 ( .A(n5645), .B(n9451), .ZN(n6089) );
  INV_X1 U6687 ( .A(n5646), .ZN(n5652) );
  XNOR2_X1 U6688 ( .A(n5647), .B(n9446), .ZN(n5724) );
  INV_X1 U6689 ( .A(n5648), .ZN(n5650) );
  XNOR2_X1 U6690 ( .A(n5649), .B(n9447), .ZN(n6072) );
  OR2_X1 U6691 ( .A1(n5650), .A2(n6072), .ZN(n5722) );
  AND2_X1 U6692 ( .A1(n5724), .A2(n5722), .ZN(n5651) );
  AND2_X1 U6693 ( .A1(n6089), .A2(n6087), .ZN(n5653) );
  INV_X1 U6694 ( .A(n5655), .ZN(n5656) );
  INV_X1 U6695 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5675) );
  INV_X1 U6696 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7960) );
  NAND2_X1 U6697 ( .A1(n5658), .A2(n5657), .ZN(n5659) );
  INV_X1 U6698 ( .A(SI_27_), .ZN(n9440) );
  NAND2_X1 U6699 ( .A1(n5660), .A2(n9440), .ZN(n5661) );
  INV_X1 U6700 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6174) );
  NOR2_X1 U6701 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n5663) );
  INV_X1 U6702 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6187) );
  INV_X1 U6703 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6111) );
  NAND4_X1 U6704 ( .A1(n6175), .A2(n5663), .A3(n6187), .A4(n6111), .ZN(n5668)
         );
  NOR2_X1 U6705 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5666) );
  NOR2_X1 U6706 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n5665) );
  NOR2_X1 U6707 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5664) );
  NAND4_X1 U6708 ( .A1(n6113), .A2(n5666), .A3(n5665), .A4(n5664), .ZN(n5667)
         );
  NAND2_X1 U6709 ( .A1(n5694), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5670) );
  INV_X1 U6710 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5669) );
  INV_X1 U6711 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5672) );
  OR2_X1 U6712 ( .A1(n8475), .A2(n5675), .ZN(n5676) );
  INV_X1 U6713 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5680) );
  INV_X1 U6714 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5682) );
  INV_X1 U6715 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9515) );
  INV_X1 U6716 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5684) );
  INV_X1 U6717 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5686) );
  INV_X1 U6718 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9418) );
  INV_X1 U6719 ( .A(n6020), .ZN(n5688) );
  INV_X1 U6720 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9502) );
  INV_X1 U6721 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5689) );
  INV_X1 U6722 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9524) );
  INV_X1 U6723 ( .A(n5708), .ZN(n5692) );
  NAND2_X1 U6724 ( .A1(n5708), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5693) );
  NAND2_X1 U6725 ( .A1(n6117), .A2(n5693), .ZN(n9033) );
  INV_X1 U6726 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5695) );
  INV_X1 U6727 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9256) );
  XNOR2_X2 U6728 ( .A(n5696), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5700) );
  XNOR2_X2 U6729 ( .A(n5697), .B(n5695), .ZN(n9262) );
  NAND2_X1 U6730 ( .A1(n9033), .A2(n6250), .ZN(n5706) );
  INV_X1 U6731 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n5703) );
  INV_X1 U6732 ( .A(n5700), .ZN(n8471) );
  NAND2_X1 U6733 ( .A1(n6252), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5702) );
  OR2_X2 U6734 ( .A1(n5700), .A2(n9262), .ZN(n5745) );
  NAND2_X1 U6735 ( .A1(n5459), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5701) );
  OAI211_X1 U6736 ( .C1(n5703), .C2(n8182), .A(n5702), .B(n5701), .ZN(n5704)
         );
  INV_X1 U6737 ( .A(n5704), .ZN(n5705) );
  NAND2_X2 U6738 ( .A1(n8740), .A2(n9041), .ZN(n8651) );
  NAND2_X1 U6739 ( .A1(n6095), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U6740 ( .A1(n5708), .A2(n5707), .ZN(n9044) );
  NAND2_X1 U6741 ( .A1(n9044), .A2(n6250), .ZN(n5714) );
  INV_X1 U6742 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U6743 ( .A1(n5459), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5710) );
  NAND2_X1 U6744 ( .A1(n6252), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5709) );
  OAI211_X1 U6745 ( .C1(n8182), .C2(n5711), .A(n5710), .B(n5709), .ZN(n5712)
         );
  INV_X1 U6746 ( .A(n5712), .ZN(n5713) );
  AND2_X1 U6747 ( .A1(n5716), .A2(n5715), .ZN(n5718) );
  NAND2_X1 U6748 ( .A1(n8288), .A2(n8473), .ZN(n5720) );
  INV_X1 U6749 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7908) );
  OR2_X1 U6750 ( .A1(n8475), .A2(n7908), .ZN(n5719) );
  NAND2_X1 U6751 ( .A1(n6086), .A2(n5721), .ZN(n5723) );
  NAND2_X1 U6752 ( .A1(n8271), .A2(n8473), .ZN(n5728) );
  INV_X1 U6753 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n5726) );
  OR2_X1 U6754 ( .A1(n8475), .A2(n5726), .ZN(n5727) );
  NAND2_X1 U6755 ( .A1(n6078), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5729) );
  NAND2_X1 U6756 ( .A1(n6093), .A2(n5729), .ZN(n9065) );
  NAND2_X1 U6757 ( .A1(n9065), .A2(n6250), .ZN(n5734) );
  INV_X1 U6758 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n9072) );
  NAND2_X1 U6759 ( .A1(n6252), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5731) );
  NAND2_X1 U6760 ( .A1(n5459), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5730) );
  OAI211_X1 U6761 ( .C1(n9072), .C2(n8182), .A(n5731), .B(n5730), .ZN(n5732)
         );
  INV_X1 U6762 ( .A(n5732), .ZN(n5733) );
  INV_X1 U6763 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6961) );
  INV_X1 U6764 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n5735) );
  INV_X1 U6765 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5736) );
  OR2_X1 U6766 ( .A1(n5760), .A2(n5736), .ZN(n5737) );
  NAND2_X1 U6767 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5738) );
  MUX2_X1 U6768 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5738), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5740) );
  INV_X1 U6769 ( .A(n6556), .ZN(n5739) );
  NAND2_X1 U6770 ( .A1(n5740), .A2(n5739), .ZN(n6564) );
  INV_X1 U6771 ( .A(n6564), .ZN(n6652) );
  NAND2_X1 U6772 ( .A1(n5742), .A2(n5213), .ZN(n5743) );
  AND2_X1 U6773 ( .A1(n5744), .A2(n5743), .ZN(n6344) );
  NAND2_X1 U6774 ( .A1(n6252), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5749) );
  INV_X1 U6775 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6893) );
  OR2_X1 U6776 ( .A1(n5930), .A2(n6893), .ZN(n5748) );
  INV_X1 U6777 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6553) );
  OR2_X1 U6778 ( .A1(n5977), .A2(n6553), .ZN(n5747) );
  INV_X1 U6779 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6920) );
  OR2_X1 U6780 ( .A1(n8182), .A2(n6920), .ZN(n5746) );
  NAND4_X1 U6781 ( .A1(n5749), .A2(n5748), .A3(n5747), .A4(n5746), .ZN(n6134)
         );
  NAND2_X1 U6782 ( .A1(n8169), .A2(SI_0_), .ZN(n5750) );
  XNOR2_X1 U6783 ( .A(n5750), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9267) );
  MUX2_X1 U6784 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9267), .S(n6306), .Z(n6135) );
  INV_X1 U6785 ( .A(n6757), .ZN(n6992) );
  NAND2_X1 U6786 ( .A1(n6991), .A2(n6992), .ZN(n6990) );
  INV_X1 U6787 ( .A(n10598), .ZN(n6997) );
  OR2_X1 U6788 ( .A1(n6754), .A2(n6997), .ZN(n5751) );
  NAND2_X1 U6789 ( .A1(n6990), .A2(n5751), .ZN(n10605) );
  NOR2_X1 U6790 ( .A1(n6556), .A2(n5672), .ZN(n5752) );
  OR2_X1 U6791 ( .A1(n8475), .A2(n5570), .ZN(n5759) );
  NAND2_X1 U6792 ( .A1(n5755), .A2(n5754), .ZN(n5757) );
  NAND2_X1 U6793 ( .A1(n5757), .A2(n5756), .ZN(n6822) );
  OR2_X1 U6794 ( .A1(n6046), .A2(n6822), .ZN(n5758) );
  OAI211_X1 U6795 ( .C1(n6306), .C2(n10503), .A(n5759), .B(n5758), .ZN(n6759)
         );
  INV_X1 U6796 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6666) );
  OR2_X1 U6797 ( .A1(n8182), .A2(n6666), .ZN(n5765) );
  NAND2_X1 U6798 ( .A1(n5459), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5764) );
  INV_X1 U6799 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5761) );
  INV_X1 U6800 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10619) );
  OR2_X1 U6801 ( .A1(n5930), .A2(n10619), .ZN(n5762) );
  INV_X1 U6802 ( .A(n10612), .ZN(n10606) );
  NAND2_X1 U6803 ( .A1(n10605), .A2(n10606), .ZN(n10604) );
  OR2_X1 U6804 ( .A1(n8905), .A2(n6759), .ZN(n5766) );
  NAND2_X1 U6805 ( .A1(n10604), .A2(n5766), .ZN(n7108) );
  NAND2_X1 U6806 ( .A1(n6252), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5772) );
  OR2_X1 U6807 ( .A1(n5930), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5771) );
  INV_X1 U6808 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5767) );
  INV_X1 U6809 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5768) );
  OR2_X1 U6810 ( .A1(n8182), .A2(n5768), .ZN(n5769) );
  NAND4_X1 U6811 ( .A1(n5772), .A2(n5771), .A3(n5770), .A4(n5769), .ZN(n10609)
         );
  NAND2_X1 U6812 ( .A1(n5774), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5773) );
  MUX2_X1 U6813 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5773), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5775) );
  OR2_X1 U6814 ( .A1(n5777), .A2(n5776), .ZN(n5778) );
  NAND2_X1 U6815 ( .A1(n5779), .A2(n5778), .ZN(n7008) );
  INV_X1 U6816 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6346) );
  OR2_X1 U6817 ( .A1(n8475), .A2(n6346), .ZN(n5780) );
  OAI211_X1 U6818 ( .C1(n6306), .C2(n6670), .A(n5781), .B(n5780), .ZN(n7116)
         );
  NAND2_X1 U6819 ( .A1(n10609), .A2(n7116), .ZN(n5782) );
  NAND2_X1 U6820 ( .A1(n7108), .A2(n5782), .ZN(n5784) );
  OR2_X1 U6821 ( .A1(n10609), .A2(n7116), .ZN(n5783) );
  INV_X2 U6822 ( .A(n8475), .ZN(n6017) );
  NAND2_X1 U6823 ( .A1(n5804), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5785) );
  XNOR2_X1 U6824 ( .A(n5785), .B(P2_IR_REG_4__SCAN_IN), .ZN(n10543) );
  AOI22_X1 U6825 ( .A1(n6017), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n6016), .B2(
        n10543), .ZN(n5791) );
  OR2_X1 U6826 ( .A1(n5787), .A2(n5786), .ZN(n5788) );
  AND2_X1 U6827 ( .A1(n5789), .A2(n5788), .ZN(n6359) );
  NAND2_X1 U6828 ( .A1(n6359), .A2(n8473), .ZN(n5790) );
  NAND2_X1 U6829 ( .A1(n5459), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5797) );
  INV_X1 U6830 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7058) );
  OR2_X1 U6831 ( .A1(n8182), .A2(n7058), .ZN(n5796) );
  NAND2_X1 U6832 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5792) );
  AND2_X1 U6833 ( .A1(n5809), .A2(n5792), .ZN(n7059) );
  OR2_X1 U6834 ( .A1(n5930), .A2(n7059), .ZN(n5795) );
  INV_X1 U6835 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5793) );
  OR2_X1 U6836 ( .A1(n5760), .A2(n5793), .ZN(n5794) );
  NAND4_X1 U6837 ( .A1(n5797), .A2(n5796), .A3(n5795), .A4(n5794), .ZN(n8904)
         );
  NOR2_X1 U6838 ( .A1(n7061), .A2(n8904), .ZN(n5799) );
  OR2_X1 U6839 ( .A1(n5801), .A2(n5800), .ZN(n5802) );
  NAND2_X1 U6840 ( .A1(n5803), .A2(n5802), .ZN(n7224) );
  OR2_X1 U6841 ( .A1(n7224), .A2(n6046), .ZN(n5807) );
  NAND2_X1 U6842 ( .A1(n5825), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5805) );
  XNOR2_X1 U6843 ( .A(n5805), .B(P2_IR_REG_5__SCAN_IN), .ZN(n10566) );
  AOI22_X1 U6844 ( .A1(n6017), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6016), .B2(
        n10566), .ZN(n5806) );
  NAND2_X1 U6845 ( .A1(n5807), .A2(n5806), .ZN(n6885) );
  NAND2_X1 U6846 ( .A1(n6252), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5815) );
  INV_X1 U6847 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5808) );
  OR2_X1 U6848 ( .A1(n5977), .A2(n5808), .ZN(n5814) );
  NAND2_X1 U6849 ( .A1(n5809), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5810) );
  AND2_X1 U6850 ( .A1(n5816), .A2(n5810), .ZN(n7041) );
  OR2_X1 U6851 ( .A1(n5930), .A2(n7041), .ZN(n5813) );
  INV_X1 U6852 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5811) );
  OR2_X1 U6853 ( .A1(n8182), .A2(n5811), .ZN(n5812) );
  NAND2_X1 U6854 ( .A1(n6252), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5821) );
  INV_X1 U6855 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6647) );
  OR2_X1 U6856 ( .A1(n5977), .A2(n6647), .ZN(n5820) );
  NAND2_X1 U6857 ( .A1(n5816), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5817) );
  AND2_X1 U6858 ( .A1(n5837), .A2(n5817), .ZN(n8856) );
  OR2_X1 U6859 ( .A1(n5930), .A2(n8856), .ZN(n5819) );
  INV_X1 U6860 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6678) );
  OR2_X1 U6861 ( .A1(n8182), .A2(n6678), .ZN(n5818) );
  NAND4_X1 U6862 ( .A1(n5821), .A2(n5820), .A3(n5819), .A4(n5818), .ZN(n8903)
         );
  OR2_X1 U6863 ( .A1(n7263), .A2(n6046), .ZN(n5828) );
  NOR2_X1 U6864 ( .A1(n5825), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5833) );
  OR2_X1 U6865 ( .A1(n5833), .A2(n5672), .ZN(n5826) );
  AOI22_X1 U6866 ( .A1(n6017), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6016), .B2(
        n6940), .ZN(n5827) );
  NAND2_X1 U6867 ( .A1(n5828), .A2(n5827), .ZN(n10670) );
  OR2_X1 U6868 ( .A1(n5830), .A2(n5829), .ZN(n5831) );
  NAND2_X1 U6869 ( .A1(n5845), .A2(n5831), .ZN(n7507) );
  OR2_X1 U6870 ( .A1(n7507), .A2(n6046), .ZN(n5835) );
  NAND2_X1 U6871 ( .A1(n5833), .A2(n5832), .ZN(n5862) );
  NAND2_X1 U6872 ( .A1(n5862), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5847) );
  XNOR2_X1 U6873 ( .A(n5847), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7143) );
  AOI22_X1 U6874 ( .A1(n6017), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6016), .B2(
        n7143), .ZN(n5834) );
  NAND2_X1 U6875 ( .A1(n6252), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5843) );
  INV_X1 U6876 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5836) );
  OR2_X1 U6877 ( .A1(n5977), .A2(n5836), .ZN(n5842) );
  NAND2_X1 U6878 ( .A1(n5837), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5838) );
  AND2_X1 U6879 ( .A1(n5851), .A2(n5838), .ZN(n7294) );
  OR2_X1 U6880 ( .A1(n5930), .A2(n7294), .ZN(n5841) );
  INV_X1 U6881 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5839) );
  OR2_X1 U6882 ( .A1(n8182), .A2(n5839), .ZN(n5840) );
  NAND4_X1 U6883 ( .A1(n5843), .A2(n5842), .A3(n5841), .A4(n5840), .ZN(n8902)
         );
  INV_X1 U6884 ( .A(n8902), .ZN(n7318) );
  OR2_X1 U6885 ( .A1(n7405), .A2(n7318), .ZN(n7358) );
  NAND2_X1 U6886 ( .A1(n7405), .A2(n7318), .ZN(n8556) );
  NAND2_X1 U6887 ( .A1(n7290), .A2(n8552), .ZN(n7289) );
  OR2_X1 U6888 ( .A1(n7405), .A2(n8902), .ZN(n7361) );
  NAND2_X1 U6889 ( .A1(n7289), .A2(n7361), .ZN(n5857) );
  NAND2_X1 U6890 ( .A1(n5847), .A2(n5282), .ZN(n5848) );
  NAND2_X1 U6891 ( .A1(n5848), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5849) );
  AOI22_X1 U6892 ( .A1(n6017), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6016), .B2(
        n7391), .ZN(n5850) );
  NAND2_X1 U6893 ( .A1(n6252), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5856) );
  INV_X1 U6894 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7149) );
  OR2_X1 U6895 ( .A1(n5977), .A2(n7149), .ZN(n5855) );
  NAND2_X1 U6896 ( .A1(n5851), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5852) );
  AND2_X1 U6897 ( .A1(n5867), .A2(n5852), .ZN(n7367) );
  OR2_X1 U6898 ( .A1(n5930), .A2(n7367), .ZN(n5854) );
  INV_X1 U6899 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7374) );
  OR2_X1 U6900 ( .A1(n8182), .A2(n7374), .ZN(n5853) );
  NAND4_X1 U6901 ( .A1(n5856), .A2(n5855), .A3(n5854), .A4(n5853), .ZN(n8901)
         );
  INV_X1 U6902 ( .A(n8901), .ZN(n7605) );
  OR2_X1 U6903 ( .A1(n10743), .A2(n7605), .ZN(n8547) );
  AND2_X1 U6904 ( .A1(n10743), .A2(n7605), .ZN(n8549) );
  INV_X1 U6905 ( .A(n8549), .ZN(n8557) );
  NAND2_X1 U6906 ( .A1(n8547), .A2(n8557), .ZN(n8491) );
  NAND2_X1 U6907 ( .A1(n5857), .A2(n8491), .ZN(n7360) );
  OR2_X1 U6908 ( .A1(n10743), .A2(n8901), .ZN(n7417) );
  XNOR2_X1 U6909 ( .A(n5858), .B(n5859), .ZN(n7543) );
  NAND2_X1 U6910 ( .A1(n7543), .A2(n8473), .ZN(n5866) );
  NAND2_X1 U6911 ( .A1(n5282), .A2(n5285), .ZN(n5861) );
  OAI21_X1 U6912 ( .B1(n5862), .B2(n5861), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5863) );
  MUX2_X1 U6913 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5863), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n5864) );
  AND2_X1 U6914 ( .A1(n5860), .A2(n5864), .ZN(n7456) );
  AOI22_X1 U6915 ( .A1(n6017), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6016), .B2(
        n7456), .ZN(n5865) );
  NAND2_X1 U6916 ( .A1(n6252), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5872) );
  INV_X1 U6917 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7382) );
  OR2_X1 U6918 ( .A1(n5977), .A2(n7382), .ZN(n5871) );
  NAND2_X1 U6919 ( .A1(n5867), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5868) );
  AND2_X1 U6920 ( .A1(n5880), .A2(n5868), .ZN(n7609) );
  OR2_X1 U6921 ( .A1(n5930), .A2(n7609), .ZN(n5870) );
  INV_X1 U6922 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7383) );
  OR2_X1 U6923 ( .A1(n8182), .A2(n7383), .ZN(n5869) );
  NAND4_X1 U6924 ( .A1(n5872), .A2(n5871), .A3(n5870), .A4(n5869), .ZN(n8900)
         );
  INV_X1 U6925 ( .A(n8900), .ZN(n7700) );
  AND2_X1 U6926 ( .A1(n7626), .A2(n7700), .ZN(n8558) );
  INV_X1 U6927 ( .A(n8558), .ZN(n5873) );
  NAND2_X1 U6928 ( .A1(n8548), .A2(n5873), .ZN(n8493) );
  NAND2_X1 U6929 ( .A1(n5162), .A2(n5874), .ZN(n5875) );
  NAND2_X1 U6930 ( .A1(n5876), .A2(n5875), .ZN(n7563) );
  OR2_X1 U6931 ( .A1(n7563), .A2(n6046), .ZN(n5879) );
  NAND2_X1 U6932 ( .A1(n5860), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5877) );
  XNOR2_X1 U6933 ( .A(n5877), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7715) );
  AOI22_X1 U6934 ( .A1(n6017), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6016), .B2(
        n7715), .ZN(n5878) );
  NAND2_X1 U6935 ( .A1(n6252), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5885) );
  INV_X1 U6936 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7457) );
  OR2_X1 U6937 ( .A1(n5977), .A2(n7457), .ZN(n5884) );
  NAND2_X1 U6938 ( .A1(n5880), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5881) );
  AND2_X1 U6939 ( .A1(n5895), .A2(n5881), .ZN(n7704) );
  OR2_X1 U6940 ( .A1(n5930), .A2(n7704), .ZN(n5883) );
  INV_X1 U6941 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7708) );
  OR2_X1 U6942 ( .A1(n8182), .A2(n7708), .ZN(n5882) );
  OR2_X1 U6943 ( .A1(n10771), .A2(n8899), .ZN(n5886) );
  NAND2_X1 U6944 ( .A1(n5887), .A2(n5886), .ZN(n7670) );
  XNOR2_X1 U6945 ( .A(n5889), .B(n5888), .ZN(n7630) );
  NAND2_X1 U6946 ( .A1(n7630), .A2(n8473), .ZN(n5892) );
  OR2_X1 U6947 ( .A1(n6183), .A2(n5672), .ZN(n5890) );
  XNOR2_X1 U6948 ( .A(n5890), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10570) );
  AOI22_X1 U6949 ( .A1(n6017), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6016), .B2(
        n10570), .ZN(n5891) );
  NAND2_X1 U6950 ( .A1(n6252), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5900) );
  INV_X1 U6951 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5893) );
  OR2_X1 U6952 ( .A1(n5977), .A2(n5893), .ZN(n5899) );
  INV_X1 U6953 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5894) );
  OR2_X1 U6954 ( .A1(n8182), .A2(n5894), .ZN(n5898) );
  NAND2_X1 U6955 ( .A1(n5895), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5896) );
  AND2_X1 U6956 ( .A1(n5913), .A2(n5896), .ZN(n7833) );
  OR2_X1 U6957 ( .A1(n5930), .A2(n7833), .ZN(n5897) );
  NAND4_X1 U6958 ( .A1(n5900), .A2(n5899), .A3(n5898), .A4(n5897), .ZN(n7889)
         );
  INV_X1 U6959 ( .A(n7889), .ZN(n7896) );
  NOR2_X1 U6960 ( .A1(n10778), .A2(n7896), .ZN(n8573) );
  INV_X1 U6961 ( .A(n8573), .ZN(n5901) );
  NAND2_X1 U6962 ( .A1(n7670), .A2(n7668), .ZN(n5903) );
  OR2_X1 U6963 ( .A1(n10778), .A2(n7889), .ZN(n5902) );
  NAND2_X1 U6964 ( .A1(n5903), .A2(n5902), .ZN(n7736) );
  NAND2_X1 U6965 ( .A1(n5905), .A2(n5904), .ZN(n5907) );
  NAND2_X1 U6966 ( .A1(n5907), .A2(n5906), .ZN(n7676) );
  OR2_X1 U6967 ( .A1(n7676), .A2(n6046), .ZN(n5911) );
  OR2_X1 U6968 ( .A1(n5908), .A2(n5672), .ZN(n5909) );
  XNOR2_X1 U6969 ( .A(n5909), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7778) );
  AOI22_X1 U6970 ( .A1(n6017), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6016), .B2(
        n7778), .ZN(n5910) );
  NAND2_X1 U6971 ( .A1(n6252), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5918) );
  INV_X1 U6972 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n5912) );
  OR2_X1 U6973 ( .A1(n5977), .A2(n5912), .ZN(n5917) );
  NAND2_X1 U6974 ( .A1(n5913), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5914) );
  AND2_X1 U6975 ( .A1(n5928), .A2(n5914), .ZN(n7901) );
  OR2_X1 U6976 ( .A1(n5930), .A2(n7901), .ZN(n5916) );
  INV_X1 U6977 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7743) );
  OR2_X1 U6978 ( .A1(n8182), .A2(n7743), .ZN(n5915) );
  NAND4_X1 U6979 ( .A1(n5918), .A2(n5917), .A3(n5916), .A4(n5915), .ZN(n8898)
         );
  NAND2_X1 U6980 ( .A1(n7903), .A2(n8898), .ZN(n7737) );
  NAND2_X1 U6981 ( .A1(n7736), .A2(n7737), .ZN(n5919) );
  OR2_X1 U6982 ( .A1(n7903), .A2(n8898), .ZN(n7738) );
  NAND2_X1 U6983 ( .A1(n5919), .A2(n7738), .ZN(n7857) );
  OR2_X1 U6984 ( .A1(n5921), .A2(n5920), .ZN(n5922) );
  NAND2_X1 U6985 ( .A1(n5923), .A2(n5922), .ZN(n7794) );
  NAND2_X1 U6986 ( .A1(n5940), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5924) );
  XNOR2_X1 U6987 ( .A(n5924), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7910) );
  AOI22_X1 U6988 ( .A1(n6017), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6016), .B2(
        n7910), .ZN(n5925) );
  NAND2_X1 U6989 ( .A1(n6252), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5934) );
  INV_X1 U6990 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5927) );
  OR2_X1 U6991 ( .A1(n5977), .A2(n5927), .ZN(n5933) );
  NAND2_X1 U6992 ( .A1(n5928), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5929) );
  AND2_X1 U6993 ( .A1(n5944), .A2(n5929), .ZN(n7952) );
  OR2_X1 U6994 ( .A1(n5930), .A2(n7952), .ZN(n5932) );
  INV_X1 U6995 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7776) );
  OR2_X1 U6996 ( .A1(n8182), .A2(n7776), .ZN(n5931) );
  NAND4_X1 U6997 ( .A1(n5934), .A2(n5933), .A3(n5932), .A4(n5931), .ZN(n7949)
         );
  INV_X1 U6998 ( .A(n7949), .ZN(n8155) );
  OR2_X1 U6999 ( .A1(n7948), .A2(n8155), .ZN(n8579) );
  NAND2_X1 U7000 ( .A1(n7948), .A2(n8155), .ZN(n8580) );
  NAND2_X1 U7001 ( .A1(n7948), .A2(n7949), .ZN(n5935) );
  OR2_X1 U7002 ( .A1(n5937), .A2(n5936), .ZN(n5938) );
  NAND2_X1 U7003 ( .A1(n5939), .A2(n5938), .ZN(n8027) );
  INV_X1 U7004 ( .A(n6003), .ZN(n5941) );
  NAND2_X1 U7005 ( .A1(n5941), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5956) );
  XNOR2_X1 U7006 ( .A(n5956), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7920) );
  AOI22_X1 U7007 ( .A1(n6017), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6016), .B2(
        n7920), .ZN(n5942) );
  NAND2_X1 U7008 ( .A1(n5944), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7009 ( .A1(n5960), .A2(n5945), .ZN(n8152) );
  NAND2_X1 U7010 ( .A1(n6250), .A2(n8152), .ZN(n5950) );
  INV_X1 U7011 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8021) );
  OR2_X1 U7012 ( .A1(n5760), .A2(n8021), .ZN(n5949) );
  INV_X1 U7013 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8024) );
  OR2_X1 U7014 ( .A1(n5977), .A2(n8024), .ZN(n5948) );
  INV_X1 U7015 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5946) );
  OR2_X1 U7016 ( .A1(n8182), .A2(n5946), .ZN(n5947) );
  NAND4_X1 U7017 ( .A1(n5950), .A2(n5949), .A3(n5948), .A4(n5947), .ZN(n8897)
         );
  NAND2_X1 U7018 ( .A1(n8578), .A2(n8897), .ZN(n8584) );
  OR2_X1 U7019 ( .A1(n5952), .A2(n5951), .ZN(n5953) );
  NAND2_X1 U7020 ( .A1(n5954), .A2(n5953), .ZN(n8032) );
  INV_X1 U7021 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U7022 ( .A1(n5956), .A2(n5955), .ZN(n5957) );
  NAND2_X1 U7023 ( .A1(n5957), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5971) );
  XNOR2_X1 U7024 ( .A(n5971), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8927) );
  AOI22_X1 U7025 ( .A1(n6017), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6016), .B2(
        n8927), .ZN(n5958) );
  NAND2_X1 U7026 ( .A1(n5960), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5961) );
  NAND2_X1 U7027 ( .A1(n5975), .A2(n5961), .ZN(n8881) );
  NAND2_X1 U7028 ( .A1(n6250), .A2(n8881), .ZN(n5966) );
  INV_X1 U7029 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8014) );
  OR2_X1 U7030 ( .A1(n5760), .A2(n8014), .ZN(n5965) );
  INV_X1 U7031 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8017) );
  OR2_X1 U7032 ( .A1(n5977), .A2(n8017), .ZN(n5964) );
  INV_X1 U7033 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n5962) );
  OR2_X1 U7034 ( .A1(n8182), .A2(n5962), .ZN(n5963) );
  NAND4_X1 U7035 ( .A1(n5966), .A2(n5965), .A3(n5964), .A4(n5963), .ZN(n8896)
         );
  INV_X1 U7036 ( .A(n8896), .ZN(n8799) );
  OR2_X1 U7037 ( .A1(n8698), .A2(n8799), .ZN(n8587) );
  NAND2_X1 U7038 ( .A1(n8698), .A2(n8799), .ZN(n8588) );
  NAND2_X1 U7039 ( .A1(n8587), .A2(n8588), .ZN(n8582) );
  NAND2_X1 U7040 ( .A1(n8698), .A2(n8896), .ZN(n5967) );
  NAND2_X1 U7041 ( .A1(n7869), .A2(n5967), .ZN(n7962) );
  XNOR2_X1 U7042 ( .A(n5969), .B(n5968), .ZN(n8125) );
  NAND2_X1 U7043 ( .A1(n8125), .A2(n8473), .ZN(n5974) );
  INV_X1 U7044 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5970) );
  NAND2_X1 U7045 ( .A1(n5971), .A2(n5970), .ZN(n5972) );
  NAND2_X1 U7046 ( .A1(n5972), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5987) );
  XNOR2_X1 U7047 ( .A(n5987), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8954) );
  AOI22_X1 U7048 ( .A1(n6017), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8954), .B2(
        n6016), .ZN(n5973) );
  NAND2_X1 U7049 ( .A1(n5975), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5976) );
  NAND2_X1 U7050 ( .A1(n5992), .A2(n5976), .ZN(n8796) );
  NAND2_X1 U7051 ( .A1(n8796), .A2(n6250), .ZN(n5982) );
  NAND2_X1 U7052 ( .A1(n6252), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5981) );
  INV_X1 U7053 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9211) );
  OR2_X1 U7054 ( .A1(n5977), .A2(n9211), .ZN(n5980) );
  INV_X1 U7055 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n5978) );
  OR2_X1 U7056 ( .A1(n8182), .A2(n5978), .ZN(n5979) );
  NAND4_X1 U7057 ( .A1(n5982), .A2(n5981), .A3(n5980), .A4(n5979), .ZN(n8895)
         );
  INV_X1 U7058 ( .A(n8895), .ZN(n8810) );
  NAND2_X1 U7059 ( .A1(n8801), .A2(n8895), .ZN(n5983) );
  XNOR2_X1 U7060 ( .A(n5985), .B(n5984), .ZN(n8210) );
  NAND2_X1 U7061 ( .A1(n8210), .A2(n8473), .ZN(n5991) );
  INV_X1 U7062 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7063 ( .A1(n5987), .A2(n5986), .ZN(n5988) );
  NAND2_X1 U7064 ( .A1(n5988), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5989) );
  XNOR2_X1 U7065 ( .A(n5989), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8984) );
  AOI22_X1 U7066 ( .A1(n8984), .A2(n6016), .B1(n6017), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7067 ( .A1(n5992), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5993) );
  NAND2_X1 U7068 ( .A1(n6007), .A2(n5993), .ZN(n8807) );
  NAND2_X1 U7069 ( .A1(n8807), .A2(n6250), .ZN(n5996) );
  AOI22_X1 U7070 ( .A1(n6252), .A2(P2_REG0_REG_17__SCAN_IN), .B1(n5459), .B2(
        P2_REG1_REG_17__SCAN_IN), .ZN(n5995) );
  INV_X1 U7071 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8957) );
  OR2_X1 U7072 ( .A1(n8182), .A2(n8957), .ZN(n5994) );
  XNOR2_X1 U7073 ( .A(n9206), .B(n9147), .ZN(n8099) );
  INV_X1 U7074 ( .A(n9147), .ZN(n8894) );
  NAND2_X1 U7075 ( .A1(n9206), .A2(n8894), .ZN(n5997) );
  NAND2_X1 U7076 ( .A1(n6000), .A2(n5999), .ZN(n8214) );
  OR2_X1 U7077 ( .A1(n8214), .A2(n6046), .ZN(n6006) );
  NOR2_X1 U7078 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n6001) );
  AND2_X1 U7079 ( .A1(n6175), .A2(n6001), .ZN(n6002) );
  NAND2_X1 U7080 ( .A1(n6003), .A2(n6002), .ZN(n6013) );
  NAND2_X1 U7081 ( .A1(n6013), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6004) );
  XNOR2_X1 U7082 ( .A(n6004), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8997) );
  AOI22_X1 U7083 ( .A1(n6017), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6016), .B2(
        n8997), .ZN(n6005) );
  INV_X1 U7084 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8995) );
  NAND2_X1 U7085 ( .A1(n6007), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6008) );
  NAND2_X1 U7086 ( .A1(n6020), .A2(n6008), .ZN(n9155) );
  NAND2_X1 U7087 ( .A1(n9155), .A2(n6250), .ZN(n6010) );
  AOI22_X1 U7088 ( .A1(n6252), .A2(P2_REG0_REG_18__SCAN_IN), .B1(n5459), .B2(
        P2_REG1_REG_18__SCAN_IN), .ZN(n6009) );
  OAI211_X1 U7089 ( .C1(n8182), .C2(n8995), .A(n6010), .B(n6009), .ZN(n8893)
         );
  OR2_X1 U7090 ( .A1(n8708), .A2(n8893), .ZN(n9131) );
  XNOR2_X1 U7091 ( .A(n6012), .B(n6011), .ZN(n8230) );
  NAND2_X1 U7092 ( .A1(n8230), .A2(n8473), .ZN(n6019) );
  INV_X1 U7093 ( .A(n6013), .ZN(n6014) );
  NAND2_X1 U7094 ( .A1(n6014), .A2(n6111), .ZN(n6015) );
  NAND2_X2 U7095 ( .A1(n6015), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6105) );
  AOI22_X1 U7096 ( .A1(n6017), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9011), .B2(
        n6016), .ZN(n6018) );
  NAND2_X1 U7097 ( .A1(n6020), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6021) );
  NAND2_X1 U7098 ( .A1(n6034), .A2(n6021), .ZN(n9140) );
  NAND2_X1 U7099 ( .A1(n9140), .A2(n6250), .ZN(n6027) );
  INV_X1 U7100 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6024) );
  NAND2_X1 U7101 ( .A1(n6252), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7102 ( .A1(n5459), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6022) );
  OAI211_X1 U7103 ( .C1(n6024), .C2(n8182), .A(n6023), .B(n6022), .ZN(n6025)
         );
  INV_X1 U7104 ( .A(n6025), .ZN(n6026) );
  NAND2_X1 U7105 ( .A1(n6027), .A2(n6026), .ZN(n8892) );
  AND2_X1 U7106 ( .A1(n9131), .A2(n9138), .ZN(n6028) );
  NAND2_X1 U7107 ( .A1(n8708), .A2(n8893), .ZN(n9132) );
  NAND2_X1 U7108 ( .A1(n8766), .A2(n8892), .ZN(n9116) );
  XNOR2_X1 U7109 ( .A(n6030), .B(n6029), .ZN(n8241) );
  NAND2_X1 U7110 ( .A1(n8241), .A2(n8473), .ZN(n6033) );
  INV_X1 U7111 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6031) );
  OR2_X1 U7112 ( .A1(n8475), .A2(n6031), .ZN(n6032) );
  NAND2_X1 U7113 ( .A1(n6034), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U7114 ( .A1(n6049), .A2(n6035), .ZN(n9124) );
  NAND2_X1 U7115 ( .A1(n9124), .A2(n6250), .ZN(n6041) );
  INV_X1 U7116 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n6038) );
  NAND2_X1 U7117 ( .A1(n6252), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U7118 ( .A1(n5459), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6036) );
  OAI211_X1 U7119 ( .C1(n6038), .C2(n8182), .A(n6037), .B(n6036), .ZN(n6039)
         );
  INV_X1 U7120 ( .A(n6039), .ZN(n6040) );
  NAND2_X1 U7121 ( .A1(n6041), .A2(n6040), .ZN(n9103) );
  INV_X1 U7122 ( .A(n9103), .ZN(n9136) );
  OR2_X1 U7123 ( .A1(n9194), .A2(n9136), .ZN(n8614) );
  NAND2_X1 U7124 ( .A1(n9194), .A2(n9136), .ZN(n8615) );
  NAND2_X1 U7125 ( .A1(n8614), .A2(n8615), .ZN(n9114) );
  NAND2_X1 U7126 ( .A1(n6044), .A2(n6043), .ZN(n6045) );
  NAND2_X1 U7127 ( .A1(n5413), .A2(n6045), .ZN(n8244) );
  INV_X1 U7128 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7629) );
  OR2_X1 U7129 ( .A1(n8475), .A2(n7629), .ZN(n6047) );
  NAND2_X1 U7130 ( .A1(n6049), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U7131 ( .A1(n6062), .A2(n6050), .ZN(n9107) );
  NAND2_X1 U7132 ( .A1(n9107), .A2(n6250), .ZN(n6055) );
  INV_X1 U7133 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9108) );
  NAND2_X1 U7134 ( .A1(n6252), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U7135 ( .A1(n5459), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6051) );
  OAI211_X1 U7136 ( .C1(n9108), .C2(n8182), .A(n6052), .B(n6051), .ZN(n6053)
         );
  INV_X1 U7137 ( .A(n6053), .ZN(n6054) );
  NAND2_X1 U7138 ( .A1(n6055), .A2(n6054), .ZN(n9085) );
  INV_X1 U7139 ( .A(n8626), .ZN(n6057) );
  INV_X1 U7140 ( .A(n8622), .ZN(n6056) );
  AOI21_X1 U7141 ( .B1(n9118), .B2(n9099), .A(n9100), .ZN(n9102) );
  XNOR2_X1 U7142 ( .A(n6059), .B(n6058), .ZN(n8253) );
  NAND2_X1 U7143 ( .A1(n8253), .A2(n8473), .ZN(n6061) );
  INV_X1 U7144 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7696) );
  OR2_X1 U7145 ( .A1(n8475), .A2(n7696), .ZN(n6060) );
  NAND2_X1 U7146 ( .A1(n6062), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U7147 ( .A1(n6076), .A2(n6063), .ZN(n9090) );
  NAND2_X1 U7148 ( .A1(n9090), .A2(n6250), .ZN(n6069) );
  INV_X1 U7149 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n6066) );
  NAND2_X1 U7150 ( .A1(n6252), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7151 ( .A1(n5459), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6064) );
  OAI211_X1 U7152 ( .C1(n6066), .C2(n8182), .A(n6065), .B(n6064), .ZN(n6067)
         );
  INV_X1 U7153 ( .A(n6067), .ZN(n6068) );
  NAND2_X1 U7154 ( .A1(n6069), .A2(n6068), .ZN(n9104) );
  NAND2_X1 U7155 ( .A1(n9184), .A2(n9104), .ZN(n8628) );
  INV_X1 U7156 ( .A(n8628), .ZN(n6070) );
  NAND2_X1 U7157 ( .A1(n6086), .A2(n6071), .ZN(n6073) );
  NAND2_X1 U7158 ( .A1(n8267), .A2(n8473), .ZN(n6075) );
  INV_X1 U7159 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7822) );
  OR2_X1 U7160 ( .A1(n8475), .A2(n7822), .ZN(n6074) );
  NAND2_X1 U7161 ( .A1(n6076), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U7162 ( .A1(n6078), .A2(n6077), .ZN(n9079) );
  NAND2_X1 U7163 ( .A1(n9079), .A2(n6250), .ZN(n6084) );
  INV_X1 U7164 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U7165 ( .A1(n6252), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7166 ( .A1(n5459), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6079) );
  OAI211_X1 U7167 ( .C1(n6081), .C2(n8182), .A(n6080), .B(n6079), .ZN(n6082)
         );
  INV_X1 U7168 ( .A(n6082), .ZN(n6083) );
  NAND2_X1 U7169 ( .A1(n8763), .A2(n9086), .ZN(n6161) );
  NAND2_X1 U7170 ( .A1(n6086), .A2(n6085), .ZN(n6088) );
  NAND2_X1 U7171 ( .A1(n8276), .A2(n8473), .ZN(n6092) );
  INV_X1 U7172 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7867) );
  OR2_X1 U7173 ( .A1(n8475), .A2(n7867), .ZN(n6091) );
  INV_X1 U7174 ( .A(n9171), .ZN(n9049) );
  NAND2_X1 U7175 ( .A1(n6093), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U7176 ( .A1(n6095), .A2(n6094), .ZN(n9056) );
  NAND2_X1 U7177 ( .A1(n9056), .A2(n6250), .ZN(n6101) );
  INV_X1 U7178 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7179 ( .A1(n6252), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7180 ( .A1(n5459), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6096) );
  OAI211_X1 U7181 ( .C1(n6098), .C2(n8182), .A(n6097), .B(n6096), .ZN(n6099)
         );
  INV_X1 U7182 ( .A(n6099), .ZN(n6100) );
  AOI21_X1 U7183 ( .B1(n8790), .B2(n9226), .A(n9039), .ZN(n6103) );
  XOR2_X1 U7184 ( .A(n8650), .B(n6237), .Z(n6133) );
  INV_X1 U7185 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6104) );
  INV_X1 U7186 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6112) );
  INV_X1 U7187 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6106) );
  OR2_X1 U7188 ( .A1(n6108), .A2(n6112), .ZN(n6109) );
  OR2_X1 U7189 ( .A1(n6746), .A2(n8675), .ZN(n6116) );
  NAND3_X1 U7190 ( .A1(n6113), .A2(n6112), .A3(n6111), .ZN(n6114) );
  OAI21_X1 U7191 ( .B1(n6013), .B2(n6114), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6115) );
  XNOR2_X1 U7192 ( .A(n6115), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8683) );
  NAND2_X1 U7193 ( .A1(n9011), .A2(n8683), .ZN(n6224) );
  NAND2_X1 U7194 ( .A1(n6116), .A2(n6224), .ZN(n10611) );
  INV_X1 U7195 ( .A(n10611), .ZN(n9145) );
  NAND2_X1 U7196 ( .A1(n6117), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6118) );
  NAND2_X1 U7197 ( .A1(n8191), .A2(n6118), .ZN(n9025) );
  NAND2_X1 U7198 ( .A1(n9025), .A2(n6250), .ZN(n6124) );
  INV_X1 U7199 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n6121) );
  NAND2_X1 U7200 ( .A1(n6252), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U7201 ( .A1(n5459), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6119) );
  OAI211_X1 U7202 ( .C1(n6121), .C2(n8182), .A(n6120), .B(n6119), .ZN(n6122)
         );
  INV_X1 U7203 ( .A(n6122), .ZN(n6123) );
  AND2_X2 U7204 ( .A1(n8516), .A2(n8683), .ZN(n8655) );
  NOR2_X1 U7205 ( .A1(n8654), .A2(n8610), .ZN(n8657) );
  INV_X1 U7206 ( .A(n8657), .ZN(n6129) );
  INV_X1 U7207 ( .A(n6126), .ZN(n8680) );
  NAND2_X1 U7208 ( .A1(n8680), .A2(n8999), .ZN(n6128) );
  NAND2_X1 U7209 ( .A1(n6306), .A2(n6128), .ZN(n6786) );
  INV_X1 U7210 ( .A(n6786), .ZN(n6785) );
  INV_X1 U7211 ( .A(n6135), .ZN(n6923) );
  INV_X1 U7212 ( .A(n6989), .ZN(n8514) );
  NAND2_X1 U7213 ( .A1(n8512), .A2(n8514), .ZN(n6137) );
  NAND2_X1 U7214 ( .A1(n6137), .A2(n6136), .ZN(n8510) );
  NAND2_X1 U7215 ( .A1(n8510), .A2(n10612), .ZN(n6138) );
  INV_X1 U7216 ( .A(n6759), .ZN(n10618) );
  OR2_X1 U7217 ( .A1(n8905), .A2(n10618), .ZN(n8523) );
  NAND2_X1 U7218 ( .A1(n6138), .A2(n8523), .ZN(n7112) );
  NAND2_X1 U7219 ( .A1(n10609), .A2(n10628), .ZN(n8535) );
  NAND2_X1 U7220 ( .A1(n7114), .A2(n8528), .ZN(n7053) );
  XNOR2_X1 U7221 ( .A(n8904), .B(n10636), .ZN(n8529) );
  INV_X1 U7222 ( .A(n8529), .ZN(n8536) );
  NAND2_X1 U7223 ( .A1(n7053), .A2(n8536), .ZN(n6139) );
  OR2_X1 U7224 ( .A1(n8904), .A2(n10636), .ZN(n8538) );
  NAND2_X1 U7225 ( .A1(n6139), .A2(n8538), .ZN(n7034) );
  NOR2_X1 U7226 ( .A1(n8854), .A2(n6885), .ZN(n8543) );
  INV_X1 U7227 ( .A(n8543), .ZN(n6140) );
  AND2_X1 U7228 ( .A1(n8854), .A2(n6885), .ZN(n8533) );
  INV_X1 U7229 ( .A(n8533), .ZN(n8537) );
  AND2_X1 U7230 ( .A1(n6140), .A2(n8537), .ZN(n7036) );
  NAND2_X1 U7231 ( .A1(n7033), .A2(n8537), .ZN(n7099) );
  AND2_X1 U7232 ( .A1(n10670), .A2(n7088), .ZN(n8532) );
  NOR2_X1 U7233 ( .A1(n10670), .A2(n7088), .ZN(n8544) );
  INV_X1 U7234 ( .A(n8544), .ZN(n8550) );
  NAND2_X1 U7235 ( .A1(n7292), .A2(n8551), .ZN(n7293) );
  NAND2_X1 U7236 ( .A1(n8547), .A2(n7358), .ZN(n8567) );
  INV_X1 U7237 ( .A(n8567), .ZN(n6141) );
  NAND2_X1 U7238 ( .A1(n7293), .A2(n6141), .ZN(n6142) );
  OR2_X1 U7239 ( .A1(n10771), .A2(n7828), .ZN(n8564) );
  NAND2_X1 U7240 ( .A1(n8564), .A2(n8548), .ZN(n8566) );
  INV_X1 U7241 ( .A(n8566), .ZN(n6143) );
  AND2_X1 U7242 ( .A1(n10771), .A2(n7828), .ZN(n8570) );
  INV_X1 U7243 ( .A(n8570), .ZN(n7666) );
  AND2_X1 U7244 ( .A1(n7666), .A2(n6145), .ZN(n6144) );
  INV_X1 U7245 ( .A(n8898), .ZN(n7830) );
  OR2_X1 U7246 ( .A1(n7903), .A2(n7830), .ZN(n8574) );
  OR2_X1 U7247 ( .A1(n8569), .A2(n8497), .ZN(n7740) );
  AND2_X1 U7248 ( .A1(n8574), .A2(n7740), .ZN(n6146) );
  NAND2_X1 U7249 ( .A1(n7903), .A2(n7830), .ZN(n8575) );
  NAND2_X1 U7250 ( .A1(n6148), .A2(n8584), .ZN(n8589) );
  NAND2_X1 U7251 ( .A1(n8578), .A2(n8695), .ZN(n6149) );
  INV_X1 U7252 ( .A(n8582), .ZN(n7874) );
  NAND2_X1 U7253 ( .A1(n7873), .A2(n8588), .ZN(n7967) );
  INV_X1 U7254 ( .A(n7967), .ZN(n6150) );
  OR2_X1 U7255 ( .A1(n8801), .A2(n8810), .ZN(n6151) );
  NAND2_X1 U7256 ( .A1(n9206), .A2(n9147), .ZN(n6152) );
  INV_X1 U7257 ( .A(n8893), .ZN(n9137) );
  NAND2_X1 U7258 ( .A1(n8708), .A2(n9137), .ZN(n6153) );
  NAND2_X1 U7259 ( .A1(n6155), .A2(n6153), .ZN(n9154) );
  INV_X1 U7260 ( .A(n8892), .ZN(n9149) );
  OR2_X1 U7261 ( .A1(n8766), .A2(n9149), .ZN(n6156) );
  INV_X1 U7262 ( .A(n9085), .ZN(n9123) );
  OR2_X1 U7263 ( .A1(n9236), .A2(n9123), .ZN(n6158) );
  INV_X1 U7264 ( .A(n9104), .ZN(n9075) );
  NOR2_X1 U7265 ( .A1(n9184), .A2(n9075), .ZN(n6160) );
  INV_X1 U7266 ( .A(n9184), .ZN(n6159) );
  NAND2_X1 U7267 ( .A1(n8634), .A2(n6161), .ZN(n9077) );
  NAND2_X1 U7268 ( .A1(n8763), .A2(n9063), .ZN(n6162) );
  NOR2_X1 U7269 ( .A1(n8819), .A2(n9076), .ZN(n8637) );
  INV_X1 U7270 ( .A(n8637), .ZN(n6163) );
  NAND2_X1 U7271 ( .A1(n9171), .A2(n9064), .ZN(n8641) );
  NAND2_X1 U7272 ( .A1(n9042), .A2(n8485), .ZN(n6164) );
  NAND2_X1 U7273 ( .A1(n8868), .A2(n8790), .ZN(n8646) );
  NAND2_X1 U7274 ( .A1(n6164), .A2(n8646), .ZN(n6165) );
  XOR2_X1 U7275 ( .A(n8650), .B(n6165), .Z(n9036) );
  INV_X1 U7276 ( .A(n8683), .ZN(n7694) );
  NAND2_X1 U7277 ( .A1(n6746), .A2(n7694), .ZN(n10650) );
  NAND2_X1 U7278 ( .A1(n8675), .A2(n8677), .ZN(n6169) );
  AND2_X1 U7279 ( .A1(n8677), .A2(n8683), .ZN(n6171) );
  INV_X1 U7280 ( .A(n6171), .ZN(n6166) );
  NAND2_X1 U7281 ( .A1(n6169), .A2(n6166), .ZN(n6167) );
  AND2_X1 U7282 ( .A1(n10650), .A2(n6167), .ZN(n6168) );
  NAND2_X1 U7283 ( .A1(n6168), .A2(n6915), .ZN(n7539) );
  OR2_X1 U7284 ( .A1(n6747), .A2(n8683), .ZN(n10767) );
  NAND2_X1 U7285 ( .A1(n7539), .A2(n10767), .ZN(n10632) );
  INV_X1 U7286 ( .A(n6169), .ZN(n6170) );
  OR2_X1 U7287 ( .A1(n8610), .A2(n6170), .ZN(n6776) );
  NAND2_X1 U7288 ( .A1(n6171), .A2(n6745), .ZN(n6172) );
  NAND2_X1 U7289 ( .A1(n8610), .A2(n6172), .ZN(n6912) );
  NAND2_X1 U7290 ( .A1(n6776), .A2(n6912), .ZN(n6907) );
  NAND3_X1 U7291 ( .A1(n6175), .A2(n6174), .A3(n6173), .ZN(n6181) );
  NOR2_X1 U7292 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n6179) );
  NOR2_X1 U7293 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n6178) );
  NOR2_X1 U7294 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n6177) );
  NOR2_X1 U7295 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n6176) );
  NAND4_X1 U7296 ( .A1(n6179), .A2(n6178), .A3(n6177), .A4(n6176), .ZN(n6180)
         );
  NOR2_X1 U7297 ( .A1(n6181), .A2(n6180), .ZN(n6182) );
  NAND2_X1 U7298 ( .A1(n6183), .A2(n6182), .ZN(n6205) );
  INV_X1 U7299 ( .A(n6205), .ZN(n6185) );
  INV_X1 U7300 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U7301 ( .A1(n6185), .A2(n6184), .ZN(n6186) );
  NAND2_X1 U7302 ( .A1(n6195), .A2(n6187), .ZN(n6191) );
  NAND2_X1 U7303 ( .A1(n6191), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6189) );
  INV_X1 U7304 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6188) );
  INV_X1 U7305 ( .A(n6195), .ZN(n6190) );
  NAND2_X1 U7306 ( .A1(n6190), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n6192) );
  XNOR2_X1 U7307 ( .A(n7866), .B(P2_B_REG_SCAN_IN), .ZN(n6193) );
  NAND2_X1 U7308 ( .A1(n7868), .A2(n6193), .ZN(n6198) );
  OAI21_X1 U7309 ( .B1(P2_IR_REG_25__SCAN_IN), .B2(P2_IR_REG_24__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7310 ( .A1(n6195), .A2(n6194), .ZN(n6197) );
  INV_X1 U7311 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6196) );
  XNOR2_X1 U7312 ( .A(n6197), .B(n6196), .ZN(n6203) );
  OR2_X1 U7313 ( .A1(n6370), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6200) );
  INV_X1 U7314 ( .A(n6203), .ZN(n7907) );
  NAND2_X1 U7315 ( .A1(n7868), .A2(n7907), .ZN(n6199) );
  NAND2_X1 U7316 ( .A1(n6200), .A2(n6199), .ZN(n6906) );
  OAI21_X1 U7317 ( .B1(n8516), .B2(n10767), .A(n6906), .ZN(n6201) );
  MUX2_X1 U7318 ( .A(n6907), .B(n6201), .S(n6748), .Z(n6220) );
  NAND2_X1 U7319 ( .A1(n6912), .A2(n6906), .ZN(n6218) );
  INV_X1 U7320 ( .A(n7866), .ZN(n6202) );
  NAND2_X1 U7321 ( .A1(n6203), .A2(n6202), .ZN(n6204) );
  OR2_X1 U7322 ( .A1(n6204), .A2(n7868), .ZN(n6775) );
  NAND2_X1 U7323 ( .A1(n6205), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6206) );
  XNOR2_X1 U7324 ( .A(n6206), .B(n6184), .ZN(n6774) );
  AND2_X1 U7325 ( .A1(n6774), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6373) );
  NAND2_X1 U7326 ( .A1(n6775), .A2(n6373), .ZN(n6788) );
  INV_X1 U7327 ( .A(n6788), .ZN(n6771) );
  NOR2_X1 U7328 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6210) );
  NOR4_X1 U7329 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6209) );
  NOR4_X1 U7330 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6208) );
  NOR4_X1 U7331 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6207) );
  NAND4_X1 U7332 ( .A1(n6210), .A2(n6209), .A3(n6208), .A4(n6207), .ZN(n6216)
         );
  NOR4_X1 U7333 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6214) );
  NOR4_X1 U7334 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6213) );
  NOR4_X1 U7335 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6212) );
  NOR4_X1 U7336 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6211) );
  NAND4_X1 U7337 ( .A1(n6214), .A2(n6213), .A3(n6212), .A4(n6211), .ZN(n6215)
         );
  NOR2_X1 U7338 ( .A1(n6216), .A2(n6215), .ZN(n6217) );
  OR2_X1 U7339 ( .A1(n6370), .A2(n6217), .ZN(n6227) );
  AND2_X1 U7340 ( .A1(n6771), .A2(n6227), .ZN(n6909) );
  NAND2_X1 U7341 ( .A1(n6218), .A2(n6909), .ZN(n6219) );
  INV_X2 U7342 ( .A(n10780), .ZN(n10781) );
  MUX2_X1 U7343 ( .A(n6221), .B(n6232), .S(n10781), .Z(n6223) );
  INV_X1 U7344 ( .A(n10650), .ZN(n10779) );
  NAND2_X1 U7345 ( .A1(n10781), .A2(n10779), .ZN(n9213) );
  NAND2_X1 U7346 ( .A1(n6223), .A2(n6222), .ZN(P2_U3486) );
  INV_X1 U7347 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6233) );
  INV_X1 U7348 ( .A(n6747), .ZN(n7859) );
  OR2_X1 U7349 ( .A1(n10650), .A2(n7859), .ZN(n10617) );
  NOR2_X1 U7350 ( .A1(n8675), .A2(n6224), .ZN(n6225) );
  NAND2_X1 U7351 ( .A1(n6746), .A2(n6225), .ZN(n6770) );
  NAND3_X1 U7352 ( .A1(n8610), .A2(n6770), .A3(n10650), .ZN(n6226) );
  NAND2_X1 U7353 ( .A1(n10617), .A2(n6226), .ZN(n6773) );
  INV_X1 U7354 ( .A(n6748), .ZN(n6905) );
  NAND3_X1 U7355 ( .A1(n6905), .A2(n6906), .A3(n6227), .ZN(n6783) );
  INV_X1 U7356 ( .A(n6783), .ZN(n6769) );
  NAND2_X1 U7357 ( .A1(n6773), .A2(n6769), .ZN(n6229) );
  INV_X1 U7358 ( .A(n6906), .ZN(n6911) );
  NAND3_X1 U7359 ( .A1(n6911), .A2(n6748), .A3(n6227), .ZN(n6789) );
  OR2_X1 U7360 ( .A1(n6789), .A2(n6770), .ZN(n6228) );
  NAND2_X1 U7361 ( .A1(n6229), .A2(n6228), .ZN(n8178) );
  NAND2_X1 U7362 ( .A1(n8178), .A2(n6771), .ZN(n6231) );
  OR2_X1 U7363 ( .A1(n6915), .A2(n6788), .ZN(n6784) );
  INV_X1 U7364 ( .A(n6784), .ZN(n8681) );
  INV_X1 U7365 ( .A(n6789), .ZN(n6767) );
  NAND2_X1 U7366 ( .A1(n8681), .A2(n6767), .ZN(n6230) );
  INV_X2 U7367 ( .A(n10782), .ZN(n10785) );
  MUX2_X1 U7368 ( .A(n6233), .B(n6232), .S(n10785), .Z(n6235) );
  OR2_X1 U7369 ( .A1(n10782), .A2(n10650), .ZN(n9252) );
  NAND2_X1 U7370 ( .A1(n8740), .A2(n9237), .ZN(n6234) );
  NAND2_X1 U7371 ( .A1(n6235), .A2(n6234), .ZN(P2_U3454) );
  NAND2_X1 U7372 ( .A1(n8740), .A2(n8890), .ZN(n6236) );
  XNOR2_X1 U7373 ( .A(n6243), .B(SI_28_), .ZN(n6246) );
  NAND2_X1 U7374 ( .A1(n8687), .A2(n8473), .ZN(n6240) );
  INV_X1 U7375 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6238) );
  OR2_X1 U7376 ( .A1(n8475), .A2(n6238), .ZN(n6239) );
  INV_X1 U7377 ( .A(n8654), .ZN(n8889) );
  NAND2_X1 U7378 ( .A1(n6242), .A2(n5552), .ZN(n6257) );
  INV_X1 U7379 ( .A(n6243), .ZN(n6244) );
  INV_X1 U7380 ( .A(SI_28_), .ZN(n9438) );
  NAND2_X1 U7381 ( .A1(n6244), .A2(n9438), .ZN(n6245) );
  INV_X1 U7382 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10405) );
  INV_X1 U7383 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9260) );
  MUX2_X1 U7384 ( .A(n10405), .B(n9260), .S(n8169), .Z(n8161) );
  NAND2_X1 U7385 ( .A1(n9664), .A2(n8473), .ZN(n6249) );
  OR2_X1 U7386 ( .A1(n8475), .A2(n9260), .ZN(n6248) );
  INV_X1 U7387 ( .A(n8191), .ZN(n6251) );
  NAND2_X1 U7388 ( .A1(n6251), .A2(n6250), .ZN(n8186) );
  INV_X1 U7389 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n9016) );
  NAND2_X1 U7390 ( .A1(n5459), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6254) );
  NAND2_X1 U7391 ( .A1(n6252), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6253) );
  OAI211_X1 U7392 ( .C1(n8182), .C2(n9016), .A(n6254), .B(n6253), .ZN(n6255)
         );
  INV_X1 U7393 ( .A(n6255), .ZN(n6256) );
  NAND2_X1 U7394 ( .A1(n8186), .A2(n6256), .ZN(n8888) );
  NAND2_X1 U7395 ( .A1(n9019), .A2(n6296), .ZN(n8667) );
  XNOR2_X1 U7396 ( .A(n6257), .B(n8505), .ZN(n6258) );
  NAND2_X1 U7397 ( .A1(n6258), .A2(n10611), .ZN(n6284) );
  INV_X1 U7398 ( .A(n6263), .ZN(n6259) );
  NAND2_X1 U7399 ( .A1(n8750), .A2(n8654), .ZN(n6260) );
  INV_X1 U7400 ( .A(n8485), .ZN(n8648) );
  OAI211_X1 U7401 ( .C1(n8648), .C2(n6264), .A(n6260), .B(n8651), .ZN(n6261)
         );
  OAI211_X1 U7402 ( .C1(n6262), .C2(n8743), .A(n6274), .B(n6261), .ZN(n6275)
         );
  INV_X1 U7403 ( .A(n6268), .ZN(n6264) );
  AND2_X1 U7404 ( .A1(n8641), .A2(n6267), .ZN(n6265) );
  NAND2_X1 U7405 ( .A1(n6266), .A2(n6265), .ZN(n6272) );
  INV_X1 U7406 ( .A(n6267), .ZN(n6270) );
  AND2_X1 U7407 ( .A1(n8485), .A2(n6268), .ZN(n6269) );
  INV_X1 U7408 ( .A(n8743), .ZN(n6273) );
  AND2_X1 U7409 ( .A1(n6306), .A2(P2_B_REG_SCAN_IN), .ZN(n6276) );
  NOR2_X1 U7410 ( .A1(n9150), .A2(n6276), .ZN(n8187) );
  INV_X1 U7411 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6280) );
  NAND2_X1 U7412 ( .A1(n5459), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6279) );
  INV_X1 U7413 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6277) );
  OR2_X1 U7414 ( .A1(n5760), .A2(n6277), .ZN(n6278) );
  OAI211_X1 U7415 ( .C1(n6280), .C2(n8182), .A(n6279), .B(n6278), .ZN(n6281)
         );
  INV_X1 U7416 ( .A(n6281), .ZN(n6282) );
  AND2_X1 U7417 ( .A1(n8186), .A2(n6282), .ZN(n8479) );
  INV_X1 U7418 ( .A(n8479), .ZN(n8887) );
  AOI22_X1 U7419 ( .A1(n8657), .A2(n6785), .B1(n8187), .B2(n8887), .ZN(n6283)
         );
  INV_X1 U7420 ( .A(n9023), .ZN(n6285) );
  INV_X1 U7421 ( .A(n10767), .ZN(n10655) );
  NOR2_X1 U7422 ( .A1(n9015), .A2(n6286), .ZN(n6294) );
  INV_X1 U7423 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6287) );
  OAI21_X1 U7424 ( .B1(n6294), .B2(n10782), .A(n6289), .ZN(P2_U3456) );
  NAND2_X1 U7425 ( .A1(n9019), .A2(n6290), .ZN(n6293) );
  INV_X1 U7426 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6291) );
  OAI21_X1 U7427 ( .B1(n6294), .B2(n10780), .A(n5553), .ZN(P2_U3488) );
  INV_X1 U7428 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6300) );
  XNOR2_X1 U7429 ( .A(n6295), .B(n8743), .ZN(n9029) );
  MUX2_X1 U7430 ( .A(n6300), .B(n6302), .S(n10781), .Z(n6301) );
  NAND2_X1 U7431 ( .A1(n6301), .A2(n5560), .ZN(P2_U3487) );
  INV_X1 U7432 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6303) );
  MUX2_X1 U7433 ( .A(n6303), .B(n6302), .S(n10785), .Z(n6304) );
  NAND2_X1 U7434 ( .A1(n6304), .A2(n5559), .ZN(P2_U3455) );
  NAND2_X1 U7435 ( .A1(n8610), .A2(n6775), .ZN(n6305) );
  NAND2_X1 U7436 ( .A1(n6305), .A2(n6774), .ZN(n6548) );
  NAND2_X1 U7437 ( .A1(n6548), .A2(n6306), .ZN(n6307) );
  NAND2_X1 U7438 ( .A1(n6307), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NAND2_X1 U7439 ( .A1(n6379), .A2(n6310), .ZN(n6397) );
  NOR2_X1 U7440 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n6313) );
  INV_X1 U7441 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6311) );
  NAND4_X1 U7442 ( .A1(n6313), .A2(n6312), .A3(n6311), .A4(n7048), .ZN(n6316)
         );
  INV_X1 U7443 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6314) );
  NAND4_X1 U7444 ( .A1(n6847), .A2(n6314), .A3(n6473), .A4(n6472), .ZN(n6315)
         );
  NOR2_X2 U7445 ( .A1(n6397), .A2(n4943), .ZN(n7067) );
  INV_X1 U7446 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6318) );
  NOR2_X1 U7447 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n6338) );
  INV_X1 U7448 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6322) );
  INV_X1 U7449 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6341) );
  NAND3_X1 U7450 ( .A1(n6338), .A2(n6322), .A3(n6341), .ZN(n6319) );
  INV_X1 U7451 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6320) );
  NAND2_X1 U7452 ( .A1(n6328), .A2(n6320), .ZN(n6331) );
  NAND2_X1 U7453 ( .A1(n6331), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6321) );
  NOR2_X1 U7454 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n6324) );
  NOR2_X1 U7455 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n6323) );
  INV_X1 U7456 ( .A(n6328), .ZN(n6329) );
  NAND2_X1 U7457 ( .A1(n6329), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6330) );
  NAND2_X1 U7458 ( .A1(n6334), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6333) );
  MUX2_X1 U7459 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6333), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n6336) );
  INV_X1 U7460 ( .A(n6335), .ZN(n6393) );
  NAND2_X1 U7461 ( .A1(n6336), .A2(n6393), .ZN(n7887) );
  NOR2_X1 U7462 ( .A1(n7882), .A2(n7887), .ZN(n6337) );
  INV_X1 U7463 ( .A(n6727), .ZN(n6616) );
  INV_X1 U7464 ( .A(n6338), .ZN(n6339) );
  NAND2_X1 U7465 ( .A1(n6339), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6340) );
  NAND2_X1 U7466 ( .A1(n6602), .A2(n6340), .ZN(n6389) );
  NAND2_X1 U7467 ( .A1(n6391), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6342) );
  XNOR2_X1 U7468 ( .A(n6342), .B(n6341), .ZN(n7771) );
  AND2_X1 U7469 ( .A1(n7771), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6414) );
  INV_X1 U7470 ( .A(n6373), .ZN(n6343) );
  INV_X2 U7471 ( .A(n8989), .ZN(P2_U3893) );
  AND2_X1 U7472 ( .A1(n8169), .A2(P2_U3151), .ZN(n7819) );
  OAI222_X1 U7473 ( .A1(n8472), .A2(n5570), .B1(n10503), .B2(P2_U3151), .C1(
        n4944), .C2(n6822), .ZN(P2_U3293) );
  INV_X1 U7474 ( .A(n6344), .ZN(n6800) );
  INV_X1 U7475 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6345) );
  INV_X1 U7476 ( .A(n8472), .ZN(n9264) );
  OAI222_X1 U7477 ( .A1(n4944), .A2(n6800), .B1(n6564), .B2(P2_U3151), .C1(
        n6345), .C2(n8472), .ZN(P2_U3294) );
  OAI222_X1 U7478 ( .A1(n4944), .A2(n7008), .B1(n6670), .B2(P2_U3151), .C1(
        n6346), .C2(n8472), .ZN(P2_U3292) );
  NAND2_X1 U7479 ( .A1(n8169), .A2(P1_U3086), .ZN(n10406) );
  INV_X1 U7480 ( .A(n10406), .ZN(n10399) );
  NAND2_X1 U7481 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6347) );
  AOI22_X1 U7482 ( .A1(n10399), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(n9973), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6348) );
  OAI21_X1 U7483 ( .B1(n6800), .B2(n10404), .A(n6348), .ZN(P1_U3354) );
  NOR2_X1 U7484 ( .A1(n6349), .A2(n10396), .ZN(n6354) );
  INV_X1 U7485 ( .A(n6354), .ZN(n6351) );
  INV_X1 U7486 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6350) );
  NAND2_X1 U7487 ( .A1(n6351), .A2(n6350), .ZN(n6355) );
  NAND2_X1 U7488 ( .A1(n6355), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6352) );
  INV_X1 U7489 ( .A(n9988), .ZN(n6353) );
  INV_X1 U7490 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7011) );
  OAI222_X1 U7491 ( .A1(P1_U3086), .A2(n6353), .B1(n10404), .B2(n7008), .C1(
        n7011), .C2(n10406), .ZN(P1_U3352) );
  NAND2_X1 U7492 ( .A1(n6354), .A2(P1_IR_REG_2__SCAN_IN), .ZN(n6356) );
  INV_X1 U7493 ( .A(n6821), .ZN(n6696) );
  INV_X1 U7494 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6825) );
  OAI222_X1 U7495 ( .A1(P1_U3086), .A2(n6696), .B1(n10404), .B2(n6822), .C1(
        n6825), .C2(n10406), .ZN(P1_U3353) );
  INV_X1 U7496 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6358) );
  NAND2_X1 U7497 ( .A1(n6911), .A2(n6771), .ZN(n6357) );
  OAI21_X1 U7498 ( .B1(n6771), .B2(n6358), .A(n6357), .ZN(P2_U3377) );
  INV_X1 U7499 ( .A(n6359), .ZN(n7189) );
  NAND2_X1 U7500 ( .A1(n6362), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6363) );
  MUX2_X1 U7501 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6363), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n6364) );
  AND2_X1 U7502 ( .A1(n6360), .A2(n6364), .ZN(n7186) );
  AOI22_X1 U7503 ( .A1(n7186), .A2(P1_STATE_REG_SCAN_IN), .B1(n10399), .B2(
        P2_DATAO_REG_4__SCAN_IN), .ZN(n6365) );
  OAI21_X1 U7504 ( .B1(n7189), .B2(n10404), .A(n6365), .ZN(P1_U3351) );
  INV_X1 U7505 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6366) );
  OAI222_X1 U7506 ( .A1(n4944), .A2(n7189), .B1(n6665), .B2(P2_U3151), .C1(
        n6366), .C2(n8472), .ZN(P2_U3291) );
  INV_X1 U7507 ( .A(n10566), .ZN(n6650) );
  INV_X1 U7508 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6367) );
  OAI222_X1 U7509 ( .A1(n4944), .A2(n7224), .B1(n6650), .B2(P2_U3151), .C1(
        n6367), .C2(n8472), .ZN(P2_U3290) );
  INV_X1 U7510 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7227) );
  NAND2_X1 U7511 ( .A1(n6360), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6368) );
  XNOR2_X1 U7512 ( .A(n6368), .B(P1_IR_REG_5__SCAN_IN), .ZN(n7223) );
  INV_X1 U7513 ( .A(n7223), .ZN(n6369) );
  OAI222_X1 U7514 ( .A1(n10406), .A2(n7227), .B1(n10404), .B2(n7224), .C1(
        n6369), .C2(P1_U3086), .ZN(P1_U3350) );
  NAND2_X1 U7515 ( .A1(n6771), .A2(n6370), .ZN(n6374) );
  INV_X1 U7516 ( .A(n6371), .ZN(n6372) );
  AOI22_X1 U7517 ( .A1(n6374), .A2(n5190), .B1(n6373), .B2(n6372), .ZN(
        P2_U3376) );
  AND2_X1 U7518 ( .A1(n6374), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U7519 ( .A1(n6374), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U7520 ( .A1(n6374), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U7521 ( .A1(n6374), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U7522 ( .A1(n6374), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U7523 ( .A1(n6374), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U7524 ( .A1(n6374), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U7525 ( .A1(n6374), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U7526 ( .A1(n6374), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U7527 ( .A1(n6374), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U7528 ( .A1(n6374), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U7529 ( .A1(n6374), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U7530 ( .A1(n6374), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U7531 ( .A1(n6374), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U7532 ( .A1(n6374), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U7533 ( .A1(n6374), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U7534 ( .A1(n6374), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U7535 ( .A1(n6374), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U7536 ( .A1(n6374), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U7537 ( .A1(n6374), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U7538 ( .A1(n6374), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U7539 ( .A1(n6374), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U7540 ( .A1(n6374), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U7541 ( .A1(n6374), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U7542 ( .A1(n6374), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U7543 ( .A1(n6374), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U7544 ( .A1(n6374), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U7545 ( .A1(n6374), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U7546 ( .A1(n6374), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U7547 ( .A1(n6374), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  INV_X1 U7548 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6454) );
  INV_X1 U7549 ( .A(n6940), .ZN(n6924) );
  OAI222_X1 U7550 ( .A1(n4944), .A2(n7263), .B1(n8472), .B2(n6454), .C1(
        P2_U3151), .C2(n6924), .ZN(P2_U3289) );
  INV_X1 U7551 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6378) );
  OR2_X1 U7552 ( .A1(n6375), .A2(n10396), .ZN(n6377) );
  XNOR2_X1 U7553 ( .A(n6377), .B(n6376), .ZN(n7265) );
  OAI222_X1 U7554 ( .A1(n10406), .A2(n6378), .B1(n10404), .B2(n7263), .C1(
        n7265), .C2(P1_U3086), .ZN(P1_U3349) );
  OR2_X1 U7555 ( .A1(n6379), .A2(n10396), .ZN(n6380) );
  XNOR2_X1 U7556 ( .A(n6380), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7508) );
  AOI22_X1 U7557 ( .A1(n7508), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10399), .ZN(n6381) );
  OAI21_X1 U7558 ( .B1(n7507), .B2(n10404), .A(n6381), .ZN(P1_U3348) );
  INV_X1 U7559 ( .A(n7143), .ZN(n7161) );
  INV_X1 U7560 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6382) );
  OAI222_X1 U7561 ( .A1(n4944), .A2(n7507), .B1(n7161), .B2(P2_U3151), .C1(
        n6382), .C2(n8472), .ZN(P2_U3288) );
  INV_X1 U7562 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6568) );
  NAND2_X1 U7563 ( .A1(n7949), .A2(P2_U3893), .ZN(n6383) );
  OAI21_X1 U7564 ( .B1(P2_U3893), .B2(n6568), .A(n6383), .ZN(P2_U3504) );
  INV_X1 U7565 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6467) );
  NAND2_X1 U7566 ( .A1(n7889), .A2(P2_U3893), .ZN(n6384) );
  OAI21_X1 U7567 ( .B1(P2_U3893), .B2(n6467), .A(n6384), .ZN(P2_U3502) );
  INV_X1 U7568 ( .A(n7771), .ZN(n6385) );
  OR2_X1 U7569 ( .A1(n6727), .A2(n6385), .ZN(n6386) );
  NAND2_X1 U7570 ( .A1(n6386), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6422) );
  INV_X1 U7571 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6601) );
  NAND2_X1 U7572 ( .A1(n6602), .A2(n6601), .ZN(n6387) );
  NAND2_X1 U7573 ( .A1(n6389), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n6390) );
  NAND2_X1 U7574 ( .A1(n6607), .A2(n9881), .ZN(n9868) );
  INV_X1 U7575 ( .A(n9868), .ZN(n6973) );
  NAND2_X1 U7576 ( .A1(n6973), .A2(n7771), .ZN(n6395) );
  INV_X1 U7577 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6426) );
  NAND2_X1 U7578 ( .A1(n6395), .A2(n6797), .ZN(n6421) );
  INV_X1 U7579 ( .A(n6421), .ZN(n6396) );
  NOR2_X1 U7580 ( .A1(n6422), .A2(n6396), .ZN(n10059) );
  NOR2_X1 U7581 ( .A1(n10059), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U7582 ( .A(n7555), .ZN(n6401) );
  NAND2_X1 U7583 ( .A1(n6398), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6399) );
  XNOR2_X1 U7584 ( .A(n6399), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7556) );
  AOI22_X1 U7585 ( .A1(n7556), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10399), .ZN(n6400) );
  OAI21_X1 U7586 ( .B1(n6401), .B2(n10404), .A(n6400), .ZN(P1_U3347) );
  INV_X1 U7587 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6402) );
  INV_X1 U7588 ( .A(n7391), .ZN(n7159) );
  OAI222_X1 U7589 ( .A1(n8472), .A2(n6402), .B1(n4944), .B2(n6401), .C1(
        P2_U3151), .C2(n7159), .ZN(P2_U3287) );
  OR2_X1 U7590 ( .A1(n6398), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6475) );
  NAND2_X1 U7591 ( .A1(n6475), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6406) );
  NAND2_X1 U7592 ( .A1(n6406), .A2(n6472), .ZN(n6403) );
  NAND2_X1 U7593 ( .A1(n6403), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6464) );
  XNOR2_X1 U7594 ( .A(n6464), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7564) );
  AOI22_X1 U7595 ( .A1(n7564), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10399), .ZN(n6404) );
  OAI21_X1 U7596 ( .B1(n7563), .B2(n10404), .A(n6404), .ZN(P1_U3345) );
  INV_X1 U7597 ( .A(n7543), .ZN(n6407) );
  INV_X1 U7598 ( .A(n7456), .ZN(n7447) );
  INV_X1 U7599 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6405) );
  OAI222_X1 U7600 ( .A1(n4944), .A2(n6407), .B1(n7447), .B2(P2_U3151), .C1(
        n6405), .C2(n8472), .ZN(P2_U3286) );
  INV_X1 U7601 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6408) );
  XNOR2_X1 U7602 ( .A(n6406), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7544) );
  INV_X1 U7603 ( .A(n7544), .ZN(n6581) );
  OAI222_X1 U7604 ( .A1(n10406), .A2(n6408), .B1(n10404), .B2(n6407), .C1(
        n6581), .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U7605 ( .A(n7715), .ZN(n7453) );
  INV_X1 U7606 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6409) );
  OAI222_X1 U7607 ( .A1(n4944), .A2(n7563), .B1(n7453), .B2(P2_U3151), .C1(
        n6409), .C2(n8472), .ZN(P2_U3285) );
  INV_X1 U7608 ( .A(n6410), .ZN(n7885) );
  NAND2_X1 U7609 ( .A1(n7885), .A2(P1_B_REG_SCAN_IN), .ZN(n6411) );
  MUX2_X1 U7610 ( .A(P1_B_REG_SCAN_IN), .B(n6411), .S(n7882), .Z(n6413) );
  INV_X1 U7611 ( .A(n7887), .ZN(n6412) );
  INV_X1 U7612 ( .A(n6723), .ZN(n6415) );
  NAND2_X1 U7613 ( .A1(n6727), .A2(n6414), .ZN(n6733) );
  INV_X1 U7614 ( .A(n6733), .ZN(n6730) );
  AND2_X1 U7615 ( .A1(n7885), .A2(n7887), .ZN(n6711) );
  NAND2_X1 U7616 ( .A1(n10408), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6416) );
  OAI21_X1 U7617 ( .B1(n10408), .B2(n6711), .A(n6416), .ZN(P1_U3440) );
  NOR2_X1 U7618 ( .A1(n8688), .A2(n10074), .ZN(n9877) );
  INV_X1 U7619 ( .A(n10074), .ZN(n6419) );
  NOR2_X1 U7620 ( .A1(n8688), .A2(n6419), .ZN(n6624) );
  AOI22_X1 U7621 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(n9877), .B1(n6624), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n6420) );
  XOR2_X1 U7622 ( .A(P1_IR_REG_0__SCAN_IN), .B(n6420), .Z(n6425) );
  NOR2_X1 U7623 ( .A1(n6422), .A2(n6421), .ZN(n6496) );
  INV_X1 U7624 ( .A(n6496), .ZN(n6424) );
  AOI22_X1 U7625 ( .A1(n10059), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n6423) );
  OAI21_X1 U7626 ( .B1(n6425), .B2(n6424), .A(n6423), .ZN(P1_U3243) );
  INV_X1 U7627 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6436) );
  INV_X1 U7628 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6427) );
  NAND2_X1 U7629 ( .A1(n6429), .A2(n6427), .ZN(n10397) );
  XNOR2_X2 U7630 ( .A(n6428), .B(P1_IR_REG_30__SCAN_IN), .ZN(n6437) );
  NAND2_X2 U7631 ( .A1(n6437), .A2(n10402), .ZN(n8218) );
  INV_X1 U7632 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n10072) );
  INV_X1 U7633 ( .A(n6437), .ZN(n8690) );
  NAND2_X1 U7634 ( .A1(n9700), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6434) );
  NAND2_X2 U7635 ( .A1(n8690), .A2(n10402), .ZN(n6815) );
  BUF_X4 U7636 ( .A(n6815), .Z(n9702) );
  INV_X1 U7637 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6432) );
  OR2_X1 U7638 ( .A1(n9702), .A2(n6432), .ZN(n6433) );
  OAI211_X1 U7639 ( .C1(n9705), .C2(n10072), .A(n6434), .B(n6433), .ZN(n10076)
         );
  NAND2_X1 U7640 ( .A1(n10076), .A2(P1_U3973), .ZN(n6435) );
  OAI21_X1 U7641 ( .B1(P1_U3973), .B2(n6436), .A(n6435), .ZN(P1_U3585) );
  INV_X1 U7642 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6565) );
  NAND2_X1 U7643 ( .A1(n7274), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6443) );
  INV_X1 U7644 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7813) );
  OR2_X1 U7645 ( .A1(n9705), .A2(n7813), .ZN(n6442) );
  NAND2_X1 U7646 ( .A1(n6431), .A2(n6437), .ZN(n6835) );
  NAND2_X1 U7647 ( .A1(n7205), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7204) );
  NAND2_X1 U7648 ( .A1(n7276), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7518) );
  INV_X1 U7649 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7517) );
  INV_X1 U7650 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7547) );
  INV_X1 U7651 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7640) );
  INV_X1 U7652 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7436) );
  NAND2_X1 U7653 ( .A1(n7643), .A2(n7436), .ZN(n6438) );
  NAND2_X1 U7654 ( .A1(n7803), .A2(n6438), .ZN(n8118) );
  OR2_X1 U7655 ( .A1(n8324), .A2(n8118), .ZN(n6441) );
  INV_X1 U7656 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n6439) );
  OR2_X1 U7657 ( .A1(n9702), .A2(n6439), .ZN(n6440) );
  NAND4_X1 U7658 ( .A1(n6443), .A2(n6442), .A3(n6441), .A4(n6440), .ZN(n8110)
         );
  NAND2_X1 U7659 ( .A1(n8110), .A2(P1_U3973), .ZN(n6444) );
  OAI21_X1 U7660 ( .B1(n6565), .B2(P1_U3973), .A(n6444), .ZN(P1_U3567) );
  NAND2_X1 U7661 ( .A1(n7274), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6452) );
  INV_X1 U7662 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6445) );
  OR2_X1 U7663 ( .A1(n8218), .A2(n6445), .ZN(n6451) );
  AND2_X1 U7664 ( .A1(n7204), .A2(n6446), .ZN(n6447) );
  OR2_X1 U7665 ( .A1(n6447), .A2(n7276), .ZN(n10695) );
  OR2_X1 U7666 ( .A1(n6835), .A2(n10695), .ZN(n6450) );
  INV_X1 U7667 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6448) );
  OR2_X1 U7668 ( .A1(n6815), .A2(n6448), .ZN(n6449) );
  NAND2_X1 U7669 ( .A1(n8200), .A2(P1_U3973), .ZN(n6453) );
  OAI21_X1 U7670 ( .B1(P1_U3973), .B2(n6454), .A(n6453), .ZN(P1_U3560) );
  NAND2_X1 U7671 ( .A1(n7274), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6461) );
  INV_X1 U7672 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n6455) );
  OR2_X1 U7673 ( .A1(n9702), .A2(n6455), .ZN(n6460) );
  INV_X1 U7674 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7802) );
  NAND2_X1 U7675 ( .A1(n8036), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8037) );
  INV_X1 U7676 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9609) );
  NAND2_X1 U7677 ( .A1(n8233), .A2(n9609), .ZN(n6457) );
  INV_X1 U7678 ( .A(n8247), .ZN(n6456) );
  NAND2_X1 U7679 ( .A1(n6457), .A2(n6456), .ZN(n10207) );
  OR2_X1 U7680 ( .A1(n8324), .A2(n10207), .ZN(n6459) );
  INV_X1 U7681 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n10208) );
  OR2_X1 U7682 ( .A1(n9705), .A2(n10208), .ZN(n6458) );
  NAND4_X1 U7683 ( .A1(n6461), .A2(n6460), .A3(n6459), .A4(n6458), .ZN(n10227)
         );
  NAND2_X1 U7684 ( .A1(n10227), .A2(P1_U3973), .ZN(n6462) );
  OAI21_X1 U7685 ( .B1(n6031), .B2(P1_U3973), .A(n6462), .ZN(P1_U3574) );
  INV_X1 U7686 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6463) );
  INV_X1 U7687 ( .A(n7630), .ZN(n6468) );
  INV_X1 U7688 ( .A(n10570), .ZN(n7720) );
  OAI222_X1 U7689 ( .A1(n8472), .A2(n6463), .B1(n4944), .B2(n6468), .C1(
        P2_U3151), .C2(n7720), .ZN(P2_U3284) );
  NAND2_X1 U7690 ( .A1(n6464), .A2(n6473), .ZN(n6465) );
  NAND2_X1 U7691 ( .A1(n6465), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6466) );
  XNOR2_X1 U7692 ( .A(n6466), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7631) );
  INV_X1 U7693 ( .A(n7631), .ZN(n6469) );
  OAI222_X1 U7694 ( .A1(P1_U3086), .A2(n6469), .B1(n10404), .B2(n6468), .C1(
        n10406), .C2(n6467), .ZN(P1_U3344) );
  INV_X1 U7695 ( .A(n7778), .ZN(n7780) );
  INV_X1 U7696 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6470) );
  OAI222_X1 U7697 ( .A1(n4944), .A2(n7676), .B1(n7780), .B2(P2_U3151), .C1(
        n6470), .C2(n8472), .ZN(P2_U3283) );
  INV_X1 U7698 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6477) );
  INV_X1 U7699 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6471) );
  NAND3_X1 U7700 ( .A1(n6473), .A2(n6472), .A3(n6471), .ZN(n6474) );
  OR2_X1 U7701 ( .A1(n6475), .A2(n6474), .ZN(n6566) );
  NAND2_X1 U7702 ( .A1(n6566), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6476) );
  XNOR2_X1 U7703 ( .A(n6476), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7677) );
  INV_X1 U7704 ( .A(n7677), .ZN(n7254) );
  OAI222_X1 U7705 ( .A1(n10406), .A2(n6477), .B1(n10404), .B2(n7676), .C1(
        n7254), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U7706 ( .A(n7265), .ZN(n6516) );
  NAND2_X1 U7707 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9971) );
  XNOR2_X1 U7708 ( .A(n6821), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n6693) );
  NOR2_X1 U7709 ( .A1(n4977), .A2(n6693), .ZN(n6692) );
  AOI21_X1 U7710 ( .B1(n6821), .B2(P1_REG1_REG_2__SCAN_IN), .A(n6692), .ZN(
        n9983) );
  XNOR2_X1 U7711 ( .A(n9988), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9982) );
  NOR2_X1 U7712 ( .A1(n9983), .A2(n9982), .ZN(n9981) );
  AOI21_X1 U7713 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n9988), .A(n9981), .ZN(
        n6590) );
  INV_X1 U7714 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7025) );
  MUX2_X1 U7715 ( .A(n7025), .B(P1_REG1_REG_4__SCAN_IN), .S(n7186), .Z(n6589)
         );
  NAND2_X1 U7716 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n7223), .ZN(n6478) );
  OAI21_X1 U7717 ( .B1(n7223), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6478), .ZN(
        n6523) );
  INV_X1 U7718 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6479) );
  MUX2_X1 U7719 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6479), .S(n7265), .Z(n6511)
         );
  NOR2_X1 U7720 ( .A1(n6512), .A2(n6511), .ZN(n6510) );
  AOI21_X1 U7721 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n6516), .A(n6510), .ZN(
        n6535) );
  OR2_X1 U7722 ( .A1(n7508), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6481) );
  NAND2_X1 U7723 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n7508), .ZN(n6480) );
  NAND2_X1 U7724 ( .A1(n6481), .A2(n6480), .ZN(n6534) );
  NOR2_X1 U7725 ( .A1(n6535), .A2(n6534), .ZN(n6533) );
  INV_X1 U7726 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6482) );
  MUX2_X1 U7727 ( .A(n6482), .B(P1_REG1_REG_8__SCAN_IN), .S(n7556), .Z(n6484)
         );
  INV_X1 U7728 ( .A(n6483), .ZN(n6486) );
  INV_X1 U7729 ( .A(n6484), .ZN(n6485) );
  AND2_X1 U7730 ( .A1(n6496), .A2(n10074), .ZN(n10024) );
  OAI21_X1 U7731 ( .B1(n6486), .B2(n6485), .A(n10024), .ZN(n6501) );
  NAND2_X1 U7732 ( .A1(n6496), .A2(n8688), .ZN(n10063) );
  INV_X1 U7733 ( .A(n10063), .ZN(n10041) );
  INV_X1 U7734 ( .A(n10059), .ZN(n10044) );
  INV_X1 U7735 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6487) );
  NAND2_X1 U7736 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7766) );
  OAI21_X1 U7737 ( .B1(n10044), .B2(n6487), .A(n7766), .ZN(n6499) );
  MUX2_X1 U7738 ( .A(n6445), .B(P1_REG2_REG_6__SCAN_IN), .S(n7265), .Z(n6488)
         );
  INV_X1 U7739 ( .A(n6488), .ZN(n6514) );
  INV_X1 U7740 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6816) );
  XNOR2_X1 U7741 ( .A(n6821), .B(n6816), .ZN(n6688) );
  INV_X1 U7742 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6736) );
  XNOR2_X1 U7743 ( .A(n9973), .B(n6736), .ZN(n9976) );
  AND2_X1 U7744 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9975) );
  NAND2_X1 U7745 ( .A1(n9976), .A2(n9975), .ZN(n9974) );
  NAND2_X1 U7746 ( .A1(n9973), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6489) );
  NAND2_X1 U7747 ( .A1(n9974), .A2(n6489), .ZN(n6687) );
  AND2_X1 U7748 ( .A1(n6688), .A2(n6687), .ZN(n6689) );
  AND2_X1 U7749 ( .A1(n6821), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6490) );
  INV_X1 U7750 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6834) );
  XNOR2_X1 U7751 ( .A(n9988), .B(n6834), .ZN(n9991) );
  NAND2_X1 U7752 ( .A1(n9990), .A2(n9991), .ZN(n9989) );
  NAND2_X1 U7753 ( .A1(n9988), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6491) );
  NAND2_X1 U7754 ( .A1(n9989), .A2(n6491), .ZN(n6586) );
  INV_X1 U7755 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6492) );
  MUX2_X1 U7756 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6492), .S(n7186), .Z(n6587)
         );
  NAND2_X1 U7757 ( .A1(n6586), .A2(n6587), .ZN(n6585) );
  INV_X1 U7758 ( .A(n6585), .ZN(n6493) );
  NAND2_X1 U7759 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n7223), .ZN(n6494) );
  OAI21_X1 U7760 ( .B1(n7223), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6494), .ZN(
        n6526) );
  NOR2_X1 U7761 ( .A1(n6527), .A2(n6526), .ZN(n6525) );
  NOR2_X1 U7762 ( .A1(n6514), .A2(n6515), .ZN(n6513) );
  AOI21_X1 U7763 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6516), .A(n6513), .ZN(
        n6538) );
  NAND2_X1 U7764 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n7508), .ZN(n6495) );
  OAI21_X1 U7765 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n7508), .A(n6495), .ZN(
        n6537) );
  NOR2_X1 U7766 ( .A1(n6538), .A2(n6537), .ZN(n6536) );
  INV_X1 U7767 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7516) );
  NAND2_X1 U7768 ( .A1(n6496), .A2(n9877), .ZN(n10037) );
  AOI211_X1 U7769 ( .C1(n6497), .C2(n5040), .A(n6575), .B(n10037), .ZN(n6498)
         );
  AOI211_X1 U7770 ( .C1(n10041), .C2(n7556), .A(n6499), .B(n6498), .ZN(n6500)
         );
  OAI21_X1 U7771 ( .B1(n6570), .B2(n6501), .A(n6500), .ZN(P1_U3251) );
  INV_X1 U7772 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6503) );
  NAND2_X1 U7773 ( .A1(n9103), .A2(P2_U3893), .ZN(n6502) );
  OAI21_X1 U7774 ( .B1(P2_U3893), .B2(n6503), .A(n6502), .ZN(P2_U3511) );
  NAND2_X1 U7775 ( .A1(n8247), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8257) );
  INV_X1 U7776 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9618) );
  OR2_X1 U7777 ( .A1(n8256), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6504) );
  NAND2_X1 U7778 ( .A1(n8256), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6702) );
  NAND2_X1 U7779 ( .A1(n6504), .A2(n6702), .ZN(n10157) );
  INV_X1 U7780 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n10158) );
  NAND2_X1 U7781 ( .A1(n8258), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6506) );
  NAND2_X1 U7782 ( .A1(n7274), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6505) );
  OAI211_X1 U7783 ( .C1(n9705), .C2(n10158), .A(n6506), .B(n6505), .ZN(n6507)
         );
  INV_X1 U7784 ( .A(n6507), .ZN(n6508) );
  OAI21_X1 U7785 ( .B1(n10157), .B2(n8324), .A(n6508), .ZN(n10326) );
  NAND2_X1 U7786 ( .A1(n10326), .A2(P1_U3973), .ZN(n6509) );
  OAI21_X1 U7787 ( .B1(P1_U3973), .B2(n7822), .A(n6509), .ZN(P1_U3577) );
  INV_X1 U7788 ( .A(n10024), .ZN(n10067) );
  AOI211_X1 U7789 ( .C1(n6512), .C2(n6511), .A(n10067), .B(n6510), .ZN(n6521)
         );
  AOI211_X1 U7790 ( .C1(n6515), .C2(n6514), .A(n6513), .B(n10037), .ZN(n6520)
         );
  INV_X1 U7791 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6518) );
  NAND2_X1 U7792 ( .A1(n10041), .A2(n6516), .ZN(n6517) );
  NAND2_X1 U7793 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7282) );
  OAI211_X1 U7794 ( .C1(n6518), .C2(n10044), .A(n6517), .B(n7282), .ZN(n6519)
         );
  OR3_X1 U7795 ( .A1(n6521), .A2(n6520), .A3(n6519), .ZN(P1_U3249) );
  AOI211_X1 U7796 ( .C1(n6524), .C2(n6523), .A(n10067), .B(n6522), .ZN(n6532)
         );
  AOI211_X1 U7797 ( .C1(n6527), .C2(n6526), .A(n6525), .B(n10037), .ZN(n6531)
         );
  INV_X1 U7798 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U7799 ( .A1(n10041), .A2(n7223), .ZN(n6528) );
  NAND2_X1 U7800 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n7238) );
  OAI211_X1 U7801 ( .C1(n6529), .C2(n10044), .A(n6528), .B(n7238), .ZN(n6530)
         );
  OR3_X1 U7802 ( .A1(n6532), .A2(n6531), .A3(n6530), .ZN(P1_U3248) );
  AOI211_X1 U7803 ( .C1(n6535), .C2(n6534), .A(n10067), .B(n6533), .ZN(n6545)
         );
  AOI211_X1 U7804 ( .C1(n6538), .C2(n6537), .A(n6536), .B(n10037), .ZN(n6544)
         );
  INV_X1 U7805 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6542) );
  NAND2_X1 U7806 ( .A1(n10041), .A2(n7508), .ZN(n6541) );
  INV_X1 U7807 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6539) );
  NOR2_X1 U7808 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6539), .ZN(n8203) );
  INV_X1 U7809 ( .A(n8203), .ZN(n6540) );
  OAI211_X1 U7810 ( .C1(n6542), .C2(n10044), .A(n6541), .B(n6540), .ZN(n6543)
         );
  OR3_X1 U7811 ( .A1(n6545), .A2(n6544), .A3(n6543), .ZN(P1_U3250) );
  NOR2_X1 U7812 ( .A1(n8679), .A2(P2_U3151), .ZN(n7936) );
  AND2_X1 U7813 ( .A1(n6548), .A2(n7936), .ZN(n6546) );
  MUX2_X1 U7814 ( .A(P2_U3893), .B(n6546), .S(n6126), .Z(n10571) );
  INV_X1 U7815 ( .A(n10571), .ZN(n10504) );
  INV_X1 U7816 ( .A(n6774), .ZN(n7820) );
  NOR2_X1 U7817 ( .A1(n6775), .A2(n7820), .ZN(n6547) );
  OR2_X1 U7818 ( .A1(P2_U3150), .A2(n6547), .ZN(n10569) );
  INV_X1 U7819 ( .A(n10569), .ZN(n10572) );
  NOR2_X1 U7820 ( .A1(n6126), .A2(P2_U3151), .ZN(n9263) );
  NAND2_X1 U7821 ( .A1(n6548), .A2(n9263), .ZN(n10486) );
  OR2_X1 U7822 ( .A1(n10486), .A2(n8999), .ZN(n10559) );
  NAND2_X1 U7823 ( .A1(n6556), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6637) );
  NAND2_X1 U7824 ( .A1(n6564), .A2(n6637), .ZN(n6551) );
  NAND2_X1 U7825 ( .A1(n5518), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6549) );
  OR2_X1 U7826 ( .A1(n6549), .A2(n6556), .ZN(n6550) );
  NAND2_X1 U7827 ( .A1(n6551), .A2(n6550), .ZN(n6636) );
  INV_X1 U7828 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6552) );
  XNOR2_X1 U7829 ( .A(n6636), .B(n6552), .ZN(n6555) );
  INV_X2 U7830 ( .A(n8999), .ZN(n8679) );
  MUX2_X1 U7831 ( .A(n6920), .B(n6553), .S(n8679), .Z(n10487) );
  AND2_X1 U7832 ( .A1(n10487), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n10489) );
  XNOR2_X1 U7833 ( .A(n6653), .B(n10489), .ZN(n6554) );
  NAND2_X1 U7834 ( .A1(P2_U3893), .A2(n6126), .ZN(n10562) );
  OAI22_X1 U7835 ( .A1(n10559), .A2(n6555), .B1(n6554), .B2(n10562), .ZN(n6562) );
  OR2_X1 U7836 ( .A1(n10486), .A2(n8679), .ZN(n10561) );
  NOR2_X1 U7837 ( .A1(n6920), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6557) );
  NAND2_X1 U7838 ( .A1(n6556), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6667) );
  OAI21_X1 U7839 ( .B1(n6564), .B2(n6557), .A(n6667), .ZN(n6559) );
  INV_X1 U7840 ( .A(n6668), .ZN(n6558) );
  AOI21_X1 U7841 ( .B1(n5735), .B2(n6559), .A(n6558), .ZN(n6560) );
  OAI22_X1 U7842 ( .A1(n10561), .A2(n6560), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6961), .ZN(n6561) );
  AOI211_X1 U7843 ( .C1(n10572), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n6562), .B(
        n6561), .ZN(n6563) );
  OAI21_X1 U7844 ( .B1(n6564), .B2(n10504), .A(n6563), .ZN(P2_U3183) );
  INV_X1 U7845 ( .A(n7910), .ZN(n7921) );
  OAI222_X1 U7846 ( .A1(n4944), .A2(n7794), .B1(n8472), .B2(n6565), .C1(
        P2_U3151), .C2(n7921), .ZN(P2_U3282) );
  NOR2_X1 U7847 ( .A1(n6566), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6632) );
  OR2_X1 U7848 ( .A1(n6632), .A2(n10396), .ZN(n6567) );
  XNOR2_X1 U7849 ( .A(n6567), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7795) );
  INV_X1 U7850 ( .A(n7795), .ZN(n6569) );
  OAI222_X1 U7851 ( .A1(P1_U3086), .A2(n6569), .B1(n10406), .B2(n6568), .C1(
        n7794), .C2(n10404), .ZN(P1_U3342) );
  INV_X1 U7852 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10754) );
  AOI22_X1 U7853 ( .A1(n7544), .A2(P1_REG1_REG_9__SCAN_IN), .B1(n10754), .B2(
        n6581), .ZN(n6571) );
  OAI21_X1 U7854 ( .B1(n6572), .B2(n6571), .A(n6868), .ZN(n6583) );
  INV_X1 U7855 ( .A(n10037), .ZN(n10065) );
  NOR2_X1 U7856 ( .A1(n7544), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6573) );
  AOI21_X1 U7857 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n7544), .A(n6573), .ZN(
        n6577) );
  AND2_X1 U7858 ( .A1(n7556), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6574) );
  NAND2_X1 U7859 ( .A1(n6577), .A2(n6576), .ZN(n6871) );
  OAI21_X1 U7860 ( .B1(n6577), .B2(n6576), .A(n6871), .ZN(n6578) );
  NAND2_X1 U7861 ( .A1(n10065), .A2(n6578), .ZN(n6580) );
  NOR2_X1 U7862 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7547), .ZN(n7846) );
  AOI21_X1 U7863 ( .B1(n10059), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7846), .ZN(
        n6579) );
  OAI211_X1 U7864 ( .C1(n10063), .C2(n6581), .A(n6580), .B(n6579), .ZN(n6582)
         );
  AOI21_X1 U7865 ( .B1(n6583), .B2(n10024), .A(n6582), .ZN(n6584) );
  INV_X1 U7866 ( .A(n6584), .ZN(P1_U3252) );
  OAI21_X1 U7867 ( .B1(n6587), .B2(n6586), .A(n6585), .ZN(n6595) );
  AOI211_X1 U7868 ( .C1(n6590), .C2(n6589), .A(n6588), .B(n10067), .ZN(n6591)
         );
  AOI21_X1 U7869 ( .B1(n10041), .B2(n7186), .A(n6591), .ZN(n6594) );
  NAND2_X1 U7870 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n7212) );
  INV_X1 U7871 ( .A(n7212), .ZN(n6592) );
  AOI21_X1 U7872 ( .B1(n10059), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6592), .ZN(
        n6593) );
  OAI211_X1 U7873 ( .C1(n10037), .C2(n6595), .A(n6594), .B(n6593), .ZN(n6625)
         );
  NAND2_X1 U7874 ( .A1(n6737), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6600) );
  INV_X1 U7875 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7309) );
  OR2_X1 U7876 ( .A1(n8218), .A2(n7309), .ZN(n6599) );
  NAND2_X1 U7877 ( .A1(n6813), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6598) );
  INV_X1 U7878 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6596) );
  NAND4_X2 U7879 ( .A1(n6600), .A2(n6599), .A3(n6598), .A4(n6597), .ZN(n9968)
         );
  XNOR2_X1 U7880 ( .A(n6602), .B(n6601), .ZN(n9879) );
  NAND2_X1 U7881 ( .A1(n6603), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6604) );
  NAND2_X1 U7882 ( .A1(n6606), .A2(n6605), .ZN(n10062) );
  NAND2_X1 U7883 ( .A1(n9879), .A2(n10062), .ZN(n6963) );
  OAI211_X2 U7884 ( .C1(n9881), .C2(n6963), .A(n6727), .B(n7350), .ZN(n8447)
         );
  INV_X2 U7885 ( .A(n8447), .ZN(n8459) );
  NAND2_X1 U7886 ( .A1(n9968), .A2(n8459), .ZN(n6613) );
  NOR2_X1 U7887 ( .A1(n8169), .A2(n6608), .ZN(n6610) );
  XNOR2_X1 U7888 ( .A(n6610), .B(n6609), .ZN(n10407) );
  AOI22_X1 U7889 ( .A1(n10592), .A2(n6806), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n6616), .ZN(n6612) );
  NAND2_X1 U7890 ( .A1(n6613), .A2(n6612), .ZN(n6619) );
  NAND2_X1 U7891 ( .A1(n9968), .A2(n6806), .ZN(n6618) );
  NAND2_X1 U7892 ( .A1(n9881), .A2(n10062), .ZN(n6964) );
  AND2_X1 U7893 ( .A1(n6964), .A2(n6614), .ZN(n6615) );
  AOI22_X1 U7894 ( .A1(n10592), .A2(n7012), .B1(P1_REG1_REG_0__SCAN_IN), .B2(
        n6616), .ZN(n6617) );
  NAND2_X1 U7895 ( .A1(n6618), .A2(n6617), .ZN(n6620) );
  NAND2_X1 U7896 ( .A1(n6620), .A2(n6619), .ZN(n6805) );
  OAI21_X1 U7897 ( .B1(n6619), .B2(n6620), .A(n6805), .ZN(n6744) );
  INV_X1 U7898 ( .A(n8688), .ZN(n6832) );
  AOI21_X1 U7899 ( .B1(n6832), .B2(P1_REG2_REG_0__SCAN_IN), .A(
        P1_IR_REG_0__SCAN_IN), .ZN(n6621) );
  NOR2_X1 U7900 ( .A1(n6621), .A2(n9975), .ZN(n6622) );
  AOI211_X1 U7901 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n8688), .A(n6624), .B(n6622), .ZN(n6623) );
  INV_X2 U7902 ( .A(P1_U3973), .ZN(n9967) );
  AOI211_X1 U7903 ( .C1(n6744), .C2(n6624), .A(n6623), .B(n9967), .ZN(n6700)
         );
  OR2_X1 U7904 ( .A1(n6625), .A2(n6700), .ZN(P1_U3247) );
  INV_X1 U7905 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6630) );
  NAND2_X1 U7906 ( .A1(n6134), .A2(n6923), .ZN(n8515) );
  AND2_X1 U7907 ( .A1(n6989), .A2(n8515), .ZN(n8511) );
  INV_X1 U7908 ( .A(n8511), .ZN(n6627) );
  OR2_X1 U7909 ( .A1(n10632), .A2(n10611), .ZN(n6626) );
  NAND2_X1 U7910 ( .A1(n6627), .A2(n6626), .ZN(n6628) );
  NAND2_X1 U7911 ( .A1(n10608), .A2(n6754), .ZN(n6919) );
  OAI211_X1 U7912 ( .C1(n10650), .C2(n6923), .A(n6628), .B(n6919), .ZN(n9218)
         );
  NAND2_X1 U7913 ( .A1(n10785), .A2(n9218), .ZN(n6629) );
  OAI21_X1 U7914 ( .B1(n10785), .B2(n6630), .A(n6629), .ZN(P2_U3390) );
  INV_X1 U7915 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6631) );
  NAND2_X1 U7916 ( .A1(n6632), .A2(n6631), .ZN(n6633) );
  NAND2_X1 U7917 ( .A1(n6633), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7046) );
  XNOR2_X1 U7918 ( .A(n7046), .B(P1_IR_REG_14__SCAN_IN), .ZN(n8063) );
  AOI22_X1 U7919 ( .A1(n8063), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n10399), .ZN(n6634) );
  OAI21_X1 U7920 ( .B1(n8027), .B2(n10404), .A(n6634), .ZN(P1_U3341) );
  INV_X1 U7921 ( .A(n10559), .ZN(n10580) );
  NAND2_X1 U7922 ( .A1(n6665), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6642) );
  INV_X1 U7923 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6635) );
  MUX2_X1 U7924 ( .A(n6635), .B(P2_REG1_REG_4__SCAN_IN), .S(n10543), .Z(n10536) );
  INV_X1 U7925 ( .A(n10503), .ZN(n6654) );
  INV_X1 U7926 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6639) );
  NAND2_X1 U7927 ( .A1(n6636), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6638) );
  NAND2_X1 U7928 ( .A1(n6638), .A2(n6637), .ZN(n10497) );
  NAND2_X1 U7929 ( .A1(n6670), .A2(n6640), .ZN(n6641) );
  NAND2_X1 U7930 ( .A1(P2_REG1_REG_3__SCAN_IN), .A2(n10517), .ZN(n10516) );
  NAND2_X1 U7931 ( .A1(n6641), .A2(n10516), .ZN(n10537) );
  NAND2_X1 U7932 ( .A1(n10536), .A2(n10537), .ZN(n10535) );
  NAND2_X1 U7933 ( .A1(n6650), .A2(n6643), .ZN(n6644) );
  MUX2_X1 U7934 ( .A(n6647), .B(P2_REG1_REG_6__SCAN_IN), .S(n6940), .Z(n6645)
         );
  NAND2_X1 U7935 ( .A1(n6646), .A2(n6645), .ZN(n6939) );
  OAI21_X1 U7936 ( .B1(n6646), .B2(n6645), .A(n6939), .ZN(n6664) );
  MUX2_X1 U7937 ( .A(n6678), .B(n6647), .S(n8679), .Z(n6649) );
  AND2_X1 U7938 ( .A1(n6649), .A2(n6940), .ZN(n6931) );
  INV_X1 U7939 ( .A(n6931), .ZN(n6648) );
  OAI21_X1 U7940 ( .B1(n6940), .B2(n6649), .A(n6648), .ZN(n6660) );
  MUX2_X1 U7941 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8679), .Z(n6651) );
  NAND2_X1 U7942 ( .A1(n6651), .A2(n6650), .ZN(n6658) );
  XNOR2_X1 U7943 ( .A(n6651), .B(n6650), .ZN(n10551) );
  MUX2_X1 U7944 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8679), .Z(n6657) );
  MUX2_X1 U7945 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8679), .Z(n6656) );
  MUX2_X1 U7946 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8679), .Z(n6655) );
  XNOR2_X1 U7947 ( .A(n6655), .B(n6654), .ZN(n10509) );
  AOI22_X1 U7948 ( .A1(n10508), .A2(n10509), .B1(n6655), .B2(n10503), .ZN(
        n10527) );
  XNOR2_X1 U7949 ( .A(n6656), .B(n10520), .ZN(n10526) );
  NAND2_X1 U7950 ( .A1(n10527), .A2(n10526), .ZN(n10525) );
  OAI21_X1 U7951 ( .B1(n6656), .B2(n6670), .A(n10525), .ZN(n10545) );
  XOR2_X1 U7952 ( .A(n10543), .B(n6657), .Z(n10546) );
  NOR2_X1 U7953 ( .A1(n6660), .A2(n6659), .ZN(n6930) );
  AOI21_X1 U7954 ( .B1(n6660), .B2(n6659), .A(n6930), .ZN(n6662) );
  NAND2_X1 U7955 ( .A1(n10572), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n6661) );
  INV_X1 U7956 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9538) );
  OR2_X1 U7957 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9538), .ZN(n8852) );
  OAI211_X1 U7958 ( .C1(n6662), .C2(n10562), .A(n6661), .B(n8852), .ZN(n6663)
         );
  AOI21_X1 U7959 ( .B1(n10580), .B2(n6664), .A(n6663), .ZN(n6685) );
  NAND2_X1 U7960 ( .A1(n6665), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6674) );
  OAI21_X1 U7961 ( .B1(n6665), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6674), .ZN(
        n10533) );
  NAND2_X1 U7962 ( .A1(n10503), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6669) );
  NOR2_X1 U7963 ( .A1(n6671), .A2(n6670), .ZN(n6672) );
  NOR2_X1 U7964 ( .A1(n6673), .A2(n10514), .ZN(n10534) );
  INV_X1 U7965 ( .A(n6674), .ZN(n6675) );
  NOR2_X1 U7966 ( .A1(n10566), .A2(n6676), .ZN(n6677) );
  INV_X1 U7967 ( .A(n6680), .ZN(n6682) );
  MUX2_X1 U7968 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6678), .S(n6940), .Z(n6679)
         );
  INV_X1 U7969 ( .A(n6679), .ZN(n6681) );
  OAI21_X1 U7970 ( .B1(n6682), .B2(n6681), .A(n6926), .ZN(n6683) );
  INV_X1 U7971 ( .A(n10561), .ZN(n10583) );
  NAND2_X1 U7972 ( .A1(n6683), .A2(n10583), .ZN(n6684) );
  OAI211_X1 U7973 ( .C1(n10504), .C2(n6924), .A(n6685), .B(n6684), .ZN(
        P2_U3188) );
  INV_X1 U7974 ( .A(n7920), .ZN(n8911) );
  INV_X1 U7975 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6686) );
  OAI222_X1 U7976 ( .A1(n4944), .A2(n8027), .B1(n8911), .B2(P2_U3151), .C1(
        n6686), .C2(n8472), .ZN(P2_U3281) );
  INV_X1 U7977 ( .A(n6687), .ZN(n6691) );
  INV_X1 U7978 ( .A(n6688), .ZN(n6690) );
  AOI211_X1 U7979 ( .C1(n6691), .C2(n6690), .A(n6689), .B(n10037), .ZN(n6699)
         );
  AOI211_X1 U7980 ( .C1(n4977), .C2(n6693), .A(n6692), .B(n10067), .ZN(n6698)
         );
  INV_X1 U7981 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6841) );
  NOR2_X1 U7982 ( .A1(n6841), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6694) );
  AOI21_X1 U7983 ( .B1(n10059), .B2(P1_ADDR_REG_2__SCAN_IN), .A(n6694), .ZN(
        n6695) );
  OAI21_X1 U7984 ( .B1(n10063), .B2(n6696), .A(n6695), .ZN(n6697) );
  OR4_X1 U7985 ( .A1(n6700), .A2(n6699), .A3(n6698), .A4(n6697), .ZN(P1_U3245)
         );
  NAND2_X1 U7986 ( .A1(n9700), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6707) );
  INV_X1 U7987 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n6701) );
  OR2_X1 U7988 ( .A1(n9702), .A2(n6701), .ZN(n6706) );
  NAND2_X1 U7989 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n6703), .ZN(n8281) );
  OAI21_X1 U7990 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n6703), .A(n8281), .ZN(
        n9601) );
  OR2_X1 U7991 ( .A1(n8324), .A2(n9601), .ZN(n6705) );
  INV_X1 U7992 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n8338) );
  OR2_X1 U7993 ( .A1(n9705), .A2(n8338), .ZN(n6704) );
  NAND4_X1 U7994 ( .A1(n6707), .A2(n6706), .A3(n6705), .A4(n6704), .ZN(n10144)
         );
  NAND2_X1 U7995 ( .A1(n10144), .A2(P1_U3973), .ZN(n6708) );
  OAI21_X1 U7996 ( .B1(n5726), .B2(P1_U3973), .A(n6708), .ZN(P1_U3578) );
  INV_X1 U7997 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6709) );
  NAND2_X1 U7998 ( .A1(n6723), .A2(n6709), .ZN(n6710) );
  NAND2_X1 U7999 ( .A1(n7882), .A2(n7887), .ZN(n10395) );
  INV_X1 U8000 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6712) );
  AOI21_X1 U8001 ( .B1(n6723), .B2(n6712), .A(n6711), .ZN(n7303) );
  NOR4_X1 U8002 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6721) );
  NOR4_X1 U8003 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6720) );
  OR4_X1 U8004 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6718) );
  NOR4_X1 U8005 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6716) );
  NOR4_X1 U8006 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6715) );
  NOR4_X1 U8007 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6714) );
  NOR4_X1 U8008 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6713) );
  NAND4_X1 U8009 ( .A1(n6716), .A2(n6715), .A3(n6714), .A4(n6713), .ZN(n6717)
         );
  NOR4_X1 U8010 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        n6718), .A4(n6717), .ZN(n6719) );
  NAND3_X1 U8011 ( .A1(n6721), .A2(n6720), .A3(n6719), .ZN(n6722) );
  NAND2_X1 U8012 ( .A1(n6723), .A2(n6722), .ZN(n7301) );
  NAND3_X1 U8013 ( .A1(n7300), .A2(n7303), .A3(n7301), .ZN(n6734) );
  NOR2_X1 U8014 ( .A1(n6734), .A2(n6733), .ZN(n6729) );
  INV_X1 U8015 ( .A(n6963), .ZN(n9945) );
  INV_X1 U8016 ( .A(n6607), .ZN(n9830) );
  INV_X1 U8017 ( .A(n9881), .ZN(n9709) );
  NAND2_X1 U8018 ( .A1(n9830), .A2(n9709), .ZN(n6965) );
  AND2_X1 U8019 ( .A1(n10820), .A2(n9868), .ZN(n6724) );
  INV_X1 U8020 ( .A(n9651), .ZN(n9632) );
  INV_X1 U8021 ( .A(n9879), .ZN(n9946) );
  NAND2_X1 U8022 ( .A1(n9946), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7426) );
  NAND2_X1 U8023 ( .A1(n10791), .A2(n7426), .ZN(n6725) );
  NAND2_X1 U8024 ( .A1(n6734), .A2(n6725), .ZN(n6728) );
  NAND2_X1 U8025 ( .A1(n6973), .A2(n6963), .ZN(n6726) );
  AND3_X1 U8026 ( .A1(n6727), .A2(n6726), .A3(n7771), .ZN(n6985) );
  NAND2_X1 U8027 ( .A1(n6728), .A2(n6985), .ZN(n7017) );
  NOR2_X1 U8028 ( .A1(n7017), .A2(P1_U3086), .ZN(n6856) );
  INV_X1 U8029 ( .A(n6856), .ZN(n6732) );
  INV_X1 U8030 ( .A(n6965), .ZN(n10593) );
  AND2_X1 U8031 ( .A1(n10593), .A2(n9946), .ZN(n7306) );
  NAND2_X1 U8032 ( .A1(n6729), .A2(n7306), .ZN(n6731) );
  NOR2_X1 U8033 ( .A1(n10257), .A2(n10062), .ZN(n6982) );
  NAND2_X1 U8034 ( .A1(n6731), .A2(n10847), .ZN(n9642) );
  AOI22_X1 U8035 ( .A1(n6732), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n10592), .B2(
        n9642), .ZN(n6743) );
  OR2_X1 U8036 ( .A1(n9868), .A2(n6963), .ZN(n7310) );
  OR2_X1 U8037 ( .A1(n6733), .A2(n7310), .ZN(n9874) );
  NOR2_X1 U8038 ( .A1(n6734), .A2(n9874), .ZN(n6833) );
  NAND2_X1 U8039 ( .A1(n6833), .A2(n8688), .ZN(n9655) );
  INV_X1 U8040 ( .A(n9655), .ZN(n9582) );
  INV_X1 U8041 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6735) );
  OR2_X1 U8042 ( .A1(n6815), .A2(n6735), .ZN(n6741) );
  OR2_X1 U8043 ( .A1(n8218), .A2(n6736), .ZN(n6740) );
  NAND2_X1 U8044 ( .A1(n6813), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6739) );
  INV_X1 U8045 ( .A(n6835), .ZN(n6737) );
  NAND4_X1 U8046 ( .A1(n6741), .A2(n6740), .A3(n6739), .A4(n6738), .ZN(n6968)
         );
  NAND2_X1 U8047 ( .A1(n9582), .A2(n10591), .ZN(n6742) );
  OAI211_X1 U8048 ( .C1(n9632), .C2(n6744), .A(n6743), .B(n6742), .ZN(P1_U3232) );
  INV_X1 U8049 ( .A(n8675), .ZN(n6745) );
  INV_X1 U8050 ( .A(n6762), .ZN(n6763) );
  XNOR2_X1 U8051 ( .A(n6751), .B(n10598), .ZN(n6755) );
  INV_X1 U8052 ( .A(n6755), .ZN(n6753) );
  INV_X1 U8053 ( .A(n6754), .ZN(n6752) );
  NAND2_X1 U8054 ( .A1(n6753), .A2(n6752), .ZN(n6758) );
  NAND2_X1 U8055 ( .A1(n6755), .A2(n6754), .ZN(n6756) );
  NAND2_X1 U8056 ( .A1(n6954), .A2(n6955), .ZN(n6953) );
  NAND2_X1 U8057 ( .A1(n6953), .A2(n6758), .ZN(n6947) );
  XNOR2_X1 U8058 ( .A(n6760), .B(n8905), .ZN(n6948) );
  XNOR2_X1 U8059 ( .A(n6751), .B(n10636), .ZN(n6764) );
  NOR2_X1 U8060 ( .A1(n6764), .A2(n8904), .ZN(n6880) );
  AOI21_X1 U8061 ( .B1(n6764), .B2(n8904), .A(n6880), .ZN(n6765) );
  OAI21_X1 U8062 ( .B1(n6766), .B2(n6765), .A(n6883), .ZN(n6795) );
  NAND3_X1 U8063 ( .A1(n8610), .A2(n10650), .A3(n6767), .ZN(n6768) );
  NAND2_X1 U8064 ( .A1(n6768), .A2(n6770), .ZN(n6772) );
  OR2_X1 U8065 ( .A1(n6770), .A2(n6769), .ZN(n6777) );
  NAND3_X1 U8066 ( .A1(n6772), .A2(n6771), .A3(n6777), .ZN(n8870) );
  INV_X1 U8067 ( .A(n8870), .ZN(n8848) );
  NAND2_X1 U8068 ( .A1(n6773), .A2(n6789), .ZN(n6779) );
  AND4_X1 U8069 ( .A1(n6777), .A2(n6776), .A3(n6775), .A4(n6774), .ZN(n6778)
         );
  NAND2_X1 U8070 ( .A1(n6779), .A2(n6778), .ZN(n6780) );
  NAND2_X1 U8071 ( .A1(n6780), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6782) );
  NAND2_X1 U8072 ( .A1(n8681), .A2(n6783), .ZN(n6781) );
  NAND2_X1 U8073 ( .A1(n6782), .A2(n6781), .ZN(n8880) );
  INV_X1 U8074 ( .A(n8880), .ZN(n7900) );
  NOR2_X1 U8075 ( .A1(n7900), .A2(n7059), .ZN(n6794) );
  NOR2_X1 U8076 ( .A1(n6784), .A2(n6783), .ZN(n6787) );
  NAND2_X1 U8077 ( .A1(n6787), .A2(n6785), .ZN(n8878) );
  NAND2_X1 U8078 ( .A1(n8876), .A2(n5079), .ZN(n6792) );
  OR2_X1 U8079 ( .A1(n10650), .A2(n6788), .ZN(n8176) );
  OR2_X1 U8080 ( .A1(n8176), .A2(n6789), .ZN(n6790) );
  NAND2_X1 U8081 ( .A1(n10620), .A2(n6790), .ZN(n8867) );
  NOR2_X1 U8082 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9523), .ZN(n10538) );
  AOI21_X1 U8083 ( .B1(n8867), .B2(n7061), .A(n10538), .ZN(n6791) );
  OAI211_X1 U8084 ( .C1(n5525), .C2(n8878), .A(n6792), .B(n6791), .ZN(n6793)
         );
  AOI211_X1 U8085 ( .C1(n6795), .C2(n8848), .A(n6794), .B(n6793), .ZN(n6796)
         );
  INV_X1 U8086 ( .A(n6796), .ZN(P2_U3170) );
  NAND2_X1 U8087 ( .A1(n10591), .A2(n6806), .ZN(n6802) );
  NAND2_X1 U8088 ( .A1(n7007), .A2(n9973), .ZN(n6798) );
  OAI211_X2 U8089 ( .C1(n7185), .C2(n6800), .A(n6799), .B(n6798), .ZN(n7347)
         );
  NAND2_X1 U8090 ( .A1(n7347), .A2(n4947), .ZN(n6801) );
  NAND2_X1 U8091 ( .A1(n6802), .A2(n6801), .ZN(n6803) );
  NAND2_X1 U8092 ( .A1(n9890), .A2(n6829), .ZN(n6804) );
  NAND2_X1 U8093 ( .A1(n6805), .A2(n6804), .ZN(n6809) );
  NAND2_X1 U8094 ( .A1(n6808), .A2(n6809), .ZN(n6851) );
  AND2_X1 U8095 ( .A1(n7347), .A2(n6806), .ZN(n6807) );
  AOI21_X1 U8096 ( .B1(n10591), .B2(n8459), .A(n6807), .ZN(n6854) );
  NAND2_X1 U8097 ( .A1(n6851), .A2(n6854), .ZN(n6812) );
  NAND2_X1 U8098 ( .A1(n6812), .A2(n6852), .ZN(n7001) );
  OR2_X1 U8099 ( .A1(n6835), .A2(n6841), .ZN(n6820) );
  NAND2_X1 U8100 ( .A1(n7274), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6819) );
  INV_X1 U8101 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6814) );
  OR2_X1 U8102 ( .A1(n9702), .A2(n6814), .ZN(n6818) );
  OR2_X1 U8103 ( .A1(n8218), .A2(n6816), .ZN(n6817) );
  NAND4_X2 U8104 ( .A1(n6820), .A2(n6819), .A3(n6818), .A4(n6817), .ZN(n9966)
         );
  NAND2_X1 U8105 ( .A1(n9966), .A2(n6806), .ZN(n6827) );
  NAND2_X1 U8106 ( .A1(n7007), .A2(n6821), .ZN(n6824) );
  OR2_X1 U8107 ( .A1(n7185), .A2(n6822), .ZN(n6823) );
  NAND2_X1 U8108 ( .A1(n7472), .A2(n4947), .ZN(n6826) );
  NAND2_X1 U8109 ( .A1(n6827), .A2(n6826), .ZN(n6830) );
  XNOR2_X1 U8110 ( .A(n6830), .B(n8460), .ZN(n7002) );
  AND2_X1 U8111 ( .A1(n7472), .A2(n6806), .ZN(n6831) );
  AOI21_X1 U8112 ( .B1(n9966), .B2(n8459), .A(n6831), .ZN(n7003) );
  XNOR2_X1 U8113 ( .A(n7002), .B(n7003), .ZN(n7000) );
  XNOR2_X1 U8114 ( .A(n7001), .B(n7000), .ZN(n6844) );
  INV_X1 U8115 ( .A(n10591), .ZN(n6979) );
  NAND2_X1 U8116 ( .A1(n6833), .A2(n6832), .ZN(n9639) );
  NAND2_X1 U8117 ( .A1(n7274), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6840) );
  OR2_X1 U8118 ( .A1(n8218), .A2(n6834), .ZN(n6839) );
  OR2_X1 U8119 ( .A1(n6835), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6838) );
  INV_X1 U8120 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6836) );
  OR2_X1 U8121 ( .A1(n6815), .A2(n6836), .ZN(n6837) );
  INV_X1 U8122 ( .A(n9965), .ZN(n6980) );
  OAI22_X1 U8123 ( .A1(n6979), .A2(n9639), .B1(n9655), .B2(n6980), .ZN(n6843)
         );
  OAI22_X1 U8124 ( .A1(n9661), .A2(n6972), .B1(n6856), .B2(n6841), .ZN(n6842)
         );
  AOI211_X1 U8125 ( .C1(n9651), .C2(n6844), .A(n6843), .B(n6842), .ZN(n6845)
         );
  INV_X1 U8126 ( .A(n6845), .ZN(P1_U3237) );
  INV_X1 U8127 ( .A(n8927), .ZN(n8936) );
  INV_X1 U8128 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6846) );
  OAI222_X1 U8129 ( .A1(n4944), .A2(n8032), .B1(n8936), .B2(P2_U3151), .C1(
        n6846), .C2(n8472), .ZN(P2_U3280) );
  INV_X1 U8130 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6850) );
  NAND2_X1 U8131 ( .A1(n7046), .A2(n6847), .ZN(n6848) );
  NAND2_X1 U8132 ( .A1(n6848), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6849) );
  XNOR2_X1 U8133 ( .A(n6849), .B(P1_IR_REG_15__SCAN_IN), .ZN(n8064) );
  INV_X1 U8134 ( .A(n8064), .ZN(n10003) );
  OAI222_X1 U8135 ( .A1(n10406), .A2(n6850), .B1(n10404), .B2(n8032), .C1(
        n10003), .C2(P1_U3086), .ZN(P1_U3340) );
  NAND2_X1 U8136 ( .A1(n6852), .A2(n6851), .ZN(n6853) );
  XOR2_X1 U8137 ( .A(n6854), .B(n6853), .Z(n6859) );
  INV_X1 U8138 ( .A(n9968), .ZN(n7177) );
  INV_X1 U8139 ( .A(n9966), .ZN(n7176) );
  OAI22_X1 U8140 ( .A1(n7177), .A2(n9639), .B1(n9655), .B2(n7176), .ZN(n6858)
         );
  INV_X1 U8141 ( .A(n7347), .ZN(n9889) );
  INV_X1 U8142 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6855) );
  OAI22_X1 U8143 ( .A1(n9661), .A2(n9889), .B1(n6856), .B2(n6855), .ZN(n6857)
         );
  AOI211_X1 U8144 ( .C1(n9651), .C2(n6859), .A(n6858), .B(n6857), .ZN(n6860)
         );
  INV_X1 U8145 ( .A(n6860), .ZN(P1_U3222) );
  INV_X1 U8146 ( .A(n8905), .ZN(n7111) );
  NAND2_X1 U8147 ( .A1(n8876), .A2(n8904), .ZN(n6862) );
  NOR2_X1 U8148 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9500), .ZN(n10518) );
  AOI21_X1 U8149 ( .B1(n8867), .B2(n7116), .A(n10518), .ZN(n6861) );
  OAI211_X1 U8150 ( .C1(n7111), .C2(n8878), .A(n6862), .B(n6861), .ZN(n6866)
         );
  AOI211_X1 U8151 ( .C1(n6864), .C2(n6863), .A(n8870), .B(n5038), .ZN(n6865)
         );
  AOI211_X1 U8152 ( .C1(n9500), .C2(n8880), .A(n6866), .B(n6865), .ZN(n6867)
         );
  INV_X1 U8153 ( .A(n6867), .ZN(P2_U3158) );
  OAI21_X1 U8154 ( .B1(n7544), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6868), .ZN(
        n6870) );
  MUX2_X1 U8155 ( .A(n10765), .B(P1_REG1_REG_10__SCAN_IN), .S(n7564), .Z(n6869) );
  NOR2_X1 U8156 ( .A1(n6870), .A2(n6869), .ZN(n7071) );
  AOI211_X1 U8157 ( .C1(n6870), .C2(n6869), .A(n7071), .B(n10067), .ZN(n6879)
         );
  OAI21_X1 U8158 ( .B1(n7544), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6871), .ZN(
        n6874) );
  NAND2_X1 U8159 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n7564), .ZN(n6872) );
  OAI21_X1 U8160 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n7564), .A(n6872), .ZN(
        n6873) );
  NOR2_X1 U8161 ( .A1(n6873), .A2(n6874), .ZN(n7074) );
  AOI211_X1 U8162 ( .C1(n6874), .C2(n6873), .A(n7074), .B(n10037), .ZN(n6878)
         );
  INV_X1 U8163 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6876) );
  NAND2_X1 U8164 ( .A1(n10041), .A2(n7564), .ZN(n6875) );
  NAND2_X1 U8165 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9310) );
  OAI211_X1 U8166 ( .C1(n6876), .C2(n10044), .A(n6875), .B(n9310), .ZN(n6877)
         );
  OR3_X1 U8167 ( .A1(n6879), .A2(n6878), .A3(n6877), .ZN(P1_U3253) );
  INV_X1 U8168 ( .A(n6880), .ZN(n6881) );
  XNOR2_X1 U8169 ( .A(n6885), .B(n6751), .ZN(n7086) );
  XNOR2_X1 U8170 ( .A(n7086), .B(n8854), .ZN(n6882) );
  AND3_X1 U8171 ( .A1(n6883), .A2(n6882), .A3(n6881), .ZN(n6884) );
  OAI21_X1 U8172 ( .B1(n7085), .B2(n6884), .A(n8848), .ZN(n6890) );
  INV_X1 U8173 ( .A(n8904), .ZN(n7110) );
  NAND2_X1 U8174 ( .A1(n8876), .A2(n8903), .ZN(n6887) );
  NOR2_X1 U8175 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5678), .ZN(n10565) );
  AOI21_X1 U8176 ( .B1(n8867), .B2(n6885), .A(n10565), .ZN(n6886) );
  OAI211_X1 U8177 ( .C1(n7110), .C2(n8878), .A(n6887), .B(n6886), .ZN(n6888)
         );
  INV_X1 U8178 ( .A(n6888), .ZN(n6889) );
  OAI211_X1 U8179 ( .C1(n7041), .C2(n7900), .A(n6890), .B(n6889), .ZN(P2_U3167) );
  NOR2_X1 U8180 ( .A1(n8880), .A2(P2_U3151), .ZN(n6962) );
  INV_X1 U8181 ( .A(n8867), .ZN(n8884) );
  OAI22_X1 U8182 ( .A1(n8884), .A2(n6923), .B1(n8511), .B2(n8870), .ZN(n6891)
         );
  AOI21_X1 U8183 ( .B1(n8876), .B2(n6754), .A(n6891), .ZN(n6892) );
  OAI21_X1 U8184 ( .B1(n6962), .B2(n6893), .A(n6892), .ZN(P2_U3172) );
  NAND2_X1 U8185 ( .A1(n8305), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6903) );
  INV_X2 U8186 ( .A(n7274), .ZN(n8307) );
  INV_X1 U8187 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6894) );
  OR2_X1 U8188 ( .A1(n8307), .A2(n6894), .ZN(n6902) );
  INV_X1 U8189 ( .A(n8281), .ZN(n6895) );
  NAND2_X1 U8190 ( .A1(n6895), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8292) );
  INV_X1 U8191 ( .A(n8292), .ZN(n6896) );
  NAND2_X1 U8192 ( .A1(n6896), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8322) );
  INV_X1 U8193 ( .A(n8322), .ZN(n6898) );
  AND2_X1 U8194 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .ZN(n6897) );
  NAND2_X1 U8195 ( .A1(n6898), .A2(n6897), .ZN(n10099) );
  OR2_X1 U8196 ( .A1(n8324), .A2(n10099), .ZN(n6901) );
  INV_X1 U8197 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6899) );
  OR2_X1 U8198 ( .A1(n9702), .A2(n6899), .ZN(n6900) );
  NAND2_X1 U8199 ( .A1(n9967), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6904) );
  OAI21_X1 U8200 ( .B1(n10280), .B2(n9967), .A(n6904), .ZN(P1_U3583) );
  MUX2_X1 U8201 ( .A(n6907), .B(n6906), .S(n6905), .Z(n6908) );
  INV_X1 U8202 ( .A(n6908), .ZN(n6914) );
  INV_X1 U8203 ( .A(n6909), .ZN(n6910) );
  AOI21_X1 U8204 ( .B1(n6912), .B2(n6911), .A(n6910), .ZN(n6913) );
  NAND2_X1 U8205 ( .A1(n6914), .A2(n6913), .ZN(n6918) );
  NOR2_X1 U8206 ( .A1(n6918), .A2(n10617), .ZN(n9111) );
  INV_X1 U8207 ( .A(n10620), .ZN(n9156) );
  INV_X1 U8208 ( .A(n6915), .ZN(n6916) );
  NOR4_X1 U8209 ( .A1(n6918), .A2(n8511), .A3(n6916), .A4(n10779), .ZN(n6917)
         );
  AOI21_X1 U8210 ( .B1(n9156), .B2(P2_REG3_REG_0__SCAN_IN), .A(n6917), .ZN(
        n6922) );
  NAND2_X2 U8211 ( .A1(n6918), .A2(n10620), .ZN(n10626) );
  MUX2_X1 U8212 ( .A(n6920), .B(n6919), .S(n10626), .Z(n6921) );
  OAI211_X1 U8213 ( .C1(n9159), .C2(n6923), .A(n6922), .B(n6921), .ZN(P2_U3233) );
  NAND2_X1 U8214 ( .A1(n6924), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6925) );
  AOI21_X1 U8215 ( .B1(n5839), .B2(n6927), .A(n7144), .ZN(n6945) );
  MUX2_X1 U8216 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8679), .Z(n6928) );
  NOR2_X1 U8217 ( .A1(n6928), .A2(n7161), .ZN(n7148) );
  AOI21_X1 U8218 ( .B1(n6928), .B2(n7161), .A(n7148), .ZN(n6929) );
  INV_X1 U8219 ( .A(n6929), .ZN(n6933) );
  NOR2_X1 U8220 ( .A1(n6931), .A2(n6930), .ZN(n6932) );
  NOR2_X1 U8221 ( .A1(n6932), .A2(n6933), .ZN(n7147) );
  AOI21_X1 U8222 ( .B1(n6933), .B2(n6932), .A(n7147), .ZN(n6935) );
  NOR2_X1 U8223 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5680), .ZN(n7091) );
  INV_X1 U8224 ( .A(n7091), .ZN(n6934) );
  OAI21_X1 U8225 ( .B1(n6935), .B2(n10562), .A(n6934), .ZN(n6938) );
  INV_X1 U8226 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6936) );
  NOR2_X1 U8227 ( .A1(n10569), .A2(n6936), .ZN(n6937) );
  AOI211_X1 U8228 ( .C1(n10571), .C2(n7143), .A(n6938), .B(n6937), .ZN(n6944)
         );
  OAI21_X1 U8229 ( .B1(P2_REG1_REG_7__SCAN_IN), .B2(n6941), .A(n7162), .ZN(
        n6942) );
  NAND2_X1 U8230 ( .A1(n6942), .A2(n10580), .ZN(n6943) );
  OAI211_X1 U8231 ( .C1(n6945), .C2(n10561), .A(n6944), .B(n6943), .ZN(
        P2_U3189) );
  OAI21_X1 U8232 ( .B1(n6948), .B2(n6947), .A(n6946), .ZN(n6949) );
  NAND2_X1 U8233 ( .A1(n6949), .A2(n8848), .ZN(n6952) );
  OAI22_X1 U8234 ( .A1(n8878), .A2(n6752), .B1(n10618), .B2(n8884), .ZN(n6950)
         );
  AOI21_X1 U8235 ( .B1(n8876), .B2(n10609), .A(n6950), .ZN(n6951) );
  OAI211_X1 U8236 ( .C1(n6962), .C2(n10619), .A(n6952), .B(n6951), .ZN(
        P2_U3177) );
  OAI21_X1 U8237 ( .B1(n6955), .B2(n6954), .A(n6953), .ZN(n6956) );
  NAND2_X1 U8238 ( .A1(n6956), .A2(n8848), .ZN(n6960) );
  INV_X1 U8239 ( .A(n6134), .ZN(n6957) );
  OAI22_X1 U8240 ( .A1(n8878), .A2(n6957), .B1(n8884), .B2(n10598), .ZN(n6958)
         );
  AOI21_X1 U8241 ( .B1(n8876), .B2(n8905), .A(n6958), .ZN(n6959) );
  OAI211_X1 U8242 ( .C1(n6962), .C2(n6961), .A(n6960), .B(n6959), .ZN(P2_U3162) );
  NAND2_X1 U8243 ( .A1(n6964), .A2(n6963), .ZN(n6966) );
  AND2_X1 U8244 ( .A1(n6966), .A2(n6965), .ZN(n6967) );
  NAND2_X1 U8245 ( .A1(n6967), .A2(n7310), .ZN(n10831) );
  OR2_X1 U8246 ( .A1(n9881), .A2(n10062), .ZN(n9831) );
  INV_X1 U8247 ( .A(n9831), .ZN(n9820) );
  NAND2_X1 U8248 ( .A1(n9820), .A2(n9879), .ZN(n10673) );
  OR2_X1 U8249 ( .A1(n10591), .A2(n7347), .ZN(n6969) );
  NAND2_X1 U8250 ( .A1(n7171), .A2(n6969), .ZN(n6970) );
  OR2_X1 U8251 ( .A1(n9966), .A2(n6972), .ZN(n9723) );
  NAND2_X1 U8252 ( .A1(n9723), .A2(n9893), .ZN(n9669) );
  NAND2_X1 U8253 ( .A1(n6970), .A2(n9669), .ZN(n7126) );
  OAI21_X1 U8254 ( .B1(n6970), .B2(n9669), .A(n7126), .ZN(n7476) );
  INV_X1 U8255 ( .A(n10257), .ZN(n10818) );
  OAI211_X1 U8256 ( .C1(n6971), .C2(n6972), .A(n7135), .B(n10818), .ZN(n7474)
         );
  OAI21_X1 U8257 ( .B1(n6972), .B2(n10820), .A(n7474), .ZN(n6981) );
  NAND2_X1 U8258 ( .A1(n6973), .A2(n8688), .ZN(n10823) );
  OR2_X1 U8259 ( .A1(n10591), .A2(n9889), .ZN(n6975) );
  NAND2_X1 U8260 ( .A1(n7174), .A2(n6975), .ZN(n9725) );
  XNOR2_X1 U8261 ( .A(n9725), .B(n9669), .ZN(n6978) );
  NAND2_X1 U8262 ( .A1(n6607), .A2(n9946), .ZN(n6977) );
  INV_X1 U8263 ( .A(n10062), .ZN(n9882) );
  NAND2_X1 U8264 ( .A1(n9881), .A2(n9882), .ZN(n6976) );
  INV_X1 U8265 ( .A(n10828), .ZN(n10794) );
  OAI222_X1 U8266 ( .A1(n10823), .A2(n6980), .B1(n10825), .B2(n6979), .C1(
        n6978), .C2(n10794), .ZN(n7471) );
  AOI211_X1 U8267 ( .C1(n10811), .C2(n7476), .A(n6981), .B(n7471), .ZN(n10603)
         );
  INV_X1 U8268 ( .A(n6982), .ZN(n6983) );
  NAND2_X1 U8269 ( .A1(n7301), .A2(n6983), .ZN(n6984) );
  OR2_X1 U8270 ( .A1(n6984), .A2(n7303), .ZN(n7121) );
  AND2_X1 U8271 ( .A1(n6985), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7302) );
  NAND2_X1 U8272 ( .A1(n7300), .A2(n7302), .ZN(n6986) );
  NAND2_X1 U8273 ( .A1(n10835), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6987) );
  OAI21_X1 U8274 ( .B1(n10603), .B2(n10835), .A(n6987), .ZN(P1_U3524) );
  INV_X1 U8275 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6988) );
  INV_X1 U8276 ( .A(n8125), .ZN(n7049) );
  INV_X1 U8277 ( .A(n8954), .ZN(n8958) );
  OAI222_X1 U8278 ( .A1(n8472), .A2(n6988), .B1(n4944), .B2(n7049), .C1(
        P2_U3151), .C2(n8958), .ZN(P2_U3279) );
  XNOR2_X1 U8279 ( .A(n8512), .B(n6989), .ZN(n10599) );
  NOR2_X1 U8280 ( .A1(n6746), .A2(n6747), .ZN(n7054) );
  NAND2_X1 U8281 ( .A1(n10626), .A2(n7054), .ZN(n9022) );
  OAI21_X1 U8282 ( .B1(n6992), .B2(n6991), .A(n6990), .ZN(n6993) );
  NAND2_X1 U8283 ( .A1(n6993), .A2(n10611), .ZN(n6995) );
  AOI22_X1 U8284 ( .A1(n10607), .A2(n6134), .B1(n10608), .B2(n8905), .ZN(n6994) );
  OAI211_X1 U8285 ( .C1(n10599), .C2(n7539), .A(n6995), .B(n6994), .ZN(n10601)
         );
  NOR2_X1 U8286 ( .A1(n10626), .A2(n5735), .ZN(n6996) );
  AOI21_X1 U8287 ( .B1(n10601), .B2(n10626), .A(n6996), .ZN(n6999) );
  AOI22_X1 U8288 ( .A1(n9111), .A2(n6997), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9156), .ZN(n6998) );
  OAI211_X1 U8289 ( .C1(n10599), .C2(n9022), .A(n6999), .B(n6998), .ZN(
        P2_U3232) );
  NAND2_X1 U8290 ( .A1(n7001), .A2(n7000), .ZN(n7006) );
  INV_X1 U8291 ( .A(n7002), .ZN(n7004) );
  NAND2_X1 U8292 ( .A1(n7004), .A2(n7003), .ZN(n7005) );
  NAND2_X1 U8293 ( .A1(n7006), .A2(n7005), .ZN(n7195) );
  NAND2_X1 U8294 ( .A1(n9965), .A2(n6806), .ZN(n7014) );
  NAND2_X1 U8295 ( .A1(n7007), .A2(n9988), .ZN(n7010) );
  OR2_X1 U8296 ( .A1(n7185), .A2(n7008), .ZN(n7009) );
  OAI211_X2 U8297 ( .C1(n7228), .C2(n7011), .A(n7010), .B(n7009), .ZN(n7331)
         );
  NAND2_X1 U8298 ( .A1(n7331), .A2(n4947), .ZN(n7013) );
  NAND2_X1 U8299 ( .A1(n7014), .A2(n7013), .ZN(n7015) );
  XNOR2_X1 U8300 ( .A(n7015), .B(n8460), .ZN(n7196) );
  AND2_X1 U8301 ( .A1(n7331), .A2(n6806), .ZN(n7016) );
  AOI21_X1 U8302 ( .B1(n9965), .B2(n8459), .A(n7016), .ZN(n7197) );
  XNOR2_X1 U8303 ( .A(n7196), .B(n7197), .ZN(n7194) );
  XNOR2_X1 U8304 ( .A(n7195), .B(n7194), .ZN(n7031) );
  OAI22_X1 U8305 ( .A1(n9639), .A2(n7176), .B1(n9654), .B2(
        P1_REG3_REG_3__SCAN_IN), .ZN(n7030) );
  INV_X1 U8306 ( .A(n7331), .ZN(n7412) );
  INV_X1 U8307 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7018) );
  OR2_X1 U8308 ( .A1(n9702), .A2(n7018), .ZN(n7024) );
  INV_X1 U8309 ( .A(n7205), .ZN(n7021) );
  INV_X1 U8310 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7409) );
  INV_X1 U8311 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n7019) );
  NAND2_X1 U8312 ( .A1(n7409), .A2(n7019), .ZN(n7020) );
  NAND2_X1 U8313 ( .A1(n7021), .A2(n7020), .ZN(n7342) );
  OR2_X1 U8314 ( .A1(n8324), .A2(n7342), .ZN(n7023) );
  NAND2_X1 U8315 ( .A1(n8305), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7022) );
  OR2_X1 U8316 ( .A1(n8307), .A2(n7025), .ZN(n7026) );
  NAND2_X2 U8317 ( .A1(n4971), .A2(n7026), .ZN(n9964) );
  NAND2_X1 U8318 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9985) );
  INV_X1 U8319 ( .A(n9985), .ZN(n7027) );
  AOI21_X1 U8320 ( .B1(n9582), .B2(n9964), .A(n7027), .ZN(n7028) );
  OAI21_X1 U8321 ( .B1(n9661), .B2(n7412), .A(n7028), .ZN(n7029) );
  AOI211_X1 U8322 ( .C1(n7031), .C2(n9651), .A(n7030), .B(n7029), .ZN(n7032)
         );
  INV_X1 U8323 ( .A(n7032), .ZN(P1_U3218) );
  OAI21_X1 U8324 ( .B1(n7034), .B2(n7036), .A(n7033), .ZN(n10654) );
  INV_X1 U8325 ( .A(n10654), .ZN(n7045) );
  INV_X1 U8326 ( .A(n7036), .ZN(n8487) );
  XNOR2_X1 U8327 ( .A(n7035), .B(n8487), .ZN(n7040) );
  AOI22_X1 U8328 ( .A1(n10607), .A2(n8904), .B1(n10608), .B2(n8903), .ZN(n7039) );
  INV_X1 U8329 ( .A(n7539), .ZN(n7037) );
  NAND2_X1 U8330 ( .A1(n10654), .A2(n7037), .ZN(n7038) );
  OAI211_X1 U8331 ( .C1(n7040), .C2(n9145), .A(n7039), .B(n7038), .ZN(n10652)
         );
  NAND2_X1 U8332 ( .A1(n10652), .A2(n10626), .ZN(n7044) );
  OAI22_X1 U8333 ( .A1(n9159), .A2(n10651), .B1(n7041), .B2(n10620), .ZN(n7042) );
  AOI21_X1 U8334 ( .B1(n9163), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7042), .ZN(
        n7043) );
  OAI211_X1 U8335 ( .C1(n7045), .C2(n9022), .A(n7044), .B(n7043), .ZN(P2_U3228) );
  INV_X1 U8336 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7050) );
  NOR2_X1 U8337 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n7047) );
  OAI21_X1 U8338 ( .B1(n7047), .B2(n10396), .A(n7046), .ZN(n7064) );
  XNOR2_X1 U8339 ( .A(n7064), .B(n7048), .ZN(n10020) );
  INV_X1 U8340 ( .A(n10020), .ZN(n10007) );
  OAI222_X1 U8341 ( .A1(n7050), .A2(n10406), .B1(P1_U3086), .B2(n10007), .C1(
        n10404), .C2(n7049), .ZN(P1_U3339) );
  INV_X1 U8342 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7051) );
  MUX2_X1 U8343 ( .A(n9063), .B(n7051), .S(n8989), .Z(n7052) );
  INV_X1 U8344 ( .A(n7052), .ZN(P2_U3514) );
  XNOR2_X1 U8345 ( .A(n7053), .B(n8529), .ZN(n10637) );
  INV_X1 U8346 ( .A(n7054), .ZN(n7055) );
  NAND2_X1 U8347 ( .A1(n7539), .A2(n7055), .ZN(n10625) );
  INV_X1 U8348 ( .A(n9161), .ZN(n9129) );
  XNOR2_X1 U8349 ( .A(n7056), .B(n8529), .ZN(n7057) );
  AOI222_X1 U8350 ( .A1(n10611), .A2(n7057), .B1(n5079), .B2(n10608), .C1(
        n10609), .C2(n10607), .ZN(n10635) );
  MUX2_X1 U8351 ( .A(n7058), .B(n10635), .S(n10626), .Z(n7063) );
  INV_X1 U8352 ( .A(n7059), .ZN(n7060) );
  AOI22_X1 U8353 ( .A1(n9111), .A2(n7061), .B1(n9156), .B2(n7060), .ZN(n7062)
         );
  OAI211_X1 U8354 ( .C1(n10637), .C2(n9129), .A(n7063), .B(n7062), .ZN(
        P2_U3229) );
  INV_X1 U8355 ( .A(n8210), .ZN(n7107) );
  OAI21_X1 U8356 ( .B1(n7064), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7065) );
  XNOR2_X1 U8357 ( .A(n7065), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10036) );
  AOI22_X1 U8358 ( .A1(n10036), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10399), .ZN(n7066) );
  OAI21_X1 U8359 ( .B1(n7107), .B2(n10404), .A(n7066), .ZN(P1_U3338) );
  INV_X1 U8360 ( .A(n7067), .ZN(n7068) );
  NAND2_X1 U8361 ( .A1(n7068), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7069) );
  XNOR2_X1 U8362 ( .A(n7069), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10040) );
  AOI22_X1 U8363 ( .A1(n10040), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10399), .ZN(n7070) );
  OAI21_X1 U8364 ( .B1(n8214), .B2(n10404), .A(n7070), .ZN(P1_U3337) );
  INV_X1 U8365 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7576) );
  MUX2_X1 U8366 ( .A(n7576), .B(P1_REG1_REG_11__SCAN_IN), .S(n7631), .Z(n7072)
         );
  AOI211_X1 U8367 ( .C1(n7073), .C2(n7072), .A(n7250), .B(n10067), .ZN(n7084)
         );
  NAND2_X1 U8368 ( .A1(n7631), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7075) );
  OAI21_X1 U8369 ( .B1(n7631), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7075), .ZN(
        n7076) );
  NOR2_X1 U8370 ( .A1(n7077), .A2(n7076), .ZN(n7246) );
  AOI211_X1 U8371 ( .C1(n7077), .C2(n7076), .A(n7246), .B(n10037), .ZN(n7083)
         );
  INV_X1 U8372 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7081) );
  NAND2_X1 U8373 ( .A1(n10041), .A2(n7631), .ZN(n7080) );
  INV_X1 U8374 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7078) );
  NOR2_X1 U8375 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7078), .ZN(n8008) );
  INV_X1 U8376 ( .A(n8008), .ZN(n7079) );
  OAI211_X1 U8377 ( .C1(n7081), .C2(n10044), .A(n7080), .B(n7079), .ZN(n7082)
         );
  OR3_X1 U8378 ( .A1(n7084), .A2(n7083), .A3(n7082), .ZN(P1_U3254) );
  XNOR2_X1 U8379 ( .A(n7405), .B(n8744), .ZN(n7317) );
  XOR2_X1 U8380 ( .A(n8902), .B(n7317), .Z(n7090) );
  XNOR2_X1 U8381 ( .A(n10670), .B(n8744), .ZN(n7087) );
  XNOR2_X1 U8382 ( .A(n7087), .B(n8903), .ZN(n8850) );
  AOI21_X1 U8383 ( .B1(n7090), .B2(n7089), .A(n7316), .ZN(n7098) );
  INV_X1 U8384 ( .A(n8878), .ZN(n8834) );
  AOI21_X1 U8385 ( .B1(n8834), .B2(n8903), .A(n7091), .ZN(n7096) );
  NAND2_X1 U8386 ( .A1(n7405), .A2(n8867), .ZN(n7095) );
  INV_X1 U8387 ( .A(n7294), .ZN(n7092) );
  NAND2_X1 U8388 ( .A1(n8880), .A2(n7092), .ZN(n7094) );
  NAND2_X1 U8389 ( .A1(n8876), .A2(n8901), .ZN(n7093) );
  AND4_X1 U8390 ( .A1(n7096), .A2(n7095), .A3(n7094), .A4(n7093), .ZN(n7097)
         );
  OAI21_X1 U8391 ( .B1(n7098), .B2(n8870), .A(n7097), .ZN(P2_U3153) );
  INV_X1 U8392 ( .A(n8532), .ZN(n8563) );
  AND2_X1 U8393 ( .A1(n8550), .A2(n8563), .ZN(n8490) );
  XOR2_X1 U8394 ( .A(n7099), .B(n8490), .Z(n10667) );
  XNOR2_X1 U8395 ( .A(n7100), .B(n8490), .ZN(n7101) );
  OAI222_X1 U8396 ( .A1(n9148), .A2(n8854), .B1(n9150), .B2(n7318), .C1(n9145), 
        .C2(n7101), .ZN(n10668) );
  NAND2_X1 U8397 ( .A1(n10668), .A2(n10626), .ZN(n7105) );
  INV_X1 U8398 ( .A(n10670), .ZN(n7102) );
  OAI22_X1 U8399 ( .A1(n9159), .A2(n7102), .B1(n8856), .B2(n10620), .ZN(n7103)
         );
  AOI21_X1 U8400 ( .B1(n9163), .B2(P2_REG2_REG_6__SCAN_IN), .A(n7103), .ZN(
        n7104) );
  OAI211_X1 U8401 ( .C1(n10667), .C2(n9129), .A(n7105), .B(n7104), .ZN(
        P2_U3227) );
  INV_X1 U8402 ( .A(n8984), .ZN(n8974) );
  INV_X1 U8403 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7106) );
  OAI222_X1 U8404 ( .A1(n4944), .A2(n7107), .B1(n8974), .B2(P2_U3151), .C1(
        n7106), .C2(n8472), .ZN(P2_U3278) );
  XNOR2_X1 U8405 ( .A(n7108), .B(n8486), .ZN(n7109) );
  OAI222_X1 U8406 ( .A1(n9148), .A2(n7111), .B1(n9150), .B2(n7110), .C1(n9145), 
        .C2(n7109), .ZN(n10629) );
  OR2_X1 U8407 ( .A1(n7112), .A2(n8486), .ZN(n7113) );
  NAND2_X1 U8408 ( .A1(n7114), .A2(n7113), .ZN(n10631) );
  NAND2_X1 U8409 ( .A1(n10631), .A2(n9161), .ZN(n7118) );
  NOR2_X1 U8410 ( .A1(n10620), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7115) );
  AOI21_X1 U8411 ( .B1(n9111), .B2(n7116), .A(n7115), .ZN(n7117) );
  OAI211_X1 U8412 ( .C1(n5768), .C2(n10626), .A(n7118), .B(n7117), .ZN(n7119)
         );
  AOI21_X1 U8413 ( .B1(n10629), .B2(n10626), .A(n7119), .ZN(n7120) );
  INV_X1 U8414 ( .A(n7120), .ZN(P2_U3230) );
  INV_X1 U8415 ( .A(n7121), .ZN(n7124) );
  INV_X1 U8416 ( .A(n7302), .ZN(n7122) );
  NOR2_X1 U8417 ( .A1(n7300), .A2(n7122), .ZN(n7123) );
  AND2_X2 U8418 ( .A1(n7124), .A2(n7123), .ZN(n10839) );
  OR2_X1 U8419 ( .A1(n9966), .A2(n7472), .ZN(n7125) );
  NAND2_X1 U8420 ( .A1(n7126), .A2(n7125), .ZN(n7127) );
  NAND2_X1 U8421 ( .A1(n7127), .A2(n7130), .ZN(n7333) );
  OAI21_X1 U8422 ( .B1(n7127), .B2(n7130), .A(n7333), .ZN(n7414) );
  INV_X1 U8423 ( .A(n7414), .ZN(n7137) );
  INV_X1 U8424 ( .A(n10831), .ZN(n10691) );
  INV_X1 U8425 ( .A(n9964), .ZN(n7239) );
  OAI22_X1 U8426 ( .A1(n7239), .A2(n10823), .B1(n7176), .B2(n10825), .ZN(n7133) );
  NAND2_X1 U8427 ( .A1(n9725), .A2(n9893), .ZN(n7128) );
  INV_X1 U8428 ( .A(n9731), .ZN(n7129) );
  NAND2_X1 U8429 ( .A1(n7129), .A2(n7130), .ZN(n7131) );
  INV_X1 U8430 ( .A(n7130), .ZN(n9667) );
  NAND2_X1 U8431 ( .A1(n9731), .A2(n9667), .ZN(n7334) );
  AOI21_X1 U8432 ( .B1(n7131), .B2(n7334), .A(n10794), .ZN(n7132) );
  AOI211_X1 U8433 ( .C1(n10691), .C2(n7414), .A(n7133), .B(n7132), .ZN(n7416)
         );
  INV_X1 U8434 ( .A(n7339), .ZN(n7134) );
  AOI211_X1 U8435 ( .C1(n7331), .C2(n7135), .A(n10257), .B(n7134), .ZN(n7408)
         );
  AOI21_X1 U8436 ( .B1(n10791), .B2(n7331), .A(n7408), .ZN(n7136) );
  OAI211_X1 U8437 ( .C1(n7137), .C2(n10673), .A(n7416), .B(n7136), .ZN(n7139)
         );
  NAND2_X1 U8438 ( .A1(n7139), .A2(n10839), .ZN(n7138) );
  OAI21_X1 U8439 ( .B1(n10839), .B2(n6836), .A(n7138), .ZN(P1_U3462) );
  INV_X2 U8440 ( .A(n10835), .ZN(n10665) );
  INV_X1 U8441 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7141) );
  NAND2_X1 U8442 ( .A1(n7139), .A2(n10665), .ZN(n7140) );
  OAI21_X1 U8443 ( .B1(n10665), .B2(n7141), .A(n7140), .ZN(P1_U3525) );
  AOI22_X1 U8444 ( .A1(n7391), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n7374), .B2(
        n7159), .ZN(n7145) );
  AOI21_X1 U8445 ( .B1(n7146), .B2(n7145), .A(n7376), .ZN(n7169) );
  NOR2_X1 U8446 ( .A1(n7148), .A2(n7147), .ZN(n7152) );
  MUX2_X1 U8447 ( .A(n7374), .B(n7149), .S(n8679), .Z(n7150) );
  NAND2_X1 U8448 ( .A1(n7150), .A2(n7391), .ZN(n7379) );
  OAI21_X1 U8449 ( .B1(n7150), .B2(n7391), .A(n7379), .ZN(n7151) );
  NOR2_X1 U8450 ( .A1(n7152), .A2(n7151), .ZN(n7381) );
  AOI21_X1 U8451 ( .B1(n7152), .B2(n7151), .A(n7381), .ZN(n7155) );
  INV_X1 U8452 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7153) );
  NOR2_X1 U8453 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7153), .ZN(n7322) );
  INV_X1 U8454 ( .A(n7322), .ZN(n7154) );
  OAI21_X1 U8455 ( .B1(n7155), .B2(n10562), .A(n7154), .ZN(n7158) );
  INV_X1 U8456 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7156) );
  NOR2_X1 U8457 ( .A1(n10569), .A2(n7156), .ZN(n7157) );
  AOI211_X1 U8458 ( .C1(n10571), .C2(n7391), .A(n7158), .B(n7157), .ZN(n7168)
         );
  AOI22_X1 U8459 ( .A1(n7391), .A2(n7149), .B1(P2_REG1_REG_8__SCAN_IN), .B2(
        n7159), .ZN(n7165) );
  NAND2_X1 U8460 ( .A1(n7161), .A2(n7160), .ZN(n7163) );
  NAND2_X1 U8461 ( .A1(n7165), .A2(n7164), .ZN(n7390) );
  OAI21_X1 U8462 ( .B1(n7165), .B2(n7164), .A(n7390), .ZN(n7166) );
  NAND2_X1 U8463 ( .A1(n7166), .A2(n10580), .ZN(n7167) );
  OAI211_X1 U8464 ( .C1(n7169), .C2(n10561), .A(n7168), .B(n7167), .ZN(
        P2_U3190) );
  INV_X1 U8465 ( .A(n7170), .ZN(n7173) );
  INV_X1 U8466 ( .A(n7171), .ZN(n7172) );
  AOI21_X1 U8467 ( .B1(n7173), .B2(n5042), .A(n7172), .ZN(n7352) );
  OAI21_X1 U8468 ( .B1(n7175), .B2(n5042), .A(n7174), .ZN(n7180) );
  OAI22_X1 U8469 ( .A1(n7177), .A2(n10825), .B1(n7176), .B2(n10823), .ZN(n7179) );
  NOR2_X1 U8470 ( .A1(n7352), .A2(n10831), .ZN(n7178) );
  AOI211_X1 U8471 ( .C1(n10828), .C2(n7180), .A(n7179), .B(n7178), .ZN(n7357)
         );
  NAND2_X1 U8472 ( .A1(n7347), .A2(n10592), .ZN(n7181) );
  NAND2_X1 U8473 ( .A1(n7181), .A2(n10818), .ZN(n7182) );
  NOR2_X1 U8474 ( .A1(n6971), .A2(n7182), .ZN(n7355) );
  AOI21_X1 U8475 ( .B1(n10791), .B2(n7347), .A(n7355), .ZN(n7183) );
  OAI211_X1 U8476 ( .C1(n7352), .C2(n10673), .A(n7357), .B(n7183), .ZN(n10377)
         );
  NAND2_X1 U8477 ( .A1(n10377), .A2(n10839), .ZN(n7184) );
  OAI21_X1 U8478 ( .B1(n10839), .B2(n6735), .A(n7184), .ZN(P1_U3456) );
  INV_X4 U8479 ( .A(n7228), .ZN(n9697) );
  NAND2_X1 U8480 ( .A1(n7264), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7188) );
  NAND2_X1 U8481 ( .A1(n7007), .A2(n7186), .ZN(n7187) );
  OAI211_X2 U8482 ( .C1(n8301), .C2(n7189), .A(n7188), .B(n7187), .ZN(n10641)
         );
  NAND2_X1 U8483 ( .A1(n10641), .A2(n4947), .ZN(n7190) );
  NAND2_X1 U8484 ( .A1(n7191), .A2(n7190), .ZN(n7192) );
  AND2_X1 U8485 ( .A1(n10641), .A2(n6806), .ZN(n7193) );
  AOI21_X1 U8486 ( .B1(n9964), .B2(n8459), .A(n7193), .ZN(n7218) );
  XNOR2_X1 U8487 ( .A(n7217), .B(n7218), .ZN(n7203) );
  INV_X1 U8488 ( .A(n7196), .ZN(n7198) );
  NAND2_X1 U8489 ( .A1(n7198), .A2(n7197), .ZN(n7199) );
  INV_X1 U8490 ( .A(n7203), .ZN(n7200) );
  INV_X1 U8491 ( .A(n7222), .ZN(n7201) );
  AOI211_X1 U8492 ( .C1(n7203), .C2(n7202), .A(n9632), .B(n7201), .ZN(n7215)
         );
  NAND2_X1 U8493 ( .A1(n7274), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7210) );
  INV_X1 U8494 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7493) );
  OR2_X1 U8495 ( .A1(n9705), .A2(n7493), .ZN(n7209) );
  OAI21_X1 U8496 ( .B1(n7205), .B2(P1_REG3_REG_5__SCAN_IN), .A(n7204), .ZN(
        n7492) );
  OR2_X1 U8497 ( .A1(n8324), .A2(n7492), .ZN(n7208) );
  INV_X1 U8498 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7206) );
  OR2_X1 U8499 ( .A1(n9702), .A2(n7206), .ZN(n7207) );
  INV_X1 U8500 ( .A(n9963), .ZN(n10681) );
  OAI22_X1 U8501 ( .A1(n9655), .A2(n10681), .B1(n9654), .B2(n7342), .ZN(n7214)
         );
  INV_X1 U8502 ( .A(n10641), .ZN(n7343) );
  INV_X1 U8503 ( .A(n9639), .ZN(n9658) );
  NAND2_X1 U8504 ( .A1(n9658), .A2(n9965), .ZN(n7211) );
  OAI211_X1 U8505 ( .C1(n9661), .C2(n7343), .A(n7212), .B(n7211), .ZN(n7213)
         );
  OR3_X1 U8506 ( .A1(n7215), .A2(n7214), .A3(n7213), .ZN(P1_U3230) );
  INV_X1 U8507 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7216) );
  INV_X1 U8508 ( .A(n8997), .ZN(n9006) );
  OAI222_X1 U8509 ( .A1(n8472), .A2(n7216), .B1(n9006), .B2(P2_U3151), .C1(
        n4944), .C2(n8214), .ZN(P2_U3277) );
  INV_X1 U8510 ( .A(n7217), .ZN(n7220) );
  INV_X1 U8511 ( .A(n7218), .ZN(n7219) );
  NAND2_X1 U8512 ( .A1(n7220), .A2(n7219), .ZN(n7221) );
  NAND2_X1 U8513 ( .A1(n7222), .A2(n7221), .ZN(n7235) );
  INV_X1 U8514 ( .A(n7235), .ZN(n7233) );
  NAND2_X1 U8515 ( .A1(n9963), .A2(n8438), .ZN(n7230) );
  NAND2_X1 U8516 ( .A1(n7007), .A2(n7223), .ZN(n7226) );
  OR2_X1 U8517 ( .A1(n8301), .A2(n7224), .ZN(n7225) );
  OAI211_X1 U8518 ( .C1(n7228), .C2(n7227), .A(n7226), .B(n7225), .ZN(n7502)
         );
  NAND2_X1 U8519 ( .A1(n7502), .A2(n4947), .ZN(n7229) );
  NAND2_X1 U8520 ( .A1(n7230), .A2(n7229), .ZN(n7231) );
  XNOR2_X1 U8521 ( .A(n7231), .B(n8460), .ZN(n7234) );
  INV_X1 U8522 ( .A(n7234), .ZN(n7232) );
  NAND2_X1 U8523 ( .A1(n7233), .A2(n7232), .ZN(n7261) );
  NAND2_X1 U8524 ( .A1(n7235), .A2(n7234), .ZN(n7260) );
  NAND2_X1 U8525 ( .A1(n7261), .A2(n7260), .ZN(n7237) );
  AND2_X1 U8526 ( .A1(n7502), .A2(n6806), .ZN(n7236) );
  AOI21_X1 U8527 ( .B1(n9963), .B2(n8459), .A(n7236), .ZN(n7259) );
  XNOR2_X1 U8528 ( .A(n7237), .B(n7259), .ZN(n7244) );
  OAI21_X1 U8529 ( .B1(n9639), .B2(n7239), .A(n7238), .ZN(n7242) );
  INV_X1 U8530 ( .A(n8200), .ZN(n7240) );
  OAI22_X1 U8531 ( .A1(n9655), .A2(n7240), .B1(n9654), .B2(n7492), .ZN(n7241)
         );
  AOI211_X1 U8532 ( .C1(n7502), .C2(n9642), .A(n7242), .B(n7241), .ZN(n7243)
         );
  OAI21_X1 U8533 ( .B1(n7244), .B2(n9632), .A(n7243), .ZN(P1_U3227) );
  NOR2_X1 U8534 ( .A1(n7677), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7245) );
  AOI21_X1 U8535 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7677), .A(n7245), .ZN(
        n7248) );
  AOI21_X1 U8536 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7631), .A(n7246), .ZN(
        n7247) );
  NAND2_X1 U8537 ( .A1(n7248), .A2(n7247), .ZN(n7428) );
  OAI21_X1 U8538 ( .B1(n7248), .B2(n7247), .A(n7428), .ZN(n7249) );
  INV_X1 U8539 ( .A(n7249), .ZN(n7258) );
  INV_X1 U8540 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10804) );
  AOI22_X1 U8541 ( .A1(n7677), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n10804), .B2(
        n7254), .ZN(n7252) );
  OAI21_X1 U8542 ( .B1(n7252), .B2(n7251), .A(n7432), .ZN(n7256) );
  AND2_X1 U8543 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8094) );
  AOI21_X1 U8544 ( .B1(n10059), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n8094), .ZN(
        n7253) );
  OAI21_X1 U8545 ( .B1(n10063), .B2(n7254), .A(n7253), .ZN(n7255) );
  AOI21_X1 U8546 ( .B1(n7256), .B2(n10024), .A(n7255), .ZN(n7257) );
  OAI21_X1 U8547 ( .B1(n7258), .B2(n10037), .A(n7257), .ZN(P1_U3255) );
  NAND2_X1 U8548 ( .A1(n7260), .A2(n7259), .ZN(n7262) );
  NAND2_X1 U8549 ( .A1(n7262), .A2(n7261), .ZN(n7750) );
  NAND2_X1 U8550 ( .A1(n8200), .A2(n6806), .ZN(n7269) );
  NAND2_X1 U8551 ( .A1(n9697), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7266) );
  NAND2_X1 U8552 ( .A1(n10698), .A2(n4947), .ZN(n7268) );
  NAND2_X1 U8553 ( .A1(n7269), .A2(n7268), .ZN(n7270) );
  XNOR2_X1 U8554 ( .A(n7270), .B(n6829), .ZN(n7272) );
  AOI22_X1 U8555 ( .A1(n8200), .A2(n8459), .B1(n6806), .B2(n10698), .ZN(n7271)
         );
  OR2_X1 U8556 ( .A1(n7272), .A2(n7271), .ZN(n7749) );
  NAND2_X1 U8557 ( .A1(n5039), .A2(n7749), .ZN(n7273) );
  XNOR2_X1 U8558 ( .A(n7750), .B(n7273), .ZN(n7288) );
  NOR2_X1 U8559 ( .A1(n9654), .A2(n10695), .ZN(n7286) );
  NAND2_X1 U8560 ( .A1(n7274), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7281) );
  INV_X1 U8561 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7275) );
  OR2_X1 U8562 ( .A1(n9702), .A2(n7275), .ZN(n7280) );
  OR2_X1 U8563 ( .A1(n7276), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7277) );
  NAND2_X1 U8564 ( .A1(n7518), .A2(n7277), .ZN(n8198) );
  OR2_X1 U8565 ( .A1(n8324), .A2(n8198), .ZN(n7279) );
  INV_X1 U8566 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7529) );
  OR2_X1 U8567 ( .A1(n9705), .A2(n7529), .ZN(n7278) );
  NAND4_X1 U8568 ( .A1(n7281), .A2(n7280), .A3(n7279), .A4(n7278), .ZN(n9962)
         );
  INV_X1 U8569 ( .A(n7282), .ZN(n7283) );
  AOI21_X1 U8570 ( .B1(n9582), .B2(n9962), .A(n7283), .ZN(n7284) );
  OAI21_X1 U8571 ( .B1(n9661), .B2(n10680), .A(n7284), .ZN(n7285) );
  AOI211_X1 U8572 ( .C1(n9658), .C2(n9963), .A(n7286), .B(n7285), .ZN(n7287)
         );
  OAI21_X1 U8573 ( .B1(n7288), .B2(n9632), .A(n7287), .ZN(P1_U3239) );
  OAI21_X1 U8574 ( .B1(n7290), .B2(n8552), .A(n7289), .ZN(n7291) );
  AOI222_X1 U8575 ( .A1(n10611), .A2(n7291), .B1(n8901), .B2(n10608), .C1(
        n8903), .C2(n10607), .ZN(n7400) );
  OR2_X1 U8576 ( .A1(n7292), .A2(n8551), .ZN(n7398) );
  NAND3_X1 U8577 ( .A1(n7398), .A2(n7397), .A3(n9161), .ZN(n7297) );
  NOR2_X1 U8578 ( .A1(n10620), .A2(n7294), .ZN(n7295) );
  AOI21_X1 U8579 ( .B1(n9111), .B2(n7405), .A(n7295), .ZN(n7296) );
  OAI211_X1 U8580 ( .C1(n5839), .C2(n10626), .A(n7297), .B(n7296), .ZN(n7298)
         );
  INV_X1 U8581 ( .A(n7298), .ZN(n7299) );
  OAI21_X1 U8582 ( .B1(n7400), .B2(n9163), .A(n7299), .ZN(P2_U3226) );
  INV_X1 U8583 ( .A(n7300), .ZN(n7304) );
  NAND4_X1 U8584 ( .A1(n7304), .A2(n7303), .A3(n7302), .A4(n7301), .ZN(n7305)
         );
  NAND2_X2 U8585 ( .A1(n7305), .A2(n10847), .ZN(n10852) );
  INV_X1 U8586 ( .A(n7306), .ZN(n7307) );
  NOR2_X2 U8587 ( .A1(n10731), .A2(n7307), .ZN(n10732) );
  AOI21_X1 U8588 ( .B1(n4942), .B2(n10593), .A(n10732), .ZN(n7315) );
  INV_X1 U8589 ( .A(n10823), .ZN(n10590) );
  NAND2_X1 U8590 ( .A1(n10852), .A2(n10590), .ZN(n10193) );
  INV_X1 U8591 ( .A(n10193), .ZN(n7585) );
  INV_X1 U8592 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7308) );
  OAI22_X1 U8593 ( .A1(n10852), .A2(n7309), .B1(n7308), .B2(n10847), .ZN(n7313) );
  INV_X1 U8594 ( .A(n10852), .ZN(n10697) );
  XNOR2_X1 U8595 ( .A(n9968), .B(n10592), .ZN(n10589) );
  INV_X1 U8596 ( .A(n7310), .ZN(n7311) );
  NOR4_X1 U8597 ( .A1(n10697), .A2(n10589), .A3(n7311), .A4(n10593), .ZN(n7312) );
  AOI211_X1 U8598 ( .C1(n7585), .C2(n10591), .A(n7313), .B(n7312), .ZN(n7314)
         );
  OAI21_X1 U8599 ( .B1(n7315), .B2(n9890), .A(n7314), .ZN(P1_U3293) );
  XNOR2_X1 U8600 ( .A(n10743), .B(n8739), .ZN(n7319) );
  AND2_X1 U8601 ( .A1(n7319), .A2(n8901), .ZN(n7610) );
  INV_X1 U8602 ( .A(n7319), .ZN(n7320) );
  NAND2_X1 U8603 ( .A1(n7320), .A2(n7605), .ZN(n7611) );
  NAND2_X1 U8604 ( .A1(n5546), .A2(n7611), .ZN(n7321) );
  XNOR2_X1 U8605 ( .A(n7612), .B(n7321), .ZN(n7329) );
  NAND2_X1 U8606 ( .A1(n10743), .A2(n8867), .ZN(n7327) );
  AOI21_X1 U8607 ( .B1(n8834), .B2(n8902), .A(n7322), .ZN(n7326) );
  INV_X1 U8608 ( .A(n7367), .ZN(n7323) );
  NAND2_X1 U8609 ( .A1(n8880), .A2(n7323), .ZN(n7325) );
  NAND2_X1 U8610 ( .A1(n8876), .A2(n8900), .ZN(n7324) );
  NAND4_X1 U8611 ( .A1(n7327), .A2(n7326), .A3(n7325), .A4(n7324), .ZN(n7328)
         );
  AOI21_X1 U8612 ( .B1(n7329), .B2(n8848), .A(n7328), .ZN(n7330) );
  INV_X1 U8613 ( .A(n7330), .ZN(P2_U3161) );
  OR2_X1 U8614 ( .A1(n9965), .A2(n7331), .ZN(n7332) );
  NAND2_X1 U8615 ( .A1(n7333), .A2(n7332), .ZN(n7481) );
  NAND2_X1 U8616 ( .A1(n9964), .A2(n7343), .ZN(n9734) );
  AND2_X2 U8617 ( .A1(n9899), .A2(n9734), .ZN(n9732) );
  XNOR2_X1 U8618 ( .A(n7481), .B(n9732), .ZN(n10645) );
  AOI21_X2 U8619 ( .B1(n10831), .B2(n7350), .A(n10731), .ZN(n10190) );
  NAND2_X1 U8620 ( .A1(n7334), .A2(n9729), .ZN(n7335) );
  OAI21_X1 U8621 ( .B1(n9732), .B2(n7335), .A(n7485), .ZN(n7336) );
  NAND2_X1 U8622 ( .A1(n7336), .A2(n10828), .ZN(n7338) );
  INV_X1 U8623 ( .A(n10825), .ZN(n10747) );
  AOI22_X1 U8624 ( .A1(n10747), .A2(n9965), .B1(n9963), .B2(n10590), .ZN(n7337) );
  AND2_X1 U8625 ( .A1(n7338), .A2(n7337), .ZN(n10648) );
  MUX2_X1 U8626 ( .A(n6492), .B(n10648), .S(n10852), .Z(n7346) );
  NAND2_X1 U8627 ( .A1(n7339), .A2(n10641), .ZN(n7340) );
  NAND2_X1 U8628 ( .A1(n7340), .A2(n10818), .ZN(n7341) );
  NOR2_X1 U8629 ( .A1(n7490), .A2(n7341), .ZN(n10643) );
  OAI22_X1 U8630 ( .A1(n10845), .A2(n7343), .B1(n10847), .B2(n7342), .ZN(n7344) );
  AOI21_X1 U8631 ( .B1(n4942), .B2(n10643), .A(n7344), .ZN(n7345) );
  OAI211_X1 U8632 ( .C1(n10645), .C2(n10265), .A(n7346), .B(n7345), .ZN(
        P1_U3289) );
  NAND2_X1 U8633 ( .A1(n10732), .A2(n7347), .ZN(n7349) );
  INV_X1 U8634 ( .A(n10847), .ZN(n10730) );
  AOI22_X1 U8635 ( .A1(n10731), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n10730), .ZN(n7348) );
  NAND2_X1 U8636 ( .A1(n7349), .A2(n7348), .ZN(n7354) );
  NOR2_X1 U8637 ( .A1(n10731), .A2(n7350), .ZN(n10843) );
  INV_X1 U8638 ( .A(n10843), .ZN(n7351) );
  NOR2_X1 U8639 ( .A1(n7352), .A2(n7351), .ZN(n7353) );
  AOI211_X1 U8640 ( .C1(n7355), .C2(n4942), .A(n7354), .B(n7353), .ZN(n7356)
         );
  OAI21_X1 U8641 ( .B1(n7357), .B2(n10697), .A(n7356), .ZN(P1_U3292) );
  NAND2_X1 U8642 ( .A1(n7397), .A2(n7358), .ZN(n7359) );
  XOR2_X1 U8643 ( .A(n8491), .B(n7359), .Z(n10740) );
  INV_X1 U8644 ( .A(n8491), .ZN(n7362) );
  NAND3_X1 U8645 ( .A1(n7289), .A2(n7362), .A3(n7361), .ZN(n7363) );
  NAND2_X1 U8646 ( .A1(n7360), .A2(n7363), .ZN(n7364) );
  NAND2_X1 U8647 ( .A1(n7364), .A2(n10611), .ZN(n7366) );
  AOI22_X1 U8648 ( .A1(n10607), .A2(n8902), .B1(n10608), .B2(n8900), .ZN(n7365) );
  NAND2_X1 U8649 ( .A1(n7366), .A2(n7365), .ZN(n10741) );
  NAND2_X1 U8650 ( .A1(n10741), .A2(n10626), .ZN(n7370) );
  OAI22_X1 U8651 ( .A1(n10626), .A2(n7374), .B1(n7367), .B2(n10620), .ZN(n7368) );
  AOI21_X1 U8652 ( .B1(n9111), .B2(n10743), .A(n7368), .ZN(n7369) );
  OAI211_X1 U8653 ( .C1(n10740), .C2(n9129), .A(n7370), .B(n7369), .ZN(
        P2_U3225) );
  INV_X1 U8654 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7371) );
  INV_X1 U8655 ( .A(n8230), .ZN(n7372) );
  OAI222_X1 U8656 ( .A1(n8472), .A2(n7371), .B1(n4944), .B2(n7372), .C1(n8677), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  INV_X1 U8657 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7373) );
  OAI222_X1 U8658 ( .A1(n10406), .A2(n7373), .B1(n10404), .B2(n7372), .C1(
        P1_U3086), .C2(n10062), .ZN(P1_U3336) );
  NOR2_X1 U8659 ( .A1(n7391), .A2(n7374), .ZN(n7375) );
  AOI21_X1 U8660 ( .B1(n7377), .B2(n7383), .A(n7444), .ZN(n7396) );
  INV_X1 U8661 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7378) );
  NOR2_X1 U8662 ( .A1(n10569), .A2(n7378), .ZN(n7389) );
  INV_X1 U8663 ( .A(n7379), .ZN(n7380) );
  NOR2_X1 U8664 ( .A1(n7381), .A2(n7380), .ZN(n7385) );
  MUX2_X1 U8665 ( .A(n7383), .B(n7382), .S(n8679), .Z(n7455) );
  XNOR2_X1 U8666 ( .A(n7455), .B(n7456), .ZN(n7384) );
  AOI21_X1 U8667 ( .B1(n7385), .B2(n7384), .A(n7454), .ZN(n7387) );
  NOR2_X1 U8668 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5682), .ZN(n7607) );
  INV_X1 U8669 ( .A(n7607), .ZN(n7386) );
  OAI21_X1 U8670 ( .B1(n7387), .B2(n10562), .A(n7386), .ZN(n7388) );
  AOI211_X1 U8671 ( .C1(n10571), .C2(n7456), .A(n7389), .B(n7388), .ZN(n7395)
         );
  XNOR2_X1 U8672 ( .A(n7448), .B(n7456), .ZN(n7392) );
  NAND2_X1 U8673 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(n7392), .ZN(n7449) );
  OAI21_X1 U8674 ( .B1(n7392), .B2(P2_REG1_REG_9__SCAN_IN), .A(n7449), .ZN(
        n7393) );
  NAND2_X1 U8675 ( .A1(n7393), .A2(n10580), .ZN(n7394) );
  OAI211_X1 U8676 ( .C1(n7396), .C2(n10561), .A(n7395), .B(n7394), .ZN(
        P2_U3191) );
  INV_X1 U8677 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7403) );
  NAND3_X1 U8678 ( .A1(n7398), .A2(n7397), .A3(n10632), .ZN(n7399) );
  NAND2_X1 U8679 ( .A1(n7400), .A2(n7399), .ZN(n7404) );
  NAND2_X1 U8680 ( .A1(n7404), .A2(n10785), .ZN(n7402) );
  INV_X1 U8681 ( .A(n9252), .ZN(n9237) );
  NAND2_X1 U8682 ( .A1(n9237), .A2(n7405), .ZN(n7401) );
  OAI211_X1 U8683 ( .C1(n7403), .C2(n10785), .A(n7402), .B(n7401), .ZN(
        P2_U3411) );
  NAND2_X1 U8684 ( .A1(n7404), .A2(n10781), .ZN(n7407) );
  NAND2_X1 U8685 ( .A1(n6290), .A2(n7405), .ZN(n7406) );
  OAI211_X1 U8686 ( .C1(n10781), .C2(n5836), .A(n7407), .B(n7406), .ZN(
        P2_U3466) );
  NAND2_X1 U8687 ( .A1(n7408), .A2(n4942), .ZN(n7411) );
  AOI22_X1 U8688 ( .A1(n10697), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10730), .B2(
        n7409), .ZN(n7410) );
  OAI211_X1 U8689 ( .C1(n7412), .C2(n10845), .A(n7411), .B(n7410), .ZN(n7413)
         );
  AOI21_X1 U8690 ( .B1(n10843), .B2(n7414), .A(n7413), .ZN(n7415) );
  OAI21_X1 U8691 ( .B1(n7416), .B2(n10697), .A(n7415), .ZN(P1_U3290) );
  NAND3_X1 U8692 ( .A1(n7360), .A2(n5467), .A3(n7417), .ZN(n7418) );
  NAND2_X1 U8693 ( .A1(n7419), .A2(n7418), .ZN(n7420) );
  AOI222_X1 U8694 ( .A1(n10611), .A2(n7420), .B1(n8901), .B2(n10607), .C1(
        n8899), .C2(n10608), .ZN(n7621) );
  INV_X1 U8695 ( .A(n10626), .ZN(n9163) );
  OAI22_X1 U8696 ( .A1(n10626), .A2(n7383), .B1(n7609), .B2(n10620), .ZN(n7421) );
  AOI21_X1 U8697 ( .B1(n7626), .B2(n9111), .A(n7421), .ZN(n7424) );
  NAND2_X1 U8698 ( .A1(n7422), .A2(n8493), .ZN(n7618) );
  NAND3_X1 U8699 ( .A1(n7619), .A2(n9161), .A3(n7618), .ZN(n7423) );
  OAI211_X1 U8700 ( .C1(n7621), .C2(n9163), .A(n7424), .B(n7423), .ZN(P2_U3224) );
  INV_X1 U8701 ( .A(n8241), .ZN(n7427) );
  NAND2_X1 U8702 ( .A1(n10399), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7425) );
  OAI211_X1 U8703 ( .C1(n7427), .C2(n10404), .A(n7426), .B(n7425), .ZN(
        P1_U3335) );
  OAI222_X1 U8704 ( .A1(n4944), .A2(n7427), .B1(n8472), .B2(n6031), .C1(n8675), 
        .C2(P2_U3151), .ZN(P2_U3275) );
  OAI21_X1 U8705 ( .B1(n7677), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7428), .ZN(
        n7431) );
  NAND2_X1 U8706 ( .A1(n7795), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7429) );
  OAI21_X1 U8707 ( .B1(n7795), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7429), .ZN(
        n7430) );
  NOR2_X1 U8708 ( .A1(n7431), .A2(n7430), .ZN(n7658) );
  AOI211_X1 U8709 ( .C1(n7431), .C2(n7430), .A(n7658), .B(n10037), .ZN(n7442)
         );
  OAI21_X1 U8710 ( .B1(n7677), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7432), .ZN(
        n7435) );
  INV_X1 U8711 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7433) );
  MUX2_X1 U8712 ( .A(n7433), .B(P1_REG1_REG_13__SCAN_IN), .S(n7795), .Z(n7434)
         );
  NOR2_X1 U8713 ( .A1(n7434), .A2(n7435), .ZN(n7654) );
  AOI211_X1 U8714 ( .C1(n7435), .C2(n7434), .A(n7654), .B(n10067), .ZN(n7441)
         );
  INV_X1 U8715 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7439) );
  NAND2_X1 U8716 ( .A1(n10041), .A2(n7795), .ZN(n7438) );
  NOR2_X1 U8717 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7436), .ZN(n8120) );
  INV_X1 U8718 ( .A(n8120), .ZN(n7437) );
  OAI211_X1 U8719 ( .C1(n7439), .C2(n10044), .A(n7438), .B(n7437), .ZN(n7440)
         );
  OR3_X1 U8720 ( .A1(n7442), .A2(n7441), .A3(n7440), .ZN(P1_U3256) );
  INV_X1 U8721 ( .A(n7443), .ZN(n7445) );
  AOI22_X1 U8722 ( .A1(n7715), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7708), .B2(
        n7453), .ZN(n7446) );
  AOI21_X1 U8723 ( .B1(n5033), .B2(n7446), .A(n7709), .ZN(n7470) );
  AOI22_X1 U8724 ( .A1(n7715), .A2(n7457), .B1(P2_REG1_REG_10__SCAN_IN), .B2(
        n7453), .ZN(n7452) );
  NAND2_X1 U8725 ( .A1(n7448), .A2(n7447), .ZN(n7450) );
  NAND2_X1 U8726 ( .A1(n7450), .A2(n7449), .ZN(n7451) );
  NAND2_X1 U8727 ( .A1(n7452), .A2(n7451), .ZN(n7714) );
  OAI21_X1 U8728 ( .B1(n7452), .B2(n7451), .A(n7714), .ZN(n7468) );
  NOR2_X1 U8729 ( .A1(n10504), .A2(n7453), .ZN(n7467) );
  INV_X1 U8730 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7465) );
  MUX2_X1 U8731 ( .A(n7708), .B(n7457), .S(n8679), .Z(n7458) );
  NOR2_X1 U8732 ( .A1(n7458), .A2(n7715), .ZN(n7721) );
  NAND2_X1 U8733 ( .A1(n7458), .A2(n7715), .ZN(n7722) );
  INV_X1 U8734 ( .A(n7722), .ZN(n7459) );
  NOR2_X1 U8735 ( .A1(n7721), .A2(n7459), .ZN(n7461) );
  INV_X1 U8736 ( .A(n10562), .ZN(n10579) );
  NAND2_X1 U8737 ( .A1(n7723), .A2(n7461), .ZN(n7460) );
  OAI211_X1 U8738 ( .C1(n7723), .C2(n7461), .A(n10579), .B(n7460), .ZN(n7464)
         );
  INV_X1 U8739 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7462) );
  NOR2_X1 U8740 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7462), .ZN(n7702) );
  INV_X1 U8741 ( .A(n7702), .ZN(n7463) );
  OAI211_X1 U8742 ( .C1(n7465), .C2(n10569), .A(n7464), .B(n7463), .ZN(n7466)
         );
  AOI211_X1 U8743 ( .C1(n7468), .C2(n10580), .A(n7467), .B(n7466), .ZN(n7469)
         );
  OAI21_X1 U8744 ( .B1(n7470), .B2(n10561), .A(n7469), .ZN(P2_U3192) );
  AOI21_X1 U8745 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n10730), .A(n7471), .ZN(
        n7478) );
  INV_X1 U8746 ( .A(n4942), .ZN(n10180) );
  AOI22_X1 U8747 ( .A1(n10732), .A2(n7472), .B1(P1_REG2_REG_2__SCAN_IN), .B2(
        n10697), .ZN(n7473) );
  OAI21_X1 U8748 ( .B1(n10180), .B2(n7474), .A(n7473), .ZN(n7475) );
  AOI21_X1 U8749 ( .B1(n10190), .B2(n7476), .A(n7475), .ZN(n7477) );
  OAI21_X1 U8750 ( .B1(n7478), .B2(n10697), .A(n7477), .ZN(P1_U3291) );
  INV_X1 U8751 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7479) );
  OAI222_X1 U8752 ( .A1(n10406), .A2(n7479), .B1(n10404), .B2(n8244), .C1(
        n9830), .C2(P1_U3086), .ZN(P1_U3334) );
  NAND2_X1 U8753 ( .A1(n9964), .A2(n10641), .ZN(n7480) );
  NAND2_X1 U8754 ( .A1(n7481), .A2(n7480), .ZN(n7483) );
  OR2_X1 U8755 ( .A1(n9964), .A2(n10641), .ZN(n7482) );
  NAND2_X1 U8756 ( .A1(n7483), .A2(n7482), .ZN(n7501) );
  NAND2_X1 U8757 ( .A1(n9963), .A2(n10660), .ZN(n9739) );
  XNOR2_X1 U8758 ( .A(n7501), .B(n10674), .ZN(n10658) );
  INV_X1 U8759 ( .A(n10658), .ZN(n7498) );
  NAND2_X1 U8760 ( .A1(n7485), .A2(n9899), .ZN(n7484) );
  INV_X1 U8761 ( .A(n10674), .ZN(n9668) );
  NAND3_X1 U8762 ( .A1(n7485), .A2(n10674), .A3(n9899), .ZN(n7486) );
  NAND2_X1 U8763 ( .A1(n10685), .A2(n7486), .ZN(n7487) );
  NAND2_X1 U8764 ( .A1(n7487), .A2(n10828), .ZN(n7489) );
  AOI22_X1 U8765 ( .A1(n10747), .A2(n9964), .B1(n8200), .B2(n10590), .ZN(n7488) );
  NAND2_X1 U8766 ( .A1(n7489), .A2(n7488), .ZN(n10662) );
  OAI21_X1 U8767 ( .B1(n7490), .B2(n10660), .A(n10818), .ZN(n7491) );
  OR2_X1 U8768 ( .A1(n7491), .A2(n10679), .ZN(n10659) );
  OAI22_X1 U8769 ( .A1(n10852), .A2(n7493), .B1(n7492), .B2(n10847), .ZN(n7494) );
  AOI21_X1 U8770 ( .B1(n10732), .B2(n7502), .A(n7494), .ZN(n7495) );
  OAI21_X1 U8771 ( .B1(n10180), .B2(n10659), .A(n7495), .ZN(n7496) );
  AOI21_X1 U8772 ( .B1(n10662), .B2(n10852), .A(n7496), .ZN(n7497) );
  OAI21_X1 U8773 ( .B1(n7498), .B2(n10265), .A(n7497), .ZN(P1_U3288) );
  OR2_X1 U8774 ( .A1(n8200), .A2(n10698), .ZN(n7503) );
  NAND2_X1 U8775 ( .A1(n7501), .A2(n7500), .ZN(n7506) );
  OR2_X1 U8776 ( .A1(n9963), .A2(n7502), .ZN(n10675) );
  OR2_X1 U8777 ( .A1(n7507), .A2(n8301), .ZN(n7510) );
  AOI22_X1 U8778 ( .A1(n9697), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7007), .B2(
        n7508), .ZN(n7509) );
  OR2_X1 U8779 ( .A1(n10720), .A2(n8204), .ZN(n9749) );
  NAND2_X1 U8780 ( .A1(n9749), .A2(n10716), .ZN(n7574) );
  XNOR2_X1 U8781 ( .A(n7575), .B(n7574), .ZN(n10707) );
  NAND2_X1 U8782 ( .A1(n9746), .A2(n10684), .ZN(n9902) );
  INV_X1 U8783 ( .A(n9902), .ZN(n7511) );
  NAND2_X1 U8784 ( .A1(n5043), .A2(n10687), .ZN(n7512) );
  NAND2_X1 U8785 ( .A1(n7512), .A2(n7574), .ZN(n7514) );
  NOR2_X1 U8786 ( .A1(n7574), .A2(n9747), .ZN(n7513) );
  NAND2_X1 U8787 ( .A1(n5043), .A2(n7513), .ZN(n10717) );
  NAND2_X1 U8788 ( .A1(n7514), .A2(n10717), .ZN(n7515) );
  NAND2_X1 U8789 ( .A1(n7515), .A2(n10828), .ZN(n7526) );
  NAND2_X1 U8790 ( .A1(n9700), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7524) );
  OR2_X1 U8791 ( .A1(n9705), .A2(n7516), .ZN(n7523) );
  NAND2_X1 U8792 ( .A1(n7518), .A2(n7517), .ZN(n7519) );
  NAND2_X1 U8793 ( .A1(n7548), .A2(n7519), .ZN(n10728) );
  OR2_X1 U8794 ( .A1(n8324), .A2(n10728), .ZN(n7522) );
  INV_X1 U8795 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7520) );
  OR2_X1 U8796 ( .A1(n9702), .A2(n7520), .ZN(n7521) );
  AOI22_X1 U8797 ( .A1(n10747), .A2(n8200), .B1(n10746), .B2(n10590), .ZN(
        n7525) );
  NAND2_X1 U8798 ( .A1(n7526), .A2(n7525), .ZN(n7527) );
  AOI21_X1 U8799 ( .B1(n10707), .B2(n10691), .A(n7527), .ZN(n10709) );
  AOI21_X1 U8800 ( .B1(n10678), .B2(n8204), .A(n10257), .ZN(n7528) );
  NAND2_X1 U8801 ( .A1(n7528), .A2(n10713), .ZN(n10705) );
  OAI22_X1 U8802 ( .A1(n10852), .A2(n7529), .B1(n8198), .B2(n10847), .ZN(n7530) );
  AOI21_X1 U8803 ( .B1(n10732), .B2(n8204), .A(n7530), .ZN(n7531) );
  OAI21_X1 U8804 ( .B1(n10705), .B2(n10180), .A(n7531), .ZN(n7532) );
  AOI21_X1 U8805 ( .B1(n10707), .B2(n10843), .A(n7532), .ZN(n7533) );
  OAI21_X1 U8806 ( .B1(n10709), .B2(n10697), .A(n7533), .ZN(P1_U3286) );
  XNOR2_X1 U8807 ( .A(n10771), .B(n7828), .ZN(n8495) );
  NAND2_X1 U8808 ( .A1(n7619), .A2(n8548), .ZN(n7534) );
  XOR2_X1 U8809 ( .A(n8495), .B(n7534), .Z(n10768) );
  XNOR2_X1 U8810 ( .A(n7535), .B(n8495), .ZN(n7536) );
  NAND2_X1 U8811 ( .A1(n7536), .A2(n10611), .ZN(n7538) );
  AOI22_X1 U8812 ( .A1(n10607), .A2(n8900), .B1(n10608), .B2(n7889), .ZN(n7537) );
  OAI211_X1 U8813 ( .C1(n10768), .C2(n7539), .A(n7538), .B(n7537), .ZN(n10769)
         );
  NAND2_X1 U8814 ( .A1(n10769), .A2(n10626), .ZN(n7542) );
  OAI22_X1 U8815 ( .A1(n10626), .A2(n7708), .B1(n7704), .B2(n10620), .ZN(n7540) );
  AOI21_X1 U8816 ( .B1(n10771), .B2(n9111), .A(n7540), .ZN(n7541) );
  OAI211_X1 U8817 ( .C1(n10768), .C2(n9022), .A(n7542), .B(n7541), .ZN(
        P2_U3223) );
  NAND2_X1 U8818 ( .A1(n7543), .A2(n9695), .ZN(n7546) );
  AOI22_X1 U8819 ( .A1(n9697), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7007), .B2(
        n7544), .ZN(n7545) );
  NAND2_X1 U8820 ( .A1(n8305), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7554) );
  OR2_X1 U8821 ( .A1(n8307), .A2(n10754), .ZN(n7553) );
  AND2_X1 U8822 ( .A1(n7548), .A2(n7547), .ZN(n7549) );
  OR2_X1 U8823 ( .A1(n7549), .A2(n7568), .ZN(n7844) );
  OR2_X1 U8824 ( .A1(n8324), .A2(n7844), .ZN(n7552) );
  INV_X1 U8825 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7550) );
  OR2_X1 U8826 ( .A1(n9702), .A2(n7550), .ZN(n7551) );
  NAND4_X1 U8827 ( .A1(n7554), .A2(n7553), .A3(n7552), .A4(n7551), .ZN(n9961)
         );
  INV_X2 U8828 ( .A(n9961), .ZN(n10757) );
  NAND2_X1 U8829 ( .A1(n7555), .A2(n9695), .ZN(n7558) );
  AOI22_X1 U8830 ( .A1(n9697), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7007), .B2(
        n7556), .ZN(n7557) );
  OR2_X1 U8831 ( .A1(n10733), .A2(n8201), .ZN(n7592) );
  INV_X1 U8832 ( .A(n9744), .ZN(n7560) );
  AND2_X1 U8833 ( .A1(n10687), .A2(n9749), .ZN(n9741) );
  INV_X1 U8834 ( .A(n9741), .ZN(n7559) );
  NOR2_X1 U8835 ( .A1(n7560), .A2(n7559), .ZN(n9901) );
  NAND2_X1 U8836 ( .A1(n10682), .A2(n9901), .ZN(n7562) );
  NAND2_X1 U8837 ( .A1(n10733), .A2(n8201), .ZN(n9751) );
  AND2_X1 U8838 ( .A1(n9751), .A2(n10716), .ZN(n9674) );
  OR2_X1 U8839 ( .A1(n7560), .A2(n9674), .ZN(n9905) );
  NAND2_X1 U8840 ( .A1(n10748), .A2(n10757), .ZN(n9758) );
  AND2_X1 U8841 ( .A1(n9905), .A2(n9758), .ZN(n7561) );
  OR2_X1 U8842 ( .A1(n7563), .A2(n8301), .ZN(n7566) );
  AOI22_X1 U8843 ( .A1(n9697), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7007), .B2(
        n7564), .ZN(n7565) );
  NAND2_X1 U8844 ( .A1(n9700), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7573) );
  INV_X1 U8845 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7567) );
  OR2_X1 U8846 ( .A1(n9702), .A2(n7567), .ZN(n7572) );
  NOR2_X1 U8847 ( .A1(n7568), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7569) );
  OR2_X1 U8848 ( .A1(n7577), .A2(n7569), .ZN(n9311) );
  OR2_X1 U8849 ( .A1(n8324), .A2(n9311), .ZN(n7571) );
  INV_X1 U8850 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7583) );
  OR2_X1 U8851 ( .A1(n9705), .A2(n7583), .ZN(n7570) );
  NAND4_X1 U8852 ( .A1(n7573), .A2(n7572), .A3(n7571), .A4(n7570), .ZN(n9960)
         );
  INV_X1 U8853 ( .A(n9904), .ZN(n9755) );
  NAND2_X1 U8854 ( .A1(n10759), .A2(n10787), .ZN(n9757) );
  NAND2_X1 U8855 ( .A1(n9755), .A2(n9757), .ZN(n9677) );
  XNOR2_X1 U8856 ( .A(n7634), .B(n9677), .ZN(n10762) );
  NAND2_X1 U8857 ( .A1(n10852), .A2(n10828), .ZN(n10202) );
  NAND2_X1 U8858 ( .A1(n9756), .A2(n9758), .ZN(n7595) );
  INV_X1 U8859 ( .A(n10748), .ZN(n7849) );
  XNOR2_X1 U8860 ( .A(n7636), .B(n7637), .ZN(n10764) );
  NAND2_X1 U8861 ( .A1(n10764), .A2(n10190), .ZN(n7591) );
  NAND2_X1 U8862 ( .A1(n10852), .A2(n10747), .ZN(n10198) );
  NAND2_X1 U8863 ( .A1(n8258), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7582) );
  OR2_X1 U8864 ( .A1(n8307), .A2(n7576), .ZN(n7581) );
  OR2_X1 U8865 ( .A1(n7577), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7578) );
  NAND2_X1 U8866 ( .A1(n7641), .A2(n7578), .ZN(n8006) );
  OR2_X1 U8867 ( .A1(n8324), .A2(n8006), .ZN(n7580) );
  INV_X1 U8868 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7639) );
  OR2_X1 U8869 ( .A1(n9705), .A2(n7639), .ZN(n7579) );
  NAND4_X1 U8870 ( .A1(n7582), .A2(n7581), .A3(n7580), .A4(n7579), .ZN(n9959)
         );
  OAI22_X1 U8871 ( .A1(n10852), .A2(n7583), .B1(n9311), .B2(n10847), .ZN(n7584) );
  AOI21_X1 U8872 ( .B1(n7585), .B2(n9959), .A(n7584), .ZN(n7586) );
  OAI21_X1 U8873 ( .B1(n10757), .B2(n10198), .A(n7586), .ZN(n7589) );
  NAND2_X1 U8874 ( .A1(n7587), .A2(n5394), .ZN(n7638) );
  OAI211_X1 U8875 ( .C1(n7587), .C2(n5394), .A(n7638), .B(n10818), .ZN(n10760)
         );
  NOR2_X1 U8876 ( .A1(n10760), .A2(n10180), .ZN(n7588) );
  AOI211_X1 U8877 ( .C1(n10732), .C2(n10759), .A(n7589), .B(n7588), .ZN(n7590)
         );
  OAI211_X1 U8878 ( .C1(n10762), .C2(n10202), .A(n7591), .B(n7590), .ZN(
        P1_U3283) );
  INV_X1 U8879 ( .A(n7592), .ZN(n7593) );
  AOI21_X1 U8880 ( .B1(n10717), .B2(n9674), .A(n7593), .ZN(n7594) );
  XNOR2_X1 U8881 ( .A(n7594), .B(n7595), .ZN(n10751) );
  XNOR2_X1 U8882 ( .A(n7596), .B(n7595), .ZN(n10753) );
  NAND2_X1 U8883 ( .A1(n10753), .A2(n10190), .ZN(n7604) );
  INV_X1 U8884 ( .A(n7844), .ZN(n7597) );
  AOI22_X1 U8885 ( .A1(n10697), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7597), .B2(
        n10730), .ZN(n7598) );
  OAI21_X1 U8886 ( .B1(n10198), .B2(n8201), .A(n7598), .ZN(n7602) );
  XNOR2_X1 U8887 ( .A(n10714), .B(n7849), .ZN(n7600) );
  AND2_X1 U8888 ( .A1(n9960), .A2(n10590), .ZN(n7599) );
  AOI21_X1 U8889 ( .B1(n7600), .B2(n10818), .A(n7599), .ZN(n10750) );
  NOR2_X1 U8890 ( .A1(n10750), .A2(n10180), .ZN(n7601) );
  AOI211_X1 U8891 ( .C1(n10732), .C2(n10748), .A(n7602), .B(n7601), .ZN(n7603)
         );
  OAI211_X1 U8892 ( .C1(n10751), .C2(n10202), .A(n7604), .B(n7603), .ZN(
        P1_U3284) );
  NOR2_X1 U8893 ( .A1(n8878), .A2(n7605), .ZN(n7606) );
  AOI211_X1 U8894 ( .C1(n8876), .C2(n8899), .A(n7607), .B(n7606), .ZN(n7608)
         );
  OAI21_X1 U8895 ( .B1(n7609), .B2(n7900), .A(n7608), .ZN(n7616) );
  XNOR2_X1 U8896 ( .A(n7626), .B(n8744), .ZN(n7697) );
  XOR2_X1 U8897 ( .A(n8900), .B(n7697), .Z(n7614) );
  AOI211_X1 U8898 ( .C1(n7614), .C2(n7613), .A(n8870), .B(n7699), .ZN(n7615)
         );
  AOI211_X1 U8899 ( .C1(n7626), .C2(n8867), .A(n7616), .B(n7615), .ZN(n7617)
         );
  INV_X1 U8900 ( .A(n7617), .ZN(P2_U3171) );
  INV_X1 U8901 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7624) );
  NAND3_X1 U8902 ( .A1(n7619), .A2(n10632), .A3(n7618), .ZN(n7620) );
  NAND2_X1 U8903 ( .A1(n7621), .A2(n7620), .ZN(n7625) );
  NAND2_X1 U8904 ( .A1(n7625), .A2(n10785), .ZN(n7623) );
  NAND2_X1 U8905 ( .A1(n7626), .A2(n9237), .ZN(n7622) );
  OAI211_X1 U8906 ( .C1(n7624), .C2(n10785), .A(n7623), .B(n7622), .ZN(
        P2_U3417) );
  NAND2_X1 U8907 ( .A1(n7625), .A2(n10781), .ZN(n7628) );
  NAND2_X1 U8908 ( .A1(n7626), .A2(n6290), .ZN(n7627) );
  OAI211_X1 U8909 ( .C1(n10781), .C2(n7382), .A(n7628), .B(n7627), .ZN(
        P2_U3468) );
  OAI222_X1 U8910 ( .A1(n4944), .A2(n8244), .B1(P2_U3151), .B2(n6746), .C1(
        n7629), .C2(n8472), .ZN(P2_U3274) );
  NAND2_X1 U8911 ( .A1(n7630), .A2(n9695), .ZN(n7633) );
  AOI22_X1 U8912 ( .A1(n9697), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7007), .B2(
        n7631), .ZN(n7632) );
  INV_X1 U8913 ( .A(n9959), .ZN(n10756) );
  OR2_X1 U8914 ( .A1(n10790), .A2(n10756), .ZN(n9772) );
  NAND2_X1 U8915 ( .A1(n10790), .A2(n10756), .ZN(n9761) );
  AND2_X1 U8916 ( .A1(n9772), .A2(n9761), .ZN(n9679) );
  XOR2_X1 U8917 ( .A(n9679), .B(n7675), .Z(n10793) );
  XOR2_X1 U8918 ( .A(n7684), .B(n9679), .Z(n10796) );
  NAND2_X1 U8919 ( .A1(n10796), .A2(n10190), .ZN(n7653) );
  INV_X1 U8920 ( .A(n7686), .ZN(n7688) );
  AOI211_X1 U8921 ( .C1(n10790), .C2(n7638), .A(n10257), .B(n7688), .ZN(n10788) );
  INV_X1 U8922 ( .A(n10790), .ZN(n8011) );
  INV_X1 U8923 ( .A(n10198), .ZN(n10172) );
  OAI22_X1 U8924 ( .A1(n10852), .A2(n7639), .B1(n8006), .B2(n10847), .ZN(n7649) );
  NAND2_X1 U8925 ( .A1(n8258), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7647) );
  OR2_X1 U8926 ( .A1(n8307), .A2(n10804), .ZN(n7646) );
  INV_X1 U8927 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7685) );
  OR2_X1 U8928 ( .A1(n9705), .A2(n7685), .ZN(n7645) );
  NAND2_X1 U8929 ( .A1(n7641), .A2(n7640), .ZN(n7642) );
  NAND2_X1 U8930 ( .A1(n7643), .A2(n7642), .ZN(n8092) );
  OR2_X1 U8931 ( .A1(n8324), .A2(n8092), .ZN(n7644) );
  NAND4_X1 U8932 ( .A1(n7647), .A2(n7646), .A3(n7645), .A4(n7644), .ZN(n9958)
         );
  NOR2_X1 U8933 ( .A1(n10193), .A2(n10786), .ZN(n7648) );
  AOI211_X1 U8934 ( .C1(n10172), .C2(n9960), .A(n7649), .B(n7648), .ZN(n7650)
         );
  OAI21_X1 U8935 ( .B1(n8011), .B2(n10845), .A(n7650), .ZN(n7651) );
  AOI21_X1 U8936 ( .B1(n10788), .B2(n4942), .A(n7651), .ZN(n7652) );
  OAI211_X1 U8937 ( .C1(n10793), .C2(n10202), .A(n7653), .B(n7652), .ZN(
        P1_U3282) );
  AOI21_X1 U8938 ( .B1(n7795), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7654), .ZN(
        n7656) );
  INV_X1 U8939 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7801) );
  MUX2_X1 U8940 ( .A(n7801), .B(P1_REG1_REG_14__SCAN_IN), .S(n8063), .Z(n7655)
         );
  NOR2_X1 U8941 ( .A1(n7656), .A2(n7655), .ZN(n8062) );
  AOI211_X1 U8942 ( .C1(n7656), .C2(n7655), .A(n8062), .B(n10067), .ZN(n7665)
         );
  NAND2_X1 U8943 ( .A1(n8063), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7657) );
  OAI21_X1 U8944 ( .B1(n8063), .B2(P1_REG2_REG_14__SCAN_IN), .A(n7657), .ZN(
        n7660) );
  NOR2_X1 U8945 ( .A1(n7659), .A2(n7660), .ZN(n8059) );
  AOI211_X1 U8946 ( .C1(n7660), .C2(n7659), .A(n8059), .B(n10037), .ZN(n7664)
         );
  INV_X1 U8947 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7662) );
  NAND2_X1 U8948 ( .A1(n10041), .A2(n8063), .ZN(n7661) );
  NAND2_X1 U8949 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9287) );
  OAI211_X1 U8950 ( .C1(n7662), .C2(n10044), .A(n7661), .B(n9287), .ZN(n7663)
         );
  OR3_X1 U8951 ( .A1(n7665), .A2(n7664), .A3(n7663), .ZN(P1_U3257) );
  NAND2_X1 U8952 ( .A1(n7667), .A2(n7666), .ZN(n7669) );
  XNOR2_X1 U8953 ( .A(n7669), .B(n7668), .ZN(n10775) );
  XNOR2_X1 U8954 ( .A(n7670), .B(n8497), .ZN(n7671) );
  OAI222_X1 U8955 ( .A1(n9150), .A2(n7830), .B1(n9148), .B2(n7828), .C1(n9145), 
        .C2(n7671), .ZN(n10776) );
  NAND2_X1 U8956 ( .A1(n10776), .A2(n10626), .ZN(n7674) );
  OAI22_X1 U8957 ( .A1(n10626), .A2(n5894), .B1(n7833), .B2(n10620), .ZN(n7672) );
  AOI21_X1 U8958 ( .B1(n10778), .B2(n9111), .A(n7672), .ZN(n7673) );
  OAI211_X1 U8959 ( .C1(n9129), .C2(n10775), .A(n7674), .B(n7673), .ZN(
        P2_U3222) );
  AOI22_X1 U8960 ( .A1(n9697), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7007), .B2(
        n7677), .ZN(n7678) );
  OR2_X1 U8961 ( .A1(n8078), .A2(n10786), .ZN(n9773) );
  NAND2_X1 U8962 ( .A1(n8078), .A2(n10786), .ZN(n9767) );
  INV_X1 U8963 ( .A(n9680), .ZN(n7680) );
  NAND3_X1 U8964 ( .A1(n7681), .A2(n9761), .A3(n7680), .ZN(n7682) );
  NAND2_X1 U8965 ( .A1(n7799), .A2(n7682), .ZN(n7683) );
  AOI222_X1 U8966 ( .A1(n10828), .A2(n7683), .B1(n8110), .B2(n10590), .C1(
        n9959), .C2(n10747), .ZN(n10800) );
  XNOR2_X1 U8967 ( .A(n7810), .B(n9680), .ZN(n10803) );
  NAND2_X1 U8968 ( .A1(n10803), .A2(n10190), .ZN(n7692) );
  OAI22_X1 U8969 ( .A1(n10852), .A2(n7685), .B1(n8092), .B2(n10847), .ZN(n7690) );
  INV_X1 U8970 ( .A(n8078), .ZN(n10801) );
  INV_X1 U8971 ( .A(n7814), .ZN(n7687) );
  OAI211_X1 U8972 ( .C1(n10801), .C2(n7688), .A(n7687), .B(n10818), .ZN(n10799) );
  NOR2_X1 U8973 ( .A1(n10799), .A2(n10180), .ZN(n7689) );
  AOI211_X1 U8974 ( .C1(n10732), .C2(n8078), .A(n7690), .B(n7689), .ZN(n7691)
         );
  OAI211_X1 U8975 ( .C1(n10697), .C2(n10800), .A(n7692), .B(n7691), .ZN(
        P1_U3281) );
  INV_X1 U8976 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7693) );
  INV_X1 U8977 ( .A(n8253), .ZN(n7695) );
  OAI222_X1 U8978 ( .A1(n10406), .A2(n7693), .B1(n10404), .B2(n7695), .C1(
        P1_U3086), .C2(n9709), .ZN(P1_U3333) );
  OAI222_X1 U8979 ( .A1(n8472), .A2(n7696), .B1(n4944), .B2(n7695), .C1(n7694), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  INV_X1 U8980 ( .A(n7697), .ZN(n7698) );
  XNOR2_X1 U8982 ( .A(n7824), .B(n10858), .ZN(n7829) );
  XNOR2_X1 U8983 ( .A(n7829), .B(n8899), .ZN(n7707) );
  NOR2_X1 U8984 ( .A1(n8878), .A2(n7700), .ZN(n7701) );
  AOI211_X1 U8985 ( .C1(n8876), .C2(n7889), .A(n7702), .B(n7701), .ZN(n7703)
         );
  OAI21_X1 U8986 ( .B1(n7704), .B2(n7900), .A(n7703), .ZN(n7705) );
  AOI21_X1 U8987 ( .B1(n10771), .B2(n8867), .A(n7705), .ZN(n7706) );
  OAI21_X1 U8988 ( .B1(n7707), .B2(n8870), .A(n7706), .ZN(P2_U3157) );
  AOI22_X1 U8989 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n7778), .B1(n7780), .B2(
        n7743), .ZN(n7712) );
  AOI21_X1 U8990 ( .B1(n7713), .B2(n7712), .A(n7774), .ZN(n7735) );
  AOI22_X1 U8991 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n7780), .B1(n7778), .B2(
        n5912), .ZN(n7719) );
  NAND2_X1 U8992 ( .A1(n7716), .A2(n7720), .ZN(n7717) );
  XNOR2_X1 U8993 ( .A(n7716), .B(n10570), .ZN(n10574) );
  NAND2_X1 U8994 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n10574), .ZN(n10573) );
  OAI21_X1 U8995 ( .B1(n7719), .B2(n7718), .A(n7777), .ZN(n7733) );
  INV_X1 U8996 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7731) );
  MUX2_X1 U8997 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8679), .Z(n7781) );
  XNOR2_X1 U8998 ( .A(n7781), .B(n7778), .ZN(n7727) );
  MUX2_X1 U8999 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8679), .Z(n7724) );
  OR2_X1 U9000 ( .A1(n7724), .A2(n7720), .ZN(n7725) );
  XNOR2_X1 U9001 ( .A(n7724), .B(n10570), .ZN(n10577) );
  NAND2_X1 U9002 ( .A1(n7725), .A2(n10575), .ZN(n7726) );
  NAND2_X1 U9003 ( .A1(n7727), .A2(n7726), .ZN(n7782) );
  OAI21_X1 U9004 ( .B1(n7727), .B2(n7726), .A(n7782), .ZN(n7729) );
  NOR2_X1 U9005 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9515), .ZN(n7898) );
  NOR2_X1 U9006 ( .A1(n10504), .A2(n7780), .ZN(n7728) );
  AOI211_X1 U9007 ( .C1(n7729), .C2(n10579), .A(n7898), .B(n7728), .ZN(n7730)
         );
  OAI21_X1 U9008 ( .B1(n10569), .B2(n7731), .A(n7730), .ZN(n7732) );
  AOI21_X1 U9009 ( .B1(n7733), .B2(n10580), .A(n7732), .ZN(n7734) );
  OAI21_X1 U9010 ( .B1(n7735), .B2(n10561), .A(n7734), .ZN(P2_U3194) );
  XNOR2_X1 U9011 ( .A(n7736), .B(n4961), .ZN(n7739) );
  OAI222_X1 U9012 ( .A1(n9148), .A2(n7896), .B1(n9150), .B2(n8155), .C1(n7739), 
        .C2(n9145), .ZN(n7850) );
  INV_X1 U9013 ( .A(n7850), .ZN(n7747) );
  AND2_X1 U9014 ( .A1(n7741), .A2(n7740), .ZN(n7742) );
  XNOR2_X1 U9015 ( .A(n7742), .B(n4961), .ZN(n7851) );
  INV_X1 U9016 ( .A(n7903), .ZN(n7856) );
  NOR2_X1 U9017 ( .A1(n7856), .A2(n9159), .ZN(n7745) );
  OAI22_X1 U9018 ( .A1(n10626), .A2(n7743), .B1(n7901), .B2(n10620), .ZN(n7744) );
  AOI211_X1 U9019 ( .C1(n7851), .C2(n9161), .A(n7745), .B(n7744), .ZN(n7746)
         );
  OAI21_X1 U9020 ( .B1(n7747), .B2(n9163), .A(n7746), .ZN(P2_U3221) );
  AND2_X1 U9021 ( .A1(n10746), .A2(n8459), .ZN(n7748) );
  AOI21_X1 U9022 ( .B1(n10733), .B2(n8438), .A(n7748), .ZN(n7764) );
  NAND2_X1 U9023 ( .A1(n8204), .A2(n6806), .ZN(n7752) );
  NAND2_X1 U9024 ( .A1(n9962), .A2(n8459), .ZN(n7751) );
  NAND2_X1 U9025 ( .A1(n7752), .A2(n7751), .ZN(n8196) );
  NAND2_X1 U9026 ( .A1(n8204), .A2(n4947), .ZN(n7754) );
  NAND2_X1 U9027 ( .A1(n9962), .A2(n6806), .ZN(n7753) );
  NAND2_X1 U9028 ( .A1(n7754), .A2(n7753), .ZN(n7755) );
  XNOR2_X1 U9029 ( .A(n7755), .B(n8460), .ZN(n8195) );
  NAND2_X1 U9030 ( .A1(n10733), .A2(n4947), .ZN(n7757) );
  NAND2_X1 U9031 ( .A1(n10746), .A2(n8438), .ZN(n7756) );
  NAND2_X1 U9032 ( .A1(n7757), .A2(n7756), .ZN(n7758) );
  XNOR2_X1 U9033 ( .A(n7758), .B(n8460), .ZN(n7761) );
  INV_X1 U9034 ( .A(n7761), .ZN(n7759) );
  NAND2_X1 U9035 ( .A1(n7760), .A2(n7759), .ZN(n7841) );
  NAND2_X1 U9036 ( .A1(n7762), .A2(n7761), .ZN(n7763) );
  OAI21_X1 U9037 ( .B1(n7764), .B2(n5035), .A(n7842), .ZN(n7765) );
  NAND2_X1 U9038 ( .A1(n7765), .A2(n9651), .ZN(n7770) );
  INV_X1 U9039 ( .A(n7766), .ZN(n7768) );
  OAI22_X1 U9040 ( .A1(n9639), .A2(n10720), .B1(n9654), .B2(n10728), .ZN(n7767) );
  AOI211_X1 U9041 ( .C1(n9582), .C2(n9961), .A(n7768), .B(n7767), .ZN(n7769)
         );
  OAI211_X1 U9042 ( .C1(n5270), .C2(n9661), .A(n7770), .B(n7769), .ZN(P1_U3221) );
  INV_X1 U9043 ( .A(n8267), .ZN(n7773) );
  OR2_X1 U9044 ( .A1(n7771), .A2(P1_U3086), .ZN(n9875) );
  INV_X1 U9045 ( .A(n9875), .ZN(n9951) );
  AOI21_X1 U9046 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n10399), .A(n9951), .ZN(
        n7772) );
  OAI21_X1 U9047 ( .B1(n7773), .B2(n10404), .A(n7772), .ZN(P1_U3332) );
  AOI21_X1 U9048 ( .B1(n7776), .B2(n7775), .A(n7911), .ZN(n7793) );
  NAND2_X1 U9049 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n7779), .ZN(n7916) );
  OAI21_X1 U9050 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n7779), .A(n7916), .ZN(
        n7791) );
  INV_X1 U9051 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7789) );
  MUX2_X1 U9052 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8679), .Z(n7922) );
  XNOR2_X1 U9053 ( .A(n7922), .B(n7910), .ZN(n7785) );
  OR2_X1 U9054 ( .A1(n7781), .A2(n7780), .ZN(n7783) );
  NAND2_X1 U9055 ( .A1(n7783), .A2(n7782), .ZN(n7784) );
  NAND2_X1 U9056 ( .A1(n7785), .A2(n7784), .ZN(n7923) );
  OAI21_X1 U9057 ( .B1(n7785), .B2(n7784), .A(n7923), .ZN(n7787) );
  NOR2_X1 U9058 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5684), .ZN(n7953) );
  NOR2_X1 U9059 ( .A1(n10504), .A2(n7921), .ZN(n7786) );
  AOI211_X1 U9060 ( .C1(n7787), .C2(n10579), .A(n7953), .B(n7786), .ZN(n7788)
         );
  OAI21_X1 U9061 ( .B1(n10569), .B2(n7789), .A(n7788), .ZN(n7790) );
  AOI21_X1 U9062 ( .B1(n7791), .B2(n10580), .A(n7790), .ZN(n7792) );
  OAI21_X1 U9063 ( .B1(n7793), .B2(n10561), .A(n7792), .ZN(P2_U3195) );
  NAND2_X1 U9064 ( .A1(n7799), .A2(n9767), .ZN(n7798) );
  AOI22_X1 U9065 ( .A1(n9697), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7007), .B2(
        n7795), .ZN(n7796) );
  INV_X1 U9066 ( .A(n8110), .ZN(n10826) );
  OR2_X1 U9067 ( .A1(n8112), .A2(n10826), .ZN(n9775) );
  NAND2_X1 U9068 ( .A1(n8112), .A2(n10826), .ZN(n9768) );
  NAND2_X1 U9069 ( .A1(n9775), .A2(n9768), .ZN(n9682) );
  INV_X1 U9070 ( .A(n9682), .ZN(n7812) );
  NAND2_X1 U9071 ( .A1(n7798), .A2(n7812), .ZN(n8044) );
  NAND3_X1 U9072 ( .A1(n7799), .A2(n9767), .A3(n9682), .ZN(n7800) );
  NAND2_X1 U9073 ( .A1(n8044), .A2(n7800), .ZN(n7809) );
  NAND2_X1 U9074 ( .A1(n8258), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7808) );
  INV_X1 U9075 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10849) );
  OR2_X1 U9076 ( .A1(n9705), .A2(n10849), .ZN(n7807) );
  OR2_X1 U9077 ( .A1(n8307), .A2(n7801), .ZN(n7806) );
  AND2_X1 U9078 ( .A1(n7803), .A2(n7802), .ZN(n7804) );
  OR2_X1 U9079 ( .A1(n7804), .A2(n8036), .ZN(n10848) );
  OR2_X1 U9080 ( .A1(n8324), .A2(n10848), .ZN(n7805) );
  NAND4_X1 U9081 ( .A1(n7808), .A2(n7807), .A3(n7806), .A4(n7805), .ZN(n10369)
         );
  AOI222_X1 U9082 ( .A1(n10828), .A2(n7809), .B1(n10369), .B2(n10590), .C1(
        n9958), .C2(n10747), .ZN(n10808) );
  AOI21_X1 U9083 ( .B1(n8078), .B2(n9958), .A(n7810), .ZN(n7811) );
  XNOR2_X1 U9084 ( .A(n8030), .B(n7812), .ZN(n10812) );
  NAND2_X1 U9085 ( .A1(n10812), .A2(n10190), .ZN(n7818) );
  OAI22_X1 U9086 ( .A1(n10852), .A2(n7813), .B1(n8118), .B2(n10847), .ZN(n7816) );
  NAND2_X1 U9087 ( .A1(n7814), .A2(n10809), .ZN(n10816) );
  OAI211_X1 U9088 ( .C1(n7814), .C2(n10809), .A(n10816), .B(n10818), .ZN(
        n10807) );
  NOR2_X1 U9089 ( .A1(n10807), .A2(n10180), .ZN(n7815) );
  AOI211_X1 U9090 ( .C1(n10732), .C2(n8112), .A(n7816), .B(n7815), .ZN(n7817)
         );
  OAI211_X1 U9091 ( .C1(n10697), .C2(n10808), .A(n7818), .B(n7817), .ZN(
        P1_U3280) );
  NAND2_X1 U9092 ( .A1(n8267), .A2(n7819), .ZN(n7821) );
  NAND2_X1 U9093 ( .A1(n7820), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8685) );
  OAI211_X1 U9094 ( .C1(n7822), .C2(n8472), .A(n7821), .B(n8685), .ZN(P2_U3272) );
  INV_X1 U9095 ( .A(n7824), .ZN(n7825) );
  NOR2_X1 U9096 ( .A1(n10858), .A2(n7825), .ZN(n7827) );
  XNOR2_X1 U9097 ( .A(n10778), .B(n8744), .ZN(n7888) );
  XOR2_X1 U9098 ( .A(n7889), .B(n7888), .Z(n7891) );
  XOR2_X1 U9099 ( .A(n7892), .B(n7891), .Z(n7836) );
  INV_X1 U9100 ( .A(n8876), .ZN(n8837) );
  INV_X1 U9101 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9533) );
  OAI22_X1 U9102 ( .A1(n8837), .A2(n7830), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9533), .ZN(n7831) );
  AOI21_X1 U9103 ( .B1(n8834), .B2(n8899), .A(n7831), .ZN(n7832) );
  OAI21_X1 U9104 ( .B1(n7833), .B2(n7900), .A(n7832), .ZN(n7834) );
  AOI21_X1 U9105 ( .B1(n10778), .B2(n8867), .A(n7834), .ZN(n7835) );
  OAI21_X1 U9106 ( .B1(n7836), .B2(n8870), .A(n7835), .ZN(P2_U3176) );
  NAND2_X1 U9107 ( .A1(n10748), .A2(n4947), .ZN(n7838) );
  NAND2_X1 U9108 ( .A1(n9961), .A2(n8438), .ZN(n7837) );
  NAND2_X1 U9109 ( .A1(n7838), .A2(n7837), .ZN(n7839) );
  XNOR2_X1 U9110 ( .A(n7839), .B(n8460), .ZN(n7978) );
  AND2_X1 U9111 ( .A1(n9961), .A2(n8459), .ZN(n7840) );
  AOI21_X1 U9112 ( .B1(n10748), .B2(n8438), .A(n7840), .ZN(n7979) );
  XNOR2_X1 U9113 ( .A(n7978), .B(n7979), .ZN(n7975) );
  NAND2_X1 U9114 ( .A1(n7977), .A2(n7975), .ZN(n7987) );
  OAI21_X1 U9115 ( .B1(n7975), .B2(n7977), .A(n7987), .ZN(n7843) );
  NAND2_X1 U9116 ( .A1(n7843), .A2(n9651), .ZN(n7848) );
  OAI22_X1 U9117 ( .A1(n9655), .A2(n10787), .B1(n9654), .B2(n7844), .ZN(n7845)
         );
  AOI211_X1 U9118 ( .C1(n9658), .C2(n10746), .A(n7846), .B(n7845), .ZN(n7847)
         );
  OAI211_X1 U9119 ( .C1(n7849), .C2(n9661), .A(n7848), .B(n7847), .ZN(P1_U3231) );
  INV_X1 U9120 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7852) );
  AOI21_X1 U9121 ( .B1(n10632), .B2(n7851), .A(n7850), .ZN(n7854) );
  MUX2_X1 U9122 ( .A(n7852), .B(n7854), .S(n10785), .Z(n7853) );
  OAI21_X1 U9123 ( .B1(n7856), .B2(n9252), .A(n7853), .ZN(P2_U3426) );
  MUX2_X1 U9124 ( .A(n5912), .B(n7854), .S(n10781), .Z(n7855) );
  OAI21_X1 U9125 ( .B1(n7856), .B2(n9213), .A(n7855), .ZN(P2_U3471) );
  XOR2_X1 U9126 ( .A(n7857), .B(n8577), .Z(n7858) );
  AOI222_X1 U9127 ( .A1(n10611), .A2(n7858), .B1(n8898), .B2(n10607), .C1(
        n8897), .C2(n10608), .ZN(n9216) );
  INV_X1 U9128 ( .A(n9216), .ZN(n7861) );
  NAND2_X1 U9129 ( .A1(n7948), .A2(n10779), .ZN(n9215) );
  OAI22_X1 U9130 ( .A1(n9215), .A2(n7859), .B1(n7952), .B2(n10620), .ZN(n7860)
         );
  OAI21_X1 U9131 ( .B1(n7861), .B2(n7860), .A(n10626), .ZN(n7865) );
  OAI21_X1 U9132 ( .B1(n8577), .B2(n7863), .A(n7862), .ZN(n9214) );
  AOI22_X1 U9133 ( .A1(n9214), .A2(n9161), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n9163), .ZN(n7864) );
  NAND2_X1 U9134 ( .A1(n7865), .A2(n7864), .ZN(P2_U3220) );
  INV_X1 U9135 ( .A(n8271), .ZN(n7881) );
  OAI222_X1 U9136 ( .A1(n4944), .A2(n7881), .B1(n8472), .B2(n5726), .C1(n7866), 
        .C2(P2_U3151), .ZN(P2_U3271) );
  INV_X1 U9137 ( .A(n8276), .ZN(n7884) );
  OAI222_X1 U9138 ( .A1(n4944), .A2(n7884), .B1(P2_U3151), .B2(n7868), .C1(
        n7867), .C2(n8472), .ZN(P2_U3270) );
  OAI211_X1 U9139 ( .C1(n7870), .C2(n8582), .A(n7869), .B(n10611), .ZN(n7872)
         );
  AOI22_X1 U9140 ( .A1(n10608), .A2(n8895), .B1(n10607), .B2(n8897), .ZN(n7871) );
  NAND2_X1 U9141 ( .A1(n7872), .A2(n7871), .ZN(n8012) );
  INV_X1 U9142 ( .A(n8012), .ZN(n7879) );
  OAI21_X1 U9143 ( .B1(n7875), .B2(n7874), .A(n7873), .ZN(n8013) );
  INV_X1 U9144 ( .A(n8698), .ZN(n8885) );
  INV_X1 U9145 ( .A(n10626), .ZN(n9157) );
  AOI22_X1 U9146 ( .A1(n9157), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n9156), .B2(
        n8881), .ZN(n7876) );
  OAI21_X1 U9147 ( .B1(n8885), .B2(n9159), .A(n7876), .ZN(n7877) );
  AOI21_X1 U9148 ( .B1(n8013), .B2(n9161), .A(n7877), .ZN(n7878) );
  OAI21_X1 U9149 ( .B1(n7879), .B2(n9163), .A(n7878), .ZN(P2_U3218) );
  INV_X1 U9150 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7880) );
  OAI222_X1 U9151 ( .A1(P1_U3086), .A2(n7882), .B1(n10404), .B2(n7881), .C1(
        n7880), .C2(n10406), .ZN(P1_U3331) );
  INV_X1 U9152 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7883) );
  OAI222_X1 U9153 ( .A1(P1_U3086), .A2(n7885), .B1(n10404), .B2(n7884), .C1(
        n7883), .C2(n10406), .ZN(P1_U3330) );
  INV_X1 U9154 ( .A(n8288), .ZN(n7906) );
  INV_X1 U9155 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7886) );
  OAI222_X1 U9156 ( .A1(P1_U3086), .A2(n7887), .B1(n10404), .B2(n7906), .C1(
        n7886), .C2(n10406), .ZN(P1_U3329) );
  INV_X1 U9157 ( .A(n7888), .ZN(n7890) );
  XNOR2_X1 U9158 ( .A(n8739), .B(n7903), .ZN(n7893) );
  NOR2_X1 U9159 ( .A1(n7893), .A2(n8898), .ZN(n7945) );
  INV_X1 U9160 ( .A(n7945), .ZN(n7894) );
  NAND2_X1 U9161 ( .A1(n7893), .A2(n8898), .ZN(n7946) );
  NAND2_X1 U9162 ( .A1(n7894), .A2(n7946), .ZN(n7895) );
  XNOR2_X1 U9163 ( .A(n7947), .B(n7895), .ZN(n7905) );
  NOR2_X1 U9164 ( .A1(n8878), .A2(n7896), .ZN(n7897) );
  AOI211_X1 U9165 ( .C1(n8876), .C2(n7949), .A(n7898), .B(n7897), .ZN(n7899)
         );
  OAI21_X1 U9166 ( .B1(n7901), .B2(n7900), .A(n7899), .ZN(n7902) );
  AOI21_X1 U9167 ( .B1(n7903), .B2(n8867), .A(n7902), .ZN(n7904) );
  OAI21_X1 U9168 ( .B1(n7905), .B2(n8870), .A(n7904), .ZN(P2_U3164) );
  OAI222_X1 U9169 ( .A1(n8472), .A2(n7908), .B1(P2_U3151), .B2(n7907), .C1(
        n4944), .C2(n7906), .ZN(P2_U3269) );
  NOR2_X1 U9170 ( .A1(n7910), .A2(n7909), .ZN(n7912) );
  NAND2_X1 U9171 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8911), .ZN(n7913) );
  OAI21_X1 U9172 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8911), .A(n7913), .ZN(
        n7914) );
  AOI21_X1 U9173 ( .B1(n5025), .B2(n7914), .A(n8906), .ZN(n7935) );
  AOI22_X1 U9174 ( .A1(n7920), .A2(n8024), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n8911), .ZN(n7919) );
  NAND2_X1 U9175 ( .A1(n7921), .A2(n7915), .ZN(n7917) );
  OAI21_X1 U9176 ( .B1(n7919), .B2(n7918), .A(n8908), .ZN(n7933) );
  INV_X1 U9177 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7931) );
  MUX2_X1 U9178 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8679), .Z(n8912) );
  XNOR2_X1 U9179 ( .A(n8912), .B(n7920), .ZN(n7926) );
  OR2_X1 U9180 ( .A1(n7922), .A2(n7921), .ZN(n7924) );
  NAND2_X1 U9181 ( .A1(n7924), .A2(n7923), .ZN(n7925) );
  NAND2_X1 U9182 ( .A1(n7926), .A2(n7925), .ZN(n8913) );
  OAI21_X1 U9183 ( .B1(n7926), .B2(n7925), .A(n8913), .ZN(n7929) );
  INV_X1 U9184 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7927) );
  NOR2_X1 U9185 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7927), .ZN(n8151) );
  NOR2_X1 U9186 ( .A1(n10504), .A2(n8911), .ZN(n7928) );
  AOI211_X1 U9187 ( .C1(n7929), .C2(n10579), .A(n8151), .B(n7928), .ZN(n7930)
         );
  OAI21_X1 U9188 ( .B1(n10569), .B2(n7931), .A(n7930), .ZN(n7932) );
  AOI21_X1 U9189 ( .B1(n7933), .B2(n10580), .A(n7932), .ZN(n7934) );
  OAI21_X1 U9190 ( .B1(n7935), .B2(n10561), .A(n7934), .ZN(P2_U3196) );
  AOI21_X1 U9191 ( .B1(n9264), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n7936), .ZN(
        n7937) );
  OAI21_X1 U9192 ( .B1(n8302), .B2(n4944), .A(n7937), .ZN(P2_U3268) );
  INV_X1 U9193 ( .A(n8578), .ZN(n8026) );
  NOR2_X1 U9194 ( .A1(n8026), .A2(n10617), .ZN(n7940) );
  INV_X1 U9195 ( .A(n8589), .ZN(n8499) );
  XNOR2_X1 U9196 ( .A(n7938), .B(n8499), .ZN(n7939) );
  OAI222_X1 U9197 ( .A1(n9148), .A2(n8155), .B1(n9150), .B2(n8799), .C1(n9145), 
        .C2(n7939), .ZN(n8019) );
  AOI211_X1 U9198 ( .C1(n9156), .C2(n8152), .A(n7940), .B(n8019), .ZN(n7944)
         );
  OAI21_X1 U9199 ( .B1(n7942), .B2(n8589), .A(n7941), .ZN(n8020) );
  AOI22_X1 U9200 ( .A1(n8020), .A2(n9161), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n9163), .ZN(n7943) );
  OAI21_X1 U9201 ( .B1(n7944), .B2(n9163), .A(n7943), .ZN(P2_U3219) );
  INV_X1 U9202 ( .A(n7948), .ZN(n7959) );
  AOI21_X1 U9203 ( .B1(n7947), .B2(n7946), .A(n7945), .ZN(n7951) );
  XNOR2_X1 U9204 ( .A(n7948), .B(n8744), .ZN(n8145) );
  XNOR2_X1 U9205 ( .A(n8145), .B(n7949), .ZN(n7950) );
  NAND2_X1 U9206 ( .A1(n7951), .A2(n7950), .ZN(n8147) );
  OAI211_X1 U9207 ( .C1(n7951), .C2(n7950), .A(n8147), .B(n8848), .ZN(n7958)
         );
  INV_X1 U9208 ( .A(n7952), .ZN(n7956) );
  AOI21_X1 U9209 ( .B1(n8834), .B2(n8898), .A(n7953), .ZN(n7954) );
  OAI21_X1 U9210 ( .B1(n8695), .B2(n8837), .A(n7954), .ZN(n7955) );
  AOI21_X1 U9211 ( .B1(n7956), .B2(n8880), .A(n7955), .ZN(n7957) );
  OAI211_X1 U9212 ( .C1(n7959), .C2(n8884), .A(n7958), .B(n7957), .ZN(P2_U3174) );
  OAI222_X1 U9213 ( .A1(n10406), .A2(n7960), .B1(n10404), .B2(n8302), .C1(
        n10074), .C2(P1_U3086), .ZN(P1_U3328) );
  OAI211_X1 U9214 ( .C1(n7962), .C2(n8594), .A(n7961), .B(n10611), .ZN(n7964)
         );
  NAND2_X1 U9215 ( .A1(n10607), .A2(n8896), .ZN(n7963) );
  OAI211_X1 U9216 ( .C1(n9147), .C2(n9150), .A(n7964), .B(n7963), .ZN(n9209)
         );
  INV_X1 U9217 ( .A(n9209), .ZN(n7971) );
  INV_X1 U9218 ( .A(n7965), .ZN(n7966) );
  AOI21_X1 U9219 ( .B1(n8594), .B2(n7967), .A(n7966), .ZN(n9210) );
  INV_X1 U9220 ( .A(n8801), .ZN(n9253) );
  AOI22_X1 U9221 ( .A1(n9157), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n9156), .B2(
        n8796), .ZN(n7968) );
  OAI21_X1 U9222 ( .B1(n9253), .B2(n9159), .A(n7968), .ZN(n7969) );
  AOI21_X1 U9223 ( .B1(n9210), .B2(n9161), .A(n7969), .ZN(n7970) );
  OAI21_X1 U9224 ( .B1(n7971), .B2(n9163), .A(n7970), .ZN(P2_U3217) );
  NAND2_X1 U9225 ( .A1(n10759), .A2(n4947), .ZN(n7973) );
  NAND2_X1 U9226 ( .A1(n9960), .A2(n8438), .ZN(n7972) );
  NAND2_X1 U9227 ( .A1(n7973), .A2(n7972), .ZN(n7974) );
  XNOR2_X1 U9228 ( .A(n7974), .B(n6829), .ZN(n7986) );
  AND2_X1 U9229 ( .A1(n7975), .A2(n7986), .ZN(n7976) );
  INV_X1 U9230 ( .A(n7986), .ZN(n7981) );
  INV_X1 U9231 ( .A(n7978), .ZN(n7980) );
  NAND2_X1 U9232 ( .A1(n7980), .A2(n7979), .ZN(n7984) );
  AND2_X1 U9233 ( .A1(n9960), .A2(n8459), .ZN(n7982) );
  AOI21_X1 U9234 ( .B1(n10759), .B2(n8438), .A(n7982), .ZN(n9308) );
  AND2_X1 U9235 ( .A1(n7989), .A2(n9308), .ZN(n7983) );
  INV_X1 U9236 ( .A(n7984), .ZN(n7985) );
  NAND2_X1 U9237 ( .A1(n4984), .A2(n7987), .ZN(n9306) );
  NAND2_X1 U9238 ( .A1(n7988), .A2(n9306), .ZN(n8002) );
  INV_X1 U9239 ( .A(n8002), .ZN(n8001) );
  INV_X1 U9240 ( .A(n9305), .ZN(n8000) );
  NAND2_X1 U9241 ( .A1(n10790), .A2(n4947), .ZN(n7992) );
  NAND2_X1 U9242 ( .A1(n9959), .A2(n8438), .ZN(n7991) );
  NAND2_X1 U9243 ( .A1(n7992), .A2(n7991), .ZN(n7993) );
  XNOR2_X1 U9244 ( .A(n7993), .B(n6829), .ZN(n7995) );
  AND2_X1 U9245 ( .A1(n9959), .A2(n8459), .ZN(n7994) );
  AOI21_X1 U9246 ( .B1(n10790), .B2(n8438), .A(n7994), .ZN(n7996) );
  NAND2_X1 U9247 ( .A1(n7995), .A2(n7996), .ZN(n8086) );
  INV_X1 U9248 ( .A(n7995), .ZN(n7998) );
  INV_X1 U9249 ( .A(n7996), .ZN(n7997) );
  NAND2_X1 U9250 ( .A1(n7998), .A2(n7997), .ZN(n7999) );
  NOR3_X1 U9251 ( .A1(n8001), .A2(n8000), .A3(n8003), .ZN(n8005) );
  NAND2_X1 U9252 ( .A1(n8002), .A2(n9305), .ZN(n8004) );
  NAND2_X1 U9253 ( .A1(n8004), .A2(n8003), .ZN(n8087) );
  INV_X1 U9254 ( .A(n8087), .ZN(n8085) );
  OAI21_X1 U9255 ( .B1(n8005), .B2(n8085), .A(n9651), .ZN(n8010) );
  OAI22_X1 U9256 ( .A1(n9639), .A2(n10787), .B1(n9654), .B2(n8006), .ZN(n8007)
         );
  AOI211_X1 U9257 ( .C1(n9582), .C2(n9958), .A(n8008), .B(n8007), .ZN(n8009)
         );
  OAI211_X1 U9258 ( .C1(n8011), .C2(n9661), .A(n8010), .B(n8009), .ZN(P1_U3236) );
  AOI21_X1 U9259 ( .B1(n10632), .B2(n8013), .A(n8012), .ZN(n8016) );
  MUX2_X1 U9260 ( .A(n8014), .B(n8016), .S(n10785), .Z(n8015) );
  OAI21_X1 U9261 ( .B1(n8885), .B2(n9252), .A(n8015), .ZN(P2_U3435) );
  MUX2_X1 U9262 ( .A(n8017), .B(n8016), .S(n10781), .Z(n8018) );
  OAI21_X1 U9263 ( .B1(n8885), .B2(n9213), .A(n8018), .ZN(P2_U3474) );
  AOI21_X1 U9264 ( .B1(n10632), .B2(n8020), .A(n8019), .ZN(n8023) );
  MUX2_X1 U9265 ( .A(n8021), .B(n8023), .S(n10785), .Z(n8022) );
  OAI21_X1 U9266 ( .B1(n8026), .B2(n9252), .A(n8022), .ZN(P2_U3432) );
  MUX2_X1 U9267 ( .A(n8024), .B(n8023), .S(n10781), .Z(n8025) );
  OAI21_X1 U9268 ( .B1(n8026), .B2(n9213), .A(n8025), .ZN(P2_U3473) );
  INV_X1 U9269 ( .A(n10369), .ZN(n8046) );
  AOI22_X1 U9270 ( .A1(n9697), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7007), .B2(
        n8063), .ZN(n8028) );
  OAI21_X1 U9271 ( .B1(n8112), .B2(n8110), .A(n8030), .ZN(n8031) );
  AOI22_X1 U9272 ( .A1(n9697), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7007), .B2(
        n8064), .ZN(n8033) );
  NAND2_X1 U9273 ( .A1(n8305), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n8043) );
  INV_X1 U9274 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n8035) );
  OR2_X1 U9275 ( .A1(n8307), .A2(n8035), .ZN(n8042) );
  OR2_X1 U9276 ( .A1(n8036), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8038) );
  NAND2_X1 U9277 ( .A1(n8038), .A2(n8037), .ZN(n9653) );
  OR2_X1 U9278 ( .A1(n8324), .A2(n9653), .ZN(n8041) );
  INV_X1 U9279 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n8039) );
  OR2_X1 U9280 ( .A1(n9702), .A2(n8039), .ZN(n8040) );
  NAND4_X1 U9281 ( .A1(n8043), .A2(n8042), .A3(n8041), .A4(n8040), .ZN(n9957)
         );
  OR2_X1 U9282 ( .A1(n9788), .A2(n10824), .ZN(n9916) );
  NAND2_X1 U9283 ( .A1(n9788), .A2(n10824), .ZN(n9913) );
  NAND2_X1 U9284 ( .A1(n9916), .A2(n9913), .ZN(n9685) );
  XNOR2_X1 U9285 ( .A(n8123), .B(n9685), .ZN(n10376) );
  INV_X1 U9286 ( .A(n10202), .ZN(n10182) );
  NAND2_X1 U9287 ( .A1(n8351), .A2(n8046), .ZN(n9912) );
  INV_X1 U9288 ( .A(n9912), .ZN(n8045) );
  OR2_X1 U9289 ( .A1(n8351), .A2(n8046), .ZN(n9911) );
  XNOR2_X1 U9290 ( .A(n8140), .B(n9685), .ZN(n10374) );
  AOI211_X1 U9291 ( .C1(n9788), .C2(n10817), .A(n10257), .B(n8128), .ZN(n10372) );
  NAND2_X1 U9292 ( .A1(n10372), .A2(n4942), .ZN(n8056) );
  NAND2_X1 U9293 ( .A1(n8258), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8051) );
  INV_X1 U9294 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n8047) );
  OR2_X1 U9295 ( .A1(n9705), .A2(n8047), .ZN(n8050) );
  INV_X1 U9296 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9998) );
  OR2_X1 U9297 ( .A1(n8307), .A2(n9998), .ZN(n8049) );
  XNOR2_X1 U9298 ( .A(P1_REG3_REG_16__SCAN_IN), .B(n8132), .ZN(n9580) );
  OR2_X1 U9299 ( .A1(n8324), .A2(n9580), .ZN(n8048) );
  NAND4_X1 U9300 ( .A1(n8051), .A2(n8050), .A3(n8049), .A4(n8048), .ZN(n10368)
         );
  INV_X1 U9301 ( .A(n10368), .ZN(n10252) );
  INV_X1 U9302 ( .A(n9653), .ZN(n8052) );
  AOI22_X1 U9303 ( .A1(n10697), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8052), .B2(
        n10730), .ZN(n8053) );
  OAI21_X1 U9304 ( .B1(n10193), .B2(n10252), .A(n8053), .ZN(n8054) );
  AOI21_X1 U9305 ( .B1(n10172), .B2(n10369), .A(n8054), .ZN(n8055) );
  OAI211_X1 U9306 ( .C1(n10371), .C2(n10845), .A(n8056), .B(n8055), .ZN(n8057)
         );
  AOI21_X1 U9307 ( .B1(n10182), .B2(n10374), .A(n8057), .ZN(n8058) );
  OAI21_X1 U9308 ( .B1(n10376), .B2(n10265), .A(n8058), .ZN(P1_U3278) );
  XOR2_X1 U9309 ( .A(n8064), .B(n10004), .Z(n8060) );
  INV_X1 U9310 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8061) );
  NAND2_X1 U9311 ( .A1(n8060), .A2(n8061), .ZN(n8072) );
  NOR2_X1 U9312 ( .A1(n8061), .A2(n8060), .ZN(n10005) );
  NOR2_X1 U9313 ( .A1(n10037), .A2(n10005), .ZN(n8071) );
  NAND2_X1 U9314 ( .A1(n8065), .A2(n8035), .ZN(n8067) );
  INV_X1 U9315 ( .A(n9996), .ZN(n8066) );
  NAND3_X1 U9316 ( .A1(n10024), .A2(n8067), .A3(n8066), .ZN(n8069) );
  AND2_X1 U9317 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9657) );
  AOI21_X1 U9318 ( .B1(n10059), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n9657), .ZN(
        n8068) );
  OAI211_X1 U9319 ( .C1(n10063), .C2(n10003), .A(n8069), .B(n8068), .ZN(n8070)
         );
  AOI21_X1 U9320 ( .B1(n8072), .B2(n8071), .A(n8070), .ZN(n8073) );
  INV_X1 U9321 ( .A(n8073), .ZN(P1_U3258) );
  INV_X1 U9322 ( .A(n8086), .ZN(n8084) );
  NAND2_X1 U9323 ( .A1(n8078), .A2(n4947), .ZN(n8075) );
  NAND2_X1 U9324 ( .A1(n9958), .A2(n8438), .ZN(n8074) );
  NAND2_X1 U9325 ( .A1(n8075), .A2(n8074), .ZN(n8076) );
  XNOR2_X1 U9326 ( .A(n8076), .B(n6829), .ZN(n8079) );
  AND2_X1 U9327 ( .A1(n9958), .A2(n8459), .ZN(n8077) );
  AOI21_X1 U9328 ( .B1(n8078), .B2(n8438), .A(n8077), .ZN(n8080) );
  NAND2_X1 U9329 ( .A1(n8079), .A2(n8080), .ZN(n8113) );
  INV_X1 U9330 ( .A(n8079), .ZN(n8082) );
  INV_X1 U9331 ( .A(n8080), .ZN(n8081) );
  NAND2_X1 U9332 ( .A1(n8082), .A2(n8081), .ZN(n8083) );
  NOR3_X1 U9333 ( .A1(n8085), .A2(n8084), .A3(n8088), .ZN(n8091) );
  NAND2_X1 U9334 ( .A1(n8087), .A2(n8086), .ZN(n8089) );
  NAND2_X1 U9335 ( .A1(n8089), .A2(n8088), .ZN(n8114) );
  INV_X1 U9336 ( .A(n8114), .ZN(n8090) );
  OAI21_X1 U9337 ( .B1(n8091), .B2(n8090), .A(n9651), .ZN(n8096) );
  OAI22_X1 U9338 ( .A1(n9655), .A2(n10826), .B1(n9654), .B2(n8092), .ZN(n8093)
         );
  AOI211_X1 U9339 ( .C1(n9658), .C2(n9959), .A(n8094), .B(n8093), .ZN(n8095)
         );
  OAI211_X1 U9340 ( .C1(n10801), .C2(n9661), .A(n8096), .B(n8095), .ZN(
        P1_U3224) );
  INV_X1 U9341 ( .A(n8099), .ZN(n8500) );
  XNOR2_X1 U9342 ( .A(n8097), .B(n8500), .ZN(n9208) );
  OAI211_X1 U9343 ( .C1(n8100), .C2(n8099), .A(n8098), .B(n10611), .ZN(n8102)
         );
  AOI22_X1 U9344 ( .A1(n8893), .A2(n10608), .B1(n10607), .B2(n8895), .ZN(n8101) );
  NAND2_X1 U9345 ( .A1(n8102), .A2(n8101), .ZN(n9205) );
  INV_X1 U9346 ( .A(n9206), .ZN(n8104) );
  AOI22_X1 U9347 ( .A1(n9157), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n9156), .B2(
        n8807), .ZN(n8103) );
  OAI21_X1 U9348 ( .B1(n8104), .B2(n9159), .A(n8103), .ZN(n8105) );
  AOI21_X1 U9349 ( .B1(n9205), .B2(n10626), .A(n8105), .ZN(n8106) );
  OAI21_X1 U9350 ( .B1(n9129), .B2(n9208), .A(n8106), .ZN(P2_U3216) );
  NAND2_X1 U9351 ( .A1(n8112), .A2(n4947), .ZN(n8108) );
  NAND2_X1 U9352 ( .A1(n8110), .A2(n8438), .ZN(n8107) );
  NAND2_X1 U9353 ( .A1(n8108), .A2(n8107), .ZN(n8109) );
  XNOR2_X1 U9354 ( .A(n8109), .B(n8460), .ZN(n8352) );
  AND2_X1 U9355 ( .A1(n8110), .A2(n8459), .ZN(n8111) );
  AOI21_X1 U9356 ( .B1(n8112), .B2(n8438), .A(n8111), .ZN(n8353) );
  XNOR2_X1 U9357 ( .A(n8352), .B(n8353), .ZN(n8116) );
  OAI21_X1 U9358 ( .B1(n8116), .B2(n8115), .A(n8356), .ZN(n8117) );
  NAND2_X1 U9359 ( .A1(n8117), .A2(n9651), .ZN(n8122) );
  OAI22_X1 U9360 ( .A1(n9639), .A2(n10786), .B1(n9654), .B2(n8118), .ZN(n8119)
         );
  AOI211_X1 U9361 ( .C1(n9582), .C2(n10369), .A(n8120), .B(n8119), .ZN(n8121)
         );
  OAI211_X1 U9362 ( .C1(n10809), .C2(n9661), .A(n8122), .B(n8121), .ZN(
        P1_U3234) );
  NAND2_X1 U9363 ( .A1(n8125), .A2(n9695), .ZN(n8127) );
  AOI22_X1 U9364 ( .A1(n9697), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7007), .B2(
        n10020), .ZN(n8126) );
  NAND2_X1 U9365 ( .A1(n10365), .A2(n10252), .ZN(n9919) );
  XNOR2_X1 U9366 ( .A(n8209), .B(n9686), .ZN(n10367) );
  INV_X1 U9367 ( .A(n8128), .ZN(n8129) );
  INV_X1 U9368 ( .A(n10365), .ZN(n9790) );
  AOI211_X1 U9369 ( .C1(n10365), .C2(n8129), .A(n10257), .B(n10254), .ZN(
        n10364) );
  NOR2_X1 U9370 ( .A1(n9790), .A2(n10845), .ZN(n8131) );
  OAI22_X1 U9371 ( .A1(n10852), .A2(n8047), .B1(n9580), .B2(n10847), .ZN(n8130) );
  AOI211_X1 U9372 ( .C1(n10364), .C2(n4942), .A(n8131), .B(n8130), .ZN(n8144)
         );
  AOI21_X1 U9373 ( .B1(P1_REG3_REG_16__SCAN_IN), .B2(n8132), .A(
        P1_REG3_REG_17__SCAN_IN), .ZN(n8133) );
  NOR2_X1 U9374 ( .A1(n8133), .A2(n8219), .ZN(n10259) );
  NAND2_X1 U9375 ( .A1(n6737), .A2(n10259), .ZN(n8139) );
  INV_X1 U9376 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10021) );
  OR2_X1 U9377 ( .A1(n8307), .A2(n10021), .ZN(n8138) );
  INV_X1 U9378 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n8134) );
  OR2_X1 U9379 ( .A1(n9702), .A2(n8134), .ZN(n8137) );
  INV_X1 U9380 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8135) );
  OR2_X1 U9381 ( .A1(n9705), .A2(n8135), .ZN(n8136) );
  NAND4_X1 U9382 ( .A1(n8139), .A2(n8138), .A3(n8137), .A4(n8136), .ZN(n9956)
         );
  INV_X1 U9383 ( .A(n9956), .ZN(n10236) );
  NAND2_X1 U9384 ( .A1(n8141), .A2(n9913), .ZN(n8313) );
  XNOR2_X1 U9385 ( .A(n8313), .B(n9686), .ZN(n8142) );
  OAI222_X1 U9386 ( .A1(n10823), .A2(n10236), .B1(n10825), .B2(n10824), .C1(
        n8142), .C2(n10794), .ZN(n10363) );
  NAND2_X1 U9387 ( .A1(n10363), .A2(n10852), .ZN(n8143) );
  OAI211_X1 U9388 ( .C1(n10367), .C2(n10265), .A(n8144), .B(n8143), .ZN(
        P1_U3277) );
  XNOR2_X1 U9389 ( .A(n8578), .B(n8744), .ZN(n8694) );
  XOR2_X1 U9390 ( .A(n8897), .B(n8694), .Z(n8150) );
  INV_X1 U9391 ( .A(n8697), .ZN(n8149) );
  AOI21_X1 U9392 ( .B1(n8150), .B2(n8148), .A(n8149), .ZN(n8158) );
  AOI21_X1 U9393 ( .B1(n8876), .B2(n8896), .A(n8151), .ZN(n8154) );
  NAND2_X1 U9394 ( .A1(n8880), .A2(n8152), .ZN(n8153) );
  OAI211_X1 U9395 ( .C1(n8155), .C2(n8878), .A(n8154), .B(n8153), .ZN(n8156)
         );
  AOI21_X1 U9396 ( .B1(n8578), .B2(n8867), .A(n8156), .ZN(n8157) );
  OAI21_X1 U9397 ( .B1(n8158), .B2(n8870), .A(n8157), .ZN(P2_U3155) );
  INV_X1 U9398 ( .A(n8159), .ZN(n8160) );
  NAND2_X1 U9399 ( .A1(n8160), .A2(SI_29_), .ZN(n8164) );
  NAND2_X1 U9400 ( .A1(n8164), .A2(n8163), .ZN(n8470) );
  INV_X1 U9401 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8691) );
  INV_X1 U9402 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8474) );
  MUX2_X1 U9403 ( .A(n8691), .B(n8474), .S(n8169), .Z(n8165) );
  INV_X1 U9404 ( .A(SI_30_), .ZN(n9433) );
  NAND2_X1 U9405 ( .A1(n8165), .A2(n9433), .ZN(n8168) );
  INV_X1 U9406 ( .A(n8165), .ZN(n8166) );
  NAND2_X1 U9407 ( .A1(n8166), .A2(SI_30_), .ZN(n8167) );
  NAND2_X1 U9408 ( .A1(n8168), .A2(n8167), .ZN(n8469) );
  MUX2_X1 U9409 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8169), .Z(n8171) );
  INV_X1 U9410 ( .A(SI_31_), .ZN(n8170) );
  XNOR2_X1 U9411 ( .A(n8171), .B(n8170), .ZN(n8172) );
  NAND2_X1 U9412 ( .A1(n9662), .A2(n8473), .ZN(n8175) );
  OR2_X1 U9413 ( .A1(n8475), .A2(n6436), .ZN(n8174) );
  INV_X1 U9414 ( .A(n8176), .ZN(n8177) );
  NAND2_X1 U9415 ( .A1(n8178), .A2(n8177), .ZN(n9221) );
  INV_X1 U9416 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8183) );
  NAND2_X1 U9417 ( .A1(n5459), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8181) );
  INV_X1 U9418 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8179) );
  OR2_X1 U9419 ( .A1(n5760), .A2(n8179), .ZN(n8180) );
  OAI211_X1 U9420 ( .C1(n8183), .C2(n8182), .A(n8181), .B(n8180), .ZN(n8184)
         );
  INV_X1 U9421 ( .A(n8184), .ZN(n8185) );
  NAND2_X1 U9422 ( .A1(n8186), .A2(n8185), .ZN(n8886) );
  NAND2_X1 U9423 ( .A1(n8886), .A2(n8187), .ZN(n8190) );
  NOR2_X1 U9424 ( .A1(n8190), .A2(n10782), .ZN(n9219) );
  AOI21_X1 U9425 ( .B1(n10782), .B2(P2_REG0_REG_31__SCAN_IN), .A(n9219), .ZN(
        n8188) );
  OAI21_X1 U9426 ( .B1(n8484), .B2(n9221), .A(n8188), .ZN(P2_U3458) );
  NOR2_X1 U9427 ( .A1(n8190), .A2(n10780), .ZN(n9165) );
  AOI21_X1 U9428 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n10780), .A(n9165), .ZN(
        n8189) );
  OAI21_X1 U9429 ( .B1(n8484), .B2(n9213), .A(n8189), .ZN(P2_U3490) );
  INV_X1 U9430 ( .A(n8190), .ZN(n8192) );
  NOR2_X1 U9431 ( .A1(n8191), .A2(n10620), .ZN(n9017) );
  NOR3_X1 U9432 ( .A1(n8192), .A2(n9163), .A3(n9017), .ZN(n9014) );
  NOR2_X1 U9433 ( .A1(n10626), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8193) );
  OAI22_X1 U9434 ( .A1(n8484), .A2(n9159), .B1(n9014), .B2(n8193), .ZN(
        P2_U3202) );
  XOR2_X1 U9435 ( .A(n8196), .B(n8195), .Z(n8197) );
  XNOR2_X1 U9436 ( .A(n8194), .B(n8197), .ZN(n8207) );
  INV_X1 U9437 ( .A(n9654), .ZN(n9590) );
  INV_X1 U9438 ( .A(n8198), .ZN(n8199) );
  AOI22_X1 U9439 ( .A1(n9658), .A2(n8200), .B1(n9590), .B2(n8199), .ZN(n8206)
         );
  NOR2_X1 U9440 ( .A1(n9655), .A2(n8201), .ZN(n8202) );
  AOI211_X1 U9441 ( .C1(n8204), .C2(n9642), .A(n8203), .B(n8202), .ZN(n8205)
         );
  OAI211_X1 U9442 ( .C1(n8207), .C2(n9632), .A(n8206), .B(n8205), .ZN(P1_U3213) );
  NAND2_X1 U9443 ( .A1(n8210), .A2(n9695), .ZN(n8212) );
  AOI22_X1 U9444 ( .A1(n9697), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7007), .B2(
        n10036), .ZN(n8211) );
  NAND2_X1 U9445 ( .A1(n10360), .A2(n9956), .ZN(n8213) );
  AOI22_X1 U9446 ( .A1(n9697), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7007), .B2(
        n10040), .ZN(n8215) );
  NAND2_X1 U9447 ( .A1(n9700), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8228) );
  INV_X1 U9448 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8217) );
  OR2_X1 U9449 ( .A1(n9705), .A2(n8217), .ZN(n8227) );
  INV_X1 U9450 ( .A(n8234), .ZN(n8223) );
  INV_X1 U9451 ( .A(n8219), .ZN(n8221) );
  INV_X1 U9452 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8220) );
  NAND2_X1 U9453 ( .A1(n8221), .A2(n8220), .ZN(n8222) );
  NAND2_X1 U9454 ( .A1(n8223), .A2(n8222), .ZN(n10240) );
  OR2_X1 U9455 ( .A1(n8324), .A2(n10240), .ZN(n8226) );
  INV_X1 U9456 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n8224) );
  OR2_X1 U9457 ( .A1(n9702), .A2(n8224), .ZN(n8225) );
  NAND4_X1 U9458 ( .A1(n8228), .A2(n8227), .A3(n8226), .A4(n8225), .ZN(n10226)
         );
  NAND2_X1 U9459 ( .A1(n10244), .A2(n10253), .ZN(n8229) );
  NAND2_X1 U9460 ( .A1(n8230), .A2(n9695), .ZN(n8232) );
  AOI22_X1 U9461 ( .A1(n9697), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9882), .B2(
        n7007), .ZN(n8231) );
  INV_X1 U9462 ( .A(n10349), .ZN(n10222) );
  NAND2_X1 U9463 ( .A1(n8258), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8239) );
  INV_X1 U9464 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10051) );
  OR2_X1 U9465 ( .A1(n8307), .A2(n10051), .ZN(n8238) );
  OAI21_X1 U9466 ( .B1(n8234), .B2(P1_REG3_REG_19__SCAN_IN), .A(n8233), .ZN(
        n10219) );
  OR2_X1 U9467 ( .A1(n8324), .A2(n10219), .ZN(n8237) );
  INV_X1 U9468 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n8235) );
  OR2_X1 U9469 ( .A1(n9705), .A2(n8235), .ZN(n8236) );
  NAND4_X1 U9470 ( .A1(n8239), .A2(n8238), .A3(n8237), .A4(n8236), .ZN(n9955)
         );
  INV_X1 U9471 ( .A(n9955), .ZN(n10237) );
  NAND2_X1 U9472 ( .A1(n8241), .A2(n9695), .ZN(n8243) );
  NAND2_X1 U9473 ( .A1(n9697), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8242) );
  NAND2_X1 U9474 ( .A1(n10345), .A2(n10335), .ZN(n10184) );
  NAND2_X1 U9475 ( .A1(n9697), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8245) );
  OAI21_X1 U9476 ( .B1(n8247), .B2(P1_REG3_REG_21__SCAN_IN), .A(n8257), .ZN(
        n10192) );
  INV_X1 U9477 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n8250) );
  NAND2_X1 U9478 ( .A1(n8258), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8249) );
  NAND2_X1 U9479 ( .A1(n9700), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n8248) );
  OAI211_X1 U9480 ( .C1(n9705), .C2(n8250), .A(n8249), .B(n8248), .ZN(n8251)
         );
  INV_X1 U9481 ( .A(n8251), .ZN(n8252) );
  OAI21_X1 U9482 ( .B1(n10192), .B2(n8324), .A(n8252), .ZN(n10325) );
  INV_X1 U9483 ( .A(n10325), .ZN(n10214) );
  NAND2_X1 U9484 ( .A1(n10339), .A2(n10214), .ZN(n9805) );
  NAND2_X1 U9485 ( .A1(n8253), .A2(n9695), .ZN(n8255) );
  NAND2_X1 U9486 ( .A1(n9697), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8254) );
  AOI21_X1 U9487 ( .B1(n8257), .B2(n9618), .A(n8256), .ZN(n10173) );
  NAND2_X1 U9488 ( .A1(n10173), .A2(n6737), .ZN(n8264) );
  INV_X1 U9489 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n8261) );
  NAND2_X1 U9490 ( .A1(n9700), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8260) );
  NAND2_X1 U9491 ( .A1(n8258), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8259) );
  OAI211_X1 U9492 ( .C1(n9705), .C2(n8261), .A(n8260), .B(n8259), .ZN(n8262)
         );
  INV_X1 U9493 ( .A(n8262), .ZN(n8263) );
  NAND2_X1 U9494 ( .A1(n8264), .A2(n8263), .ZN(n10161) );
  OR2_X1 U9495 ( .A1(n10178), .A2(n10336), .ZN(n9714) );
  NAND2_X1 U9496 ( .A1(n10178), .A2(n10336), .ZN(n9713) );
  NAND2_X1 U9497 ( .A1(n10167), .A2(n9689), .ZN(n8266) );
  INV_X1 U9498 ( .A(n10178), .ZN(n10329) );
  NAND2_X1 U9499 ( .A1(n10329), .A2(n10336), .ZN(n8265) );
  NAND2_X1 U9500 ( .A1(n9697), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8268) );
  NOR2_X1 U9501 ( .A1(n10321), .A2(n10326), .ZN(n8270) );
  NAND2_X1 U9502 ( .A1(n10321), .A2(n10326), .ZN(n8269) );
  NAND2_X1 U9503 ( .A1(n9697), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8272) );
  NOR2_X1 U9504 ( .A1(n8337), .A2(n10318), .ZN(n8275) );
  NAND2_X1 U9505 ( .A1(n8337), .A2(n10318), .ZN(n8274) );
  NAND2_X1 U9506 ( .A1(n9697), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8277) );
  NAND2_X1 U9507 ( .A1(n8305), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8287) );
  INV_X1 U9508 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n8279) );
  OR2_X1 U9509 ( .A1(n8307), .A2(n8279), .ZN(n8286) );
  INV_X1 U9510 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8280) );
  NAND2_X1 U9511 ( .A1(n8281), .A2(n8280), .ZN(n8282) );
  NAND2_X1 U9512 ( .A1(n8292), .A2(n8282), .ZN(n10140) );
  OR2_X1 U9513 ( .A1(n8324), .A2(n10140), .ZN(n8285) );
  INV_X1 U9514 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n8283) );
  OR2_X1 U9515 ( .A1(n9702), .A2(n8283), .ZN(n8284) );
  NAND4_X1 U9516 ( .A1(n8287), .A2(n8286), .A3(n8285), .A4(n8284), .ZN(n10297)
         );
  NAND2_X1 U9517 ( .A1(n9697), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8289) );
  NAND2_X1 U9518 ( .A1(n8305), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8298) );
  INV_X1 U9519 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n8291) );
  OR2_X1 U9520 ( .A1(n8307), .A2(n8291), .ZN(n8297) );
  INV_X1 U9521 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9637) );
  NAND2_X1 U9522 ( .A1(n8292), .A2(n9637), .ZN(n8293) );
  NAND2_X1 U9523 ( .A1(n8322), .A2(n8293), .ZN(n10126) );
  OR2_X1 U9524 ( .A1(n8324), .A2(n10126), .ZN(n8296) );
  INV_X1 U9525 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n8294) );
  OR2_X1 U9526 ( .A1(n9702), .A2(n8294), .ZN(n8295) );
  NAND4_X1 U9527 ( .A1(n8298), .A2(n8297), .A3(n8296), .A4(n8295), .ZN(n9954)
         );
  NOR2_X1 U9528 ( .A1(n5262), .A2(n10305), .ZN(n8300) );
  NAND2_X1 U9529 ( .A1(n9697), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8303) );
  NAND2_X1 U9530 ( .A1(n8305), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8312) );
  INV_X1 U9531 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8306) );
  OR2_X1 U9532 ( .A1(n8307), .A2(n8306), .ZN(n8311) );
  INV_X1 U9533 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9274) );
  XNOR2_X1 U9534 ( .A(n8322), .B(n9274), .ZN(n9275) );
  OR2_X1 U9535 ( .A1(n8324), .A2(n9275), .ZN(n8310) );
  INV_X1 U9536 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n8308) );
  OR2_X1 U9537 ( .A1(n9702), .A2(n8308), .ZN(n8309) );
  NAND4_X1 U9538 ( .A1(n8312), .A2(n8311), .A3(n8310), .A4(n8309), .ZN(n10296)
         );
  XNOR2_X1 U9539 ( .A(n10091), .B(n10089), .ZN(n10295) );
  NAND2_X1 U9540 ( .A1(n10360), .A2(n10236), .ZN(n9720) );
  INV_X1 U9541 ( .A(n9720), .ZN(n8314) );
  OR2_X1 U9542 ( .A1(n10360), .A2(n10236), .ZN(n9922) );
  OR2_X1 U9543 ( .A1(n10355), .A2(n10253), .ZN(n9719) );
  INV_X1 U9544 ( .A(n9719), .ZN(n8315) );
  AND2_X1 U9545 ( .A1(n10355), .A2(n10253), .ZN(n9718) );
  INV_X1 U9546 ( .A(n9718), .ZN(n9721) );
  OR2_X1 U9547 ( .A1(n10349), .A2(n10237), .ZN(n9717) );
  NAND2_X1 U9548 ( .A1(n10349), .A2(n10237), .ZN(n9925) );
  NAND2_X1 U9549 ( .A1(n9717), .A2(n9925), .ZN(n9688) );
  NAND2_X1 U9550 ( .A1(n10224), .A2(n10225), .ZN(n10223) );
  INV_X1 U9551 ( .A(n9930), .ZN(n8316) );
  NAND2_X1 U9552 ( .A1(n9805), .A2(n10184), .ZN(n8317) );
  NAND2_X1 U9553 ( .A1(n8317), .A2(n9930), .ZN(n9855) );
  INV_X1 U9554 ( .A(n9713), .ZN(n8318) );
  INV_X1 U9555 ( .A(n10326), .ZN(n10176) );
  NAND2_X1 U9556 ( .A1(n9809), .A2(n9838), .ZN(n10153) );
  INV_X1 U9557 ( .A(n9838), .ZN(n8319) );
  NAND2_X1 U9558 ( .A1(n10314), .A2(n10318), .ZN(n9857) );
  NOR2_X1 U9559 ( .A1(n10308), .A2(n9638), .ZN(n9812) );
  INV_X1 U9560 ( .A(n9812), .ZN(n9844) );
  NAND2_X1 U9561 ( .A1(n10131), .A2(n10305), .ZN(n9816) );
  NAND2_X1 U9562 ( .A1(n8320), .A2(n10089), .ZN(n10087) );
  OAI21_X1 U9563 ( .B1(n8320), .B2(n10089), .A(n10087), .ZN(n10292) );
  INV_X1 U9564 ( .A(n10291), .ZN(n8449) );
  AOI211_X1 U9565 ( .C1(n10291), .C2(n10125), .A(n10257), .B(n10070), .ZN(
        n10289) );
  NAND2_X1 U9566 ( .A1(n10289), .A2(n4942), .ZN(n8333) );
  NAND2_X1 U9567 ( .A1(n9700), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8328) );
  INV_X1 U9568 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n8321) );
  OR2_X1 U9569 ( .A1(n9702), .A2(n8321), .ZN(n8327) );
  INV_X1 U9570 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8465) );
  OAI21_X1 U9571 ( .B1(n8322), .B2(n9274), .A(n8465), .ZN(n8323) );
  NAND2_X1 U9572 ( .A1(n8323), .A2(n10099), .ZN(n10114) );
  OR2_X1 U9573 ( .A1(n8324), .A2(n10114), .ZN(n8326) );
  INV_X1 U9574 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n10115) );
  OR2_X1 U9575 ( .A1(n9705), .A2(n10115), .ZN(n8325) );
  NAND4_X1 U9576 ( .A1(n8328), .A2(n8327), .A3(n8326), .A4(n8325), .ZN(n10093)
         );
  INV_X1 U9577 ( .A(n9275), .ZN(n8329) );
  AOI22_X1 U9578 ( .A1(n10697), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n8329), .B2(
        n10730), .ZN(n8330) );
  OAI21_X1 U9579 ( .B1(n10193), .B2(n10288), .A(n8330), .ZN(n8331) );
  AOI21_X1 U9580 ( .B1(n10172), .B2(n9954), .A(n8331), .ZN(n8332) );
  OAI211_X1 U9581 ( .C1(n8449), .C2(n10845), .A(n8333), .B(n8332), .ZN(n8334)
         );
  AOI21_X1 U9582 ( .B1(n10292), .B2(n10182), .A(n8334), .ZN(n8335) );
  OAI21_X1 U9583 ( .B1(n10295), .B2(n10265), .A(n8335), .ZN(P1_U3266) );
  INV_X1 U9584 ( .A(n9811), .ZN(n9691) );
  XNOR2_X1 U9585 ( .A(n8336), .B(n9691), .ZN(n10316) );
  AOI211_X1 U9586 ( .C1(n10314), .C2(n10155), .A(n10257), .B(n10139), .ZN(
        n10313) );
  NOR2_X1 U9587 ( .A1(n8337), .A2(n10845), .ZN(n8340) );
  OAI22_X1 U9588 ( .A1(n10852), .A2(n8338), .B1(n9601), .B2(n10847), .ZN(n8339) );
  AOI211_X1 U9589 ( .C1(n10313), .C2(n4942), .A(n8340), .B(n8339), .ZN(n8346)
         );
  OAI211_X1 U9590 ( .C1(n8342), .C2(n9811), .A(n8341), .B(n10828), .ZN(n8344)
         );
  AOI22_X1 U9591 ( .A1(n10326), .A2(n10747), .B1(n10590), .B2(n10297), .ZN(
        n8343) );
  NAND2_X1 U9592 ( .A1(n8344), .A2(n8343), .ZN(n10312) );
  NAND2_X1 U9593 ( .A1(n10312), .A2(n10852), .ZN(n8345) );
  OAI211_X1 U9594 ( .C1(n10316), .C2(n10265), .A(n8346), .B(n8345), .ZN(
        P1_U3269) );
  NAND2_X1 U9595 ( .A1(n8351), .A2(n4947), .ZN(n8348) );
  NAND2_X1 U9596 ( .A1(n10369), .A2(n8438), .ZN(n8347) );
  NAND2_X1 U9597 ( .A1(n8348), .A2(n8347), .ZN(n8349) );
  XNOR2_X1 U9598 ( .A(n8349), .B(n6829), .ZN(n9283) );
  AND2_X1 U9599 ( .A1(n10369), .A2(n8459), .ZN(n8350) );
  AOI21_X1 U9600 ( .B1(n8351), .B2(n8438), .A(n8350), .ZN(n9282) );
  INV_X1 U9601 ( .A(n8352), .ZN(n8354) );
  AND2_X1 U9602 ( .A1(n8354), .A2(n8353), .ZN(n9280) );
  AOI21_X1 U9603 ( .B1(n9283), .B2(n9282), .A(n9280), .ZN(n8355) );
  INV_X1 U9604 ( .A(n9283), .ZN(n8358) );
  INV_X1 U9605 ( .A(n9282), .ZN(n8357) );
  NAND2_X1 U9606 ( .A1(n9788), .A2(n4947), .ZN(n8360) );
  NAND2_X1 U9607 ( .A1(n9957), .A2(n8438), .ZN(n8359) );
  NAND2_X1 U9608 ( .A1(n8360), .A2(n8359), .ZN(n8361) );
  XNOR2_X1 U9609 ( .A(n8361), .B(n8460), .ZN(n8367) );
  AND2_X2 U9610 ( .A1(n8366), .A2(n8367), .ZN(n9652) );
  NAND2_X1 U9611 ( .A1(n10365), .A2(n4947), .ZN(n8363) );
  NAND2_X1 U9612 ( .A1(n10368), .A2(n8438), .ZN(n8362) );
  NAND2_X1 U9613 ( .A1(n8363), .A2(n8362), .ZN(n8364) );
  XNOR2_X1 U9614 ( .A(n8364), .B(n6829), .ZN(n8373) );
  AND2_X1 U9615 ( .A1(n10368), .A2(n8459), .ZN(n8365) );
  AOI21_X1 U9616 ( .B1(n10365), .B2(n8438), .A(n8365), .ZN(n8372) );
  XNOR2_X1 U9617 ( .A(n8373), .B(n8372), .ZN(n9576) );
  INV_X1 U9618 ( .A(n8366), .ZN(n8369) );
  AND2_X1 U9619 ( .A1(n9957), .A2(n8459), .ZN(n8370) );
  AOI21_X1 U9620 ( .B1(n9788), .B2(n8438), .A(n8370), .ZN(n9648) );
  NAND2_X1 U9621 ( .A1(n10360), .A2(n4947), .ZN(n8376) );
  NAND2_X1 U9622 ( .A1(n9956), .A2(n8438), .ZN(n8375) );
  NAND2_X1 U9623 ( .A1(n8376), .A2(n8375), .ZN(n8377) );
  XNOR2_X1 U9624 ( .A(n8377), .B(n6829), .ZN(n8380) );
  AND2_X1 U9625 ( .A1(n9956), .A2(n8459), .ZN(n8378) );
  AOI21_X1 U9626 ( .B1(n10360), .B2(n8438), .A(n8378), .ZN(n8379) );
  NOR2_X1 U9627 ( .A1(n8380), .A2(n8379), .ZN(n9587) );
  NAND2_X1 U9628 ( .A1(n8380), .A2(n8379), .ZN(n9585) );
  AOI22_X1 U9629 ( .A1(n10355), .A2(n4947), .B1(n8438), .B2(n10226), .ZN(n8381) );
  XNOR2_X1 U9630 ( .A(n8381), .B(n8460), .ZN(n8382) );
  NOR2_X1 U9631 ( .A1(n8383), .A2(n8382), .ZN(n9626) );
  OAI22_X1 U9632 ( .A1(n10244), .A2(n8448), .B1(n10253), .B2(n8447), .ZN(n9627) );
  NAND2_X1 U9633 ( .A1(n8383), .A2(n8382), .ZN(n9624) );
  OAI21_X1 U9634 ( .B1(n9626), .B2(n9627), .A(n9624), .ZN(n9549) );
  NAND2_X1 U9635 ( .A1(n10349), .A2(n4947), .ZN(n8385) );
  NAND2_X1 U9636 ( .A1(n9955), .A2(n8438), .ZN(n8384) );
  NAND2_X1 U9637 ( .A1(n8385), .A2(n8384), .ZN(n8386) );
  XNOR2_X1 U9638 ( .A(n8386), .B(n6829), .ZN(n9551) );
  AND2_X1 U9639 ( .A1(n9955), .A2(n8459), .ZN(n8387) );
  INV_X1 U9640 ( .A(n9551), .ZN(n8389) );
  INV_X1 U9641 ( .A(n9550), .ZN(n8388) );
  NAND2_X1 U9642 ( .A1(n10345), .A2(n4947), .ZN(n8392) );
  NAND2_X1 U9643 ( .A1(n10227), .A2(n8438), .ZN(n8391) );
  NAND2_X1 U9644 ( .A1(n8392), .A2(n8391), .ZN(n8393) );
  XNOR2_X1 U9645 ( .A(n8393), .B(n8460), .ZN(n8398) );
  AOI22_X1 U9646 ( .A1(n10345), .A2(n8438), .B1(n8459), .B2(n10227), .ZN(n8399) );
  XNOR2_X1 U9647 ( .A(n8398), .B(n8399), .ZN(n9607) );
  NAND2_X1 U9648 ( .A1(n10339), .A2(n4947), .ZN(n8395) );
  NAND2_X1 U9649 ( .A1(n10325), .A2(n8438), .ZN(n8394) );
  NAND2_X1 U9650 ( .A1(n8395), .A2(n8394), .ZN(n8396) );
  XNOR2_X1 U9651 ( .A(n8396), .B(n8460), .ZN(n8402) );
  AND2_X1 U9652 ( .A1(n10325), .A2(n8459), .ZN(n8397) );
  XNOR2_X1 U9653 ( .A(n8402), .B(n8403), .ZN(n9560) );
  INV_X1 U9654 ( .A(n8398), .ZN(n8400) );
  NAND2_X1 U9655 ( .A1(n8400), .A2(n8399), .ZN(n9561) );
  NAND2_X1 U9656 ( .A1(n9559), .A2(n8405), .ZN(n9296) );
  NAND2_X1 U9657 ( .A1(n10321), .A2(n4947), .ZN(n8407) );
  NAND2_X1 U9658 ( .A1(n10326), .A2(n8438), .ZN(n8406) );
  NAND2_X1 U9659 ( .A1(n8407), .A2(n8406), .ZN(n8408) );
  XNOR2_X1 U9660 ( .A(n8408), .B(n6829), .ZN(n8418) );
  AND2_X1 U9661 ( .A1(n10326), .A2(n8459), .ZN(n8409) );
  AOI21_X1 U9662 ( .B1(n10321), .B2(n8438), .A(n8409), .ZN(n8419) );
  NAND2_X1 U9663 ( .A1(n8418), .A2(n8419), .ZN(n9293) );
  NAND2_X1 U9664 ( .A1(n10178), .A2(n4947), .ZN(n8411) );
  NAND2_X1 U9665 ( .A1(n10161), .A2(n8438), .ZN(n8410) );
  NAND2_X1 U9666 ( .A1(n8411), .A2(n8410), .ZN(n8412) );
  NAND2_X1 U9667 ( .A1(n10178), .A2(n8438), .ZN(n8414) );
  NAND2_X1 U9668 ( .A1(n10161), .A2(n8459), .ZN(n8413) );
  NAND2_X1 U9669 ( .A1(n9296), .A2(n8417), .ZN(n8432) );
  INV_X1 U9670 ( .A(n8418), .ZN(n8421) );
  INV_X1 U9671 ( .A(n8419), .ZN(n8420) );
  AOI21_X1 U9672 ( .B1(n9295), .B2(n9617), .A(n9292), .ZN(n8422) );
  NAND2_X1 U9673 ( .A1(n10314), .A2(n4947), .ZN(n8424) );
  NAND2_X1 U9674 ( .A1(n10144), .A2(n8438), .ZN(n8423) );
  NAND2_X1 U9675 ( .A1(n8424), .A2(n8423), .ZN(n8425) );
  XNOR2_X1 U9676 ( .A(n8425), .B(n8460), .ZN(n8429) );
  NAND2_X1 U9677 ( .A1(n10314), .A2(n8438), .ZN(n8427) );
  NAND2_X1 U9678 ( .A1(n10144), .A2(n8459), .ZN(n8426) );
  NAND2_X1 U9679 ( .A1(n8427), .A2(n8426), .ZN(n8428) );
  AOI21_X1 U9680 ( .B1(n8429), .B2(n8428), .A(n8433), .ZN(n9595) );
  INV_X1 U9681 ( .A(n8433), .ZN(n8434) );
  NAND2_X1 U9682 ( .A1(n10308), .A2(n4947), .ZN(n8436) );
  NAND2_X1 U9683 ( .A1(n10297), .A2(n8438), .ZN(n8435) );
  NAND2_X1 U9684 ( .A1(n8436), .A2(n8435), .ZN(n8437) );
  XNOR2_X1 U9685 ( .A(n8437), .B(n8460), .ZN(n8443) );
  AOI22_X1 U9686 ( .A1(n10308), .A2(n8438), .B1(n8459), .B2(n10297), .ZN(n8444) );
  XNOR2_X1 U9687 ( .A(n8443), .B(n8444), .ZN(n9569) );
  NAND2_X1 U9688 ( .A1(n10131), .A2(n4947), .ZN(n8440) );
  NAND2_X1 U9689 ( .A1(n9954), .A2(n8438), .ZN(n8439) );
  NAND2_X1 U9690 ( .A1(n8440), .A2(n8439), .ZN(n8441) );
  XNOR2_X1 U9691 ( .A(n8441), .B(n8460), .ZN(n8454) );
  AND2_X1 U9692 ( .A1(n9954), .A2(n8459), .ZN(n8442) );
  AOI21_X1 U9693 ( .B1(n10131), .B2(n8438), .A(n8442), .ZN(n8452) );
  XNOR2_X1 U9694 ( .A(n8454), .B(n8452), .ZN(n9634) );
  INV_X1 U9695 ( .A(n8443), .ZN(n8445) );
  NAND2_X1 U9696 ( .A1(n8445), .A2(n8444), .ZN(n9635) );
  AOI22_X1 U9697 ( .A1(n10291), .A2(n4947), .B1(n8438), .B2(n10296), .ZN(n8446) );
  XOR2_X1 U9698 ( .A(n8460), .B(n8446), .Z(n8451) );
  OAI22_X1 U9699 ( .A1(n8449), .A2(n8448), .B1(n10281), .B2(n8447), .ZN(n8450)
         );
  NOR2_X1 U9700 ( .A1(n8451), .A2(n8450), .ZN(n8456) );
  AOI21_X1 U9701 ( .B1(n8451), .B2(n8450), .A(n8456), .ZN(n9270) );
  INV_X1 U9702 ( .A(n8452), .ZN(n8453) );
  NAND2_X1 U9703 ( .A1(n8454), .A2(n8453), .ZN(n9271) );
  NAND2_X1 U9704 ( .A1(n9269), .A2(n8455), .ZN(n9268) );
  NAND2_X1 U9705 ( .A1(n9697), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8457) );
  AOI22_X1 U9706 ( .A1(n10284), .A2(n4947), .B1(n8438), .B2(n10093), .ZN(n8463) );
  AOI22_X1 U9707 ( .A1(n10284), .A2(n8438), .B1(n8459), .B2(n10093), .ZN(n8461) );
  XNOR2_X1 U9708 ( .A(n8461), .B(n8460), .ZN(n8462) );
  XOR2_X1 U9709 ( .A(n8463), .B(n8462), .Z(n8464) );
  OAI22_X1 U9710 ( .A1(n9639), .A2(n10281), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8465), .ZN(n8467) );
  OAI22_X1 U9711 ( .A1(n9655), .A2(n10280), .B1(n9654), .B2(n10114), .ZN(n8466) );
  AOI211_X1 U9712 ( .C1(n10284), .C2(n9642), .A(n8467), .B(n8466), .ZN(n8468)
         );
  INV_X1 U9713 ( .A(n9696), .ZN(n8692) );
  OAI222_X1 U9714 ( .A1(n8472), .A2(n8474), .B1(n4944), .B2(n8692), .C1(
        P2_U3151), .C2(n8471), .ZN(P2_U3265) );
  NAND2_X1 U9715 ( .A1(n9696), .A2(n8473), .ZN(n8477) );
  OR2_X1 U9716 ( .A1(n8475), .A2(n8474), .ZN(n8476) );
  INV_X1 U9717 ( .A(n8478), .ZN(n8663) );
  NOR2_X1 U9718 ( .A1(n8480), .A2(n8479), .ZN(n8664) );
  INV_X1 U9719 ( .A(n8664), .ZN(n8669) );
  NAND2_X1 U9720 ( .A1(n8669), .A2(n8886), .ZN(n8482) );
  NAND2_X1 U9721 ( .A1(n8482), .A2(n8481), .ZN(n8483) );
  NOR2_X1 U9722 ( .A1(n8484), .A2(n8886), .ZN(n8674) );
  NAND2_X1 U9723 ( .A1(n8485), .A2(n8646), .ZN(n9043) );
  NAND2_X1 U9724 ( .A1(n8642), .A2(n8641), .ZN(n8638) );
  AND2_X1 U9725 ( .A1(n8631), .A2(n8628), .ZN(n9089) );
  NAND4_X1 U9726 ( .A1(n8486), .A2(n8511), .A3(n8512), .A4(n10612), .ZN(n8488)
         );
  NOR3_X1 U9727 ( .A1(n8488), .A2(n8487), .A3(n8529), .ZN(n8489) );
  NAND3_X1 U9728 ( .A1(n8551), .A2(n8490), .A3(n8489), .ZN(n8492) );
  OR3_X1 U9729 ( .A1(n8493), .A2(n8492), .A3(n8491), .ZN(n8494) );
  NOR2_X1 U9730 ( .A1(n8495), .A2(n8494), .ZN(n8496) );
  NAND4_X1 U9731 ( .A1(n8577), .A2(n8497), .A3(n8496), .A4(n4961), .ZN(n8498)
         );
  NAND4_X1 U9732 ( .A1(n9100), .A2(n4975), .A3(n5059), .A4(n8500), .ZN(n8501)
         );
  NOR4_X1 U9733 ( .A1(n9138), .A2(n9089), .A3(n8501), .A4(n9114), .ZN(n8502)
         );
  NAND4_X1 U9734 ( .A1(n5237), .A2(n8502), .A3(n9060), .A4(n9077), .ZN(n8503)
         );
  NOR4_X1 U9735 ( .A1(n8743), .A2(n9043), .A3(n8650), .A4(n8503), .ZN(n8504)
         );
  NAND4_X1 U9736 ( .A1(n8505), .A2(n8669), .A3(n8504), .A4(n8668), .ZN(n8506)
         );
  NOR3_X1 U9737 ( .A1(n8674), .A2(n8507), .A3(n8506), .ZN(n8508) );
  AOI21_X1 U9738 ( .B1(n8512), .B2(n8511), .A(n8510), .ZN(n8521) );
  AOI211_X1 U9739 ( .C1(n8516), .C2(n8515), .A(n8514), .B(n8513), .ZN(n8519)
         );
  NOR2_X1 U9740 ( .A1(n8519), .A2(n8518), .ZN(n8520) );
  NAND2_X1 U9741 ( .A1(n8905), .A2(n10618), .ZN(n8522) );
  NAND2_X1 U9742 ( .A1(n8535), .A2(n8522), .ZN(n8525) );
  NAND2_X1 U9743 ( .A1(n8528), .A2(n8523), .ZN(n8524) );
  MUX2_X1 U9744 ( .A(n8525), .B(n8524), .S(n8610), .Z(n8526) );
  INV_X1 U9745 ( .A(n8528), .ZN(n8530) );
  NOR3_X1 U9746 ( .A1(n8540), .A2(n8530), .A3(n8529), .ZN(n8531) );
  AOI211_X1 U9747 ( .C1(n10636), .C2(n8904), .A(n8543), .B(n8531), .ZN(n8534)
         );
  NOR3_X1 U9748 ( .A1(n8534), .A2(n8533), .A3(n8532), .ZN(n8542) );
  NAND2_X1 U9749 ( .A1(n8536), .A2(n8535), .ZN(n8539) );
  OAI211_X1 U9750 ( .C1(n8540), .C2(n8539), .A(n8538), .B(n8537), .ZN(n8541)
         );
  MUX2_X1 U9751 ( .A(n8542), .B(n8541), .S(n8610), .Z(n8546) );
  OAI21_X1 U9752 ( .B1(n8544), .B2(n8543), .A(n8610), .ZN(n8545) );
  NAND2_X1 U9753 ( .A1(n8546), .A2(n8545), .ZN(n8555) );
  NOR2_X1 U9754 ( .A1(n8550), .A2(n8610), .ZN(n8553) );
  NOR3_X1 U9755 ( .A1(n8565), .A2(n8553), .A3(n8552), .ZN(n8554) );
  NOR3_X1 U9756 ( .A1(n8559), .A2(n8558), .A3(n8570), .ZN(n8560) );
  OAI21_X1 U9757 ( .B1(n8655), .B2(n8563), .A(n8562), .ZN(n8572) );
  INV_X1 U9758 ( .A(n8565), .ZN(n8568) );
  AOI21_X1 U9759 ( .B1(n8568), .B2(n8567), .A(n8566), .ZN(n8571) );
  MUX2_X1 U9760 ( .A(n8575), .B(n8574), .S(n8610), .Z(n8576) );
  MUX2_X1 U9761 ( .A(n8897), .B(n8578), .S(n8610), .Z(n8590) );
  INV_X1 U9762 ( .A(n8579), .ZN(n8581) );
  MUX2_X1 U9763 ( .A(n8581), .B(n5275), .S(n8610), .Z(n8583) );
  AOI211_X1 U9764 ( .C1(n8590), .C2(n8584), .A(n8583), .B(n8582), .ZN(n8585)
         );
  NAND2_X1 U9765 ( .A1(n8586), .A2(n8585), .ZN(n8601) );
  OAI21_X1 U9766 ( .B1(n8610), .B2(n8896), .A(n8698), .ZN(n8596) );
  OAI21_X1 U9767 ( .B1(n8655), .B2(n8799), .A(n8885), .ZN(n8595) );
  INV_X1 U9768 ( .A(n8587), .ZN(n8592) );
  INV_X1 U9769 ( .A(n8588), .ZN(n8591) );
  NOR4_X1 U9770 ( .A1(n8592), .A2(n8591), .A3(n8590), .A4(n8589), .ZN(n8593)
         );
  AOI211_X1 U9771 ( .C1(n8596), .C2(n8595), .A(n8594), .B(n8593), .ZN(n8600)
         );
  NOR2_X1 U9772 ( .A1(n8801), .A2(n8610), .ZN(n8598) );
  NOR2_X1 U9773 ( .A1(n9253), .A2(n8655), .ZN(n8597) );
  MUX2_X1 U9774 ( .A(n8598), .B(n8597), .S(n8810), .Z(n8599) );
  AOI21_X1 U9775 ( .B1(n8601), .B2(n8600), .A(n8599), .ZN(n8609) );
  MUX2_X1 U9776 ( .A(n8894), .B(n9206), .S(n8610), .Z(n8605) );
  NOR2_X1 U9777 ( .A1(n9147), .A2(n8655), .ZN(n8602) );
  AOI21_X1 U9778 ( .B1(n6154), .B2(n8605), .A(n8606), .ZN(n8608) );
  OAI21_X1 U9779 ( .B1(n8655), .B2(n8893), .A(n8708), .ZN(n8604) );
  INV_X1 U9780 ( .A(n8708), .ZN(n9247) );
  OAI21_X1 U9781 ( .B1(n9137), .B2(n8610), .A(n9247), .ZN(n8603) );
  AOI22_X1 U9782 ( .A1(n8606), .A2(n8605), .B1(n8604), .B2(n8603), .ZN(n8607)
         );
  OAI211_X1 U9783 ( .C1(n8609), .C2(n8608), .A(n8607), .B(n8709), .ZN(n8620)
         );
  NOR2_X1 U9784 ( .A1(n9149), .A2(n8655), .ZN(n8612) );
  NOR2_X1 U9785 ( .A1(n8892), .A2(n8610), .ZN(n8611) );
  MUX2_X1 U9786 ( .A(n8612), .B(n8611), .S(n8766), .Z(n8613) );
  NOR2_X1 U9787 ( .A1(n9114), .A2(n8613), .ZN(n8619) );
  INV_X1 U9788 ( .A(n8614), .ZN(n8617) );
  INV_X1 U9789 ( .A(n8615), .ZN(n8616) );
  MUX2_X1 U9790 ( .A(n8617), .B(n8616), .S(n8610), .Z(n8618) );
  AOI21_X1 U9791 ( .B1(n8620), .B2(n8619), .A(n8618), .ZN(n8623) );
  INV_X1 U9792 ( .A(n8623), .ZN(n8625) );
  MUX2_X1 U9793 ( .A(n9236), .B(n9085), .S(n8610), .Z(n8621) );
  AOI21_X1 U9794 ( .B1(n8623), .B2(n8622), .A(n8621), .ZN(n8624) );
  AOI21_X1 U9795 ( .B1(n8626), .B2(n8625), .A(n8624), .ZN(n8629) );
  INV_X1 U9796 ( .A(n8629), .ZN(n8632) );
  MUX2_X1 U9797 ( .A(n9184), .B(n9104), .S(n8610), .Z(n8627) );
  OAI21_X1 U9798 ( .B1(n8632), .B2(n8631), .A(n8630), .ZN(n8635) );
  INV_X1 U9799 ( .A(n8763), .ZN(n9232) );
  MUX2_X1 U9800 ( .A(n9063), .B(n9232), .S(n8610), .Z(n8633) );
  AOI22_X1 U9801 ( .A1(n8635), .A2(n9077), .B1(n8634), .B2(n8633), .ZN(n8640)
         );
  NOR2_X1 U9802 ( .A1(n9179), .A2(n9051), .ZN(n8636) );
  MUX2_X1 U9803 ( .A(n8637), .B(n8636), .S(n8610), .Z(n8639) );
  INV_X1 U9804 ( .A(n8641), .ZN(n8644) );
  INV_X1 U9805 ( .A(n8642), .ZN(n8643) );
  MUX2_X1 U9806 ( .A(n8644), .B(n8643), .S(n8610), .Z(n8645) );
  INV_X1 U9807 ( .A(n8646), .ZN(n8647) );
  MUX2_X1 U9808 ( .A(n8648), .B(n8647), .S(n8610), .Z(n8649) );
  INV_X1 U9809 ( .A(n8651), .ZN(n8652) );
  MUX2_X1 U9810 ( .A(n8652), .B(n6264), .S(n8610), .Z(n8653) );
  MUX2_X1 U9811 ( .A(n9027), .B(n8654), .S(n8610), .Z(n8658) );
  NOR2_X1 U9812 ( .A1(n9027), .A2(n8655), .ZN(n8656) );
  NAND2_X1 U9813 ( .A1(n8659), .A2(n8658), .ZN(n8661) );
  NOR3_X1 U9814 ( .A1(n8671), .A2(n8664), .A3(n8663), .ZN(n8666) );
  NAND2_X1 U9815 ( .A1(n8668), .A2(n8667), .ZN(n8670) );
  OAI21_X1 U9816 ( .B1(n8671), .B2(n8670), .A(n8669), .ZN(n8672) );
  XNOR2_X1 U9817 ( .A(n8678), .B(n8677), .ZN(n8686) );
  NAND3_X1 U9818 ( .A1(n8681), .A2(n8680), .A3(n8679), .ZN(n8682) );
  OAI211_X1 U9819 ( .C1(n8683), .C2(n8685), .A(n8682), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8684) );
  OAI21_X1 U9820 ( .B1(n8686), .B2(n8685), .A(n8684), .ZN(P2_U3296) );
  INV_X1 U9821 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8689) );
  INV_X1 U9822 ( .A(n8687), .ZN(n9266) );
  OAI222_X1 U9823 ( .A1(n10406), .A2(n8689), .B1(n10404), .B2(n9266), .C1(
        P1_U3086), .C2(n8688), .ZN(P1_U3327) );
  OAI222_X1 U9824 ( .A1(P1_U3086), .A2(n8690), .B1(n10404), .B2(n8692), .C1(
        n8691), .C2(n10406), .ZN(P1_U3325) );
  NAND2_X1 U9825 ( .A1(n8694), .A2(n8695), .ZN(n8696) );
  XNOR2_X1 U9826 ( .A(n8698), .B(n8744), .ZN(n8700) );
  XOR2_X1 U9827 ( .A(n8896), .B(n8700), .Z(n8872) );
  INV_X1 U9828 ( .A(n8872), .ZN(n8699) );
  INV_X1 U9829 ( .A(n8700), .ZN(n8701) );
  NAND2_X1 U9830 ( .A1(n8701), .A2(n8896), .ZN(n8702) );
  NAND2_X1 U9831 ( .A1(n8874), .A2(n8702), .ZN(n8795) );
  XNOR2_X1 U9832 ( .A(n8801), .B(n8744), .ZN(n8703) );
  XNOR2_X1 U9833 ( .A(n8703), .B(n8895), .ZN(n8794) );
  NAND2_X1 U9834 ( .A1(n8795), .A2(n8794), .ZN(n8705) );
  NAND2_X1 U9835 ( .A1(n8705), .A2(n8704), .ZN(n8804) );
  XNOR2_X1 U9836 ( .A(n9206), .B(n8744), .ZN(n8805) );
  NOR2_X1 U9837 ( .A1(n8805), .A2(n9147), .ZN(n8707) );
  INV_X1 U9838 ( .A(n8805), .ZN(n8706) );
  OAI22_X1 U9839 ( .A1(n8804), .A2(n8707), .B1(n8706), .B2(n8894), .ZN(n8767)
         );
  INV_X1 U9840 ( .A(n8767), .ZN(n8710) );
  XNOR2_X1 U9841 ( .A(n8708), .B(n8744), .ZN(n8711) );
  XOR2_X1 U9842 ( .A(n8893), .B(n8711), .Z(n8841) );
  XNOR2_X1 U9843 ( .A(n8709), .B(n8744), .ZN(n8772) );
  INV_X1 U9844 ( .A(n8711), .ZN(n8712) );
  NAND2_X1 U9845 ( .A1(n8712), .A2(n8893), .ZN(n8768) );
  OR2_X1 U9846 ( .A1(n8713), .A2(n8768), .ZN(n8769) );
  NAND2_X1 U9847 ( .A1(n8713), .A2(n8892), .ZN(n8714) );
  XNOR2_X1 U9848 ( .A(n9194), .B(n8744), .ZN(n8719) );
  XOR2_X1 U9849 ( .A(n9103), .B(n8719), .Z(n8825) );
  XNOR2_X1 U9850 ( .A(n9236), .B(n8744), .ZN(n8716) );
  NAND2_X1 U9851 ( .A1(n8716), .A2(n9123), .ZN(n8720) );
  INV_X1 U9852 ( .A(n8720), .ZN(n8717) );
  XNOR2_X1 U9853 ( .A(n8716), .B(n9085), .ZN(n8780) );
  NOR2_X1 U9854 ( .A1(n8717), .A2(n8780), .ZN(n8722) );
  OR2_X1 U9855 ( .A1(n8825), .A2(n8722), .ZN(n8718) );
  NAND2_X1 U9856 ( .A1(n8719), .A2(n9136), .ZN(n8778) );
  AND2_X1 U9857 ( .A1(n8778), .A2(n8720), .ZN(n8721) );
  OR2_X1 U9858 ( .A1(n8722), .A2(n8721), .ZN(n8723) );
  XOR2_X1 U9859 ( .A(n8744), .B(n9184), .Z(n8725) );
  INV_X1 U9860 ( .A(n8725), .ZN(n8724) );
  XNOR2_X1 U9861 ( .A(n8724), .B(n9104), .ZN(n8832) );
  NOR2_X1 U9862 ( .A1(n8725), .A2(n9104), .ZN(n8726) );
  XNOR2_X1 U9863 ( .A(n8763), .B(n8744), .ZN(n8727) );
  XNOR2_X1 U9864 ( .A(n8729), .B(n8727), .ZN(n8759) );
  NAND2_X1 U9865 ( .A1(n8759), .A2(n9063), .ZN(n8731) );
  INV_X1 U9866 ( .A(n8727), .ZN(n8728) );
  NAND2_X1 U9867 ( .A1(n8731), .A2(n8730), .ZN(n8814) );
  XNOR2_X1 U9868 ( .A(n8819), .B(n6751), .ZN(n8732) );
  XNOR2_X1 U9869 ( .A(n8732), .B(n9051), .ZN(n8815) );
  NAND2_X1 U9870 ( .A1(n8814), .A2(n8815), .ZN(n8734) );
  NAND2_X1 U9871 ( .A1(n8732), .A2(n9076), .ZN(n8733) );
  XNOR2_X1 U9872 ( .A(n9171), .B(n8744), .ZN(n8735) );
  XNOR2_X1 U9873 ( .A(n8735), .B(n8891), .ZN(n8787) );
  NAND2_X1 U9874 ( .A1(n8786), .A2(n8787), .ZN(n8737) );
  NAND2_X1 U9875 ( .A1(n8735), .A2(n9064), .ZN(n8736) );
  NAND2_X1 U9876 ( .A1(n8737), .A2(n8736), .ZN(n8862) );
  XNOR2_X1 U9877 ( .A(n8868), .B(n6751), .ZN(n8738) );
  XNOR2_X1 U9878 ( .A(n8738), .B(n9052), .ZN(n8863) );
  XNOR2_X1 U9879 ( .A(n8740), .B(n8739), .ZN(n8741) );
  NAND2_X1 U9880 ( .A1(n8741), .A2(n8890), .ZN(n8742) );
  OAI21_X1 U9881 ( .B1(n8741), .B2(n8890), .A(n8742), .ZN(n8753) );
  XOR2_X1 U9882 ( .A(n8744), .B(n8743), .Z(n8745) );
  XNOR2_X1 U9883 ( .A(n8746), .B(n8745), .ZN(n8752) );
  NAND2_X1 U9884 ( .A1(n8888), .A2(n8876), .ZN(n8748) );
  AOI22_X1 U9885 ( .A1(n9025), .A2(n8880), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8747) );
  OAI211_X1 U9886 ( .C1(n9041), .C2(n8878), .A(n8748), .B(n8747), .ZN(n8749)
         );
  AOI21_X1 U9887 ( .B1(n8750), .B2(n8867), .A(n8749), .ZN(n8751) );
  OAI21_X1 U9888 ( .B1(n8752), .B2(n8870), .A(n8751), .ZN(P2_U3160) );
  AOI22_X1 U9889 ( .A1(n9033), .A2(n8880), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8755) );
  OAI21_X1 U9890 ( .B1(n8790), .B2(n8878), .A(n8755), .ZN(n8756) );
  AOI21_X1 U9891 ( .B1(n8889), .B2(n8876), .A(n8756), .ZN(n8757) );
  OAI211_X1 U9892 ( .C1(n5048), .C2(n8884), .A(n8758), .B(n8757), .ZN(P2_U3154) );
  XNOR2_X1 U9893 ( .A(n8759), .B(n9086), .ZN(n8765) );
  AOI22_X1 U9894 ( .A1(n9104), .A2(n8834), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8761) );
  NAND2_X1 U9895 ( .A1(n9079), .A2(n8880), .ZN(n8760) );
  OAI211_X1 U9896 ( .C1(n9076), .C2(n8837), .A(n8761), .B(n8760), .ZN(n8762)
         );
  AOI21_X1 U9897 ( .B1(n8763), .B2(n8867), .A(n8762), .ZN(n8764) );
  OAI21_X1 U9898 ( .B1(n8765), .B2(n8870), .A(n8764), .ZN(P2_U3156) );
  INV_X1 U9899 ( .A(n8766), .ZN(n9243) );
  NAND2_X1 U9900 ( .A1(n8842), .A2(n8768), .ZN(n8773) );
  AND2_X1 U9901 ( .A1(n8770), .A2(n8769), .ZN(n8771) );
  OAI211_X1 U9902 ( .C1(n8773), .C2(n8772), .A(n8771), .B(n8848), .ZN(n8777)
         );
  NOR2_X1 U9903 ( .A1(n9502), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9003) );
  AOI21_X1 U9904 ( .B1(n9103), .B2(n8876), .A(n9003), .ZN(n8774) );
  OAI21_X1 U9905 ( .B1(n9137), .B2(n8878), .A(n8774), .ZN(n8775) );
  AOI21_X1 U9906 ( .B1(n9140), .B2(n8880), .A(n8775), .ZN(n8776) );
  OAI211_X1 U9907 ( .C1(n9243), .C2(n8884), .A(n8777), .B(n8776), .ZN(P2_U3159) );
  OR2_X1 U9908 ( .A1(n8824), .A2(n8825), .ZN(n8822) );
  NAND2_X1 U9909 ( .A1(n8822), .A2(n8778), .ZN(n8779) );
  XOR2_X1 U9910 ( .A(n8780), .B(n8779), .Z(n8785) );
  AOI22_X1 U9911 ( .A1(n9104), .A2(n8876), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8782) );
  NAND2_X1 U9912 ( .A1(n9107), .A2(n8880), .ZN(n8781) );
  OAI211_X1 U9913 ( .C1(n9136), .C2(n8878), .A(n8782), .B(n8781), .ZN(n8783)
         );
  AOI21_X1 U9914 ( .B1(n9236), .B2(n8867), .A(n8783), .ZN(n8784) );
  OAI21_X1 U9915 ( .B1(n8785), .B2(n8870), .A(n8784), .ZN(P2_U3163) );
  XOR2_X1 U9916 ( .A(n8787), .B(n8786), .Z(n8793) );
  AOI22_X1 U9917 ( .A1(n9051), .A2(n8834), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8789) );
  NAND2_X1 U9918 ( .A1(n9056), .A2(n8880), .ZN(n8788) );
  OAI211_X1 U9919 ( .C1(n8790), .C2(n8837), .A(n8789), .B(n8788), .ZN(n8791)
         );
  AOI21_X1 U9920 ( .B1(n9171), .B2(n8867), .A(n8791), .ZN(n8792) );
  OAI21_X1 U9921 ( .B1(n8793), .B2(n8870), .A(n8792), .ZN(P2_U3165) );
  XNOR2_X1 U9922 ( .A(n8795), .B(n8794), .ZN(n8803) );
  INV_X1 U9923 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9399) );
  NOR2_X1 U9924 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9399), .ZN(n8943) );
  AOI21_X1 U9925 ( .B1(n8876), .B2(n8894), .A(n8943), .ZN(n8798) );
  NAND2_X1 U9926 ( .A1(n8880), .A2(n8796), .ZN(n8797) );
  OAI211_X1 U9927 ( .C1(n8799), .C2(n8878), .A(n8798), .B(n8797), .ZN(n8800)
         );
  AOI21_X1 U9928 ( .B1(n8801), .B2(n8867), .A(n8800), .ZN(n8802) );
  OAI21_X1 U9929 ( .B1(n8803), .B2(n8870), .A(n8802), .ZN(P2_U3166) );
  XNOR2_X1 U9930 ( .A(n8805), .B(n8894), .ZN(n8806) );
  XNOR2_X1 U9931 ( .A(n8804), .B(n8806), .ZN(n8813) );
  NOR2_X1 U9932 ( .A1(n9418), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8966) );
  AOI21_X1 U9933 ( .B1(n8876), .B2(n8893), .A(n8966), .ZN(n8809) );
  NAND2_X1 U9934 ( .A1(n8880), .A2(n8807), .ZN(n8808) );
  OAI211_X1 U9935 ( .C1(n8810), .C2(n8878), .A(n8809), .B(n8808), .ZN(n8811)
         );
  AOI21_X1 U9936 ( .B1(n9206), .B2(n8867), .A(n8811), .ZN(n8812) );
  OAI21_X1 U9937 ( .B1(n8813), .B2(n8870), .A(n8812), .ZN(P2_U3168) );
  XOR2_X1 U9938 ( .A(n8815), .B(n8814), .Z(n8821) );
  OAI22_X1 U9939 ( .A1(n9063), .A2(n8878), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9524), .ZN(n8816) );
  AOI21_X1 U9940 ( .B1(n9065), .B2(n8880), .A(n8816), .ZN(n8817) );
  OAI21_X1 U9941 ( .B1(n9064), .B2(n8837), .A(n8817), .ZN(n8818) );
  AOI21_X1 U9942 ( .B1(n8819), .B2(n8867), .A(n8818), .ZN(n8820) );
  OAI21_X1 U9943 ( .B1(n8821), .B2(n8870), .A(n8820), .ZN(P2_U3169) );
  INV_X1 U9944 ( .A(n8822), .ZN(n8823) );
  AOI21_X1 U9945 ( .B1(n8825), .B2(n8824), .A(n8823), .ZN(n8830) );
  AOI22_X1 U9946 ( .A1(n9085), .A2(n8876), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8827) );
  NAND2_X1 U9947 ( .A1(n8880), .A2(n9124), .ZN(n8826) );
  OAI211_X1 U9948 ( .C1(n9149), .C2(n8878), .A(n8827), .B(n8826), .ZN(n8828)
         );
  AOI21_X1 U9949 ( .B1(n9194), .B2(n8867), .A(n8828), .ZN(n8829) );
  OAI21_X1 U9950 ( .B1(n8830), .B2(n8870), .A(n8829), .ZN(P2_U3173) );
  XOR2_X1 U9951 ( .A(n8832), .B(n8831), .Z(n8840) );
  AOI22_X1 U9952 ( .A1(n9085), .A2(n8834), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8836) );
  NAND2_X1 U9953 ( .A1(n9090), .A2(n8880), .ZN(n8835) );
  OAI211_X1 U9954 ( .C1(n9063), .C2(n8837), .A(n8836), .B(n8835), .ZN(n8838)
         );
  AOI21_X1 U9955 ( .B1(n9184), .B2(n8867), .A(n8838), .ZN(n8839) );
  OAI21_X1 U9956 ( .B1(n8840), .B2(n8870), .A(n8839), .ZN(P2_U3175) );
  AOI21_X1 U9957 ( .B1(n8767), .B2(n8841), .A(n8870), .ZN(n8843) );
  NAND2_X1 U9958 ( .A1(n8843), .A2(n8842), .ZN(n8847) );
  INV_X1 U9959 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9536) );
  NOR2_X1 U9960 ( .A1(n9536), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8990) );
  AOI21_X1 U9961 ( .B1(n8876), .B2(n8892), .A(n8990), .ZN(n8844) );
  OAI21_X1 U9962 ( .B1(n9147), .B2(n8878), .A(n8844), .ZN(n8845) );
  AOI21_X1 U9963 ( .B1(n9155), .B2(n8880), .A(n8845), .ZN(n8846) );
  OAI211_X1 U9964 ( .C1(n9247), .C2(n8884), .A(n8847), .B(n8846), .ZN(P2_U3178) );
  OAI211_X1 U9965 ( .C1(n8851), .C2(n8850), .A(n8849), .B(n8848), .ZN(n8861)
         );
  NAND2_X1 U9966 ( .A1(n8876), .A2(n8902), .ZN(n8853) );
  OAI211_X1 U9967 ( .C1(n8854), .C2(n8878), .A(n8853), .B(n8852), .ZN(n8855)
         );
  INV_X1 U9968 ( .A(n8855), .ZN(n8860) );
  INV_X1 U9969 ( .A(n8856), .ZN(n8857) );
  NAND2_X1 U9970 ( .A1(n8880), .A2(n8857), .ZN(n8859) );
  NAND2_X1 U9971 ( .A1(n8867), .A2(n10670), .ZN(n8858) );
  NAND4_X1 U9972 ( .A1(n8861), .A2(n8860), .A3(n8859), .A4(n8858), .ZN(
        P2_U3179) );
  XOR2_X1 U9973 ( .A(n8863), .B(n8862), .Z(n8871) );
  NAND2_X1 U9974 ( .A1(n8890), .A2(n8876), .ZN(n8865) );
  AOI22_X1 U9975 ( .A1(n9044), .A2(n8880), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8864) );
  OAI211_X1 U9976 ( .C1(n9064), .C2(n8878), .A(n8865), .B(n8864), .ZN(n8866)
         );
  AOI21_X1 U9977 ( .B1(n8868), .B2(n8867), .A(n8866), .ZN(n8869) );
  OAI21_X1 U9978 ( .B1(n8871), .B2(n8870), .A(n8869), .ZN(P2_U3180) );
  AOI21_X1 U9979 ( .B1(n8873), .B2(n8872), .A(n8870), .ZN(n8875) );
  NAND2_X1 U9980 ( .A1(n8875), .A2(n8874), .ZN(n8883) );
  AND2_X1 U9981 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8918) );
  AOI21_X1 U9982 ( .B1(n8876), .B2(n8895), .A(n8918), .ZN(n8877) );
  OAI21_X1 U9983 ( .B1(n8695), .B2(n8878), .A(n8877), .ZN(n8879) );
  AOI21_X1 U9984 ( .B1(n8881), .B2(n8880), .A(n8879), .ZN(n8882) );
  OAI211_X1 U9985 ( .C1(n8885), .C2(n8884), .A(n8883), .B(n8882), .ZN(P2_U3181) );
  MUX2_X1 U9986 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8886), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9987 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8887), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9988 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8888), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9989 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8889), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9990 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8890), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9991 ( .A(n9052), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8989), .Z(
        P2_U3517) );
  MUX2_X1 U9992 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8891), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9993 ( .A(n9051), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8989), .Z(
        P2_U3515) );
  MUX2_X1 U9994 ( .A(n9104), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8989), .Z(
        P2_U3513) );
  MUX2_X1 U9995 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9085), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9996 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8892), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9997 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8893), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9998 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8894), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9999 ( .A(n8895), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8989), .Z(
        P2_U3507) );
  MUX2_X1 U10000 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8896), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10001 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8897), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U10002 ( .A(n8898), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8989), .Z(
        P2_U3503) );
  MUX2_X1 U10003 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8899), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10004 ( .A(n8900), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8989), .Z(
        P2_U3500) );
  MUX2_X1 U10005 ( .A(n8901), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8989), .Z(
        P2_U3499) );
  MUX2_X1 U10006 ( .A(n8902), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8989), .Z(
        P2_U3498) );
  MUX2_X1 U10007 ( .A(n8903), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8989), .Z(
        P2_U3497) );
  MUX2_X1 U10008 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n5079), .S(P2_U3893), .Z(
        P2_U3496) );
  MUX2_X1 U10009 ( .A(n8904), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8989), .Z(
        P2_U3495) );
  MUX2_X1 U10010 ( .A(n10609), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8989), .Z(
        P2_U3494) );
  MUX2_X1 U10011 ( .A(n8905), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8989), .Z(
        P2_U3493) );
  MUX2_X1 U10012 ( .A(n6754), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8989), .Z(
        P2_U3492) );
  MUX2_X1 U10013 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n6134), .S(P2_U3893), .Z(
        P2_U3491) );
  AOI21_X1 U10014 ( .B1(n5962), .B2(n8907), .A(n8928), .ZN(n8925) );
  NAND2_X1 U10015 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8911), .ZN(n8909) );
  NAND2_X1 U10016 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8910), .ZN(n8932) );
  OAI21_X1 U10017 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n8910), .A(n8932), .ZN(
        n8923) );
  INV_X1 U10018 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8921) );
  MUX2_X1 U10019 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8679), .Z(n8937) );
  XNOR2_X1 U10020 ( .A(n8937), .B(n8927), .ZN(n8916) );
  OR2_X1 U10021 ( .A1(n8912), .A2(n8911), .ZN(n8914) );
  NAND2_X1 U10022 ( .A1(n8914), .A2(n8913), .ZN(n8915) );
  NAND2_X1 U10023 ( .A1(n8916), .A2(n8915), .ZN(n8938) );
  OAI21_X1 U10024 ( .B1(n8916), .B2(n8915), .A(n8938), .ZN(n8919) );
  NOR2_X1 U10025 ( .A1(n10504), .A2(n8936), .ZN(n8917) );
  AOI211_X1 U10026 ( .C1(n8919), .C2(n10579), .A(n8918), .B(n8917), .ZN(n8920)
         );
  OAI21_X1 U10027 ( .B1(n10569), .B2(n8921), .A(n8920), .ZN(n8922) );
  AOI21_X1 U10028 ( .B1(n8923), .B2(n10580), .A(n8922), .ZN(n8924) );
  OAI21_X1 U10029 ( .B1(n8925), .B2(n10561), .A(n8924), .ZN(P2_U3197) );
  NOR2_X1 U10030 ( .A1(n8927), .A2(n8926), .ZN(n8929) );
  AOI22_X1 U10031 ( .A1(n8954), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n5978), .B2(
        n8958), .ZN(n8930) );
  AOI21_X1 U10032 ( .B1(n5026), .B2(n8930), .A(n8951), .ZN(n8950) );
  AOI22_X1 U10033 ( .A1(n8954), .A2(n9211), .B1(P2_REG1_REG_16__SCAN_IN), .B2(
        n8958), .ZN(n8935) );
  NAND2_X1 U10034 ( .A1(n8936), .A2(n8931), .ZN(n8933) );
  OAI21_X1 U10035 ( .B1(n8935), .B2(n8934), .A(n8953), .ZN(n8948) );
  INV_X1 U10036 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8946) );
  MUX2_X1 U10037 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8679), .Z(n8959) );
  XNOR2_X1 U10038 ( .A(n8954), .B(n8959), .ZN(n8941) );
  OR2_X1 U10039 ( .A1(n8937), .A2(n8936), .ZN(n8939) );
  NAND2_X1 U10040 ( .A1(n8939), .A2(n8938), .ZN(n8940) );
  NAND2_X1 U10041 ( .A1(n8941), .A2(n8940), .ZN(n8960) );
  OAI21_X1 U10042 ( .B1(n8941), .B2(n8940), .A(n8960), .ZN(n8944) );
  NOR2_X1 U10043 ( .A1(n10504), .A2(n8958), .ZN(n8942) );
  AOI211_X1 U10044 ( .C1(n8944), .C2(n10579), .A(n8943), .B(n8942), .ZN(n8945)
         );
  OAI21_X1 U10045 ( .B1(n10569), .B2(n8946), .A(n8945), .ZN(n8947) );
  AOI21_X1 U10046 ( .B1(n8948), .B2(n10580), .A(n8947), .ZN(n8949) );
  OAI21_X1 U10047 ( .B1(n8950), .B2(n10561), .A(n8949), .ZN(P2_U3198) );
  AOI21_X1 U10048 ( .B1(n8957), .B2(n8952), .A(n8977), .ZN(n8972) );
  NAND2_X1 U10049 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n8955), .ZN(n8975) );
  OAI21_X1 U10050 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8955), .A(n8975), .ZN(
        n8970) );
  INV_X1 U10051 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8956) );
  MUX2_X1 U10052 ( .A(n8957), .B(n8956), .S(n8679), .Z(n8983) );
  XNOR2_X1 U10053 ( .A(n8974), .B(n8983), .ZN(n8963) );
  OR2_X1 U10054 ( .A1(n8959), .A2(n8958), .ZN(n8961) );
  NAND2_X1 U10055 ( .A1(n8961), .A2(n8960), .ZN(n8962) );
  OAI21_X1 U10056 ( .B1(n8963), .B2(n8962), .A(n8982), .ZN(n8964) );
  INV_X1 U10057 ( .A(n8964), .ZN(n8968) );
  NOR2_X1 U10058 ( .A1(n10504), .A2(n8974), .ZN(n8965) );
  AOI211_X1 U10059 ( .C1(n10572), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n8966), .B(
        n8965), .ZN(n8967) );
  OAI21_X1 U10060 ( .B1(n8968), .B2(n10562), .A(n8967), .ZN(n8969) );
  AOI21_X1 U10061 ( .B1(n8970), .B2(n10580), .A(n8969), .ZN(n8971) );
  OAI21_X1 U10062 ( .B1(n8972), .B2(n10561), .A(n8971), .ZN(P2_U3199) );
  XNOR2_X1 U10063 ( .A(n8997), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n9007) );
  NAND2_X1 U10064 ( .A1(n8974), .A2(n8973), .ZN(n8976) );
  NAND2_X1 U10065 ( .A1(n8976), .A2(n8975), .ZN(n9008) );
  XOR2_X1 U10066 ( .A(n9007), .B(n9008), .Z(n8993) );
  MUX2_X1 U10067 ( .A(n8995), .B(P2_REG2_REG_18__SCAN_IN), .S(n8997), .Z(n8980) );
  NOR2_X1 U10068 ( .A1(n8984), .A2(n5019), .ZN(n8978) );
  OAI21_X1 U10069 ( .B1(n8980), .B2(n8979), .A(n8994), .ZN(n8981) );
  NAND2_X1 U10070 ( .A1(n8981), .A2(n10583), .ZN(n8992) );
  MUX2_X1 U10071 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8679), .Z(n8985) );
  INV_X1 U10072 ( .A(n8998), .ZN(n8987) );
  NAND2_X1 U10073 ( .A1(n8986), .A2(n8985), .ZN(n8996) );
  NAND2_X1 U10074 ( .A1(n8987), .A2(n8996), .ZN(n8988) );
  OAI211_X1 U10075 ( .C1(n10559), .C2(n8993), .A(n8992), .B(n8991), .ZN(
        P2_U3200) );
  MUX2_X1 U10076 ( .A(n6024), .B(P2_REG2_REG_19__SCAN_IN), .S(n9011), .Z(n9000) );
  OAI21_X1 U10077 ( .B1(n8998), .B2(n8997), .A(n8996), .ZN(n9002) );
  XNOR2_X1 U10078 ( .A(n9011), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n9009) );
  MUX2_X1 U10079 ( .A(n9009), .B(n9000), .S(n8999), .Z(n9001) );
  XNOR2_X1 U10080 ( .A(n9002), .B(n9001), .ZN(n9005) );
  AOI21_X1 U10081 ( .B1(n10572), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n9003), .ZN(
        n9004) );
  OAI21_X1 U10082 ( .B1(n10562), .B2(n9005), .A(n9004), .ZN(n9010) );
  NOR2_X1 U10083 ( .A1(n10626), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9013) );
  OAI22_X1 U10084 ( .A1(n9222), .A2(n9159), .B1(n9014), .B2(n9013), .ZN(
        P2_U3203) );
  NAND2_X1 U10085 ( .A1(n9015), .A2(n10626), .ZN(n9021) );
  NOR2_X1 U10086 ( .A1(n10626), .A2(n9016), .ZN(n9018) );
  AOI211_X1 U10087 ( .C1(n9019), .C2(n9111), .A(n9018), .B(n9017), .ZN(n9020)
         );
  OAI211_X1 U10088 ( .C1(n9023), .C2(n9022), .A(n9021), .B(n9020), .ZN(
        P2_U3204) );
  INV_X1 U10089 ( .A(n9024), .ZN(n9031) );
  AOI22_X1 U10090 ( .A1(n9025), .A2(n9156), .B1(n9157), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n9026) );
  OAI21_X1 U10091 ( .B1(n9027), .B2(n9159), .A(n9026), .ZN(n9028) );
  AOI21_X1 U10092 ( .B1(n9029), .B2(n9161), .A(n9028), .ZN(n9030) );
  OAI21_X1 U10093 ( .B1(n9031), .B2(n9163), .A(n9030), .ZN(P2_U3205) );
  INV_X1 U10094 ( .A(n9032), .ZN(n9038) );
  AOI22_X1 U10095 ( .A1(n9033), .A2(n9156), .B1(n9157), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n9034) );
  OAI21_X1 U10096 ( .B1(n5048), .B2(n9159), .A(n9034), .ZN(n9035) );
  AOI21_X1 U10097 ( .B1(n9036), .B2(n9161), .A(n9035), .ZN(n9037) );
  OAI21_X1 U10098 ( .B1(n9038), .B2(n9163), .A(n9037), .ZN(P2_U3206) );
  XOR2_X1 U10099 ( .A(n9043), .B(n9039), .Z(n9040) );
  OAI222_X1 U10100 ( .A1(n9148), .A2(n9064), .B1(n9150), .B2(n9041), .C1(n9145), .C2(n9040), .ZN(n9167) );
  INV_X1 U10101 ( .A(n9167), .ZN(n9048) );
  XOR2_X1 U10102 ( .A(n9043), .B(n9042), .Z(n9168) );
  AOI22_X1 U10103 ( .A1(n9044), .A2(n9156), .B1(n9157), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n9045) );
  OAI21_X1 U10104 ( .B1(n9226), .B2(n9159), .A(n9045), .ZN(n9046) );
  AOI21_X1 U10105 ( .B1(n9168), .B2(n9161), .A(n9046), .ZN(n9047) );
  OAI21_X1 U10106 ( .B1(n9048), .B2(n9163), .A(n9047), .ZN(P2_U3207) );
  NOR2_X1 U10107 ( .A1(n9049), .A2(n10617), .ZN(n9055) );
  XNOR2_X1 U10108 ( .A(n9050), .B(n5237), .ZN(n9053) );
  AOI222_X1 U10109 ( .A1(n10611), .A2(n9053), .B1(n9052), .B2(n10608), .C1(
        n9051), .C2(n10607), .ZN(n9174) );
  INV_X1 U10110 ( .A(n9174), .ZN(n9054) );
  AOI211_X1 U10111 ( .C1(n9156), .C2(n9056), .A(n9055), .B(n9054), .ZN(n9059)
         );
  XNOR2_X1 U10112 ( .A(n9057), .B(n5237), .ZN(n9172) );
  AOI22_X1 U10113 ( .A1(n9172), .A2(n9161), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n9163), .ZN(n9058) );
  OAI21_X1 U10114 ( .B1(n9059), .B2(n9163), .A(n9058), .ZN(P2_U3208) );
  AOI21_X1 U10115 ( .B1(n9061), .B2(n9060), .A(n5015), .ZN(n9062) );
  OAI222_X1 U10116 ( .A1(n9150), .A2(n9064), .B1(n9148), .B2(n9063), .C1(n9145), .C2(n9062), .ZN(n9175) );
  INV_X1 U10117 ( .A(n9065), .ZN(n9066) );
  OAI22_X1 U10118 ( .A1(n9179), .A2(n10617), .B1(n9066), .B2(n10620), .ZN(
        n9067) );
  OAI21_X1 U10119 ( .B1(n9175), .B2(n9067), .A(n10626), .ZN(n9071) );
  NAND2_X1 U10120 ( .A1(n9069), .A2(n5492), .ZN(n9176) );
  NAND3_X1 U10121 ( .A1(n9068), .A2(n9176), .A3(n9161), .ZN(n9070) );
  OAI211_X1 U10122 ( .C1(n10626), .C2(n9072), .A(n9071), .B(n9070), .ZN(
        P2_U3209) );
  XNOR2_X1 U10123 ( .A(n9073), .B(n9077), .ZN(n9074) );
  OAI222_X1 U10124 ( .A1(n9150), .A2(n9076), .B1(n9148), .B2(n9075), .C1(n9074), .C2(n9145), .ZN(n9180) );
  INV_X1 U10125 ( .A(n9180), .ZN(n9083) );
  XNOR2_X1 U10126 ( .A(n9078), .B(n9077), .ZN(n9181) );
  AOI22_X1 U10127 ( .A1(n9079), .A2(n9156), .B1(n9157), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n9080) );
  OAI21_X1 U10128 ( .B1(n9232), .B2(n9159), .A(n9080), .ZN(n9081) );
  AOI21_X1 U10129 ( .B1(n9181), .B2(n9161), .A(n9081), .ZN(n9082) );
  OAI21_X1 U10130 ( .B1(n9083), .B2(n9163), .A(n9082), .ZN(P2_U3210) );
  XOR2_X1 U10131 ( .A(n9089), .B(n9084), .Z(n9087) );
  AOI222_X1 U10132 ( .A1(n10611), .A2(n9087), .B1(n9086), .B2(n10608), .C1(
        n9085), .C2(n10607), .ZN(n9187) );
  XNOR2_X1 U10133 ( .A(n9088), .B(n9089), .ZN(n9185) );
  NAND2_X1 U10134 ( .A1(n9184), .A2(n9111), .ZN(n9092) );
  AOI22_X1 U10135 ( .A1(n9157), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9090), .B2(
        n9156), .ZN(n9091) );
  NAND2_X1 U10136 ( .A1(n9092), .A2(n9091), .ZN(n9093) );
  AOI21_X1 U10137 ( .B1(n9185), .B2(n9161), .A(n9093), .ZN(n9094) );
  OAI21_X1 U10138 ( .B1(n9187), .B2(n9163), .A(n9094), .ZN(P2_U3211) );
  NAND2_X1 U10139 ( .A1(n9096), .A2(n9095), .ZN(n9097) );
  NAND2_X1 U10140 ( .A1(n9098), .A2(n9097), .ZN(n9188) );
  AND3_X1 U10141 ( .A1(n9118), .A2(n9100), .A3(n9099), .ZN(n9101) );
  OAI21_X1 U10142 ( .B1(n9102), .B2(n9101), .A(n10611), .ZN(n9106) );
  AOI22_X1 U10143 ( .A1(n9104), .A2(n10608), .B1(n10607), .B2(n9103), .ZN(
        n9105) );
  NAND2_X1 U10144 ( .A1(n9106), .A2(n9105), .ZN(n9190) );
  NAND2_X1 U10145 ( .A1(n9190), .A2(n10626), .ZN(n9113) );
  INV_X1 U10146 ( .A(n9107), .ZN(n9109) );
  OAI22_X1 U10147 ( .A1(n9109), .A2(n10620), .B1(n10626), .B2(n9108), .ZN(
        n9110) );
  AOI21_X1 U10148 ( .B1(n9236), .B2(n9111), .A(n9110), .ZN(n9112) );
  OAI211_X1 U10149 ( .C1(n9188), .C2(n9129), .A(n9113), .B(n9112), .ZN(
        P2_U3212) );
  INV_X1 U10150 ( .A(n9114), .ZN(n9121) );
  XNOR2_X1 U10151 ( .A(n9115), .B(n9121), .ZN(n9196) );
  NAND2_X1 U10152 ( .A1(n9117), .A2(n9116), .ZN(n9120) );
  INV_X1 U10153 ( .A(n9118), .ZN(n9119) );
  AOI21_X1 U10154 ( .B1(n9121), .B2(n9120), .A(n9119), .ZN(n9122) );
  OAI222_X1 U10155 ( .A1(n9150), .A2(n9123), .B1(n9148), .B2(n9149), .C1(n9145), .C2(n9122), .ZN(n9193) );
  INV_X1 U10156 ( .A(n9194), .ZN(n9126) );
  AOI22_X1 U10157 ( .A1(n9157), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9156), .B2(
        n9124), .ZN(n9125) );
  OAI21_X1 U10158 ( .B1(n9126), .B2(n9159), .A(n9125), .ZN(n9127) );
  AOI21_X1 U10159 ( .B1(n9193), .B2(n10626), .A(n9127), .ZN(n9128) );
  OAI21_X1 U10160 ( .B1(n9196), .B2(n9129), .A(n9128), .ZN(P2_U3213) );
  NAND2_X1 U10161 ( .A1(n9130), .A2(n9131), .ZN(n9133) );
  NAND2_X1 U10162 ( .A1(n9133), .A2(n9132), .ZN(n9134) );
  XNOR2_X1 U10163 ( .A(n9134), .B(n9138), .ZN(n9135) );
  OAI222_X1 U10164 ( .A1(n9148), .A2(n9137), .B1(n9150), .B2(n9136), .C1(n9145), .C2(n9135), .ZN(n9197) );
  INV_X1 U10165 ( .A(n9197), .ZN(n9144) );
  XNOR2_X1 U10166 ( .A(n9139), .B(n9138), .ZN(n9198) );
  AOI22_X1 U10167 ( .A1(n9157), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n9156), .B2(
        n9140), .ZN(n9141) );
  OAI21_X1 U10168 ( .B1(n9243), .B2(n9159), .A(n9141), .ZN(n9142) );
  AOI21_X1 U10169 ( .B1(n9198), .B2(n9161), .A(n9142), .ZN(n9143) );
  OAI21_X1 U10170 ( .B1(n9144), .B2(n9163), .A(n9143), .ZN(P2_U3214) );
  XNOR2_X1 U10171 ( .A(n9130), .B(n9154), .ZN(n9146) );
  OAI222_X1 U10172 ( .A1(n9150), .A2(n9149), .B1(n9148), .B2(n9147), .C1(n9146), .C2(n9145), .ZN(n9201) );
  INV_X1 U10173 ( .A(n9201), .ZN(n9164) );
  INV_X1 U10174 ( .A(n9151), .ZN(n9152) );
  AOI21_X1 U10175 ( .B1(n9154), .B2(n9153), .A(n9152), .ZN(n9202) );
  AOI22_X1 U10176 ( .A1(n9157), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9156), .B2(
        n9155), .ZN(n9158) );
  OAI21_X1 U10177 ( .B1(n9247), .B2(n9159), .A(n9158), .ZN(n9160) );
  AOI21_X1 U10178 ( .B1(n9202), .B2(n9161), .A(n9160), .ZN(n9162) );
  OAI21_X1 U10179 ( .B1(n9164), .B2(n9163), .A(n9162), .ZN(P2_U3215) );
  AOI21_X1 U10180 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n10780), .A(n9165), .ZN(
        n9166) );
  OAI21_X1 U10181 ( .B1(n9222), .B2(n9213), .A(n9166), .ZN(P2_U3489) );
  INV_X1 U10182 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9169) );
  AOI21_X1 U10183 ( .B1(n9168), .B2(n10632), .A(n9167), .ZN(n9223) );
  MUX2_X1 U10184 ( .A(n9169), .B(n9223), .S(n10781), .Z(n9170) );
  OAI21_X1 U10185 ( .B1(n9226), .B2(n9213), .A(n9170), .ZN(P2_U3485) );
  AOI22_X1 U10186 ( .A1(n9172), .A2(n10632), .B1(n10779), .B2(n9171), .ZN(
        n9173) );
  NAND2_X1 U10187 ( .A1(n9174), .A2(n9173), .ZN(n9227) );
  MUX2_X1 U10188 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9227), .S(n10781), .Z(
        P2_U3484) );
  INV_X1 U10189 ( .A(n9175), .ZN(n9178) );
  NAND3_X1 U10190 ( .A1(n9068), .A2(n9176), .A3(n10632), .ZN(n9177) );
  OAI211_X1 U10191 ( .C1(n9179), .C2(n10650), .A(n9178), .B(n9177), .ZN(n9228)
         );
  MUX2_X1 U10192 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9228), .S(n10781), .Z(
        P2_U3483) );
  INV_X1 U10193 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9182) );
  AOI21_X1 U10194 ( .B1(n10632), .B2(n9181), .A(n9180), .ZN(n9229) );
  MUX2_X1 U10195 ( .A(n9182), .B(n9229), .S(n10781), .Z(n9183) );
  OAI21_X1 U10196 ( .B1(n9232), .B2(n9213), .A(n9183), .ZN(P2_U3482) );
  AOI22_X1 U10197 ( .A1(n9185), .A2(n10632), .B1(n10779), .B2(n9184), .ZN(
        n9186) );
  NAND2_X1 U10198 ( .A1(n9187), .A2(n9186), .ZN(n9233) );
  MUX2_X1 U10199 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9233), .S(n10781), .Z(
        P2_U3481) );
  INV_X1 U10200 ( .A(n10632), .ZN(n10774) );
  NOR2_X1 U10201 ( .A1(n9188), .A2(n10774), .ZN(n9189) );
  OR2_X1 U10202 ( .A1(n9190), .A2(n9189), .ZN(n9234) );
  MUX2_X1 U10203 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9234), .S(n10781), .Z(
        n9191) );
  AOI21_X1 U10204 ( .B1(n6290), .B2(n9236), .A(n9191), .ZN(n9192) );
  INV_X1 U10205 ( .A(n9192), .ZN(P2_U3480) );
  AOI21_X1 U10206 ( .B1(n10779), .B2(n9194), .A(n9193), .ZN(n9195) );
  OAI21_X1 U10207 ( .B1(n10774), .B2(n9196), .A(n9195), .ZN(n9239) );
  MUX2_X1 U10208 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9239), .S(n10781), .Z(
        P2_U3479) );
  INV_X1 U10209 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9199) );
  AOI21_X1 U10210 ( .B1(n9198), .B2(n10632), .A(n9197), .ZN(n9240) );
  MUX2_X1 U10211 ( .A(n9199), .B(n9240), .S(n10781), .Z(n9200) );
  OAI21_X1 U10212 ( .B1(n9243), .B2(n9213), .A(n9200), .ZN(P2_U3478) );
  INV_X1 U10213 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9203) );
  AOI21_X1 U10214 ( .B1(n9202), .B2(n10632), .A(n9201), .ZN(n9244) );
  MUX2_X1 U10215 ( .A(n9203), .B(n9244), .S(n10781), .Z(n9204) );
  OAI21_X1 U10216 ( .B1(n9247), .B2(n9213), .A(n9204), .ZN(P2_U3477) );
  AOI21_X1 U10217 ( .B1(n10779), .B2(n9206), .A(n9205), .ZN(n9207) );
  OAI21_X1 U10218 ( .B1(n10774), .B2(n9208), .A(n9207), .ZN(n9248) );
  MUX2_X1 U10219 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9248), .S(n10781), .Z(
        P2_U3476) );
  AOI21_X1 U10220 ( .B1(n9210), .B2(n10632), .A(n9209), .ZN(n9249) );
  MUX2_X1 U10221 ( .A(n9211), .B(n9249), .S(n10781), .Z(n9212) );
  OAI21_X1 U10222 ( .B1(n9253), .B2(n9213), .A(n9212), .ZN(P2_U3475) );
  INV_X1 U10223 ( .A(n9214), .ZN(n9217) );
  OAI211_X1 U10224 ( .C1(n10774), .C2(n9217), .A(n9216), .B(n9215), .ZN(n9254)
         );
  MUX2_X1 U10225 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9254), .S(n10781), .Z(
        P2_U3472) );
  MUX2_X1 U10226 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n9218), .S(n10781), .Z(
        P2_U3459) );
  AOI21_X1 U10227 ( .B1(n10782), .B2(P2_REG0_REG_30__SCAN_IN), .A(n9219), .ZN(
        n9220) );
  OAI21_X1 U10228 ( .B1(n9222), .B2(n9221), .A(n9220), .ZN(P2_U3457) );
  INV_X1 U10229 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9224) );
  MUX2_X1 U10230 ( .A(n9224), .B(n9223), .S(n10785), .Z(n9225) );
  OAI21_X1 U10231 ( .B1(n9226), .B2(n9252), .A(n9225), .ZN(P2_U3453) );
  MUX2_X1 U10232 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9227), .S(n10785), .Z(
        P2_U3452) );
  MUX2_X1 U10233 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9228), .S(n10785), .Z(
        P2_U3451) );
  INV_X1 U10234 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9230) );
  MUX2_X1 U10235 ( .A(n9230), .B(n9229), .S(n10785), .Z(n9231) );
  OAI21_X1 U10236 ( .B1(n9232), .B2(n9252), .A(n9231), .ZN(P2_U3450) );
  MUX2_X1 U10237 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9233), .S(n10785), .Z(
        P2_U3449) );
  MUX2_X1 U10238 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9234), .S(n10785), .Z(
        n9235) );
  AOI21_X1 U10239 ( .B1(n9237), .B2(n9236), .A(n9235), .ZN(n9238) );
  INV_X1 U10240 ( .A(n9238), .ZN(P2_U3448) );
  MUX2_X1 U10241 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9239), .S(n10785), .Z(
        P2_U3447) );
  INV_X1 U10242 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9241) );
  MUX2_X1 U10243 ( .A(n9241), .B(n9240), .S(n10785), .Z(n9242) );
  OAI21_X1 U10244 ( .B1(n9243), .B2(n9252), .A(n9242), .ZN(P2_U3446) );
  INV_X1 U10245 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9245) );
  MUX2_X1 U10246 ( .A(n9245), .B(n9244), .S(n10785), .Z(n9246) );
  OAI21_X1 U10247 ( .B1(n9247), .B2(n9252), .A(n9246), .ZN(P2_U3444) );
  MUX2_X1 U10248 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9248), .S(n10785), .Z(
        P2_U3441) );
  INV_X1 U10249 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9250) );
  MUX2_X1 U10250 ( .A(n9250), .B(n9249), .S(n10785), .Z(n9251) );
  OAI21_X1 U10251 ( .B1(n9253), .B2(n9252), .A(n9251), .ZN(P2_U3438) );
  MUX2_X1 U10252 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n9254), .S(n10785), .Z(
        P2_U3429) );
  INV_X1 U10253 ( .A(n9662), .ZN(n10401) );
  NAND3_X1 U10254 ( .A1(n9256), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n9257) );
  OAI22_X1 U10255 ( .A1(n9255), .A2(n9257), .B1(n6436), .B2(n8472), .ZN(n9258)
         );
  INV_X1 U10256 ( .A(n9258), .ZN(n9259) );
  OAI21_X1 U10257 ( .B1(n10401), .B2(n4944), .A(n9259), .ZN(P2_U3264) );
  INV_X1 U10258 ( .A(n9664), .ZN(n10403) );
  OAI222_X1 U10259 ( .A1(n4944), .A2(n10403), .B1(n9262), .B2(P2_U3151), .C1(
        n9260), .C2(n8472), .ZN(P2_U3266) );
  AOI21_X1 U10260 ( .B1(n9264), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n9263), .ZN(
        n9265) );
  OAI21_X1 U10261 ( .B1(n9266), .B2(n4944), .A(n9265), .ZN(P2_U3267) );
  MUX2_X1 U10262 ( .A(n9267), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10263 ( .A(n9268), .ZN(n9273) );
  AOI21_X1 U10264 ( .B1(n9269), .B2(n9271), .A(n9270), .ZN(n9272) );
  OAI21_X1 U10265 ( .B1(n9273), .B2(n9272), .A(n9651), .ZN(n9279) );
  OAI22_X1 U10266 ( .A1(n9639), .A2(n10305), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9274), .ZN(n9277) );
  OAI22_X1 U10267 ( .A1(n9654), .A2(n9275), .B1(n10288), .B2(n9655), .ZN(n9276) );
  AOI211_X1 U10268 ( .C1(n10291), .C2(n9642), .A(n9277), .B(n9276), .ZN(n9278)
         );
  NAND2_X1 U10269 ( .A1(n9279), .A2(n9278), .ZN(P1_U3214) );
  INV_X1 U10270 ( .A(n8356), .ZN(n9281) );
  NOR2_X1 U10271 ( .A1(n9281), .A2(n9280), .ZN(n9285) );
  XNOR2_X1 U10272 ( .A(n9283), .B(n9282), .ZN(n9284) );
  XNOR2_X1 U10273 ( .A(n9285), .B(n9284), .ZN(n9286) );
  NAND2_X1 U10274 ( .A1(n9286), .A2(n9651), .ZN(n9291) );
  INV_X1 U10275 ( .A(n9287), .ZN(n9289) );
  OAI22_X1 U10276 ( .A1(n9639), .A2(n10826), .B1(n9654), .B2(n10848), .ZN(
        n9288) );
  AOI211_X1 U10277 ( .C1(n9582), .C2(n9957), .A(n9289), .B(n9288), .ZN(n9290)
         );
  OAI211_X1 U10278 ( .C1(n10846), .C2(n9661), .A(n9291), .B(n9290), .ZN(
        P1_U3215) );
  INV_X1 U10279 ( .A(n10321), .ZN(n10163) );
  OR2_X1 U10280 ( .A1(n9296), .A2(n9295), .ZN(n9615) );
  NAND2_X1 U10281 ( .A1(n9615), .A2(n9617), .ZN(n9298) );
  INV_X1 U10282 ( .A(n9292), .ZN(n9294) );
  AND2_X1 U10283 ( .A1(n9294), .A2(n9293), .ZN(n9297) );
  NAND2_X1 U10284 ( .A1(n9296), .A2(n9295), .ZN(n9614) );
  NAND3_X1 U10285 ( .A1(n9298), .A2(n9297), .A3(n9614), .ZN(n9598) );
  INV_X1 U10286 ( .A(n9598), .ZN(n9300) );
  AOI21_X1 U10287 ( .B1(n9298), .B2(n9614), .A(n9297), .ZN(n9299) );
  OAI21_X1 U10288 ( .B1(n9300), .B2(n9299), .A(n9651), .ZN(n9304) );
  NOR2_X1 U10289 ( .A1(n9655), .A2(n10318), .ZN(n9302) );
  OAI22_X1 U10290 ( .A1(n9639), .A2(n10336), .B1(n9654), .B2(n10157), .ZN(
        n9301) );
  AOI211_X1 U10291 ( .C1(P1_REG3_REG_23__SCAN_IN), .C2(P1_U3086), .A(n9302), 
        .B(n9301), .ZN(n9303) );
  OAI211_X1 U10292 ( .C1(n10163), .C2(n9661), .A(n9304), .B(n9303), .ZN(
        P1_U3216) );
  AND2_X1 U10293 ( .A1(n9306), .A2(n9305), .ZN(n9307) );
  OAI21_X1 U10294 ( .B1(n9308), .B2(n9307), .A(n8002), .ZN(n9309) );
  NAND2_X1 U10295 ( .A1(n9309), .A2(n9651), .ZN(n9315) );
  INV_X1 U10296 ( .A(n9310), .ZN(n9313) );
  OAI22_X1 U10297 ( .A1(n9639), .A2(n10757), .B1(n9654), .B2(n9311), .ZN(n9312) );
  AOI211_X1 U10298 ( .C1(n9582), .C2(n9959), .A(n9313), .B(n9312), .ZN(n9314)
         );
  OAI211_X1 U10299 ( .C1(n5394), .C2(n9661), .A(n9315), .B(n9314), .ZN(
        P1_U3217) );
  INV_X1 U10300 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9316) );
  OAI22_X1 U10301 ( .A1(n9316), .A2(keyinput_62), .B1(keyinput_61), .B2(
        P2_REG3_REG_6__SCAN_IN), .ZN(n9319) );
  INV_X1 U10302 ( .A(keyinput_62), .ZN(n9317) );
  NOR2_X1 U10303 ( .A1(n9317), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n9318) );
  AOI211_X1 U10304 ( .C1(P2_REG3_REG_6__SCAN_IN), .C2(keyinput_61), .A(n9319), 
        .B(n9318), .ZN(n9548) );
  OAI22_X1 U10305 ( .A1(n6893), .A2(keyinput_54), .B1(keyinput_55), .B2(
        P2_REG3_REG_20__SCAN_IN), .ZN(n9320) );
  AOI221_X1 U10306 ( .B1(n6893), .B2(keyinput_54), .C1(P2_REG3_REG_20__SCAN_IN), .C2(keyinput_55), .A(n9320), .ZN(n9408) );
  OAI22_X1 U10307 ( .A1(n5678), .A2(keyinput_49), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(keyinput_50), .ZN(n9321) );
  AOI221_X1 U10308 ( .B1(n5678), .B2(keyinput_49), .C1(keyinput_50), .C2(
        P2_REG3_REG_17__SCAN_IN), .A(n9321), .ZN(n9397) );
  INV_X1 U10309 ( .A(keyinput_47), .ZN(n9395) );
  INV_X1 U10310 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9517) );
  INV_X1 U10311 ( .A(keyinput_46), .ZN(n9393) );
  INV_X1 U10312 ( .A(keyinput_42), .ZN(n9385) );
  INV_X1 U10313 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9506) );
  INV_X1 U10314 ( .A(keyinput_41), .ZN(n9383) );
  INV_X1 U10315 ( .A(keyinput_40), .ZN(n9381) );
  AOI22_X1 U10316 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_37), .B1(
        P2_REG3_REG_23__SCAN_IN), .B2(keyinput_38), .ZN(n9322) );
  OAI221_X1 U10317 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_37), .C1(
        P2_REG3_REG_23__SCAN_IN), .C2(keyinput_38), .A(n9322), .ZN(n9378) );
  INV_X1 U10318 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9376) );
  OAI22_X1 U10319 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_34), .B1(
        keyinput_35), .B2(P2_REG3_REG_7__SCAN_IN), .ZN(n9323) );
  AOI221_X1 U10320 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_34), .C1(
        P2_REG3_REG_7__SCAN_IN), .C2(keyinput_35), .A(n9323), .ZN(n9374) );
  INV_X1 U10321 ( .A(keyinput_23), .ZN(n9358) );
  INV_X1 U10322 ( .A(SI_12_), .ZN(n9423) );
  OAI22_X1 U10323 ( .A1(n9423), .A2(keyinput_20), .B1(keyinput_21), .B2(SI_11_), .ZN(n9324) );
  AOI221_X1 U10324 ( .B1(n9423), .B2(keyinput_20), .C1(SI_11_), .C2(
        keyinput_21), .A(n9324), .ZN(n9354) );
  INV_X1 U10325 ( .A(keyinput_12), .ZN(n9343) );
  INV_X1 U10326 ( .A(SI_21_), .ZN(n9457) );
  INV_X1 U10327 ( .A(keyinput_11), .ZN(n9341) );
  INV_X1 U10328 ( .A(keyinput_10), .ZN(n9339) );
  OAI22_X1 U10329 ( .A1(n9451), .A2(keyinput_7), .B1(n9446), .B2(keyinput_8), 
        .ZN(n9325) );
  AOI221_X1 U10330 ( .B1(n9451), .B2(keyinput_7), .C1(keyinput_8), .C2(n9446), 
        .A(n9325), .ZN(n9336) );
  INV_X1 U10331 ( .A(keyinput_6), .ZN(n9334) );
  INV_X1 U10332 ( .A(keyinput_5), .ZN(n9332) );
  INV_X1 U10333 ( .A(SI_29_), .ZN(n9432) );
  OAI22_X1 U10334 ( .A1(n9432), .A2(keyinput_3), .B1(n9433), .B2(keyinput_2), 
        .ZN(n9326) );
  AOI221_X1 U10335 ( .B1(n9432), .B2(keyinput_3), .C1(keyinput_2), .C2(n9433), 
        .A(n9326), .ZN(n9329) );
  AOI22_X1 U10336 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_0), .B1(SI_31_), .B2(
        keyinput_1), .ZN(n9327) );
  OAI221_X1 U10337 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_0), .C1(SI_31_), 
        .C2(keyinput_1), .A(n9327), .ZN(n9328) );
  AOI22_X1 U10338 ( .A1(keyinput_4), .A2(n9438), .B1(n9329), .B2(n9328), .ZN(
        n9330) );
  OAI21_X1 U10339 ( .B1(n9438), .B2(keyinput_4), .A(n9330), .ZN(n9331) );
  OAI221_X1 U10340 ( .B1(SI_27_), .B2(n9332), .C1(n9440), .C2(keyinput_5), .A(
        n9331), .ZN(n9333) );
  OAI221_X1 U10341 ( .B1(SI_26_), .B2(n9334), .C1(n9444), .C2(keyinput_6), .A(
        n9333), .ZN(n9335) );
  OAI211_X1 U10342 ( .C1(SI_23_), .C2(keyinput_9), .A(n9336), .B(n9335), .ZN(
        n9337) );
  AOI21_X1 U10343 ( .B1(SI_23_), .B2(keyinput_9), .A(n9337), .ZN(n9338) );
  AOI221_X1 U10344 ( .B1(SI_22_), .B2(keyinput_10), .C1(n9453), .C2(n9339), 
        .A(n9338), .ZN(n9340) );
  AOI221_X1 U10345 ( .B1(SI_21_), .B2(keyinput_11), .C1(n9457), .C2(n9341), 
        .A(n9340), .ZN(n9342) );
  AOI221_X1 U10346 ( .B1(SI_20_), .B2(n9343), .C1(n9459), .C2(keyinput_12), 
        .A(n9342), .ZN(n9348) );
  AOI22_X1 U10347 ( .A1(n9427), .A2(keyinput_16), .B1(n9428), .B2(keyinput_14), 
        .ZN(n9344) );
  OAI221_X1 U10348 ( .B1(n9427), .B2(keyinput_16), .C1(n9428), .C2(keyinput_14), .A(n9344), .ZN(n9347) );
  AOI22_X1 U10349 ( .A1(SI_17_), .A2(keyinput_15), .B1(SI_19_), .B2(
        keyinput_13), .ZN(n9345) );
  OAI221_X1 U10350 ( .B1(SI_17_), .B2(keyinput_15), .C1(SI_19_), .C2(
        keyinput_13), .A(n9345), .ZN(n9346) );
  NOR3_X1 U10351 ( .A1(n9348), .A2(n9347), .A3(n9346), .ZN(n9351) );
  AOI22_X1 U10352 ( .A1(SI_15_), .A2(keyinput_17), .B1(n9425), .B2(keyinput_18), .ZN(n9349) );
  OAI221_X1 U10353 ( .B1(SI_15_), .B2(keyinput_17), .C1(n9425), .C2(
        keyinput_18), .A(n9349), .ZN(n9350) );
  AOI211_X1 U10354 ( .C1(n9467), .C2(keyinput_19), .A(n9351), .B(n9350), .ZN(
        n9352) );
  OAI21_X1 U10355 ( .B1(n9467), .B2(keyinput_19), .A(n9352), .ZN(n9353) );
  AOI22_X1 U10356 ( .A1(keyinput_22), .A2(n9356), .B1(n9354), .B2(n9353), .ZN(
        n9355) );
  OAI21_X1 U10357 ( .B1(n9356), .B2(keyinput_22), .A(n9355), .ZN(n9357) );
  OAI221_X1 U10358 ( .B1(SI_9_), .B2(keyinput_23), .C1(n9472), .C2(n9358), .A(
        n9357), .ZN(n9366) );
  OAI22_X1 U10359 ( .A1(n9475), .A2(keyinput_24), .B1(n9476), .B2(keyinput_25), 
        .ZN(n9359) );
  AOI221_X1 U10360 ( .B1(n9475), .B2(keyinput_24), .C1(keyinput_25), .C2(n9476), .A(n9359), .ZN(n9365) );
  AOI22_X1 U10361 ( .A1(SI_5_), .A2(keyinput_27), .B1(SI_6_), .B2(keyinput_26), 
        .ZN(n9360) );
  OAI221_X1 U10362 ( .B1(SI_5_), .B2(keyinput_27), .C1(SI_6_), .C2(keyinput_26), .A(n9360), .ZN(n9364) );
  XNOR2_X1 U10363 ( .A(SI_3_), .B(keyinput_29), .ZN(n9362) );
  XNOR2_X1 U10364 ( .A(SI_4_), .B(keyinput_28), .ZN(n9361) );
  NAND2_X1 U10365 ( .A1(n9362), .A2(n9361), .ZN(n9363) );
  AOI211_X1 U10366 ( .C1(n9366), .C2(n9365), .A(n9364), .B(n9363), .ZN(n9372)
         );
  XNOR2_X1 U10367 ( .A(SI_2_), .B(keyinput_30), .ZN(n9368) );
  XNOR2_X1 U10368 ( .A(SI_1_), .B(keyinput_31), .ZN(n9367) );
  NAND2_X1 U10369 ( .A1(n9368), .A2(n9367), .ZN(n9371) );
  OAI22_X1 U10370 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput_33), .B1(keyinput_32), 
        .B2(SI_0_), .ZN(n9369) );
  AOI221_X1 U10371 ( .B1(P2_RD_REG_SCAN_IN), .B2(keyinput_33), .C1(SI_0_), 
        .C2(keyinput_32), .A(n9369), .ZN(n9370) );
  OAI21_X1 U10372 ( .B1(n9372), .B2(n9371), .A(n9370), .ZN(n9373) );
  AOI22_X1 U10373 ( .A1(n9374), .A2(n9373), .B1(keyinput_36), .B2(n9376), .ZN(
        n9375) );
  OAI21_X1 U10374 ( .B1(keyinput_36), .B2(n9376), .A(n9375), .ZN(n9377) );
  OAI22_X1 U10375 ( .A1(n9378), .A2(n9377), .B1(keyinput_39), .B2(
        P2_REG3_REG_10__SCAN_IN), .ZN(n9379) );
  AOI21_X1 U10376 ( .B1(keyinput_39), .B2(P2_REG3_REG_10__SCAN_IN), .A(n9379), 
        .ZN(n9380) );
  AOI221_X1 U10377 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n9381), .C1(n9500), .C2(
        keyinput_40), .A(n9380), .ZN(n9382) );
  AOI221_X1 U10378 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(n9383), .C1(n9502), 
        .C2(keyinput_41), .A(n9382), .ZN(n9384) );
  AOI221_X1 U10379 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(n9385), .C1(n9506), 
        .C2(keyinput_42), .A(n9384), .ZN(n9390) );
  XNOR2_X1 U10380 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_44), .ZN(n9388) );
  XNOR2_X1 U10381 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_43), .ZN(n9387) );
  NAND2_X1 U10382 ( .A1(keyinput_45), .A2(n5689), .ZN(n9386) );
  NAND3_X1 U10383 ( .A1(n9388), .A2(n9387), .A3(n9386), .ZN(n9389) );
  NOR2_X1 U10384 ( .A1(n9390), .A2(n9389), .ZN(n9391) );
  OAI21_X1 U10385 ( .B1(n5689), .B2(keyinput_45), .A(n9391), .ZN(n9392) );
  OAI221_X1 U10386 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(n9393), .C1(n9515), 
        .C2(keyinput_46), .A(n9392), .ZN(n9394) );
  OAI221_X1 U10387 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(n9395), .C1(n9517), 
        .C2(keyinput_47), .A(n9394), .ZN(n9396) );
  OAI211_X1 U10388 ( .C1(n9399), .C2(keyinput_48), .A(n9397), .B(n9396), .ZN(
        n9398) );
  AOI21_X1 U10389 ( .B1(n9399), .B2(keyinput_48), .A(n9398), .ZN(n9402) );
  AOI22_X1 U10390 ( .A1(n5682), .A2(keyinput_53), .B1(keyinput_52), .B2(n9523), 
        .ZN(n9400) );
  OAI221_X1 U10391 ( .B1(n5682), .B2(keyinput_53), .C1(n9523), .C2(keyinput_52), .A(n9400), .ZN(n9401) );
  AOI211_X1 U10392 ( .C1(P2_REG3_REG_24__SCAN_IN), .C2(keyinput_51), .A(n9402), 
        .B(n9401), .ZN(n9403) );
  OAI21_X1 U10393 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_51), .A(n9403), 
        .ZN(n9407) );
  INV_X1 U10394 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9405) );
  AOI22_X1 U10395 ( .A1(n9405), .A2(keyinput_57), .B1(keyinput_56), .B2(n5684), 
        .ZN(n9404) );
  OAI221_X1 U10396 ( .B1(n9405), .B2(keyinput_57), .C1(n5684), .C2(keyinput_56), .A(n9404), .ZN(n9406) );
  AOI21_X1 U10397 ( .B1(n9408), .B2(n9407), .A(n9406), .ZN(n9414) );
  XOR2_X1 U10398 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_58), .Z(n9413) );
  INV_X1 U10399 ( .A(keyinput_60), .ZN(n9411) );
  AOI22_X1 U10400 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_59), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_60), .ZN(n9409) );
  OAI21_X1 U10401 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_59), .A(n9409), 
        .ZN(n9410) );
  AOI21_X1 U10402 ( .B1(n9536), .B2(n9411), .A(n9410), .ZN(n9412) );
  OAI21_X1 U10403 ( .B1(n9414), .B2(n9413), .A(n9412), .ZN(n9547) );
  INV_X1 U10404 ( .A(keyinput_122), .ZN(n9534) );
  INV_X1 U10405 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9416) );
  OAI22_X1 U10406 ( .A1(n9416), .A2(keyinput_119), .B1(n6893), .B2(
        keyinput_118), .ZN(n9415) );
  AOI221_X1 U10407 ( .B1(n9416), .B2(keyinput_119), .C1(keyinput_118), .C2(
        n6893), .A(n9415), .ZN(n9531) );
  OAI22_X1 U10408 ( .A1(n9418), .A2(keyinput_114), .B1(keyinput_112), .B2(
        P2_REG3_REG_16__SCAN_IN), .ZN(n9417) );
  AOI221_X1 U10409 ( .B1(n9418), .B2(keyinput_114), .C1(
        P2_REG3_REG_16__SCAN_IN), .C2(keyinput_112), .A(n9417), .ZN(n9520) );
  INV_X1 U10410 ( .A(keyinput_111), .ZN(n9518) );
  INV_X1 U10411 ( .A(keyinput_110), .ZN(n9514) );
  INV_X1 U10412 ( .A(keyinput_106), .ZN(n9505) );
  INV_X1 U10413 ( .A(keyinput_105), .ZN(n9503) );
  INV_X1 U10414 ( .A(keyinput_104), .ZN(n9499) );
  INV_X1 U10415 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9420) );
  AOI22_X1 U10416 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_101), .B1(n9420), .B2(keyinput_102), .ZN(n9419) );
  OAI221_X1 U10417 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_101), .C1(
        n9420), .C2(keyinput_102), .A(n9419), .ZN(n9496) );
  AOI22_X1 U10418 ( .A1(n5680), .A2(keyinput_99), .B1(P2_U3151), .B2(
        keyinput_98), .ZN(n9421) );
  OAI221_X1 U10419 ( .B1(n5680), .B2(keyinput_99), .C1(P2_U3151), .C2(
        keyinput_98), .A(n9421), .ZN(n9494) );
  INV_X1 U10420 ( .A(keyinput_87), .ZN(n9473) );
  AOI22_X1 U10421 ( .A1(SI_11_), .A2(keyinput_85), .B1(n9423), .B2(keyinput_84), .ZN(n9422) );
  OAI221_X1 U10422 ( .B1(SI_11_), .B2(keyinput_85), .C1(n9423), .C2(
        keyinput_84), .A(n9422), .ZN(n9469) );
  OAI22_X1 U10423 ( .A1(n9425), .A2(keyinput_82), .B1(SI_15_), .B2(keyinput_81), .ZN(n9424) );
  AOI221_X1 U10424 ( .B1(n9425), .B2(keyinput_82), .C1(keyinput_81), .C2(
        SI_15_), .A(n9424), .ZN(n9465) );
  OAI22_X1 U10425 ( .A1(n9428), .A2(keyinput_78), .B1(n9427), .B2(keyinput_80), 
        .ZN(n9426) );
  AOI221_X1 U10426 ( .B1(n9428), .B2(keyinput_78), .C1(keyinput_80), .C2(n9427), .A(n9426), .ZN(n9463) );
  OAI22_X1 U10427 ( .A1(n9430), .A2(keyinput_77), .B1(SI_17_), .B2(keyinput_79), .ZN(n9429) );
  AOI221_X1 U10428 ( .B1(n9430), .B2(keyinput_77), .C1(keyinput_79), .C2(
        SI_17_), .A(n9429), .ZN(n9462) );
  INV_X1 U10429 ( .A(keyinput_76), .ZN(n9460) );
  INV_X1 U10430 ( .A(keyinput_75), .ZN(n9456) );
  INV_X1 U10431 ( .A(keyinput_74), .ZN(n9454) );
  INV_X1 U10432 ( .A(keyinput_70), .ZN(n9443) );
  INV_X1 U10433 ( .A(keyinput_69), .ZN(n9441) );
  AOI22_X1 U10434 ( .A1(n9433), .A2(keyinput_66), .B1(n9432), .B2(keyinput_67), 
        .ZN(n9431) );
  OAI221_X1 U10435 ( .B1(n9433), .B2(keyinput_66), .C1(n9432), .C2(keyinput_67), .A(n9431), .ZN(n9436) );
  OAI22_X1 U10436 ( .A1(SI_31_), .A2(keyinput_65), .B1(P2_WR_REG_SCAN_IN), 
        .B2(keyinput_64), .ZN(n9434) );
  AOI221_X1 U10437 ( .B1(SI_31_), .B2(keyinput_65), .C1(keyinput_64), .C2(
        P2_WR_REG_SCAN_IN), .A(n9434), .ZN(n9435) );
  OAI22_X1 U10438 ( .A1(keyinput_68), .A2(n9438), .B1(n9436), .B2(n9435), .ZN(
        n9437) );
  AOI21_X1 U10439 ( .B1(keyinput_68), .B2(n9438), .A(n9437), .ZN(n9439) );
  AOI221_X1 U10440 ( .B1(SI_27_), .B2(n9441), .C1(n9440), .C2(keyinput_69), 
        .A(n9439), .ZN(n9442) );
  AOI221_X1 U10441 ( .B1(SI_26_), .B2(keyinput_70), .C1(n9444), .C2(n9443), 
        .A(n9442), .ZN(n9449) );
  AOI22_X1 U10442 ( .A1(n9447), .A2(keyinput_73), .B1(n9446), .B2(keyinput_72), 
        .ZN(n9445) );
  OAI221_X1 U10443 ( .B1(n9447), .B2(keyinput_73), .C1(n9446), .C2(keyinput_72), .A(n9445), .ZN(n9448) );
  AOI211_X1 U10444 ( .C1(n9451), .C2(keyinput_71), .A(n9449), .B(n9448), .ZN(
        n9450) );
  OAI21_X1 U10445 ( .B1(n9451), .B2(keyinput_71), .A(n9450), .ZN(n9452) );
  OAI221_X1 U10446 ( .B1(SI_22_), .B2(n9454), .C1(n9453), .C2(keyinput_74), 
        .A(n9452), .ZN(n9455) );
  OAI221_X1 U10447 ( .B1(SI_21_), .B2(keyinput_75), .C1(n9457), .C2(n9456), 
        .A(n9455), .ZN(n9458) );
  OAI221_X1 U10448 ( .B1(SI_20_), .B2(n9460), .C1(n9459), .C2(keyinput_76), 
        .A(n9458), .ZN(n9461) );
  NAND3_X1 U10449 ( .A1(n9463), .A2(n9462), .A3(n9461), .ZN(n9464) );
  OAI211_X1 U10450 ( .C1(n9467), .C2(keyinput_83), .A(n9465), .B(n9464), .ZN(
        n9466) );
  AOI21_X1 U10451 ( .B1(n9467), .B2(keyinput_83), .A(n9466), .ZN(n9468) );
  OAI22_X1 U10452 ( .A1(n9469), .A2(n9468), .B1(keyinput_86), .B2(SI_10_), 
        .ZN(n9470) );
  AOI21_X1 U10453 ( .B1(keyinput_86), .B2(SI_10_), .A(n9470), .ZN(n9471) );
  AOI221_X1 U10454 ( .B1(SI_9_), .B2(n9473), .C1(n9472), .C2(keyinput_87), .A(
        n9471), .ZN(n9480) );
  AOI22_X1 U10455 ( .A1(n9476), .A2(keyinput_89), .B1(n9475), .B2(keyinput_88), 
        .ZN(n9474) );
  OAI221_X1 U10456 ( .B1(n9476), .B2(keyinput_89), .C1(n9475), .C2(keyinput_88), .A(n9474), .ZN(n9479) );
  OAI22_X1 U10457 ( .A1(SI_5_), .A2(keyinput_91), .B1(keyinput_93), .B2(SI_3_), 
        .ZN(n9477) );
  AOI221_X1 U10458 ( .B1(SI_5_), .B2(keyinput_91), .C1(SI_3_), .C2(keyinput_93), .A(n9477), .ZN(n9478) );
  OAI21_X1 U10459 ( .B1(n9480), .B2(n9479), .A(n9478), .ZN(n9487) );
  AOI22_X1 U10460 ( .A1(n9483), .A2(keyinput_92), .B1(n9482), .B2(keyinput_90), 
        .ZN(n9481) );
  OAI221_X1 U10461 ( .B1(n9483), .B2(keyinput_92), .C1(n9482), .C2(keyinput_90), .A(n9481), .ZN(n9486) );
  XOR2_X1 U10462 ( .A(SI_2_), .B(keyinput_94), .Z(n9485) );
  XNOR2_X1 U10463 ( .A(SI_1_), .B(keyinput_95), .ZN(n9484) );
  OAI211_X1 U10464 ( .C1(n9487), .C2(n9486), .A(n9485), .B(n9484), .ZN(n9488)
         );
  INV_X1 U10465 ( .A(n9488), .ZN(n9491) );
  AOI22_X1 U10466 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput_97), .B1(n6608), .B2(
        keyinput_96), .ZN(n9489) );
  OAI221_X1 U10467 ( .B1(P2_RD_REG_SCAN_IN), .B2(keyinput_97), .C1(n6608), 
        .C2(keyinput_96), .A(n9489), .ZN(n9490) );
  NOR2_X1 U10468 ( .A1(n9491), .A2(n9490), .ZN(n9493) );
  NAND2_X1 U10469 ( .A1(keyinput_100), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n9492) );
  OAI221_X1 U10470 ( .B1(n9494), .B2(n9493), .C1(keyinput_100), .C2(
        P2_REG3_REG_27__SCAN_IN), .A(n9492), .ZN(n9495) );
  OAI22_X1 U10471 ( .A1(n9496), .A2(n9495), .B1(keyinput_103), .B2(
        P2_REG3_REG_10__SCAN_IN), .ZN(n9497) );
  AOI21_X1 U10472 ( .B1(keyinput_103), .B2(P2_REG3_REG_10__SCAN_IN), .A(n9497), 
        .ZN(n9498) );
  AOI221_X1 U10473 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_104), .C1(n9500), .C2(n9499), .A(n9498), .ZN(n9501) );
  AOI221_X1 U10474 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(n9503), .C1(n9502), 
        .C2(keyinput_105), .A(n9501), .ZN(n9504) );
  AOI221_X1 U10475 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_106), .C1(
        n9506), .C2(n9505), .A(n9504), .ZN(n9511) );
  XNOR2_X1 U10476 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_108), .ZN(n9509)
         );
  XNOR2_X1 U10477 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_107), .ZN(n9508)
         );
  NAND2_X1 U10478 ( .A1(keyinput_109), .A2(n5689), .ZN(n9507) );
  NAND3_X1 U10479 ( .A1(n9509), .A2(n9508), .A3(n9507), .ZN(n9510) );
  NOR2_X1 U10480 ( .A1(n9511), .A2(n9510), .ZN(n9512) );
  OAI21_X1 U10481 ( .B1(n5689), .B2(keyinput_109), .A(n9512), .ZN(n9513) );
  OAI221_X1 U10482 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_110), .C1(
        n9515), .C2(n9514), .A(n9513), .ZN(n9516) );
  OAI221_X1 U10483 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(n9518), .C1(n9517), 
        .C2(keyinput_111), .A(n9516), .ZN(n9519) );
  OAI211_X1 U10484 ( .C1(P2_REG3_REG_5__SCAN_IN), .C2(keyinput_113), .A(n9520), 
        .B(n9519), .ZN(n9521) );
  AOI21_X1 U10485 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_113), .A(n9521), 
        .ZN(n9526) );
  AOI22_X1 U10486 ( .A1(n9524), .A2(keyinput_115), .B1(keyinput_116), .B2(
        n9523), .ZN(n9522) );
  OAI221_X1 U10487 ( .B1(n9524), .B2(keyinput_115), .C1(n9523), .C2(
        keyinput_116), .A(n9522), .ZN(n9525) );
  AOI211_X1 U10488 ( .C1(n5682), .C2(keyinput_117), .A(n9526), .B(n9525), .ZN(
        n9527) );
  OAI21_X1 U10489 ( .B1(n5682), .B2(keyinput_117), .A(n9527), .ZN(n9530) );
  AOI22_X1 U10490 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput_120), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput_121), .ZN(n9528) );
  OAI221_X1 U10491 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_120), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_121), .A(n9528), .ZN(n9529) );
  AOI21_X1 U10492 ( .B1(n9531), .B2(n9530), .A(n9529), .ZN(n9532) );
  AOI221_X1 U10493 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(n9534), .C1(n9533), 
        .C2(keyinput_122), .A(n9532), .ZN(n9541) );
  AOI22_X1 U10494 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_123), .B1(n9536), 
        .B2(keyinput_124), .ZN(n9535) );
  OAI221_X1 U10495 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_123), .C1(n9536), .C2(keyinput_124), .A(n9535), .ZN(n9540) );
  OAI22_X1 U10496 ( .A1(n9538), .A2(keyinput_125), .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_126), .ZN(n9537) );
  AOI221_X1 U10497 ( .B1(n9538), .B2(keyinput_125), .C1(keyinput_126), .C2(
        P2_REG3_REG_26__SCAN_IN), .A(n9537), .ZN(n9539) );
  OAI21_X1 U10498 ( .B1(n9541), .B2(n9540), .A(n9539), .ZN(n9543) );
  AOI21_X1 U10499 ( .B1(keyinput_127), .B2(n9543), .A(keyinput_63), .ZN(n9545)
         );
  INV_X1 U10500 ( .A(keyinput_127), .ZN(n9542) );
  AOI21_X1 U10501 ( .B1(n9543), .B2(n9542), .A(P2_REG3_REG_15__SCAN_IN), .ZN(
        n9544) );
  AOI22_X1 U10502 ( .A1(n9545), .A2(P2_REG3_REG_15__SCAN_IN), .B1(n9544), .B2(
        keyinput_63), .ZN(n9546) );
  AOI21_X1 U10503 ( .B1(n9548), .B2(n9547), .A(n9546), .ZN(n9558) );
  XNOR2_X1 U10504 ( .A(n9551), .B(n9550), .ZN(n9552) );
  XNOR2_X1 U10505 ( .A(n9549), .B(n9552), .ZN(n9556) );
  NAND2_X1 U10506 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n10061)
         );
  OAI21_X1 U10507 ( .B1(n9655), .B2(n10335), .A(n10061), .ZN(n9554) );
  OAI22_X1 U10508 ( .A1(n9639), .A2(n10253), .B1(n9654), .B2(n10219), .ZN(
        n9553) );
  AOI211_X1 U10509 ( .C1(n10349), .C2(n9642), .A(n9554), .B(n9553), .ZN(n9555)
         );
  OAI21_X1 U10510 ( .B1(n9556), .B2(n9632), .A(n9555), .ZN(n9557) );
  XOR2_X1 U10511 ( .A(n9558), .B(n9557), .Z(P1_U3219) );
  NAND2_X1 U10512 ( .A1(n9559), .A2(n9651), .ZN(n9567) );
  AOI21_X1 U10513 ( .B1(n9606), .B2(n9561), .A(n9560), .ZN(n9566) );
  INV_X1 U10514 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9562) );
  OAI22_X1 U10515 ( .A1(n9639), .A2(n10335), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9562), .ZN(n9564) );
  OAI22_X1 U10516 ( .A1(n9655), .A2(n10336), .B1(n9654), .B2(n10192), .ZN(
        n9563) );
  AOI211_X1 U10517 ( .C1(n10339), .C2(n9642), .A(n9564), .B(n9563), .ZN(n9565)
         );
  OAI21_X1 U10518 ( .B1(n9567), .B2(n9566), .A(n9565), .ZN(P1_U3223) );
  OAI21_X1 U10519 ( .B1(n9569), .B2(n9568), .A(n9636), .ZN(n9570) );
  NAND2_X1 U10520 ( .A1(n9570), .A2(n9651), .ZN(n9574) );
  NOR2_X1 U10521 ( .A1(n9655), .A2(n10305), .ZN(n9572) );
  OAI22_X1 U10522 ( .A1(n9639), .A2(n10318), .B1(n9654), .B2(n10140), .ZN(
        n9571) );
  AOI211_X1 U10523 ( .C1(P1_REG3_REG_25__SCAN_IN), .C2(P1_U3086), .A(n9572), 
        .B(n9571), .ZN(n9573) );
  OAI211_X1 U10524 ( .C1(n10146), .C2(n9661), .A(n9574), .B(n9573), .ZN(
        P1_U3225) );
  INV_X1 U10525 ( .A(n9575), .ZN(n9646) );
  OAI21_X1 U10526 ( .B1(n9646), .B2(n9652), .A(n9576), .ZN(n9577) );
  INV_X1 U10527 ( .A(n9577), .ZN(n9578) );
  OAI21_X1 U10528 ( .B1(n9579), .B2(n9578), .A(n9651), .ZN(n9584) );
  AND2_X1 U10529 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10001) );
  OAI22_X1 U10530 ( .A1(n9639), .A2(n10824), .B1(n9654), .B2(n9580), .ZN(n9581) );
  AOI211_X1 U10531 ( .C1(n9582), .C2(n9956), .A(n10001), .B(n9581), .ZN(n9583)
         );
  OAI211_X1 U10532 ( .C1(n9790), .C2(n9661), .A(n9584), .B(n9583), .ZN(
        P1_U3226) );
  INV_X1 U10533 ( .A(n9585), .ZN(n9586) );
  NOR2_X1 U10534 ( .A1(n9587), .A2(n9586), .ZN(n9588) );
  XNOR2_X1 U10535 ( .A(n9589), .B(n9588), .ZN(n9594) );
  AOI22_X1 U10536 ( .A1(n9658), .A2(n10368), .B1(n9590), .B2(n10259), .ZN(
        n9591) );
  NAND2_X1 U10537 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10026)
         );
  OAI211_X1 U10538 ( .C1(n10253), .C2(n9655), .A(n9591), .B(n10026), .ZN(n9592) );
  AOI21_X1 U10539 ( .B1(n10360), .B2(n9642), .A(n9592), .ZN(n9593) );
  OAI21_X1 U10540 ( .B1(n9594), .B2(n9632), .A(n9593), .ZN(P1_U3228) );
  NOR2_X1 U10541 ( .A1(n9595), .A2(n8416), .ZN(n9599) );
  INV_X1 U10542 ( .A(n9596), .ZN(n9597) );
  AOI21_X1 U10543 ( .B1(n9599), .B2(n9598), .A(n9597), .ZN(n9605) );
  INV_X1 U10544 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9600) );
  OAI22_X1 U10545 ( .A1(n9655), .A2(n9638), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9600), .ZN(n9603) );
  OAI22_X1 U10546 ( .A1(n10176), .A2(n9639), .B1(n9654), .B2(n9601), .ZN(n9602) );
  AOI211_X1 U10547 ( .C1(n10314), .C2(n9642), .A(n9603), .B(n9602), .ZN(n9604)
         );
  OAI21_X1 U10548 ( .B1(n9605), .B2(n9632), .A(n9604), .ZN(P1_U3229) );
  OAI21_X1 U10549 ( .B1(n9607), .B2(n4964), .A(n9606), .ZN(n9608) );
  NAND2_X1 U10550 ( .A1(n9608), .A2(n9651), .ZN(n9613) );
  OAI22_X1 U10551 ( .A1(n9655), .A2(n10214), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9609), .ZN(n9611) );
  OAI22_X1 U10552 ( .A1(n9639), .A2(n10237), .B1(n9654), .B2(n10207), .ZN(
        n9610) );
  AOI211_X1 U10553 ( .C1(n10345), .C2(n9642), .A(n9611), .B(n9610), .ZN(n9612)
         );
  NAND2_X1 U10554 ( .A1(n9613), .A2(n9612), .ZN(P1_U3233) );
  NAND2_X1 U10555 ( .A1(n9615), .A2(n9614), .ZN(n9616) );
  XOR2_X1 U10556 ( .A(n9617), .B(n9616), .Z(n9623) );
  OAI22_X1 U10557 ( .A1(n10176), .A2(n9655), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9618), .ZN(n9621) );
  INV_X1 U10558 ( .A(n10173), .ZN(n9619) );
  OAI22_X1 U10559 ( .A1(n9639), .A2(n10214), .B1(n9654), .B2(n9619), .ZN(n9620) );
  AOI211_X1 U10560 ( .C1(n10178), .C2(n9642), .A(n9621), .B(n9620), .ZN(n9622)
         );
  OAI21_X1 U10561 ( .B1(n9623), .B2(n9632), .A(n9622), .ZN(P1_U3235) );
  INV_X1 U10562 ( .A(n9624), .ZN(n9625) );
  NOR2_X1 U10563 ( .A1(n9626), .A2(n9625), .ZN(n9628) );
  XNOR2_X1 U10564 ( .A(n9628), .B(n9627), .ZN(n9633) );
  NAND2_X1 U10565 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10042)
         );
  OAI21_X1 U10566 ( .B1(n9655), .B2(n10237), .A(n10042), .ZN(n9630) );
  OAI22_X1 U10567 ( .A1(n9639), .A2(n10236), .B1(n9654), .B2(n10240), .ZN(
        n9629) );
  AOI211_X1 U10568 ( .C1(n10355), .C2(n9642), .A(n9630), .B(n9629), .ZN(n9631)
         );
  OAI21_X1 U10569 ( .B1(n9633), .B2(n9632), .A(n9631), .ZN(P1_U3238) );
  NAND2_X1 U10570 ( .A1(n9269), .A2(n9651), .ZN(n9645) );
  AOI21_X1 U10571 ( .B1(n9636), .B2(n9635), .A(n9634), .ZN(n9644) );
  OAI22_X1 U10572 ( .A1(n9639), .A2(n9638), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9637), .ZN(n9641) );
  OAI22_X1 U10573 ( .A1(n9655), .A2(n10281), .B1(n9654), .B2(n10126), .ZN(
        n9640) );
  AOI211_X1 U10574 ( .C1(n10131), .C2(n9642), .A(n9641), .B(n9640), .ZN(n9643)
         );
  OAI21_X1 U10575 ( .B1(n9645), .B2(n9644), .A(n9643), .ZN(P1_U3240) );
  INV_X1 U10576 ( .A(n9647), .ZN(n9649) );
  OAI21_X1 U10577 ( .B1(n9649), .B2(n9652), .A(n9648), .ZN(n9650) );
  OAI211_X1 U10578 ( .C1(n9575), .C2(n9652), .A(n9651), .B(n9650), .ZN(n9660)
         );
  OAI22_X1 U10579 ( .A1(n9655), .A2(n10252), .B1(n9654), .B2(n9653), .ZN(n9656) );
  AOI211_X1 U10580 ( .C1(n9658), .C2(n10369), .A(n9657), .B(n9656), .ZN(n9659)
         );
  OAI211_X1 U10581 ( .C1(n10371), .C2(n9661), .A(n9660), .B(n9659), .ZN(
        P1_U3241) );
  INV_X1 U10582 ( .A(n10076), .ZN(n9663) );
  INV_X1 U10583 ( .A(n9942), .ZN(n9832) );
  NAND2_X1 U10584 ( .A1(n9664), .A2(n9695), .ZN(n9666) );
  NAND2_X1 U10585 ( .A1(n9697), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n9665) );
  NAND2_X1 U10586 ( .A1(n10272), .A2(n10280), .ZN(n9934) );
  INV_X1 U10587 ( .A(n10188), .ZN(n10186) );
  NAND4_X1 U10588 ( .A1(n9668), .A2(n9667), .A3(n10589), .A4(n9830), .ZN(n9673) );
  INV_X1 U10589 ( .A(n9669), .ZN(n9671) );
  NAND4_X1 U10590 ( .A1(n9671), .A2(n9732), .A3(n9746), .A4(n5042), .ZN(n9672)
         );
  NOR2_X1 U10591 ( .A1(n9673), .A2(n9672), .ZN(n9675) );
  NAND3_X1 U10592 ( .A1(n9675), .A2(n9674), .A3(n9758), .ZN(n9676) );
  NOR2_X1 U10593 ( .A1(n9677), .A2(n9676), .ZN(n9678) );
  NAND4_X1 U10594 ( .A1(n9680), .A2(n9901), .A3(n9679), .A4(n9678), .ZN(n9681)
         );
  NOR2_X1 U10595 ( .A1(n9682), .A2(n9681), .ZN(n9683) );
  NAND2_X1 U10596 ( .A1(n10821), .A2(n9683), .ZN(n9684) );
  OR3_X1 U10597 ( .A1(n9686), .A2(n9685), .A3(n9684), .ZN(n9687) );
  XNOR2_X1 U10598 ( .A(n10355), .B(n10253), .ZN(n10234) );
  AND2_X1 U10599 ( .A1(n9922), .A2(n9720), .ZN(n10248) );
  INV_X1 U10600 ( .A(n10248), .ZN(n10249) );
  OR4_X1 U10601 ( .A1(n9688), .A2(n9687), .A3(n10234), .A4(n10249), .ZN(n9690)
         );
  OR4_X1 U10602 ( .A1(n10186), .A2(n9690), .A3(n9689), .A4(n10211), .ZN(n9692)
         );
  OR4_X1 U10603 ( .A1(n9692), .A2(n10137), .A3(n9691), .A4(n10153), .ZN(n9693)
         );
  NOR2_X1 U10604 ( .A1(n10123), .A2(n9693), .ZN(n9694) );
  NAND4_X1 U10605 ( .A1(n5417), .A2(n10089), .A3(n10109), .A4(n9694), .ZN(
        n9708) );
  NAND2_X1 U10606 ( .A1(n9696), .A2(n9695), .ZN(n9699) );
  NAND2_X1 U10607 ( .A1(n9697), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9698) );
  INV_X1 U10608 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n10081) );
  NAND2_X1 U10609 ( .A1(n9700), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n9704) );
  INV_X1 U10610 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9701) );
  OR2_X1 U10611 ( .A1(n9702), .A2(n9701), .ZN(n9703) );
  OAI211_X1 U10612 ( .C1(n9705), .C2(n10081), .A(n9704), .B(n9703), .ZN(n10098) );
  INV_X1 U10613 ( .A(n10098), .ZN(n9706) );
  OR2_X1 U10614 ( .A1(n10084), .A2(n9706), .ZN(n9937) );
  NAND2_X1 U10615 ( .A1(n10084), .A2(n9706), .ZN(n9933) );
  NAND2_X1 U10616 ( .A1(n9937), .A2(n9933), .ZN(n9707) );
  AOI211_X1 U10617 ( .C1(n6607), .C2(n9709), .A(n10062), .B(n9837), .ZN(n9886)
         );
  INV_X1 U10618 ( .A(n9862), .ZN(n10088) );
  INV_X1 U10619 ( .A(n9850), .ZN(n9710) );
  MUX2_X1 U10620 ( .A(n10088), .B(n9710), .S(n9820), .Z(n9826) );
  AND2_X1 U10621 ( .A1(n9954), .A2(n9820), .ZN(n9712) );
  OAI21_X1 U10622 ( .B1(n9820), .B2(n9954), .A(n10131), .ZN(n9711) );
  OAI21_X1 U10623 ( .B1(n9712), .B2(n10131), .A(n9711), .ZN(n9823) );
  NAND2_X1 U10624 ( .A1(n9838), .A2(n9713), .ZN(n9854) );
  NAND2_X1 U10625 ( .A1(n9809), .A2(n9714), .ZN(n9839) );
  NAND2_X1 U10626 ( .A1(n9929), .A2(n9717), .ZN(n9716) );
  NAND2_X1 U10627 ( .A1(n10184), .A2(n9925), .ZN(n9715) );
  MUX2_X1 U10628 ( .A(n9716), .B(n9715), .S(n9831), .Z(n9804) );
  NAND2_X1 U10629 ( .A1(n9717), .A2(n9719), .ZN(n9927) );
  MUX2_X1 U10630 ( .A(n9718), .B(n9927), .S(n9831), .Z(n9801) );
  AND2_X1 U10631 ( .A1(n9719), .A2(n9922), .ZN(n9722) );
  AND2_X1 U10632 ( .A1(n9721), .A2(n9720), .ZN(n9887) );
  MUX2_X1 U10633 ( .A(n9722), .B(n9887), .S(n9831), .Z(n9798) );
  INV_X1 U10634 ( .A(n9723), .ZN(n9724) );
  OAI211_X1 U10635 ( .C1(n9725), .C2(n9724), .A(n9894), .B(n9893), .ZN(n9726)
         );
  NAND2_X1 U10636 ( .A1(n9726), .A2(n9729), .ZN(n9727) );
  NAND3_X1 U10637 ( .A1(n9727), .A2(n9732), .A3(n9739), .ZN(n9728) );
  NAND2_X1 U10638 ( .A1(n9728), .A2(n10684), .ZN(n9738) );
  INV_X1 U10639 ( .A(n9729), .ZN(n9730) );
  OR2_X1 U10640 ( .A1(n9731), .A2(n9730), .ZN(n9896) );
  NAND2_X1 U10641 ( .A1(n9896), .A2(n9894), .ZN(n9733) );
  NAND2_X1 U10642 ( .A1(n9733), .A2(n9732), .ZN(n9736) );
  AND2_X1 U10643 ( .A1(n9739), .A2(n9734), .ZN(n9897) );
  INV_X1 U10644 ( .A(n10684), .ZN(n9735) );
  AOI21_X1 U10645 ( .B1(n9736), .B2(n9897), .A(n9735), .ZN(n9737) );
  MUX2_X1 U10646 ( .A(n9738), .B(n9737), .S(n9820), .Z(n9748) );
  INV_X1 U10647 ( .A(n9739), .ZN(n9740) );
  OAI21_X1 U10648 ( .B1(n9740), .B2(n9899), .A(n9746), .ZN(n9742) );
  OAI21_X1 U10649 ( .B1(n9748), .B2(n9742), .A(n9741), .ZN(n9743) );
  NAND3_X1 U10650 ( .A1(n9743), .A2(n10718), .A3(n10716), .ZN(n9745) );
  NAND2_X1 U10651 ( .A1(n9745), .A2(n9744), .ZN(n9754) );
  OAI211_X1 U10652 ( .C1(n9748), .C2(n9747), .A(n9746), .B(n10716), .ZN(n9750)
         );
  NAND3_X1 U10653 ( .A1(n9750), .A2(n10718), .A3(n9749), .ZN(n9752) );
  NAND3_X1 U10654 ( .A1(n9752), .A2(n9758), .A3(n9751), .ZN(n9753) );
  MUX2_X1 U10655 ( .A(n9754), .B(n9753), .S(n9820), .Z(n9771) );
  OAI211_X1 U10656 ( .C1(n5442), .C2(n9756), .A(n9772), .B(n9755), .ZN(n9759)
         );
  OAI211_X1 U10657 ( .C1(n9904), .C2(n9758), .A(n9761), .B(n9757), .ZN(n9907)
         );
  MUX2_X1 U10658 ( .A(n9759), .B(n9907), .S(n9831), .Z(n9769) );
  INV_X1 U10659 ( .A(n9769), .ZN(n9760) );
  OAI21_X1 U10660 ( .B1(n9771), .B2(n5442), .A(n9760), .ZN(n9762) );
  NAND3_X1 U10661 ( .A1(n9762), .A2(n9767), .A3(n9761), .ZN(n9763) );
  NAND3_X1 U10662 ( .A1(n9763), .A2(n9773), .A3(n9775), .ZN(n9764) );
  NAND2_X1 U10663 ( .A1(n9764), .A2(n9768), .ZN(n9766) );
  NAND4_X1 U10664 ( .A1(n9919), .A2(n9820), .A3(n9913), .A4(n9912), .ZN(n9765)
         );
  AOI21_X1 U10665 ( .B1(n9766), .B2(n10821), .A(n9765), .ZN(n9796) );
  NAND2_X1 U10666 ( .A1(n9768), .A2(n9767), .ZN(n9909) );
  NOR2_X1 U10667 ( .A1(n9909), .A2(n9769), .ZN(n9770) );
  OAI21_X1 U10668 ( .B1(n9771), .B2(n9904), .A(n9770), .ZN(n9777) );
  AND2_X1 U10669 ( .A1(n9773), .A2(n9772), .ZN(n9774) );
  OR2_X1 U10670 ( .A1(n9909), .A2(n9774), .ZN(n9776) );
  AND2_X1 U10671 ( .A1(n9776), .A2(n9775), .ZN(n9888) );
  INV_X1 U10672 ( .A(n10821), .ZN(n10814) );
  AOI21_X1 U10673 ( .B1(n9777), .B2(n9888), .A(n10814), .ZN(n9794) );
  NAND4_X1 U10674 ( .A1(n9921), .A2(n9831), .A3(n9911), .A4(n9916), .ZN(n9793)
         );
  NAND3_X1 U10675 ( .A1(n9788), .A2(n10824), .A3(n9831), .ZN(n9778) );
  OR2_X1 U10676 ( .A1(n10368), .A2(n9820), .ZN(n9779) );
  NAND2_X1 U10677 ( .A1(n9778), .A2(n9779), .ZN(n9785) );
  INV_X1 U10678 ( .A(n9779), .ZN(n9780) );
  NAND2_X1 U10679 ( .A1(n9780), .A2(n10824), .ZN(n9781) );
  NAND2_X1 U10680 ( .A1(n9788), .A2(n9781), .ZN(n9784) );
  NAND2_X1 U10681 ( .A1(n10368), .A2(n9820), .ZN(n9786) );
  NOR2_X1 U10682 ( .A1(n9786), .A2(n10824), .ZN(n9782) );
  OR2_X1 U10683 ( .A1(n9788), .A2(n9782), .ZN(n9783) );
  AOI22_X1 U10684 ( .A1(n10365), .A2(n9785), .B1(n9784), .B2(n9783), .ZN(n9792) );
  NAND2_X1 U10685 ( .A1(n9957), .A2(n9820), .ZN(n9787) );
  OAI21_X1 U10686 ( .B1(n9788), .B2(n9787), .A(n9786), .ZN(n9789) );
  NAND2_X1 U10687 ( .A1(n9790), .A2(n9789), .ZN(n9791) );
  OAI211_X1 U10688 ( .C1(n9794), .C2(n9793), .A(n9792), .B(n9791), .ZN(n9795)
         );
  OAI21_X1 U10689 ( .B1(n9796), .B2(n9795), .A(n10248), .ZN(n9797) );
  NAND2_X1 U10690 ( .A1(n9798), .A2(n9797), .ZN(n9799) );
  NAND2_X1 U10691 ( .A1(n9799), .A2(n9925), .ZN(n9800) );
  NOR2_X1 U10692 ( .A1(n9801), .A2(n9800), .ZN(n9803) );
  MUX2_X1 U10693 ( .A(n10184), .B(n9929), .S(n9831), .Z(n9802) );
  OAI211_X1 U10694 ( .C1(n9804), .C2(n9803), .A(n10188), .B(n9802), .ZN(n9807)
         );
  MUX2_X1 U10695 ( .A(n9805), .B(n9930), .S(n9820), .Z(n9806) );
  NAND2_X1 U10696 ( .A1(n9807), .A2(n9806), .ZN(n9808) );
  MUX2_X1 U10697 ( .A(n9838), .B(n9809), .S(n9831), .Z(n9810) );
  OAI211_X1 U10698 ( .C1(n9814), .C2(n9813), .A(n9831), .B(n9846), .ZN(n9822)
         );
  AND2_X1 U10699 ( .A1(n9816), .A2(n9815), .ZN(n9845) );
  NAND3_X1 U10700 ( .A1(n9818), .A2(n9817), .A3(n9841), .ZN(n9819) );
  NAND3_X1 U10701 ( .A1(n9845), .A2(n9820), .A3(n9819), .ZN(n9821) );
  NAND4_X1 U10702 ( .A1(n10089), .A2(n9823), .A3(n9822), .A4(n9821), .ZN(n9825) );
  MUX2_X1 U10703 ( .A(n10086), .B(n9847), .S(n9831), .Z(n9824) );
  MUX2_X1 U10704 ( .A(n9934), .B(n9853), .S(n9831), .Z(n9827) );
  NOR2_X1 U10705 ( .A1(n9829), .A2(n10270), .ZN(n9836) );
  AND2_X1 U10706 ( .A1(n10098), .A2(n10076), .ZN(n9864) );
  OAI211_X1 U10707 ( .C1(n10084), .C2(n9831), .A(n10078), .B(n9864), .ZN(n9835) );
  AOI211_X1 U10708 ( .C1(n9831), .C2(n10084), .A(n9864), .B(n9939), .ZN(n9828)
         );
  OAI211_X1 U10709 ( .C1(n9836), .C2(n9829), .A(n9828), .B(n9942), .ZN(n9834)
         );
  AOI21_X1 U10710 ( .B1(n9832), .B2(n9831), .A(n9830), .ZN(n9833) );
  OAI211_X1 U10711 ( .C1(n9836), .C2(n9835), .A(n9834), .B(n9833), .ZN(n9885)
         );
  INV_X1 U10712 ( .A(n9837), .ZN(n9873) );
  NAND2_X1 U10713 ( .A1(n9839), .A2(n9838), .ZN(n9840) );
  NAND2_X1 U10714 ( .A1(n9841), .A2(n9840), .ZN(n9842) );
  NAND2_X1 U10715 ( .A1(n9842), .A2(n9857), .ZN(n9843) );
  AND2_X1 U10716 ( .A1(n9844), .A2(n9843), .ZN(n9848) );
  INV_X1 U10717 ( .A(n9845), .ZN(n9859) );
  OAI211_X1 U10718 ( .C1(n9848), .C2(n9859), .A(n9847), .B(n9846), .ZN(n9849)
         );
  NAND3_X1 U10719 ( .A1(n9862), .A2(n10086), .A3(n9849), .ZN(n9851) );
  AND2_X1 U10720 ( .A1(n9851), .A2(n9850), .ZN(n9852) );
  NAND2_X1 U10721 ( .A1(n9853), .A2(n9852), .ZN(n9936) );
  INV_X1 U10722 ( .A(n9854), .ZN(n9856) );
  NAND3_X1 U10723 ( .A1(n9857), .A2(n9856), .A3(n9855), .ZN(n9858) );
  NOR2_X1 U10724 ( .A1(n9859), .A2(n9858), .ZN(n9860) );
  AND2_X1 U10725 ( .A1(n10086), .A2(n9860), .ZN(n9861) );
  NAND2_X1 U10726 ( .A1(n9862), .A2(n9861), .ZN(n9932) );
  NOR2_X1 U10727 ( .A1(n9932), .A2(n9863), .ZN(n9867) );
  INV_X1 U10728 ( .A(n9864), .ZN(n9865) );
  NAND2_X1 U10729 ( .A1(n10084), .A2(n9865), .ZN(n9866) );
  OAI211_X1 U10730 ( .C1(n9936), .C2(n9867), .A(n9934), .B(n9866), .ZN(n9871)
         );
  INV_X1 U10731 ( .A(n9937), .ZN(n9869) );
  AOI21_X1 U10732 ( .B1(n9869), .B2(n10078), .A(n9868), .ZN(n9870) );
  OAI211_X1 U10733 ( .C1(n9939), .C2(n9871), .A(n9870), .B(n9942), .ZN(n9872)
         );
  AOI21_X1 U10734 ( .B1(n9873), .B2(n9872), .A(n9882), .ZN(n9880) );
  INV_X1 U10735 ( .A(n9874), .ZN(n9878) );
  OAI21_X1 U10736 ( .B1(n9875), .B2(n9881), .A(P1_B_REG_SCAN_IN), .ZN(n9876)
         );
  AOI21_X1 U10737 ( .B1(n9878), .B2(n9877), .A(n9876), .ZN(n9950) );
  OR3_X1 U10738 ( .A1(n9880), .A2(n9950), .A3(n9879), .ZN(n9884) );
  AOI211_X1 U10739 ( .C1(n9882), .C2(n9939), .A(n9881), .B(n9885), .ZN(n9883)
         );
  AOI211_X1 U10740 ( .C1(n9886), .C2(n9885), .A(n9884), .B(n9883), .ZN(n9953)
         );
  INV_X1 U10741 ( .A(n9887), .ZN(n9924) );
  INV_X1 U10742 ( .A(n9888), .ZN(n9915) );
  NAND2_X1 U10743 ( .A1(n10591), .A2(n9889), .ZN(n9892) );
  NAND2_X1 U10744 ( .A1(n9968), .A2(n9890), .ZN(n9891) );
  AND4_X1 U10745 ( .A1(n9893), .A2(n6607), .A3(n9892), .A4(n9891), .ZN(n9895)
         );
  OAI21_X1 U10746 ( .B1(n9896), .B2(n9895), .A(n9894), .ZN(n9900) );
  INV_X1 U10747 ( .A(n9897), .ZN(n9898) );
  AOI21_X1 U10748 ( .B1(n9900), .B2(n9899), .A(n9898), .ZN(n9903) );
  OAI21_X1 U10749 ( .B1(n9903), .B2(n9902), .A(n9901), .ZN(n9906) );
  AOI21_X1 U10750 ( .B1(n9906), .B2(n9905), .A(n9904), .ZN(n9908) );
  OR3_X1 U10751 ( .A1(n9909), .A2(n9908), .A3(n9907), .ZN(n9910) );
  NAND2_X1 U10752 ( .A1(n9911), .A2(n9910), .ZN(n9914) );
  OAI211_X1 U10753 ( .C1(n9915), .C2(n9914), .A(n9913), .B(n9912), .ZN(n9917)
         );
  NAND2_X1 U10754 ( .A1(n9917), .A2(n9916), .ZN(n9918) );
  NAND2_X1 U10755 ( .A1(n9919), .A2(n9918), .ZN(n9920) );
  AND3_X1 U10756 ( .A1(n9922), .A2(n9921), .A3(n9920), .ZN(n9923) );
  NOR2_X1 U10757 ( .A1(n9924), .A2(n9923), .ZN(n9926) );
  OAI21_X1 U10758 ( .B1(n9927), .B2(n9926), .A(n9925), .ZN(n9928) );
  AND3_X1 U10759 ( .A1(n9930), .A2(n9929), .A3(n9928), .ZN(n9931) );
  NOR2_X1 U10760 ( .A1(n9932), .A2(n9931), .ZN(n9935) );
  OAI211_X1 U10761 ( .C1(n9936), .C2(n9935), .A(n9934), .B(n9933), .ZN(n9938)
         );
  NAND2_X1 U10762 ( .A1(n9938), .A2(n9937), .ZN(n9941) );
  INV_X1 U10763 ( .A(n9939), .ZN(n9940) );
  NAND2_X1 U10764 ( .A1(n9941), .A2(n9940), .ZN(n9943) );
  NAND2_X1 U10765 ( .A1(n9943), .A2(n9942), .ZN(n9947) );
  INV_X1 U10766 ( .A(n9950), .ZN(n9944) );
  NAND3_X1 U10767 ( .A1(n9947), .A2(n9945), .A3(n9944), .ZN(n9949) );
  OR4_X1 U10768 ( .A1(n9947), .A2(n9950), .A3(n9946), .A4(n10062), .ZN(n9948)
         );
  OAI211_X1 U10769 ( .C1(n9951), .C2(n9950), .A(n9949), .B(n9948), .ZN(n9952)
         );
  NOR2_X1 U10770 ( .A1(n9953), .A2(n9952), .ZN(P1_U3242) );
  MUX2_X1 U10771 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n10098), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10772 ( .A(n10093), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9967), .Z(
        P1_U3582) );
  MUX2_X1 U10773 ( .A(n10296), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9967), .Z(
        P1_U3581) );
  MUX2_X1 U10774 ( .A(n9954), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9967), .Z(
        P1_U3580) );
  MUX2_X1 U10775 ( .A(n10297), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9967), .Z(
        P1_U3579) );
  MUX2_X1 U10776 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n10161), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10777 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n10325), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10778 ( .A(n9955), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9967), .Z(
        P1_U3573) );
  MUX2_X1 U10779 ( .A(n10226), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9967), .Z(
        P1_U3572) );
  MUX2_X1 U10780 ( .A(n9956), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9967), .Z(
        P1_U3571) );
  MUX2_X1 U10781 ( .A(n10368), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9967), .Z(
        P1_U3570) );
  MUX2_X1 U10782 ( .A(n9957), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9967), .Z(
        P1_U3569) );
  MUX2_X1 U10783 ( .A(n10369), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9967), .Z(
        P1_U3568) );
  MUX2_X1 U10784 ( .A(n9958), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9967), .Z(
        P1_U3566) );
  MUX2_X1 U10785 ( .A(n9959), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9967), .Z(
        P1_U3565) );
  MUX2_X1 U10786 ( .A(n9960), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9967), .Z(
        P1_U3564) );
  MUX2_X1 U10787 ( .A(n9961), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9967), .Z(
        P1_U3563) );
  MUX2_X1 U10788 ( .A(n10746), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9967), .Z(
        P1_U3562) );
  MUX2_X1 U10789 ( .A(n9962), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9967), .Z(
        P1_U3561) );
  MUX2_X1 U10790 ( .A(n9963), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9967), .Z(
        P1_U3559) );
  MUX2_X1 U10791 ( .A(n9964), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9967), .Z(
        P1_U3558) );
  MUX2_X1 U10792 ( .A(n9965), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9967), .Z(
        P1_U3557) );
  MUX2_X1 U10793 ( .A(n9966), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9967), .Z(
        P1_U3556) );
  MUX2_X1 U10794 ( .A(n10591), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9967), .Z(
        P1_U3555) );
  MUX2_X1 U10795 ( .A(n9968), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9967), .Z(
        P1_U3554) );
  AOI211_X1 U10796 ( .C1(n9971), .C2(n9970), .A(n9969), .B(n10067), .ZN(n9972)
         );
  INV_X1 U10797 ( .A(n9972), .ZN(n9980) );
  AOI22_X1 U10798 ( .A1(n10059), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9979) );
  NAND2_X1 U10799 ( .A1(n10041), .A2(n9973), .ZN(n9978) );
  OAI211_X1 U10800 ( .C1(n9976), .C2(n9975), .A(n10065), .B(n9974), .ZN(n9977)
         );
  NAND4_X1 U10801 ( .A1(n9980), .A2(n9979), .A3(n9978), .A4(n9977), .ZN(
        P1_U3244) );
  AOI211_X1 U10802 ( .C1(n9983), .C2(n9982), .A(n9981), .B(n10067), .ZN(n9984)
         );
  INV_X1 U10803 ( .A(n9984), .ZN(n9994) );
  INV_X1 U10804 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9986) );
  OAI21_X1 U10805 ( .B1(n10044), .B2(n9986), .A(n9985), .ZN(n9987) );
  AOI21_X1 U10806 ( .B1(n9988), .B2(n10041), .A(n9987), .ZN(n9993) );
  OAI211_X1 U10807 ( .C1(n9991), .C2(n9990), .A(n10065), .B(n9989), .ZN(n9992)
         );
  NAND3_X1 U10808 ( .A1(n9994), .A2(n9993), .A3(n9992), .ZN(P1_U3246) );
  NOR2_X1 U10809 ( .A1(n9995), .A2(n10003), .ZN(n9997) );
  NOR2_X1 U10810 ( .A1(n9997), .A2(n9996), .ZN(n10000) );
  AOI22_X1 U10811 ( .A1(n10020), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9998), 
        .B2(n10007), .ZN(n9999) );
  NAND2_X1 U10812 ( .A1(n9999), .A2(n10000), .ZN(n10019) );
  OAI21_X1 U10813 ( .B1(n10000), .B2(n9999), .A(n10019), .ZN(n10012) );
  AOI21_X1 U10814 ( .B1(n10059), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n10001), 
        .ZN(n10002) );
  OAI21_X1 U10815 ( .B1(n10063), .B2(n10007), .A(n10002), .ZN(n10011) );
  NOR2_X1 U10816 ( .A1(n10004), .A2(n10003), .ZN(n10006) );
  AOI22_X1 U10817 ( .A1(n10020), .A2(n8047), .B1(P1_REG2_REG_16__SCAN_IN), 
        .B2(n10007), .ZN(n10008) );
  NOR2_X1 U10818 ( .A1(n10009), .A2(n10008), .ZN(n10015) );
  AOI211_X1 U10819 ( .C1(n10009), .C2(n10008), .A(n10015), .B(n10037), .ZN(
        n10010) );
  AOI211_X1 U10820 ( .C1(n10024), .C2(n10012), .A(n10011), .B(n10010), .ZN(
        n10013) );
  INV_X1 U10821 ( .A(n10013), .ZN(P1_U3259) );
  NOR2_X1 U10822 ( .A1(n10036), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n10014) );
  AOI21_X1 U10823 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n10036), .A(n10014), 
        .ZN(n10017) );
  NAND2_X1 U10824 ( .A1(n10017), .A2(n10016), .ZN(n10035) );
  OAI21_X1 U10825 ( .B1(n10017), .B2(n10016), .A(n10035), .ZN(n10018) );
  INV_X1 U10826 ( .A(n10018), .ZN(n10031) );
  OAI21_X1 U10827 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n10020), .A(n10019), 
        .ZN(n10023) );
  XNOR2_X1 U10828 ( .A(n10036), .B(n10021), .ZN(n10022) );
  NAND2_X1 U10829 ( .A1(n10022), .A2(n10023), .ZN(n10032) );
  OAI21_X1 U10830 ( .B1(n10023), .B2(n10022), .A(n10032), .ZN(n10025) );
  NAND2_X1 U10831 ( .A1(n10025), .A2(n10024), .ZN(n10030) );
  INV_X1 U10832 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10027) );
  OAI21_X1 U10833 ( .B1(n10044), .B2(n10027), .A(n10026), .ZN(n10028) );
  AOI21_X1 U10834 ( .B1(n10036), .B2(n10041), .A(n10028), .ZN(n10029) );
  OAI211_X1 U10835 ( .C1(n10031), .C2(n10037), .A(n10030), .B(n10029), .ZN(
        P1_U3260) );
  NAND2_X1 U10836 ( .A1(n10040), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n10048) );
  OAI21_X1 U10837 ( .B1(n10040), .B2(P1_REG1_REG_18__SCAN_IN), .A(n10048), 
        .ZN(n10034) );
  OAI21_X1 U10838 ( .B1(n10036), .B2(P1_REG1_REG_17__SCAN_IN), .A(n10032), 
        .ZN(n10033) );
  NOR2_X1 U10839 ( .A1(n10033), .A2(n10034), .ZN(n10050) );
  AOI211_X1 U10840 ( .C1(n10034), .C2(n10033), .A(n10050), .B(n10067), .ZN(
        n10047) );
  OAI21_X1 U10841 ( .B1(n10036), .B2(P1_REG2_REG_17__SCAN_IN), .A(n10035), 
        .ZN(n10039) );
  NAND2_X1 U10842 ( .A1(n10040), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n10054) );
  OAI21_X1 U10843 ( .B1(n10040), .B2(P1_REG2_REG_18__SCAN_IN), .A(n10054), 
        .ZN(n10038) );
  NOR2_X1 U10844 ( .A1(n10038), .A2(n10039), .ZN(n10056) );
  AOI211_X1 U10845 ( .C1(n10039), .C2(n10038), .A(n10056), .B(n10037), .ZN(
        n10046) );
  INV_X1 U10846 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10479) );
  NAND2_X1 U10847 ( .A1(n10041), .A2(n10040), .ZN(n10043) );
  OAI211_X1 U10848 ( .C1(n10479), .C2(n10044), .A(n10043), .B(n10042), .ZN(
        n10045) );
  OR3_X1 U10849 ( .A1(n10047), .A2(n10046), .A3(n10045), .ZN(P1_U3261) );
  INV_X1 U10850 ( .A(n10048), .ZN(n10049) );
  NOR2_X1 U10851 ( .A1(n10050), .A2(n10049), .ZN(n10053) );
  XNOR2_X1 U10852 ( .A(n10062), .B(n10051), .ZN(n10052) );
  XNOR2_X1 U10853 ( .A(n10053), .B(n10052), .ZN(n10068) );
  MUX2_X1 U10854 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n8235), .S(n10062), .Z(
        n10058) );
  INV_X1 U10855 ( .A(n10054), .ZN(n10055) );
  NOR2_X1 U10856 ( .A1(n10056), .A2(n10055), .ZN(n10057) );
  NAND2_X1 U10857 ( .A1(n10059), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n10060) );
  OAI211_X1 U10858 ( .C1(n10063), .C2(n10062), .A(n10061), .B(n10060), .ZN(
        n10064) );
  OAI21_X1 U10859 ( .B1(n10068), .B2(n10067), .A(n10066), .ZN(P1_U3262) );
  NAND2_X1 U10860 ( .A1(n10270), .A2(n10096), .ZN(n10080) );
  XNOR2_X1 U10861 ( .A(n10267), .B(n10080), .ZN(n10071) );
  NAND2_X1 U10862 ( .A1(n10071), .A2(n10818), .ZN(n10266) );
  NOR2_X1 U10863 ( .A1(n10852), .A2(n10072), .ZN(n10077) );
  INV_X1 U10864 ( .A(P1_B_REG_SCAN_IN), .ZN(n10073) );
  NOR2_X1 U10865 ( .A1(n10074), .A2(n10073), .ZN(n10075) );
  NOR2_X1 U10866 ( .A1(n10823), .A2(n10075), .ZN(n10097) );
  NAND2_X1 U10867 ( .A1(n10076), .A2(n10097), .ZN(n10268) );
  NOR2_X1 U10868 ( .A1(n10731), .A2(n10268), .ZN(n10082) );
  AOI211_X1 U10869 ( .C1(n10078), .C2(n10732), .A(n10077), .B(n10082), .ZN(
        n10079) );
  OAI21_X1 U10870 ( .B1(n10266), .B2(n10180), .A(n10079), .ZN(P1_U3263) );
  OAI211_X1 U10871 ( .C1(n10270), .C2(n10096), .A(n10818), .B(n10080), .ZN(
        n10269) );
  NOR2_X1 U10872 ( .A1(n10852), .A2(n10081), .ZN(n10083) );
  AOI211_X1 U10873 ( .C1(n10084), .C2(n10732), .A(n10083), .B(n10082), .ZN(
        n10085) );
  OAI21_X1 U10874 ( .B1(n10269), .B2(n10180), .A(n10085), .ZN(P1_U3264) );
  NAND2_X1 U10875 ( .A1(n10087), .A2(n10086), .ZN(n10108) );
  INV_X1 U10876 ( .A(n10277), .ZN(n10106) );
  NAND2_X1 U10877 ( .A1(n10069), .A2(n10288), .ZN(n10092) );
  NAND2_X1 U10878 ( .A1(n10284), .A2(n10093), .ZN(n10094) );
  NAND2_X1 U10879 ( .A1(n10271), .A2(n10190), .ZN(n10105) );
  NAND2_X1 U10880 ( .A1(n10272), .A2(n10732), .ZN(n10102) );
  NAND2_X1 U10881 ( .A1(n10098), .A2(n10097), .ZN(n10273) );
  OAI22_X1 U10882 ( .A1(n10697), .A2(n10273), .B1(n10099), .B2(n10847), .ZN(
        n10100) );
  AOI21_X1 U10883 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(n10731), .A(n10100), 
        .ZN(n10101) );
  OAI211_X1 U10884 ( .C1(n10288), .C2(n10198), .A(n10102), .B(n10101), .ZN(
        n10103) );
  AOI21_X1 U10885 ( .B1(n10276), .B2(n4942), .A(n10103), .ZN(n10104) );
  OAI211_X1 U10886 ( .C1(n10202), .C2(n10106), .A(n10105), .B(n10104), .ZN(
        P1_U3356) );
  XNOR2_X1 U10887 ( .A(n10108), .B(n10107), .ZN(n10287) );
  XNOR2_X1 U10888 ( .A(n10110), .B(n10109), .ZN(n10279) );
  NAND2_X1 U10889 ( .A1(n10279), .A2(n10190), .ZN(n10121) );
  INV_X1 U10890 ( .A(n10111), .ZN(n10112) );
  OAI22_X1 U10891 ( .A1(n10852), .A2(n10115), .B1(n10114), .B2(n10847), .ZN(
        n10117) );
  NOR2_X1 U10892 ( .A1(n10193), .A2(n10280), .ZN(n10116) );
  AOI211_X1 U10893 ( .C1(n10172), .C2(n10296), .A(n10117), .B(n10116), .ZN(
        n10118) );
  OAI21_X1 U10894 ( .B1(n10069), .B2(n10845), .A(n10118), .ZN(n10119) );
  AOI21_X1 U10895 ( .B1(n10282), .B2(n4942), .A(n10119), .ZN(n10120) );
  OAI211_X1 U10896 ( .C1(n10287), .C2(n10202), .A(n10121), .B(n10120), .ZN(
        P1_U3265) );
  XNOR2_X1 U10897 ( .A(n10122), .B(n10123), .ZN(n10303) );
  XNOR2_X1 U10898 ( .A(n10124), .B(n10123), .ZN(n10301) );
  OAI211_X1 U10899 ( .C1(n4948), .C2(n5262), .A(n10818), .B(n10125), .ZN(
        n10299) );
  NAND2_X1 U10900 ( .A1(n10172), .A2(n10297), .ZN(n10129) );
  INV_X1 U10901 ( .A(n10126), .ZN(n10127) );
  AOI22_X1 U10902 ( .A1(n10697), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n10127), 
        .B2(n10730), .ZN(n10128) );
  OAI211_X1 U10903 ( .C1(n10281), .C2(n10193), .A(n10129), .B(n10128), .ZN(
        n10130) );
  AOI21_X1 U10904 ( .B1(n10131), .B2(n10732), .A(n10130), .ZN(n10132) );
  OAI21_X1 U10905 ( .B1(n10299), .B2(n10180), .A(n10132), .ZN(n10133) );
  AOI21_X1 U10906 ( .B1(n10301), .B2(n10182), .A(n10133), .ZN(n10134) );
  OAI21_X1 U10907 ( .B1(n10303), .B2(n10265), .A(n10134), .ZN(P1_U3267) );
  AOI21_X1 U10908 ( .B1(n10136), .B2(n10137), .A(n10135), .ZN(n10311) );
  XNOR2_X1 U10909 ( .A(n10138), .B(n10137), .ZN(n10304) );
  NAND2_X1 U10910 ( .A1(n10304), .A2(n10190), .ZN(n10149) );
  AOI211_X1 U10911 ( .C1(n10308), .C2(n5264), .A(n10257), .B(n4948), .ZN(
        n10306) );
  INV_X1 U10912 ( .A(n10140), .ZN(n10141) );
  AOI22_X1 U10913 ( .A1(n10697), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n10141), 
        .B2(n10730), .ZN(n10142) );
  OAI21_X1 U10914 ( .B1(n10193), .B2(n10305), .A(n10142), .ZN(n10143) );
  AOI21_X1 U10915 ( .B1(n10172), .B2(n10144), .A(n10143), .ZN(n10145) );
  OAI21_X1 U10916 ( .B1(n10146), .B2(n10845), .A(n10145), .ZN(n10147) );
  AOI21_X1 U10917 ( .B1(n10306), .B2(n4942), .A(n10147), .ZN(n10148) );
  OAI211_X1 U10918 ( .C1(n10311), .C2(n10202), .A(n10149), .B(n10148), .ZN(
        P1_U3268) );
  AOI21_X1 U10919 ( .B1(n10151), .B2(n10153), .A(n10150), .ZN(n10324) );
  XNOR2_X1 U10920 ( .A(n10152), .B(n10153), .ZN(n10317) );
  NAND2_X1 U10921 ( .A1(n10317), .A2(n10190), .ZN(n10166) );
  INV_X1 U10922 ( .A(n10155), .ZN(n10156) );
  AOI211_X1 U10923 ( .C1(n10321), .C2(n10171), .A(n10257), .B(n10156), .ZN(
        n10319) );
  OAI22_X1 U10924 ( .A1(n10852), .A2(n10158), .B1(n10157), .B2(n10847), .ZN(
        n10160) );
  NOR2_X1 U10925 ( .A1(n10193), .A2(n10318), .ZN(n10159) );
  AOI211_X1 U10926 ( .C1(n10172), .C2(n10161), .A(n10160), .B(n10159), .ZN(
        n10162) );
  OAI21_X1 U10927 ( .B1(n10163), .B2(n10845), .A(n10162), .ZN(n10164) );
  AOI21_X1 U10928 ( .B1(n10319), .B2(n4942), .A(n10164), .ZN(n10165) );
  OAI211_X1 U10929 ( .C1(n10324), .C2(n10202), .A(n10166), .B(n10165), .ZN(
        P1_U3270) );
  XNOR2_X1 U10930 ( .A(n10167), .B(n10168), .ZN(n10333) );
  XNOR2_X1 U10931 ( .A(n10169), .B(n10168), .ZN(n10331) );
  INV_X1 U10932 ( .A(n10170), .ZN(n10191) );
  OAI211_X1 U10933 ( .C1(n10329), .C2(n10191), .A(n10818), .B(n10171), .ZN(
        n10328) );
  NAND2_X1 U10934 ( .A1(n10172), .A2(n10325), .ZN(n10175) );
  AOI22_X1 U10935 ( .A1(n10697), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n10173), 
        .B2(n10730), .ZN(n10174) );
  OAI211_X1 U10936 ( .C1(n10176), .C2(n10193), .A(n10175), .B(n10174), .ZN(
        n10177) );
  AOI21_X1 U10937 ( .B1(n10178), .B2(n10732), .A(n10177), .ZN(n10179) );
  OAI21_X1 U10938 ( .B1(n10328), .B2(n10180), .A(n10179), .ZN(n10181) );
  AOI21_X1 U10939 ( .B1(n10331), .B2(n10182), .A(n10181), .ZN(n10183) );
  OAI21_X1 U10940 ( .B1(n10333), .B2(n10265), .A(n10183), .ZN(P1_U3271) );
  NAND2_X1 U10941 ( .A1(n10185), .A2(n10184), .ZN(n10187) );
  XNOR2_X1 U10942 ( .A(n10187), .B(n10186), .ZN(n10342) );
  XNOR2_X1 U10943 ( .A(n10189), .B(n10188), .ZN(n10334) );
  NAND2_X1 U10944 ( .A1(n10334), .A2(n10190), .ZN(n10201) );
  AOI211_X1 U10945 ( .C1(n10339), .C2(n10204), .A(n10257), .B(n10191), .ZN(
        n10337) );
  NAND2_X1 U10946 ( .A1(n10339), .A2(n10732), .ZN(n10197) );
  NOR2_X1 U10947 ( .A1(n10192), .A2(n10847), .ZN(n10195) );
  NOR2_X1 U10948 ( .A1(n10193), .A2(n10336), .ZN(n10194) );
  AOI211_X1 U10949 ( .C1(n10697), .C2(P1_REG2_REG_21__SCAN_IN), .A(n10195), 
        .B(n10194), .ZN(n10196) );
  OAI211_X1 U10950 ( .C1(n10335), .C2(n10198), .A(n10197), .B(n10196), .ZN(
        n10199) );
  AOI21_X1 U10951 ( .B1(n10337), .B2(n4942), .A(n10199), .ZN(n10200) );
  OAI211_X1 U10952 ( .C1(n10342), .C2(n10202), .A(n10201), .B(n10200), .ZN(
        P1_U3272) );
  XOR2_X1 U10953 ( .A(n10211), .B(n10203), .Z(n10347) );
  INV_X1 U10954 ( .A(n10204), .ZN(n10205) );
  AOI211_X1 U10955 ( .C1(n10345), .C2(n5269), .A(n10257), .B(n10205), .ZN(
        n10344) );
  NOR2_X1 U10956 ( .A1(n10206), .A2(n10845), .ZN(n10210) );
  OAI22_X1 U10957 ( .A1(n10852), .A2(n10208), .B1(n10207), .B2(n10847), .ZN(
        n10209) );
  AOI211_X1 U10958 ( .C1(n10344), .C2(n4942), .A(n10210), .B(n10209), .ZN(
        n10216) );
  XNOR2_X1 U10959 ( .A(n10212), .B(n10211), .ZN(n10213) );
  OAI222_X1 U10960 ( .A1(n10823), .A2(n10214), .B1(n10825), .B2(n10237), .C1(
        n10213), .C2(n10794), .ZN(n10343) );
  NAND2_X1 U10961 ( .A1(n10343), .A2(n10852), .ZN(n10215) );
  OAI211_X1 U10962 ( .C1(n10347), .C2(n10265), .A(n10216), .B(n10215), .ZN(
        P1_U3273) );
  XNOR2_X1 U10963 ( .A(n10217), .B(n10225), .ZN(n10352) );
  AOI211_X1 U10964 ( .C1(n10349), .C2(n10238), .A(n10257), .B(n10218), .ZN(
        n10348) );
  INV_X1 U10965 ( .A(n10219), .ZN(n10220) );
  AOI22_X1 U10966 ( .A1(n10697), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n10220), 
        .B2(n10730), .ZN(n10221) );
  OAI21_X1 U10967 ( .B1(n10222), .B2(n10845), .A(n10221), .ZN(n10230) );
  OAI21_X1 U10968 ( .B1(n10225), .B2(n10224), .A(n10223), .ZN(n10228) );
  AOI222_X1 U10969 ( .A1(n10828), .A2(n10228), .B1(n10227), .B2(n10590), .C1(
        n10226), .C2(n10747), .ZN(n10351) );
  NOR2_X1 U10970 ( .A1(n10351), .A2(n10697), .ZN(n10229) );
  AOI211_X1 U10971 ( .C1(n10348), .C2(n4942), .A(n10230), .B(n10229), .ZN(
        n10231) );
  OAI21_X1 U10972 ( .B1(n10352), .B2(n10265), .A(n10231), .ZN(P1_U3274) );
  XNOR2_X1 U10973 ( .A(n10232), .B(n10234), .ZN(n10357) );
  XOR2_X1 U10974 ( .A(n10233), .B(n10234), .Z(n10235) );
  OAI222_X1 U10975 ( .A1(n10823), .A2(n10237), .B1(n10825), .B2(n10236), .C1(
        n10235), .C2(n10794), .ZN(n10353) );
  INV_X1 U10976 ( .A(n10238), .ZN(n10239) );
  AOI211_X1 U10977 ( .C1(n10355), .C2(n10255), .A(n10257), .B(n10239), .ZN(
        n10354) );
  NAND2_X1 U10978 ( .A1(n10354), .A2(n4942), .ZN(n10243) );
  INV_X1 U10979 ( .A(n10240), .ZN(n10241) );
  AOI22_X1 U10980 ( .A1(n10697), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n10241), 
        .B2(n10730), .ZN(n10242) );
  OAI211_X1 U10981 ( .C1(n10244), .C2(n10845), .A(n10243), .B(n10242), .ZN(
        n10245) );
  AOI21_X1 U10982 ( .B1(n10353), .B2(n10852), .A(n10245), .ZN(n10246) );
  OAI21_X1 U10983 ( .B1(n10357), .B2(n10265), .A(n10246), .ZN(P1_U3275) );
  XNOR2_X1 U10984 ( .A(n10247), .B(n10248), .ZN(n10362) );
  XNOR2_X1 U10985 ( .A(n10250), .B(n10249), .ZN(n10251) );
  OAI222_X1 U10986 ( .A1(n10823), .A2(n10253), .B1(n10825), .B2(n10252), .C1(
        n10251), .C2(n10794), .ZN(n10358) );
  INV_X1 U10987 ( .A(n10254), .ZN(n10258) );
  INV_X1 U10988 ( .A(n10255), .ZN(n10256) );
  AOI211_X1 U10989 ( .C1(n10360), .C2(n10258), .A(n10257), .B(n10256), .ZN(
        n10359) );
  NAND2_X1 U10990 ( .A1(n10359), .A2(n4942), .ZN(n10261) );
  AOI22_X1 U10991 ( .A1(n10697), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n10259), 
        .B2(n10730), .ZN(n10260) );
  OAI211_X1 U10992 ( .C1(n10262), .C2(n10845), .A(n10261), .B(n10260), .ZN(
        n10263) );
  AOI21_X1 U10993 ( .B1(n10358), .B2(n10852), .A(n10263), .ZN(n10264) );
  OAI21_X1 U10994 ( .B1(n10362), .B2(n10265), .A(n10264), .ZN(P1_U3276) );
  OAI211_X1 U10995 ( .C1(n10267), .C2(n10820), .A(n10266), .B(n10268), .ZN(
        n10378) );
  MUX2_X1 U10996 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10378), .S(n10665), .Z(
        P1_U3553) );
  OAI211_X1 U10997 ( .C1(n10270), .C2(n10820), .A(n10269), .B(n10268), .ZN(
        n10379) );
  MUX2_X1 U10998 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10379), .S(n10665), .Z(
        P1_U3552) );
  NAND2_X1 U10999 ( .A1(n10271), .A2(n10811), .ZN(n10278) );
  NAND2_X1 U11000 ( .A1(n10272), .A2(n10791), .ZN(n10274) );
  OAI211_X1 U11001 ( .C1(n10288), .C2(n10825), .A(n10274), .B(n10273), .ZN(
        n10275) );
  MUX2_X1 U11002 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10380), .S(n10665), .Z(
        P1_U3551) );
  NAND2_X1 U11003 ( .A1(n10279), .A2(n10811), .ZN(n10286) );
  OAI22_X1 U11004 ( .A1(n10281), .A2(n10825), .B1(n10280), .B2(n10823), .ZN(
        n10283) );
  AOI211_X1 U11005 ( .C1(n10791), .C2(n10284), .A(n10283), .B(n10282), .ZN(
        n10285) );
  OAI211_X1 U11006 ( .C1(n10794), .C2(n10287), .A(n10286), .B(n10285), .ZN(
        n10381) );
  MUX2_X1 U11007 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10381), .S(n10665), .Z(
        P1_U3550) );
  INV_X1 U11008 ( .A(n10811), .ZN(n10644) );
  OAI22_X1 U11009 ( .A1(n10305), .A2(n10825), .B1(n10288), .B2(n10823), .ZN(
        n10290) );
  AOI211_X1 U11010 ( .C1(n10791), .C2(n10291), .A(n10290), .B(n10289), .ZN(
        n10294) );
  NAND2_X1 U11011 ( .A1(n10292), .A2(n10828), .ZN(n10293) );
  OAI211_X1 U11012 ( .C1(n10295), .C2(n10644), .A(n10294), .B(n10293), .ZN(
        n10382) );
  MUX2_X1 U11013 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10382), .S(n10665), .Z(
        P1_U3549) );
  AOI22_X1 U11014 ( .A1(n10747), .A2(n10297), .B1(n10296), .B2(n10590), .ZN(
        n10298) );
  OAI211_X1 U11015 ( .C1(n5262), .C2(n10820), .A(n10299), .B(n10298), .ZN(
        n10300) );
  AOI21_X1 U11016 ( .B1(n10301), .B2(n10828), .A(n10300), .ZN(n10302) );
  OAI21_X1 U11017 ( .B1(n10303), .B2(n10644), .A(n10302), .ZN(n10383) );
  MUX2_X1 U11018 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10383), .S(n10665), .Z(
        P1_U3548) );
  NAND2_X1 U11019 ( .A1(n10304), .A2(n10811), .ZN(n10310) );
  OAI22_X1 U11020 ( .A1(n10318), .A2(n10825), .B1(n10305), .B2(n10823), .ZN(
        n10307) );
  AOI211_X1 U11021 ( .C1(n10791), .C2(n10308), .A(n10307), .B(n10306), .ZN(
        n10309) );
  OAI211_X1 U11022 ( .C1(n10794), .C2(n10311), .A(n10310), .B(n10309), .ZN(
        n10384) );
  MUX2_X1 U11023 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10384), .S(n10665), .Z(
        P1_U3547) );
  AOI211_X1 U11024 ( .C1(n10791), .C2(n10314), .A(n10313), .B(n10312), .ZN(
        n10315) );
  OAI21_X1 U11025 ( .B1(n10316), .B2(n10644), .A(n10315), .ZN(n10385) );
  MUX2_X1 U11026 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10385), .S(n10665), .Z(
        P1_U3546) );
  NAND2_X1 U11027 ( .A1(n10317), .A2(n10811), .ZN(n10323) );
  OAI22_X1 U11028 ( .A1(n10336), .A2(n10825), .B1(n10318), .B2(n10823), .ZN(
        n10320) );
  AOI211_X1 U11029 ( .C1(n10791), .C2(n10321), .A(n10320), .B(n10319), .ZN(
        n10322) );
  OAI211_X1 U11030 ( .C1(n10794), .C2(n10324), .A(n10323), .B(n10322), .ZN(
        n10386) );
  MUX2_X1 U11031 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10386), .S(n10665), .Z(
        P1_U3545) );
  AOI22_X1 U11032 ( .A1(n10326), .A2(n10590), .B1(n10747), .B2(n10325), .ZN(
        n10327) );
  OAI211_X1 U11033 ( .C1(n10329), .C2(n10820), .A(n10328), .B(n10327), .ZN(
        n10330) );
  AOI21_X1 U11034 ( .B1(n10331), .B2(n10828), .A(n10330), .ZN(n10332) );
  OAI21_X1 U11035 ( .B1(n10333), .B2(n10644), .A(n10332), .ZN(n10387) );
  MUX2_X1 U11036 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10387), .S(n10665), .Z(
        P1_U3544) );
  NAND2_X1 U11037 ( .A1(n10334), .A2(n10811), .ZN(n10341) );
  OAI22_X1 U11038 ( .A1(n10336), .A2(n10823), .B1(n10335), .B2(n10825), .ZN(
        n10338) );
  AOI211_X1 U11039 ( .C1(n10791), .C2(n10339), .A(n10338), .B(n10337), .ZN(
        n10340) );
  OAI211_X1 U11040 ( .C1(n10794), .C2(n10342), .A(n10341), .B(n10340), .ZN(
        n10388) );
  MUX2_X1 U11041 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10388), .S(n10665), .Z(
        P1_U3543) );
  AOI211_X1 U11042 ( .C1(n10791), .C2(n10345), .A(n10344), .B(n10343), .ZN(
        n10346) );
  OAI21_X1 U11043 ( .B1(n10347), .B2(n10644), .A(n10346), .ZN(n10389) );
  MUX2_X1 U11044 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10389), .S(n10665), .Z(
        P1_U3542) );
  AOI21_X1 U11045 ( .B1(n10791), .B2(n10349), .A(n10348), .ZN(n10350) );
  OAI211_X1 U11046 ( .C1(n10352), .C2(n10644), .A(n10351), .B(n10350), .ZN(
        n10390) );
  MUX2_X1 U11047 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10390), .S(n10665), .Z(
        P1_U3541) );
  AOI211_X1 U11048 ( .C1(n10791), .C2(n10355), .A(n10354), .B(n10353), .ZN(
        n10356) );
  OAI21_X1 U11049 ( .B1(n10357), .B2(n10644), .A(n10356), .ZN(n10391) );
  MUX2_X1 U11050 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10391), .S(n10665), .Z(
        P1_U3540) );
  AOI211_X1 U11051 ( .C1(n10791), .C2(n10360), .A(n10359), .B(n10358), .ZN(
        n10361) );
  OAI21_X1 U11052 ( .B1(n10362), .B2(n10644), .A(n10361), .ZN(n10392) );
  MUX2_X1 U11053 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10392), .S(n10665), .Z(
        P1_U3539) );
  AOI211_X1 U11054 ( .C1(n10791), .C2(n10365), .A(n10364), .B(n10363), .ZN(
        n10366) );
  OAI21_X1 U11055 ( .B1(n10367), .B2(n10644), .A(n10366), .ZN(n10393) );
  MUX2_X1 U11056 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10393), .S(n10665), .Z(
        P1_U3538) );
  AOI22_X1 U11057 ( .A1(n10747), .A2(n10369), .B1(n10368), .B2(n10590), .ZN(
        n10370) );
  OAI21_X1 U11058 ( .B1(n10371), .B2(n10820), .A(n10370), .ZN(n10373) );
  AOI211_X1 U11059 ( .C1(n10828), .C2(n10374), .A(n10373), .B(n10372), .ZN(
        n10375) );
  OAI21_X1 U11060 ( .B1(n10376), .B2(n10644), .A(n10375), .ZN(n10394) );
  MUX2_X1 U11061 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10394), .S(n10665), .Z(
        P1_U3537) );
  MUX2_X1 U11062 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10377), .S(n10665), .Z(
        P1_U3523) );
  MUX2_X1 U11063 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10378), .S(n10839), .Z(
        P1_U3521) );
  MUX2_X1 U11064 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10379), .S(n10839), .Z(
        P1_U3520) );
  MUX2_X1 U11065 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10380), .S(n10839), .Z(
        P1_U3519) );
  MUX2_X1 U11066 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10381), .S(n10839), .Z(
        P1_U3518) );
  MUX2_X1 U11067 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10382), .S(n10839), .Z(
        P1_U3517) );
  MUX2_X1 U11068 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10383), .S(n10839), .Z(
        P1_U3516) );
  MUX2_X1 U11069 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10384), .S(n10839), .Z(
        P1_U3515) );
  MUX2_X1 U11070 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10385), .S(n10839), .Z(
        P1_U3514) );
  MUX2_X1 U11071 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10386), .S(n10839), .Z(
        P1_U3513) );
  MUX2_X1 U11072 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10387), .S(n10839), .Z(
        P1_U3512) );
  MUX2_X1 U11073 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10388), .S(n10839), .Z(
        P1_U3511) );
  MUX2_X1 U11074 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10389), .S(n10839), .Z(
        P1_U3510) );
  MUX2_X1 U11075 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10390), .S(n10839), .Z(
        P1_U3509) );
  MUX2_X1 U11076 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10391), .S(n10839), .Z(
        P1_U3507) );
  MUX2_X1 U11077 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10392), .S(n10839), .Z(
        P1_U3504) );
  MUX2_X1 U11078 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10393), .S(n10839), .Z(
        P1_U3501) );
  MUX2_X1 U11079 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10394), .S(n10839), .Z(
        P1_U3498) );
  MUX2_X1 U11080 ( .A(n10395), .B(P1_D_REG_0__SCAN_IN), .S(n10408), .Z(
        P1_U3439) );
  NOR4_X1 U11081 ( .A1(n10397), .A2(P1_IR_REG_30__SCAN_IN), .A3(n10396), .A4(
        P1_U3086), .ZN(n10398) );
  AOI21_X1 U11082 ( .B1(n10399), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10398), 
        .ZN(n10400) );
  OAI21_X1 U11083 ( .B1(n10401), .B2(n10404), .A(n10400), .ZN(P1_U3324) );
  OAI222_X1 U11084 ( .A1(n10406), .A2(n10405), .B1(n10404), .B2(n10403), .C1(
        n10402), .C2(P1_U3086), .ZN(P1_U3326) );
  MUX2_X1 U11085 ( .A(n10407), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AND2_X1 U11086 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10408), .ZN(P1_U3323) );
  AND2_X1 U11087 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10408), .ZN(P1_U3322) );
  AND2_X1 U11088 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10408), .ZN(P1_U3321) );
  AND2_X1 U11089 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10408), .ZN(P1_U3320) );
  AND2_X1 U11090 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10408), .ZN(P1_U3319) );
  AND2_X1 U11091 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10408), .ZN(P1_U3318) );
  AND2_X1 U11092 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10408), .ZN(P1_U3317) );
  AND2_X1 U11093 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10408), .ZN(P1_U3316) );
  AND2_X1 U11094 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10408), .ZN(P1_U3315) );
  AND2_X1 U11095 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10408), .ZN(P1_U3314) );
  AND2_X1 U11096 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10408), .ZN(P1_U3313) );
  AND2_X1 U11097 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10408), .ZN(P1_U3312) );
  AND2_X1 U11098 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10408), .ZN(P1_U3311) );
  AND2_X1 U11099 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10408), .ZN(P1_U3310) );
  AND2_X1 U11100 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10408), .ZN(P1_U3309) );
  AND2_X1 U11101 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10408), .ZN(P1_U3308) );
  AND2_X1 U11102 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10408), .ZN(P1_U3307) );
  AND2_X1 U11103 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10408), .ZN(P1_U3306) );
  AND2_X1 U11104 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10408), .ZN(P1_U3305) );
  AND2_X1 U11105 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10408), .ZN(P1_U3304) );
  AND2_X1 U11106 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10408), .ZN(P1_U3303) );
  AND2_X1 U11107 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10408), .ZN(P1_U3302) );
  AND2_X1 U11108 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10408), .ZN(P1_U3301) );
  AND2_X1 U11109 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10408), .ZN(P1_U3300) );
  AND2_X1 U11110 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10408), .ZN(P1_U3299) );
  AND2_X1 U11111 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10408), .ZN(P1_U3298) );
  AND2_X1 U11112 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10408), .ZN(P1_U3297) );
  AND2_X1 U11113 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10408), .ZN(P1_U3296) );
  AND2_X1 U11114 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10408), .ZN(P1_U3295) );
  AND2_X1 U11115 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10408), .ZN(P1_U3294) );
  NAND2_X1 U11116 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .ZN(n10412) );
  OAI21_X1 U11117 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(n10412), .ZN(n10409) );
  INV_X1 U11118 ( .A(n10409), .ZN(ADD_1068_U46) );
  INV_X1 U11119 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10410) );
  NAND2_X1 U11120 ( .A1(n10410), .A2(n10412), .ZN(n10413) );
  OAI21_X1 U11121 ( .B1(n10410), .B2(n10412), .A(n10413), .ZN(n10411) );
  XNOR2_X1 U11122 ( .A(n10411), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(ADD_1068_U5)
         );
  INV_X1 U11123 ( .A(n10412), .ZN(n10414) );
  AOI22_X1 U11124 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n10414), .B1(
        P2_ADDR_REG_1__SCAN_IN), .B2(n10413), .ZN(n10417) );
  NAND2_X1 U11125 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10415) );
  OAI21_X1 U11126 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10415), .ZN(n10416) );
  NOR2_X1 U11127 ( .A1(n10417), .A2(n10416), .ZN(n10418) );
  AOI21_X1 U11128 ( .B1(n10417), .B2(n10416), .A(n10418), .ZN(ADD_1068_U54) );
  AOI21_X1 U11129 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10418), .ZN(n10421) );
  NAND2_X1 U11130 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n10419) );
  OAI21_X1 U11131 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10419), .ZN(n10420) );
  NOR2_X1 U11132 ( .A1(n10421), .A2(n10420), .ZN(n10422) );
  AOI21_X1 U11133 ( .B1(n10421), .B2(n10420), .A(n10422), .ZN(ADD_1068_U53) );
  AOI21_X1 U11134 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10422), .ZN(n10425) );
  NOR2_X1 U11135 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10423) );
  AOI21_X1 U11136 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n10423), .ZN(n10424) );
  NAND2_X1 U11137 ( .A1(n10425), .A2(n10424), .ZN(n10427) );
  OAI21_X1 U11138 ( .B1(n10425), .B2(n10424), .A(n10427), .ZN(ADD_1068_U52) );
  NOR2_X1 U11139 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10426) );
  AOI21_X1 U11140 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10426), .ZN(n10429) );
  OAI21_X1 U11141 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10427), .ZN(n10428) );
  NAND2_X1 U11142 ( .A1(n10429), .A2(n10428), .ZN(n10431) );
  OAI21_X1 U11143 ( .B1(n10429), .B2(n10428), .A(n10431), .ZN(ADD_1068_U51) );
  NOR2_X1 U11144 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10430) );
  AOI21_X1 U11145 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n10430), .ZN(n10433) );
  OAI21_X1 U11146 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10431), .ZN(n10432) );
  NAND2_X1 U11147 ( .A1(n10433), .A2(n10432), .ZN(n10435) );
  OAI21_X1 U11148 ( .B1(n10433), .B2(n10432), .A(n10435), .ZN(ADD_1068_U50) );
  NOR2_X1 U11149 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10434) );
  AOI21_X1 U11150 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n10434), .ZN(n10437) );
  OAI21_X1 U11151 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10435), .ZN(n10436) );
  NAND2_X1 U11152 ( .A1(n10437), .A2(n10436), .ZN(n10439) );
  OAI21_X1 U11153 ( .B1(n10437), .B2(n10436), .A(n10439), .ZN(ADD_1068_U49) );
  NOR2_X1 U11154 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10438) );
  AOI21_X1 U11155 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n10438), .ZN(n10441) );
  OAI21_X1 U11156 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10439), .ZN(n10440) );
  NAND2_X1 U11157 ( .A1(n10441), .A2(n10440), .ZN(n10443) );
  OAI21_X1 U11158 ( .B1(n10441), .B2(n10440), .A(n10443), .ZN(ADD_1068_U48) );
  NOR2_X1 U11159 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10442) );
  AOI21_X1 U11160 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n10442), .ZN(n10445) );
  OAI21_X1 U11161 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10443), .ZN(n10444) );
  NAND2_X1 U11162 ( .A1(n10445), .A2(n10444), .ZN(n10447) );
  OAI21_X1 U11163 ( .B1(n10445), .B2(n10444), .A(n10447), .ZN(ADD_1068_U47) );
  NOR2_X1 U11164 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10446) );
  AOI21_X1 U11165 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10446), .ZN(n10449) );
  OAI21_X1 U11166 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10447), .ZN(n10448) );
  NAND2_X1 U11167 ( .A1(n10449), .A2(n10448), .ZN(n10451) );
  OAI21_X1 U11168 ( .B1(n10449), .B2(n10448), .A(n10451), .ZN(ADD_1068_U63) );
  NOR2_X1 U11169 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10450) );
  AOI21_X1 U11170 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10450), .ZN(n10453) );
  OAI21_X1 U11171 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10451), .ZN(n10452) );
  NAND2_X1 U11172 ( .A1(n10453), .A2(n10452), .ZN(n10455) );
  OAI21_X1 U11173 ( .B1(n10453), .B2(n10452), .A(n10455), .ZN(ADD_1068_U62) );
  NOR2_X1 U11174 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10454) );
  AOI21_X1 U11175 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10454), .ZN(n10457) );
  OAI21_X1 U11176 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10455), .ZN(n10456) );
  NAND2_X1 U11177 ( .A1(n10457), .A2(n10456), .ZN(n10459) );
  OAI21_X1 U11178 ( .B1(n10457), .B2(n10456), .A(n10459), .ZN(ADD_1068_U61) );
  NOR2_X1 U11179 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10458) );
  AOI21_X1 U11180 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10458), .ZN(n10461) );
  OAI21_X1 U11181 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10459), .ZN(n10460) );
  NAND2_X1 U11182 ( .A1(n10461), .A2(n10460), .ZN(n10463) );
  OAI21_X1 U11183 ( .B1(n10461), .B2(n10460), .A(n10463), .ZN(ADD_1068_U60) );
  NOR2_X1 U11184 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10462) );
  AOI21_X1 U11185 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10462), .ZN(n10465) );
  OAI21_X1 U11186 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10463), .ZN(n10464) );
  NAND2_X1 U11187 ( .A1(n10465), .A2(n10464), .ZN(n10467) );
  OAI21_X1 U11188 ( .B1(n10465), .B2(n10464), .A(n10467), .ZN(ADD_1068_U59) );
  NOR2_X1 U11189 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10466) );
  AOI21_X1 U11190 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10466), .ZN(n10469) );
  OAI21_X1 U11191 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10467), .ZN(n10468) );
  NAND2_X1 U11192 ( .A1(n10469), .A2(n10468), .ZN(n10471) );
  OAI21_X1 U11193 ( .B1(n10469), .B2(n10468), .A(n10471), .ZN(ADD_1068_U58) );
  NOR2_X1 U11194 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10470) );
  AOI21_X1 U11195 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10470), .ZN(n10473) );
  OAI21_X1 U11196 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10471), .ZN(n10472) );
  NAND2_X1 U11197 ( .A1(n10473), .A2(n10472), .ZN(n10475) );
  OAI21_X1 U11198 ( .B1(n10473), .B2(n10472), .A(n10475), .ZN(ADD_1068_U57) );
  NOR2_X1 U11199 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10474) );
  AOI21_X1 U11200 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10474), .ZN(n10477) );
  OAI21_X1 U11201 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10475), .ZN(n10476) );
  NAND2_X1 U11202 ( .A1(n10477), .A2(n10476), .ZN(n10480) );
  OAI21_X1 U11203 ( .B1(n10477), .B2(n10476), .A(n10480), .ZN(ADD_1068_U56) );
  INV_X1 U11204 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10478) );
  AOI22_X1 U11205 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P1_ADDR_REG_18__SCAN_IN), 
        .B1(n10479), .B2(n10478), .ZN(n10482) );
  OAI21_X1 U11206 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10480), .ZN(n10481) );
  NAND2_X1 U11207 ( .A1(n10482), .A2(n10481), .ZN(n10483) );
  OAI21_X1 U11208 ( .B1(n10482), .B2(n10481), .A(n10483), .ZN(ADD_1068_U55) );
  OAI21_X1 U11209 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10483), .ZN(n10485) );
  XOR2_X1 U11210 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n10484) );
  XNOR2_X1 U11211 ( .A(n10485), .B(n10484), .ZN(ADD_1068_U4) );
  AOI22_X1 U11212 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(n10571), .B1(n10572), .B2(
        P2_ADDR_REG_0__SCAN_IN), .ZN(n10492) );
  INV_X1 U11213 ( .A(n10486), .ZN(n10490) );
  NOR2_X1 U11214 ( .A1(n10487), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n10488) );
  OAI22_X1 U11215 ( .A1(n10490), .A2(n10579), .B1(n10489), .B2(n10488), .ZN(
        n10491) );
  OAI211_X1 U11216 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6893), .A(n10492), .B(
        n10491), .ZN(P2_U3182) );
  INV_X1 U11217 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10513) );
  OAI21_X1 U11218 ( .B1(n10495), .B2(n10494), .A(n10493), .ZN(n10507) );
  INV_X1 U11219 ( .A(n10496), .ZN(n10499) );
  INV_X1 U11220 ( .A(n10497), .ZN(n10498) );
  NAND2_X1 U11221 ( .A1(n10499), .A2(n10498), .ZN(n10500) );
  AND2_X1 U11222 ( .A1(n10501), .A2(n10500), .ZN(n10502) );
  OAI22_X1 U11223 ( .A1(n10559), .A2(n10502), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10619), .ZN(n10506) );
  NOR2_X1 U11224 ( .A1(n10504), .A2(n10503), .ZN(n10505) );
  AOI211_X1 U11225 ( .C1(n10583), .C2(n10507), .A(n10506), .B(n10505), .ZN(
        n10512) );
  XOR2_X1 U11226 ( .A(n10509), .B(n10508), .Z(n10510) );
  NAND2_X1 U11227 ( .A1(n10510), .A2(n10579), .ZN(n10511) );
  OAI211_X1 U11228 ( .C1(n10513), .C2(n10569), .A(n10512), .B(n10511), .ZN(
        P2_U3184) );
  INV_X1 U11229 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10531) );
  AOI21_X1 U11230 ( .B1(n10515), .B2(n5768), .A(n10514), .ZN(n10523) );
  OAI21_X1 U11231 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n10517), .A(n10516), .ZN(
        n10519) );
  AOI21_X1 U11232 ( .B1(n10580), .B2(n10519), .A(n10518), .ZN(n10522) );
  NAND2_X1 U11233 ( .A1(n10571), .A2(n10520), .ZN(n10521) );
  OAI211_X1 U11234 ( .C1(n10523), .C2(n10561), .A(n10522), .B(n10521), .ZN(
        n10524) );
  INV_X1 U11235 ( .A(n10524), .ZN(n10530) );
  OAI21_X1 U11236 ( .B1(n10527), .B2(n10526), .A(n10525), .ZN(n10528) );
  NAND2_X1 U11237 ( .A1(n10528), .A2(n10579), .ZN(n10529) );
  OAI211_X1 U11238 ( .C1(n10531), .C2(n10569), .A(n10530), .B(n10529), .ZN(
        P2_U3185) );
  INV_X1 U11239 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10550) );
  AOI21_X1 U11240 ( .B1(n10534), .B2(n10533), .A(n10532), .ZN(n10541) );
  OAI21_X1 U11241 ( .B1(n10537), .B2(n10536), .A(n10535), .ZN(n10539) );
  AOI21_X1 U11242 ( .B1(n10580), .B2(n10539), .A(n10538), .ZN(n10540) );
  OAI21_X1 U11243 ( .B1(n10541), .B2(n10561), .A(n10540), .ZN(n10542) );
  AOI21_X1 U11244 ( .B1(n10543), .B2(n10571), .A(n10542), .ZN(n10549) );
  AOI211_X1 U11245 ( .C1(n10546), .C2(n10545), .A(n10562), .B(n10544), .ZN(
        n10547) );
  INV_X1 U11246 ( .A(n10547), .ZN(n10548) );
  OAI211_X1 U11247 ( .C1(n10550), .C2(n10569), .A(n10549), .B(n10548), .ZN(
        P2_U3186) );
  INV_X1 U11248 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10568) );
  XNOR2_X1 U11249 ( .A(n10552), .B(n10551), .ZN(n10563) );
  AOI21_X1 U11250 ( .B1(n5811), .B2(n10554), .A(n10553), .ZN(n10560) );
  OAI21_X1 U11251 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(n10556), .A(n10555), .ZN(
        n10557) );
  INV_X1 U11252 ( .A(n10557), .ZN(n10558) );
  OAI222_X1 U11253 ( .A1(n10563), .A2(n10562), .B1(n10561), .B2(n10560), .C1(
        n10559), .C2(n10558), .ZN(n10564) );
  AOI211_X1 U11254 ( .C1(n10566), .C2(n10571), .A(n10565), .B(n10564), .ZN(
        n10567) );
  OAI21_X1 U11255 ( .B1(n10569), .B2(n10568), .A(n10567), .ZN(P2_U3187) );
  AOI22_X1 U11256 ( .A1(n10572), .A2(P2_ADDR_REG_11__SCAN_IN), .B1(n10571), 
        .B2(n10570), .ZN(n10588) );
  OAI21_X1 U11257 ( .B1(n10574), .B2(P2_REG1_REG_11__SCAN_IN), .A(n10573), 
        .ZN(n10581) );
  OAI21_X1 U11258 ( .B1(n10577), .B2(n10576), .A(n10575), .ZN(n10578) );
  AOI22_X1 U11259 ( .A1(n10581), .A2(n10580), .B1(n10579), .B2(n10578), .ZN(
        n10587) );
  NAND2_X1 U11260 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3151), .ZN(n10586)
         );
  XNOR2_X1 U11261 ( .A(n10582), .B(n5894), .ZN(n10584) );
  NAND2_X1 U11262 ( .A1(n10584), .A2(n10583), .ZN(n10585) );
  NAND4_X1 U11263 ( .A1(n10588), .A2(n10587), .A3(n10586), .A4(n10585), .ZN(
        P2_U3193) );
  XNOR2_X1 U11264 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11265 ( .A(n10589), .ZN(n10595) );
  NAND2_X1 U11266 ( .A1(n10644), .A2(n10794), .ZN(n10594) );
  AOI222_X1 U11267 ( .A1(n10595), .A2(n10594), .B1(n10593), .B2(n10592), .C1(
        n10591), .C2(n10590), .ZN(n10597) );
  INV_X1 U11268 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10596) );
  AOI22_X1 U11269 ( .A1(n10665), .A2(n10597), .B1(n10596), .B2(n10835), .ZN(
        P1_U3522) );
  AOI22_X1 U11270 ( .A1(n10839), .A2(n10597), .B1(n6596), .B2(n10836), .ZN(
        P1_U3453) );
  OAI22_X1 U11271 ( .A1(n10599), .A2(n10767), .B1(n10598), .B2(n10650), .ZN(
        n10600) );
  NOR2_X1 U11272 ( .A1(n10601), .A2(n10600), .ZN(n10602) );
  AOI22_X1 U11273 ( .A1(n10781), .A2(n10602), .B1(n6552), .B2(n10780), .ZN(
        P2_U3460) );
  AOI22_X1 U11274 ( .A1(n10785), .A2(n10602), .B1(n5736), .B2(n10782), .ZN(
        P2_U3393) );
  AOI22_X1 U11275 ( .A1(n10839), .A2(n10603), .B1(n6814), .B2(n10836), .ZN(
        P1_U3459) );
  OAI21_X1 U11276 ( .B1(n10606), .B2(n10605), .A(n10604), .ZN(n10610) );
  AOI222_X1 U11277 ( .A1(n10611), .A2(n10610), .B1(n10609), .B2(n10608), .C1(
        n6754), .C2(n10607), .ZN(n10621) );
  XNOR2_X1 U11278 ( .A(n8510), .B(n10612), .ZN(n10624) );
  NAND2_X1 U11279 ( .A1(n10624), .A2(n10632), .ZN(n10613) );
  OAI211_X1 U11280 ( .C1(n10618), .C2(n10650), .A(n10621), .B(n10613), .ZN(
        n10615) );
  OAI22_X1 U11281 ( .A1(n10780), .A2(n10615), .B1(P2_REG1_REG_2__SCAN_IN), 
        .B2(n10781), .ZN(n10614) );
  INV_X1 U11282 ( .A(n10614), .ZN(P2_U3461) );
  OAI22_X1 U11283 ( .A1(n10782), .A2(n10615), .B1(P2_REG0_REG_2__SCAN_IN), 
        .B2(n10785), .ZN(n10616) );
  INV_X1 U11284 ( .A(n10616), .ZN(P2_U3396) );
  OAI22_X1 U11285 ( .A1(n10620), .A2(n10619), .B1(n10618), .B2(n10617), .ZN(
        n10623) );
  INV_X1 U11286 ( .A(n10621), .ZN(n10622) );
  AOI211_X1 U11287 ( .C1(n10625), .C2(n10624), .A(n10623), .B(n10622), .ZN(
        n10627) );
  AOI22_X1 U11288 ( .A1(n9163), .A2(n6666), .B1(n10627), .B2(n10626), .ZN(
        P2_U3231) );
  NOR2_X1 U11289 ( .A1(n10650), .A2(n10628), .ZN(n10630) );
  AOI211_X1 U11290 ( .C1(n10632), .C2(n10631), .A(n10630), .B(n10629), .ZN(
        n10634) );
  AOI22_X1 U11291 ( .A1(n10781), .A2(n10634), .B1(n5767), .B2(n10780), .ZN(
        P2_U3462) );
  INV_X1 U11292 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10633) );
  AOI22_X1 U11293 ( .A1(n10785), .A2(n10634), .B1(n10633), .B2(n10782), .ZN(
        P2_U3399) );
  INV_X1 U11294 ( .A(n10635), .ZN(n10639) );
  OAI22_X1 U11295 ( .A1(n10637), .A2(n10774), .B1(n10636), .B2(n10650), .ZN(
        n10638) );
  NOR2_X1 U11296 ( .A1(n10639), .A2(n10638), .ZN(n10640) );
  AOI22_X1 U11297 ( .A1(n10781), .A2(n10640), .B1(n6635), .B2(n10780), .ZN(
        P2_U3463) );
  AOI22_X1 U11298 ( .A1(n10785), .A2(n10640), .B1(n5793), .B2(n10782), .ZN(
        P2_U3402) );
  AND2_X1 U11299 ( .A1(n10641), .A2(n10791), .ZN(n10642) );
  NOR2_X1 U11300 ( .A1(n10643), .A2(n10642), .ZN(n10647) );
  OR2_X1 U11301 ( .A1(n10645), .A2(n10644), .ZN(n10646) );
  AND3_X1 U11302 ( .A1(n10648), .A2(n10647), .A3(n10646), .ZN(n10649) );
  AOI22_X1 U11303 ( .A1(n10665), .A2(n10649), .B1(n7025), .B2(n10835), .ZN(
        P1_U3526) );
  AOI22_X1 U11304 ( .A1(n10839), .A2(n10649), .B1(n7018), .B2(n10836), .ZN(
        P1_U3465) );
  NOR2_X1 U11305 ( .A1(n10651), .A2(n10650), .ZN(n10653) );
  AOI211_X1 U11306 ( .C1(n10655), .C2(n10654), .A(n10653), .B(n10652), .ZN(
        n10657) );
  AOI22_X1 U11307 ( .A1(n10781), .A2(n10657), .B1(n5808), .B2(n10780), .ZN(
        P2_U3464) );
  INV_X1 U11308 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10656) );
  AOI22_X1 U11309 ( .A1(n10785), .A2(n10657), .B1(n10656), .B2(n10782), .ZN(
        P2_U3405) );
  AND2_X1 U11310 ( .A1(n10658), .A2(n10811), .ZN(n10663) );
  OAI21_X1 U11311 ( .B1(n10660), .B2(n10820), .A(n10659), .ZN(n10661) );
  NOR3_X1 U11312 ( .A1(n10663), .A2(n10662), .A3(n10661), .ZN(n10666) );
  INV_X1 U11313 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10664) );
  AOI22_X1 U11314 ( .A1(n10665), .A2(n10666), .B1(n10664), .B2(n10835), .ZN(
        P1_U3527) );
  AOI22_X1 U11315 ( .A1(n10839), .A2(n10666), .B1(n7206), .B2(n10836), .ZN(
        P1_U3468) );
  NOR2_X1 U11316 ( .A1(n10667), .A2(n10774), .ZN(n10669) );
  AOI211_X1 U11317 ( .C1(n10779), .C2(n10670), .A(n10669), .B(n10668), .ZN(
        n10672) );
  AOI22_X1 U11318 ( .A1(n10781), .A2(n10672), .B1(n6647), .B2(n10780), .ZN(
        P2_U3465) );
  INV_X1 U11319 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10671) );
  AOI22_X1 U11320 ( .A1(n10785), .A2(n10672), .B1(n10671), .B2(n10782), .ZN(
        P2_U3408) );
  INV_X1 U11321 ( .A(n10673), .ZN(n10834) );
  NAND2_X1 U11322 ( .A1(n7501), .A2(n10674), .ZN(n10676) );
  NAND2_X1 U11323 ( .A1(n10676), .A2(n10675), .ZN(n10677) );
  XNOR2_X1 U11324 ( .A(n10677), .B(n10683), .ZN(n10701) );
  OAI211_X1 U11325 ( .C1(n10679), .C2(n10680), .A(n10818), .B(n10678), .ZN(
        n10699) );
  OAI21_X1 U11326 ( .B1(n10680), .B2(n10820), .A(n10699), .ZN(n10693) );
  OAI22_X1 U11327 ( .A1(n10720), .A2(n10823), .B1(n10681), .B2(n10825), .ZN(
        n10690) );
  INV_X1 U11328 ( .A(n5043), .ZN(n10688) );
  AOI21_X1 U11329 ( .B1(n10685), .B2(n10684), .A(n7499), .ZN(n10686) );
  AOI211_X1 U11330 ( .C1(n10688), .C2(n10687), .A(n10794), .B(n10686), .ZN(
        n10689) );
  AOI211_X1 U11331 ( .C1(n10691), .C2(n10701), .A(n10690), .B(n10689), .ZN(
        n10704) );
  INV_X1 U11332 ( .A(n10704), .ZN(n10692) );
  AOI211_X1 U11333 ( .C1(n10834), .C2(n10701), .A(n10693), .B(n10692), .ZN(
        n10694) );
  AOI22_X1 U11334 ( .A1(n10665), .A2(n10694), .B1(n6479), .B2(n10835), .ZN(
        P1_U3528) );
  AOI22_X1 U11335 ( .A1(n10839), .A2(n10694), .B1(n6448), .B2(n10836), .ZN(
        P1_U3471) );
  INV_X1 U11336 ( .A(n10695), .ZN(n10696) );
  AOI222_X1 U11337 ( .A1(n10698), .A2(n10732), .B1(P1_REG2_REG_6__SCAN_IN), 
        .B2(n10697), .C1(n10730), .C2(n10696), .ZN(n10703) );
  INV_X1 U11338 ( .A(n10699), .ZN(n10700) );
  AOI22_X1 U11339 ( .A1(n10701), .A2(n10843), .B1(n4942), .B2(n10700), .ZN(
        n10702) );
  OAI211_X1 U11340 ( .C1(n10697), .C2(n10704), .A(n10703), .B(n10702), .ZN(
        P1_U3287) );
  OAI21_X1 U11341 ( .B1(n5271), .B2(n10820), .A(n10705), .ZN(n10706) );
  AOI21_X1 U11342 ( .B1(n10707), .B2(n10834), .A(n10706), .ZN(n10708) );
  AND2_X1 U11343 ( .A1(n10709), .A2(n10708), .ZN(n10711) );
  INV_X1 U11344 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10710) );
  AOI22_X1 U11345 ( .A1(n10665), .A2(n10711), .B1(n10710), .B2(n10835), .ZN(
        P1_U3529) );
  AOI22_X1 U11346 ( .A1(n10839), .A2(n10711), .B1(n7275), .B2(n10836), .ZN(
        P1_U3474) );
  XOR2_X1 U11347 ( .A(n10712), .B(n10718), .Z(n10721) );
  INV_X1 U11348 ( .A(n10721), .ZN(n10736) );
  INV_X1 U11349 ( .A(n10713), .ZN(n10715) );
  OAI211_X1 U11350 ( .C1(n10715), .C2(n5270), .A(n10818), .B(n10714), .ZN(
        n10734) );
  OAI21_X1 U11351 ( .B1(n5270), .B2(n10820), .A(n10734), .ZN(n10726) );
  NAND2_X1 U11352 ( .A1(n10717), .A2(n10716), .ZN(n10719) );
  XNOR2_X1 U11353 ( .A(n10719), .B(n10718), .ZN(n10724) );
  OAI22_X1 U11354 ( .A1(n10720), .A2(n10825), .B1(n10757), .B2(n10823), .ZN(
        n10723) );
  NOR2_X1 U11355 ( .A1(n10721), .A2(n10831), .ZN(n10722) );
  AOI211_X1 U11356 ( .C1(n10724), .C2(n10828), .A(n10723), .B(n10722), .ZN(
        n10739) );
  INV_X1 U11357 ( .A(n10739), .ZN(n10725) );
  AOI211_X1 U11358 ( .C1(n10834), .C2(n10736), .A(n10726), .B(n10725), .ZN(
        n10727) );
  AOI22_X1 U11359 ( .A1(n10665), .A2(n10727), .B1(n6482), .B2(n10835), .ZN(
        P1_U3530) );
  AOI22_X1 U11360 ( .A1(n10839), .A2(n10727), .B1(n7520), .B2(n10836), .ZN(
        P1_U3477) );
  INV_X1 U11361 ( .A(n10728), .ZN(n10729) );
  AOI222_X1 U11362 ( .A1(n10733), .A2(n10732), .B1(P1_REG2_REG_8__SCAN_IN), 
        .B2(n10731), .C1(n10730), .C2(n10729), .ZN(n10738) );
  INV_X1 U11363 ( .A(n10734), .ZN(n10735) );
  AOI22_X1 U11364 ( .A1(n10736), .A2(n10843), .B1(n4942), .B2(n10735), .ZN(
        n10737) );
  OAI211_X1 U11365 ( .C1(n10697), .C2(n10739), .A(n10738), .B(n10737), .ZN(
        P1_U3285) );
  NOR2_X1 U11366 ( .A1(n10740), .A2(n10774), .ZN(n10742) );
  AOI211_X1 U11367 ( .C1(n10779), .C2(n10743), .A(n10742), .B(n10741), .ZN(
        n10745) );
  AOI22_X1 U11368 ( .A1(n10781), .A2(n10745), .B1(n7149), .B2(n10780), .ZN(
        P2_U3467) );
  INV_X1 U11369 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10744) );
  AOI22_X1 U11370 ( .A1(n10785), .A2(n10745), .B1(n10744), .B2(n10782), .ZN(
        P2_U3414) );
  AOI22_X1 U11371 ( .A1(n10748), .A2(n10791), .B1(n10747), .B2(n10746), .ZN(
        n10749) );
  OAI211_X1 U11372 ( .C1(n10751), .C2(n10794), .A(n10750), .B(n10749), .ZN(
        n10752) );
  AOI21_X1 U11373 ( .B1(n10753), .B2(n10811), .A(n10752), .ZN(n10755) );
  AOI22_X1 U11374 ( .A1(n10665), .A2(n10755), .B1(n10754), .B2(n10835), .ZN(
        P1_U3531) );
  AOI22_X1 U11375 ( .A1(n10839), .A2(n10755), .B1(n7550), .B2(n10836), .ZN(
        P1_U3480) );
  OAI22_X1 U11376 ( .A1(n10757), .A2(n10825), .B1(n10756), .B2(n10823), .ZN(
        n10758) );
  AOI21_X1 U11377 ( .B1(n10759), .B2(n10791), .A(n10758), .ZN(n10761) );
  OAI211_X1 U11378 ( .C1(n10762), .C2(n10794), .A(n10761), .B(n10760), .ZN(
        n10763) );
  AOI21_X1 U11379 ( .B1(n10764), .B2(n10811), .A(n10763), .ZN(n10766) );
  INV_X1 U11380 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10765) );
  AOI22_X1 U11381 ( .A1(n10665), .A2(n10766), .B1(n10765), .B2(n10835), .ZN(
        P1_U3532) );
  AOI22_X1 U11382 ( .A1(n10839), .A2(n10766), .B1(n7567), .B2(n10836), .ZN(
        P1_U3483) );
  NOR2_X1 U11383 ( .A1(n10768), .A2(n10767), .ZN(n10770) );
  AOI211_X1 U11384 ( .C1(n10779), .C2(n10771), .A(n10770), .B(n10769), .ZN(
        n10773) );
  AOI22_X1 U11385 ( .A1(n10781), .A2(n10773), .B1(n7457), .B2(n10780), .ZN(
        P2_U3469) );
  INV_X1 U11386 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U11387 ( .A1(n10785), .A2(n10773), .B1(n10772), .B2(n10782), .ZN(
        P2_U3420) );
  NOR2_X1 U11388 ( .A1(n10775), .A2(n10774), .ZN(n10777) );
  AOI211_X1 U11389 ( .C1(n10779), .C2(n10778), .A(n10777), .B(n10776), .ZN(
        n10784) );
  AOI22_X1 U11390 ( .A1(n10781), .A2(n10784), .B1(n5893), .B2(n10780), .ZN(
        P2_U3470) );
  INV_X1 U11391 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10783) );
  AOI22_X1 U11392 ( .A1(n10785), .A2(n10784), .B1(n10783), .B2(n10782), .ZN(
        P2_U3423) );
  OAI22_X1 U11393 ( .A1(n10787), .A2(n10825), .B1(n10786), .B2(n10823), .ZN(
        n10789) );
  AOI211_X1 U11394 ( .C1(n10791), .C2(n10790), .A(n10789), .B(n10788), .ZN(
        n10792) );
  OAI21_X1 U11395 ( .B1(n10794), .B2(n10793), .A(n10792), .ZN(n10795) );
  AOI21_X1 U11396 ( .B1(n10796), .B2(n10811), .A(n10795), .ZN(n10798) );
  AOI22_X1 U11397 ( .A1(n10665), .A2(n10798), .B1(n7576), .B2(n10835), .ZN(
        P1_U3533) );
  INV_X1 U11398 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10797) );
  AOI22_X1 U11399 ( .A1(n10839), .A2(n10798), .B1(n10797), .B2(n10836), .ZN(
        P1_U3486) );
  OAI211_X1 U11400 ( .C1(n10801), .C2(n10820), .A(n10800), .B(n10799), .ZN(
        n10802) );
  AOI21_X1 U11401 ( .B1(n10803), .B2(n10811), .A(n10802), .ZN(n10806) );
  AOI22_X1 U11402 ( .A1(n10665), .A2(n10806), .B1(n10804), .B2(n10835), .ZN(
        P1_U3534) );
  INV_X1 U11403 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10805) );
  AOI22_X1 U11404 ( .A1(n10839), .A2(n10806), .B1(n10805), .B2(n10836), .ZN(
        P1_U3489) );
  OAI211_X1 U11405 ( .C1(n10809), .C2(n10820), .A(n10808), .B(n10807), .ZN(
        n10810) );
  AOI21_X1 U11406 ( .B1(n10812), .B2(n10811), .A(n10810), .ZN(n10813) );
  AOI22_X1 U11407 ( .A1(n10665), .A2(n10813), .B1(n7433), .B2(n10835), .ZN(
        P1_U3535) );
  AOI22_X1 U11408 ( .A1(n10839), .A2(n10813), .B1(n6439), .B2(n10836), .ZN(
        P1_U3492) );
  XNOR2_X1 U11409 ( .A(n10815), .B(n10814), .ZN(n10832) );
  INV_X1 U11410 ( .A(n10832), .ZN(n10844) );
  INV_X1 U11411 ( .A(n10816), .ZN(n10819) );
  OAI211_X1 U11412 ( .C1(n10819), .C2(n10846), .A(n10818), .B(n10817), .ZN(
        n10840) );
  OAI21_X1 U11413 ( .B1(n10846), .B2(n10820), .A(n10840), .ZN(n10833) );
  XNOR2_X1 U11414 ( .A(n10822), .B(n10821), .ZN(n10829) );
  OAI22_X1 U11415 ( .A1(n10826), .A2(n10825), .B1(n10824), .B2(n10823), .ZN(
        n10827) );
  AOI21_X1 U11416 ( .B1(n10829), .B2(n10828), .A(n10827), .ZN(n10830) );
  OAI21_X1 U11417 ( .B1(n10832), .B2(n10831), .A(n10830), .ZN(n10853) );
  AOI211_X1 U11418 ( .C1(n10834), .C2(n10844), .A(n10833), .B(n10853), .ZN(
        n10838) );
  AOI22_X1 U11419 ( .A1(n10665), .A2(n10838), .B1(n7801), .B2(n10835), .ZN(
        P1_U3536) );
  INV_X1 U11420 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10837) );
  AOI22_X1 U11421 ( .A1(n10839), .A2(n10838), .B1(n10837), .B2(n10836), .ZN(
        P1_U3495) );
  INV_X1 U11422 ( .A(n10840), .ZN(n10841) );
  AOI22_X1 U11423 ( .A1(n10844), .A2(n10843), .B1(n4942), .B2(n10841), .ZN(
        n10855) );
  NOR2_X1 U11424 ( .A1(n10846), .A2(n10845), .ZN(n10851) );
  OAI22_X1 U11425 ( .A1(n10852), .A2(n10849), .B1(n10848), .B2(n10847), .ZN(
        n10850) );
  AOI211_X1 U11426 ( .C1(n10853), .C2(n10852), .A(n10851), .B(n10850), .ZN(
        n10854) );
  NAND2_X1 U11427 ( .A1(n10855), .A2(n10854), .ZN(P1_U3279) );
  XNOR2_X1 U11428 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  CLKBUF_X1 U5018 ( .A(n5745), .Z(n5977) );
  NAND2_X1 U6300 ( .A1(n6306), .A2(n8169), .ZN(n6046) );
  BUF_X1 U5216 ( .A(n7185), .Z(n8301) );
  INV_X1 U5012 ( .A(n8301), .ZN(n9695) );
  CLKBUF_X1 U5181 ( .A(n5700), .Z(n5699) );
  XOR2_X1 U6537 ( .A(n10771), .B(n8744), .Z(n10858) );
endmodule

