

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput127, keyinput126,
         keyinput125, keyinput124, keyinput123, keyinput122, keyinput121,
         keyinput120, keyinput119, keyinput118, keyinput117, keyinput116,
         keyinput115, keyinput114, keyinput113, keyinput112, keyinput111,
         keyinput110, keyinput109, keyinput108, keyinput107, keyinput106,
         keyinput105, keyinput104, keyinput103, keyinput102, keyinput101,
         keyinput100, keyinput99, keyinput98, keyinput97, keyinput96,
         keyinput95, keyinput94, keyinput93, keyinput92, keyinput91,
         keyinput90, keyinput89, keyinput88, keyinput87, keyinput86,
         keyinput85, keyinput84, keyinput83, keyinput82, keyinput81,
         keyinput80, keyinput79, keyinput78, keyinput77, keyinput76,
         keyinput75, keyinput74, keyinput73, keyinput72, keyinput71,
         keyinput70, keyinput69, keyinput68, keyinput67, keyinput66,
         keyinput65, keyinput64, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858;

  CLKBUF_X2 U3549 ( .A(n4143), .Z(n3121) );
  CLKBUF_X2 U3550 ( .A(n3285), .Z(n4151) );
  CLKBUF_X2 U3551 ( .A(n3309), .Z(n4150) );
  BUF_X1 U3552 ( .A(n3279), .Z(n4148) );
  CLKBUF_X2 U3553 ( .A(n3106), .Z(n3422) );
  AND2_X1 U3554 ( .A1(n4510), .A2(n3224), .ZN(n3285) );
  AND2_X1 U3555 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4606) );
  INV_X1 U3556 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4586) );
  OAI21_X1 U3557 ( .B1(n4496), .B2(STATE2_REG_0__SCAN_IN), .A(n3454), .ZN(
        n3460) );
  AOI22_X1 U3558 ( .A1(n6553), .A2(keyinput124), .B1(n4308), .B2(keyinput16), 
        .ZN(n6552) );
  NAND2_X1 U3559 ( .A1(n3366), .A2(n3293), .ZN(n3330) );
  AND2_X1 U3560 ( .A1(n4557), .A2(n5282), .ZN(n4352) );
  NAND2_X1 U3561 ( .A1(n3522), .A2(n3521), .ZN(n3523) );
  OAI221_X1 U3562 ( .B1(n6553), .B2(keyinput124), .C1(n4308), .C2(keyinput16), 
        .A(n6552), .ZN(n6554) );
  INV_X1 U3564 ( .A(n3365), .ZN(n4387) );
  NAND2_X1 U3565 ( .A1(n3333), .A2(n3706), .ZN(n3339) );
  INV_X1 U3566 ( .A(n4548), .ZN(n4557) );
  NAND2_X1 U3567 ( .A1(n3407), .A2(n3130), .ZN(n3707) );
  NAND2_X1 U3568 ( .A1(n3516), .A2(n3515), .ZN(n4689) );
  INV_X1 U3569 ( .A(n3349), .ZN(n3701) );
  INV_X1 U3570 ( .A(n3101), .ZN(n4695) );
  XNOR2_X1 U3571 ( .A(n4180), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4459)
         );
  INV_X1 U3572 ( .A(n5704), .ZN(n5693) );
  NAND2_X2 U3573 ( .A1(n3762), .A2(n3761), .ZN(n4820) );
  XNOR2_X1 U3574 ( .A(n3525), .B(n4689), .ZN(n3725) );
  NAND2_X2 U3575 ( .A1(n5021), .A2(n5020), .ZN(n5973) );
  NAND2_X2 U3576 ( .A1(n3189), .A2(n3188), .ZN(n5021) );
  AND2_X4 U3577 ( .A1(n4616), .A2(n3748), .ZN(n3101) );
  NAND2_X4 U3578 ( .A1(n3241), .A2(n3240), .ZN(n3333) );
  AND2_X2 U3579 ( .A1(n4505), .A2(n3224), .ZN(n3271) );
  NAND4_X2 U3580 ( .A1(n3101), .A2(n3195), .A3(n4820), .A4(n4768), .ZN(n4766)
         );
  BUF_X4 U3583 ( .A(n4256), .Z(n5282) );
  NAND2_X4 U3584 ( .A1(n3610), .A2(n3609), .ZN(n5704) );
  NOR2_X1 U3585 ( .A1(n4696), .A2(n4759), .ZN(n3195) );
  INV_X2 U3586 ( .A(n5903), .ZN(n5892) );
  XNOR2_X1 U3587 ( .A(n3569), .B(n3570), .ZN(n3731) );
  BUF_X1 U3589 ( .A(n4594), .Z(n3122) );
  NAND2_X1 U3590 ( .A1(n5204), .A2(n4220), .ZN(n4482) );
  NAND2_X1 U3593 ( .A1(n3374), .A2(n3365), .ZN(n4480) );
  INV_X1 U3594 ( .A(n3332), .ZN(n3374) );
  INV_X2 U3595 ( .A(n3294), .ZN(n4417) );
  AND4_X1 U3596 ( .A1(n3317), .A2(n3316), .A3(n3315), .A4(n3314), .ZN(n3328)
         );
  AND4_X1 U3597 ( .A1(n3325), .A2(n3324), .A3(n3323), .A4(n3322), .ZN(n3326)
         );
  BUF_X2 U3598 ( .A(n4122), .Z(n4041) );
  BUF_X2 U3599 ( .A(n3271), .Z(n3109) );
  CLKBUF_X2 U3600 ( .A(n3269), .Z(n4142) );
  BUF_X2 U3601 ( .A(n3278), .Z(n4123) );
  BUF_X2 U3602 ( .A(n3792), .Z(n4087) );
  BUF_X2 U3603 ( .A(n3872), .Z(n3980) );
  AND2_X1 U3604 ( .A1(n4585), .A2(n3219), .ZN(n3309) );
  NOR2_X1 U3605 ( .A1(n4207), .A2(n4206), .ZN(n5413) );
  NOR2_X1 U3606 ( .A1(n4381), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4382)
         );
  OR2_X1 U3607 ( .A1(n5339), .A2(n4178), .ZN(n4381) );
  NAND2_X1 U3608 ( .A1(n4193), .A2(n4192), .ZN(n5584) );
  AOI21_X1 U3609 ( .B1(n4209), .B2(n4192), .A(n4216), .ZN(n5653) );
  OR2_X1 U3610 ( .A1(n4191), .A2(n3135), .ZN(n4193) );
  NAND2_X1 U3611 ( .A1(n3632), .A2(n3170), .ZN(n3169) );
  OAI21_X1 U3612 ( .B1(n5264), .B2(n5263), .A(n5358), .ZN(n5625) );
  INV_X1 U3613 ( .A(n3183), .ZN(n3182) );
  AOI21_X1 U3614 ( .B1(n3190), .B2(n3192), .A(n3131), .ZN(n3188) );
  AOI21_X1 U3615 ( .B1(n3619), .B2(n3186), .A(n3140), .ZN(n3185) );
  AND2_X1 U3616 ( .A1(n3620), .A2(n3187), .ZN(n3186) );
  AND2_X2 U3617 ( .A1(n4698), .A2(n4699), .ZN(n4616) );
  AND2_X1 U3618 ( .A1(n5972), .A2(n3618), .ZN(n3619) );
  NAND2_X1 U3619 ( .A1(n3720), .A2(n4555), .ZN(n4703) );
  XNOR2_X1 U3620 ( .A(n3610), .B(n3597), .ZN(n3757) );
  CLKBUF_X3 U3621 ( .A(n3725), .Z(n3114) );
  NOR2_X1 U3622 ( .A1(n4182), .A2(n4181), .ZN(n4183) );
  CLKBUF_X1 U3623 ( .A(n4624), .Z(n4825) );
  INV_X1 U3624 ( .A(n4241), .ZN(n4971) );
  XNOR2_X1 U3625 ( .A(n3406), .B(n3405), .ZN(n3464) );
  AND2_X1 U3626 ( .A1(n4482), .A2(n4476), .ZN(n6518) );
  OAI21_X1 U3627 ( .B1(n4884), .B2(n3472), .A(n3480), .ZN(n4513) );
  OAI22_X1 U3628 ( .A1(n4594), .A2(STATE2_REG_0__SCAN_IN), .B1(n3517), .B2(
        n3607), .ZN(n3406) );
  INV_X1 U3629 ( .A(n3460), .ZN(n3486) );
  NAND2_X1 U3630 ( .A1(n3477), .A2(n3476), .ZN(n4884) );
  NAND2_X2 U3631 ( .A1(n3686), .A2(n3685), .ZN(n5204) );
  OAI21_X1 U3632 ( .B1(n3707), .B2(STATE2_REG_0__SCAN_IN), .A(n3474), .ZN(
        n3439) );
  AOI21_X1 U3633 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6525), .A(n3680), 
        .ZN(n3681) );
  INV_X1 U3634 ( .A(n3391), .ZN(n3177) );
  NAND2_X1 U3635 ( .A1(n3503), .A2(n3502), .ZN(n6182) );
  AND2_X1 U3636 ( .A1(n3371), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3377) );
  OAI21_X1 U3637 ( .B1(n3148), .B2(n3654), .A(n3684), .ZN(n3659) );
  AND2_X1 U3638 ( .A1(n5195), .A2(n3375), .ZN(n3376) );
  AND3_X1 U3639 ( .A1(n3356), .A2(n3355), .A3(n3354), .ZN(n3361) );
  OAI211_X1 U3640 ( .C1(n3298), .C2(n4368), .A(n3297), .B(n3296), .ZN(n3373)
         );
  NOR2_X1 U3641 ( .A1(n4503), .A2(n6525), .ZN(n4138) );
  INV_X1 U3642 ( .A(n3107), .ZN(n3108) );
  AND2_X2 U3643 ( .A1(n3607), .A2(n3504), .ZN(n3682) );
  NAND2_X1 U3644 ( .A1(n4387), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3504) );
  OR2_X1 U3646 ( .A1(n3432), .A2(n3431), .ZN(n3489) );
  NAND2_X2 U3647 ( .A1(n3365), .A2(n3332), .ZN(n4548) );
  AND2_X1 U3648 ( .A1(n3365), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3652) );
  NOR2_X1 U3649 ( .A1(n3332), .A2(n3365), .ZN(n5203) );
  AND4_X1 U3650 ( .A1(n3284), .A2(n3283), .A3(n3282), .A4(n3281), .ZN(n3213)
         );
  OR2_X2 U3651 ( .A1(n3308), .A2(n3307), .ZN(n3365) );
  AND4_X1 U3652 ( .A1(n3289), .A2(n3288), .A3(n3287), .A4(n3286), .ZN(n3290)
         );
  AND4_X1 U3653 ( .A1(n3259), .A2(n3258), .A3(n3257), .A4(n3256), .ZN(n3260)
         );
  AND4_X1 U3654 ( .A1(n3268), .A2(n3267), .A3(n3266), .A4(n3265), .ZN(n3277)
         );
  AND4_X1 U3655 ( .A1(n3275), .A2(n3274), .A3(n3273), .A4(n3272), .ZN(n3276)
         );
  AND4_X1 U3656 ( .A1(n3321), .A2(n3320), .A3(n3319), .A4(n3318), .ZN(n3327)
         );
  AND4_X1 U3657 ( .A1(n3313), .A2(n3312), .A3(n3311), .A4(n3310), .ZN(n3329)
         );
  AND4_X1 U3658 ( .A1(n3239), .A2(n3238), .A3(n3237), .A4(n3236), .ZN(n3240)
         );
  AND4_X1 U3659 ( .A1(n3223), .A2(n3222), .A3(n3221), .A4(n3220), .ZN(n3231)
         );
  CLKBUF_X2 U3660 ( .A(n3410), .Z(n3103) );
  BUF_X2 U3661 ( .A(n3855), .Z(n4149) );
  BUF_X1 U3662 ( .A(n3410), .Z(n3102) );
  AND2_X2 U3663 ( .A1(n3225), .A2(n4606), .ZN(n3119) );
  AND2_X2 U3664 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4504) );
  NOR2_X1 U3665 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3219) );
  AND2_X2 U3666 ( .A1(n3144), .A2(n4495), .ZN(n4505) );
  BUF_X4 U3667 ( .A(n3443), .Z(n3106) );
  NAND2_X2 U3668 ( .A1(n3231), .A2(n3230), .ZN(n3338) );
  AND2_X1 U3669 ( .A1(n4582), .A2(n4504), .ZN(n3415) );
  AND2_X1 U3670 ( .A1(n4582), .A2(n4504), .ZN(n3115) );
  AND2_X2 U3671 ( .A1(n4582), .A2(n4504), .ZN(n3116) );
  AND2_X2 U3672 ( .A1(n4510), .A2(n4606), .ZN(n3270) );
  BUF_X4 U3673 ( .A(n3410), .Z(n3104) );
  AND2_X2 U3674 ( .A1(n4505), .A2(n4581), .ZN(n4143) );
  INV_X1 U3675 ( .A(n5203), .ZN(n3107) );
  AND2_X2 U3676 ( .A1(n3143), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4581)
         );
  AOI21_X2 U3677 ( .B1(n3363), .B2(n3344), .A(n3210), .ZN(n3408) );
  AND2_X2 U3678 ( .A1(n4581), .A2(n4504), .ZN(n3278) );
  AND2_X1 U3680 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4585) );
  BUF_X1 U3681 ( .A(n4208), .Z(n4216) );
  AND2_X1 U3682 ( .A1(n4510), .A2(n3224), .ZN(n3112) );
  INV_X2 U3683 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3144) );
  XNOR2_X1 U3684 ( .A(n4572), .B(n6182), .ZN(n4578) );
  AND2_X2 U3685 ( .A1(n3402), .A2(n3333), .ZN(n3357) );
  NAND2_X2 U3686 ( .A1(n3384), .A2(n3383), .ZN(n3441) );
  NAND2_X1 U3687 ( .A1(n3402), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3607) );
  OAI21_X2 U3688 ( .B1(n5681), .B2(n3139), .A(n3631), .ZN(n3632) );
  OAI21_X2 U3689 ( .B1(n5708), .B2(n3622), .A(n3621), .ZN(n5390) );
  NAND2_X2 U3690 ( .A1(n3180), .A2(n3179), .ZN(n5708) );
  INV_X2 U3691 ( .A(n5233), .ZN(n4079) );
  NOR2_X4 U3692 ( .A1(n5298), .A2(n5299), .ZN(n5290) );
  NAND2_X2 U3693 ( .A1(n3724), .A2(n3723), .ZN(n4698) );
  NAND2_X2 U3694 ( .A1(n5113), .A2(n3199), .ZN(n5298) );
  NAND2_X2 U3695 ( .A1(n5085), .A2(n3852), .ZN(n5113) );
  AND2_X2 U3696 ( .A1(n5262), .A2(n5357), .ZN(n5243) );
  NOR2_X2 U3697 ( .A1(n5260), .A2(n5259), .ZN(n5262) );
  AND2_X2 U3698 ( .A1(n3652), .A2(n3338), .ZN(n3677) );
  AND2_X2 U3699 ( .A1(n4394), .A2(n3364), .ZN(n4386) );
  AND2_X1 U3700 ( .A1(n4585), .A2(n3219), .ZN(n3117) );
  AND2_X1 U3701 ( .A1(n4585), .A2(n3219), .ZN(n3118) );
  AND2_X4 U3702 ( .A1(n3224), .A2(n4504), .ZN(n3279) );
  AND2_X2 U3703 ( .A1(n3143), .A2(n4586), .ZN(n3224) );
  INV_X2 U3704 ( .A(n3338), .ZN(n3402) );
  AND2_X2 U3705 ( .A1(n3225), .A2(n4606), .ZN(n3120) );
  AND2_X2 U3706 ( .A1(n3225), .A2(n4606), .ZN(n3854) );
  AND2_X1 U3707 ( .A1(n3349), .A2(n3402), .ZN(n3331) );
  OR2_X2 U3708 ( .A1(n3251), .A2(n3250), .ZN(n3349) );
  OAI211_X1 U3709 ( .C1(n3178), .C2(n3177), .A(n3176), .B(n3174), .ZN(n4594)
         );
  OR2_X1 U3710 ( .A1(n3682), .A2(n3582), .ZN(n3584) );
  INV_X1 U3711 ( .A(n3185), .ZN(n3184) );
  NAND2_X1 U3712 ( .A1(n4100), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4119)
         );
  INV_X1 U3713 ( .A(n3750), .ZN(n4141) );
  AND2_X1 U3714 ( .A1(n3350), .A2(n3332), .ZN(n4256) );
  NAND2_X1 U3715 ( .A1(n3571), .A2(n3134), .ZN(n3610) );
  OAI21_X1 U3716 ( .B1(n3126), .B2(n3184), .A(n5501), .ZN(n3183) );
  INV_X1 U3717 ( .A(n5433), .ZN(n3170) );
  AND2_X1 U3718 ( .A1(n5256), .A2(n5447), .ZN(n3161) );
  NOR2_X1 U3719 ( .A1(n3165), .A2(n5295), .ZN(n3164) );
  INV_X1 U3720 ( .A(n5285), .ZN(n3165) );
  AND2_X1 U3721 ( .A1(n6426), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3690) );
  AND2_X1 U3722 ( .A1(n5317), .A2(n4374), .ZN(n5932) );
  INV_X1 U3723 ( .A(n5317), .ZN(n5931) );
  INV_X1 U3724 ( .A(n3585), .ZN(n3561) );
  AND2_X1 U3725 ( .A1(n3656), .A2(n3657), .ZN(n3147) );
  NAND2_X1 U3726 ( .A1(n3637), .A2(n3636), .ZN(n3672) );
  NAND2_X1 U3727 ( .A1(n3548), .A2(n3547), .ZN(n3569) );
  NAND2_X1 U3728 ( .A1(n3560), .A2(n3559), .ZN(n3570) );
  OR2_X1 U3729 ( .A1(n3581), .A2(n3580), .ZN(n3599) );
  INV_X1 U3730 ( .A(n3684), .ZN(n3679) );
  OR3_X1 U3731 ( .A1(n3643), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(n6113), 
        .ZN(n4221) );
  INV_X1 U3732 ( .A(n5112), .ZN(n3203) );
  NAND2_X1 U3733 ( .A1(n3701), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4136) );
  INV_X1 U3734 ( .A(n5091), .ZN(n3187) );
  INV_X1 U3735 ( .A(n3191), .ZN(n3190) );
  OAI21_X1 U3736 ( .B1(n5989), .B2(n3192), .A(n3616), .ZN(n3191) );
  INV_X1 U3737 ( .A(n3615), .ZN(n3192) );
  NOR2_X2 U3738 ( .A1(n4548), .A2(n5282), .ZN(n4341) );
  BUF_X1 U3739 ( .A(n4257), .Z(n4346) );
  INV_X1 U3740 ( .A(n4681), .ZN(n3168) );
  INV_X1 U3741 ( .A(n5282), .ZN(n4461) );
  AOI21_X1 U3742 ( .B1(n4556), .B2(n4557), .A(n4261), .ZN(n4748) );
  OAI21_X1 U3743 ( .B1(n4394), .B2(n4480), .A(n4421), .ZN(n3353) );
  NOR2_X1 U3744 ( .A1(n3352), .A2(n4422), .ZN(n3355) );
  OR2_X1 U3745 ( .A1(n5760), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3696) );
  NAND2_X1 U3746 ( .A1(n5622), .A2(n3212), .ZN(n5597) );
  NAND2_X1 U3747 ( .A1(n5820), .A2(n6832), .ZN(n5799) );
  NOR2_X1 U3748 ( .A1(n5182), .A2(n5282), .ZN(n4353) );
  NAND2_X1 U3749 ( .A1(n4461), .A2(n4346), .ZN(n4529) );
  INV_X1 U3750 ( .A(n4536), .ZN(n5966) );
  AND2_X1 U3751 ( .A1(n3197), .A2(n5276), .ZN(n3196) );
  NAND2_X1 U3752 ( .A1(n3804), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3807)
         );
  AND2_X1 U3753 ( .A1(n4742), .A2(n4617), .ZN(n3748) );
  OR2_X1 U3754 ( .A1(n4354), .A2(n4356), .ZN(n5182) );
  NAND2_X1 U3755 ( .A1(n5448), .A2(n3141), .ZN(n5252) );
  INV_X1 U3756 ( .A(n5249), .ZN(n3160) );
  NOR2_X1 U3757 ( .A1(n3124), .A2(n5265), .ZN(n5448) );
  OR2_X1 U3758 ( .A1(n5312), .A2(n5305), .ZN(n5294) );
  AND2_X1 U3759 ( .A1(n4311), .A2(n4310), .ZN(n5295) );
  NAND2_X1 U3760 ( .A1(n5310), .A2(n5309), .ZN(n5312) );
  OR2_X1 U3761 ( .A1(n5704), .A2(n6052), .ZN(n3618) );
  NOR2_X1 U3762 ( .A1(n4681), .A2(n3166), .ZN(n5036) );
  NAND2_X1 U3763 ( .A1(n3123), .A2(n3127), .ZN(n3166) );
  NAND2_X1 U3764 ( .A1(n4404), .A2(n6436), .ZN(n4426) );
  AND2_X1 U3765 ( .A1(n5204), .A2(n4405), .ZN(n6417) );
  NOR2_X1 U3766 ( .A1(n5219), .A2(n5916), .ZN(n3145) );
  AND2_X1 U3767 ( .A1(n4249), .A2(n4248), .ZN(n4250) );
  NAND2_X1 U3768 ( .A1(n4371), .A2(n4536), .ZN(n5317) );
  OAI21_X1 U3769 ( .B1(n4485), .B2(n4369), .A(n6436), .ZN(n4371) );
  AOI21_X1 U3770 ( .B1(n6022), .B2(n5579), .A(n4195), .ZN(n4196) );
  INV_X1 U3771 ( .A(n6045), .ZN(n6022) );
  AND2_X1 U3772 ( .A1(n6417), .A2(n6436), .ZN(n6040) );
  INV_X1 U3773 ( .A(n6040), .ZN(n5773) );
  NOR2_X1 U3774 ( .A1(n3169), .A2(n3207), .ZN(n4179) );
  AND2_X1 U3775 ( .A1(n3690), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6436) );
  NOR2_X1 U3776 ( .A1(n3332), .A2(n4237), .ZN(n3370) );
  OR2_X1 U3777 ( .A1(n3607), .A2(n3455), .ZN(n3454) );
  AND2_X1 U3778 ( .A1(n6183), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3649)
         );
  CLKBUF_X2 U3779 ( .A(n3270), .Z(n3889) );
  OR2_X1 U3780 ( .A1(n3682), .A2(n3561), .ZN(n3537) );
  OR2_X1 U3781 ( .A1(n3535), .A2(n3534), .ZN(n3585) );
  OR2_X1 U3782 ( .A1(n3401), .A2(n3400), .ZN(n3403) );
  OR2_X1 U3783 ( .A1(n3514), .A2(n3513), .ZN(n3538) );
  NAND2_X1 U3784 ( .A1(n3477), .A2(n3209), .ZN(n3485) );
  NOR2_X1 U3785 ( .A1(n3687), .A2(n3689), .ZN(n4398) );
  AOI21_X1 U3786 ( .B1(n3339), .B2(n3350), .A(n3701), .ZN(n3296) );
  OR2_X1 U3787 ( .A1(n4240), .A2(n4239), .ZN(n5208) );
  INV_X1 U3788 ( .A(n3333), .ZN(n3366) );
  NOR2_X1 U3789 ( .A1(n3350), .A2(n3294), .ZN(n4367) );
  INV_X1 U3790 ( .A(n4209), .ZN(n3204) );
  NOR2_X1 U3791 ( .A1(n3206), .A2(n5235), .ZN(n3205) );
  INV_X1 U3792 ( .A(n3135), .ZN(n3206) );
  INV_X1 U3793 ( .A(n5371), .ZN(n3972) );
  NOR2_X1 U3794 ( .A1(n3198), .A2(n5278), .ZN(n3197) );
  INV_X1 U3795 ( .A(n5292), .ZN(n3198) );
  NAND2_X1 U3796 ( .A1(n3830), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3835)
         );
  AOI21_X1 U3797 ( .B1(n5519), .B2(n3877), .A(n4174), .ZN(n3720) );
  NOR2_X1 U3798 ( .A1(n3625), .A2(n3194), .ZN(n3193) );
  AND2_X1 U3799 ( .A1(n5704), .A2(n6579), .ZN(n3625) );
  INV_X1 U3800 ( .A(n3624), .ZN(n3194) );
  INV_X1 U3801 ( .A(n4352), .ZN(n4349) );
  NAND2_X1 U3802 ( .A1(n5704), .A2(n3613), .ZN(n3614) );
  INV_X1 U3803 ( .A(n4752), .ZN(n3167) );
  INV_X1 U3804 ( .A(n4680), .ZN(n4275) );
  NAND2_X1 U3805 ( .A1(n3151), .A2(n3149), .ZN(n4261) );
  NAND2_X1 U3806 ( .A1(n4341), .A2(n4921), .ZN(n3151) );
  AND2_X1 U3807 ( .A1(n3333), .A2(n3332), .ZN(n3644) );
  INV_X1 U3808 ( .A(n3606), .ZN(n3611) );
  OR2_X1 U3809 ( .A1(n3339), .A2(n3688), .ZN(n4503) );
  AND2_X2 U3810 ( .A1(n4586), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4582)
         );
  AOI21_X1 U3811 ( .B1(n3263), .B2(INSTQUEUE_REG_10__2__SCAN_IN), .A(n3264), 
        .ZN(n3268) );
  AND2_X1 U3812 ( .A1(n3119), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3264) );
  AND2_X1 U3813 ( .A1(n3103), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3280) );
  AOI21_X1 U3814 ( .B1(n6521), .B2(n4807), .A(n5118), .ZN(n4622) );
  OR2_X1 U3815 ( .A1(n6116), .A2(n4626), .ZN(n4688) );
  OAI21_X1 U3816 ( .B1(n3677), .B2(n4221), .A(n3676), .ZN(n3678) );
  NAND2_X1 U3817 ( .A1(n3642), .A2(n3641), .ZN(n4226) );
  OR2_X1 U3818 ( .A1(n3643), .A2(n3640), .ZN(n3642) );
  AND2_X1 U3819 ( .A1(n6113), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3640)
         );
  AND2_X1 U3820 ( .A1(n3677), .A2(n3644), .ZN(n3684) );
  INV_X1 U3821 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5807) );
  INV_X1 U3822 ( .A(n5208), .ZN(n5207) );
  NAND2_X1 U3823 ( .A1(n5207), .A2(REIP_REG_1__SCAN_IN), .ZN(n5009) );
  AND2_X1 U3824 ( .A1(n5238), .A2(n5228), .ZN(n5229) );
  NAND2_X1 U3825 ( .A1(n4322), .A2(n3164), .ZN(n3163) );
  OR2_X1 U3826 ( .A1(n5204), .A2(n5196), .ZN(n4551) );
  INV_X1 U3827 ( .A(n4136), .ZN(n4175) );
  OR2_X1 U3828 ( .A1(n4119), .A2(n3695), .ZN(n4182) );
  NAND2_X1 U3829 ( .A1(n3974), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3993)
         );
  OR2_X1 U3830 ( .A1(n3993), .A2(n3992), .ZN(n4038) );
  CLKBUF_X1 U3831 ( .A(n5260), .Z(n5261) );
  OR2_X1 U3832 ( .A1(n3940), .A2(n5633), .ZN(n3956) );
  NOR2_X1 U3833 ( .A1(n3956), .A2(n5373), .ZN(n3974) );
  NOR2_X1 U3834 ( .A1(n3912), .A2(n5791), .ZN(n3926) );
  NOR2_X1 U3835 ( .A1(n3884), .A2(n5807), .ZN(n3898) );
  CLKBUF_X1 U3836 ( .A(n5290), .Z(n5291) );
  NAND2_X1 U3837 ( .A1(n3881), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3884)
         );
  NOR2_X1 U3838 ( .A1(n3202), .A2(n3200), .ZN(n3199) );
  INV_X1 U3839 ( .A(n5303), .ZN(n3200) );
  AND2_X1 U3840 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n3853), .ZN(n3881)
         );
  NOR2_X1 U3841 ( .A1(n3835), .A2(n3693), .ZN(n3853) );
  INV_X1 U3842 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6553) );
  NOR2_X1 U3843 ( .A1(n6553), .A2(n3807), .ZN(n3830) );
  CLKBUF_X1 U3844 ( .A(n4928), .Z(n4929) );
  NOR2_X1 U3845 ( .A1(n3779), .A2(n3692), .ZN(n3804) );
  OR2_X1 U3846 ( .A1(n3763), .A2(n5874), .ZN(n3779) );
  CLKBUF_X1 U3847 ( .A(n4766), .Z(n4767) );
  NOR2_X1 U3848 ( .A1(n3749), .A2(n3691), .ZN(n3758) );
  NAND2_X1 U3849 ( .A1(n3758), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3763)
         );
  INV_X1 U3850 ( .A(n3760), .ZN(n3761) );
  AOI21_X1 U3851 ( .B1(n3756), .B2(n3877), .A(n3755), .ZN(n4696) );
  OR2_X1 U3852 ( .A1(n3754), .A2(n3753), .ZN(n3755) );
  NAND2_X1 U3853 ( .A1(n3742), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3749)
         );
  INV_X1 U3854 ( .A(n3734), .ZN(n3735) );
  NAND2_X1 U3855 ( .A1(n3731), .A2(n3877), .ZN(n3736) );
  OAI21_X1 U3856 ( .B1(n4136), .B2(n3733), .A(n3732), .ZN(n3734) );
  NOR2_X1 U3857 ( .A1(n6550), .A2(n3743), .ZN(n3742) );
  INV_X1 U3858 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6550) );
  NAND2_X1 U3859 ( .A1(n3726), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3743)
         );
  INV_X1 U3860 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6822) );
  NOR2_X1 U3861 ( .A1(n5252), .A2(n5237), .ZN(n5238) );
  AND2_X1 U3862 ( .A1(n5448), .A2(n5447), .ZN(n5449) );
  OAI21_X1 U3863 ( .B1(n5384), .B2(n5382), .A(n5380), .ZN(n5376) );
  AND3_X1 U3864 ( .A1(n4433), .A2(n5479), .A3(n4432), .ZN(n5460) );
  AOI21_X1 U3865 ( .B1(n3182), .B2(n3184), .A(n3132), .ZN(n3179) );
  OR2_X1 U3866 ( .A1(n4436), .A2(n4435), .ZN(n5747) );
  NOR2_X1 U3867 ( .A1(n5114), .A2(n5115), .ZN(n5310) );
  NAND2_X1 U3868 ( .A1(n3153), .A2(n3152), .ZN(n5114) );
  INV_X1 U3869 ( .A(n5087), .ZN(n3152) );
  INV_X1 U3870 ( .A(n5099), .ZN(n3153) );
  NAND2_X1 U3871 ( .A1(n3155), .A2(n3154), .ZN(n5099) );
  INV_X1 U3872 ( .A(n5096), .ZN(n3154) );
  INV_X1 U3873 ( .A(n5097), .ZN(n3155) );
  NOR3_X1 U3874 ( .A1(n6095), .A2(n4431), .A3(n4678), .ZN(n5102) );
  AND2_X1 U3875 ( .A1(n4289), .A2(n4288), .ZN(n5034) );
  NAND2_X1 U3876 ( .A1(n5987), .A2(n5989), .ZN(n5988) );
  NAND2_X1 U3877 ( .A1(n3168), .A2(n3123), .ZN(n5880) );
  NAND2_X1 U3878 ( .A1(n3168), .A2(n4275), .ZN(n4753) );
  NAND2_X1 U3879 ( .A1(n4655), .A2(n4271), .ZN(n4681) );
  AND2_X1 U3880 ( .A1(n5747), .A2(n5503), .ZN(n5029) );
  AND2_X1 U3881 ( .A1(n4677), .A2(n4676), .ZN(n6104) );
  OAI21_X1 U3882 ( .B1(n3345), .B2(n3347), .A(n3332), .ZN(n3356) );
  NAND2_X1 U3883 ( .A1(n3390), .A2(n3389), .ZN(n3391) );
  INV_X1 U3884 ( .A(n4628), .ZN(n5049) );
  AND2_X1 U3885 ( .A1(n6255), .A2(n6154), .ZN(n6188) );
  NOR2_X1 U3886 ( .A1(n6116), .A2(n4689), .ZN(n6255) );
  OR2_X1 U3887 ( .A1(n6334), .A2(n4825), .ZN(n4873) );
  INV_X1 U3888 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6412) );
  NOR2_X1 U3889 ( .A1(n4688), .A2(n4825), .ZN(n4885) );
  AND2_X1 U3890 ( .A1(n4825), .A2(n4884), .ZN(n6217) );
  NOR2_X1 U3891 ( .A1(n4622), .A2(n4621), .ZN(n4661) );
  INV_X1 U3892 ( .A(n4688), .ZN(n4826) );
  OR2_X1 U3893 ( .A1(n5201), .A2(n6434), .ZN(n4476) );
  OAI211_X1 U3894 ( .C1(n5320), .C2(n5902), .A(n5215), .B(n3158), .ZN(n3157)
         );
  OR2_X1 U3895 ( .A1(n5216), .A2(n5217), .ZN(n3158) );
  NAND2_X1 U3896 ( .A1(n5793), .A2(n3142), .ZN(n5639) );
  INV_X1 U3897 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5791) );
  NAND2_X1 U3898 ( .A1(n5899), .A2(n3215), .ZN(n5872) );
  INV_X1 U3899 ( .A(n5893), .ZN(n5904) );
  NOR2_X1 U3900 ( .A1(n5909), .A2(n6467), .ZN(n5899) );
  NAND2_X1 U3901 ( .A1(n4946), .A2(REIP_REG_4__SCAN_IN), .ZN(n5909) );
  INV_X1 U3902 ( .A(n5891), .ZN(n5916) );
  AND2_X1 U3903 ( .A1(n4247), .A2(n4918), .ZN(n5908) );
  NOR2_X1 U3904 ( .A1(n4971), .A2(n5768), .ZN(n5907) );
  INV_X1 U3905 ( .A(n5908), .ZN(n5897) );
  OAI21_X1 U3906 ( .B1(n4462), .B2(n5181), .A(n5184), .ZN(n4464) );
  OR2_X1 U3907 ( .A1(n5928), .A2(n5932), .ZN(n5335) );
  INV_X1 U3908 ( .A(n5335), .ZN(n5089) );
  OR2_X1 U3909 ( .A1(n4808), .A2(n5960), .ZN(n5957) );
  INV_X1 U3910 ( .A(n6520), .ZN(n5960) );
  NAND2_X1 U3911 ( .A1(n4806), .A2(n4805), .ZN(n5965) );
  NAND2_X1 U3912 ( .A1(n5163), .A2(n4804), .ZN(n4806) );
  INV_X2 U3913 ( .A(n5957), .ZN(n5962) );
  OR2_X1 U3914 ( .A1(n4482), .A2(n4481), .ZN(n5968) );
  OR2_X1 U3915 ( .A1(n4482), .A2(n3332), .ZN(n5163) );
  OR2_X1 U3916 ( .A1(n4482), .A2(n4370), .ZN(n4536) );
  INV_X1 U3917 ( .A(n5968), .ZN(n4547) );
  OR2_X1 U3918 ( .A1(n6040), .A2(n3697), .ZN(n5393) );
  NAND2_X1 U3919 ( .A1(n5393), .A2(n4514), .ZN(n6045) );
  INV_X1 U3920 ( .A(n5393), .ZN(n6036) );
  OR2_X1 U3921 ( .A1(n5436), .A2(n5424), .ZN(n5414) );
  INV_X1 U3922 ( .A(n3632), .ZN(n5434) );
  NAND2_X1 U3923 ( .A1(n5448), .A2(n3161), .ZN(n5250) );
  NOR2_X1 U3924 ( .A1(n5294), .A2(n3162), .ZN(n5271) );
  INV_X1 U3925 ( .A(n3164), .ZN(n3162) );
  NAND2_X1 U3926 ( .A1(n5973), .A2(n3126), .ZN(n3181) );
  OAI21_X1 U3927 ( .B1(n5973), .B2(n3620), .A(n3619), .ZN(n5090) );
  OR2_X1 U3928 ( .A1(n4426), .A2(n5196), .ZN(n6095) );
  OR2_X1 U3929 ( .A1(n4426), .A2(n4412), .ZN(n5733) );
  OAI21_X1 U3930 ( .B1(n3402), .B2(n4406), .A(n4407), .ZN(n4408) );
  OR2_X1 U3931 ( .A1(n4426), .A2(n4599), .ZN(n5503) );
  INV_X1 U3932 ( .A(n5733), .ZN(n6099) );
  INV_X1 U3933 ( .A(n4825), .ZN(n6154) );
  INV_X1 U3934 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4866) );
  CLKBUF_X1 U3935 ( .A(n4623), .Z(n6116) );
  INV_X1 U3936 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6113) );
  AND2_X2 U3937 ( .A1(n4495), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4510)
         );
  INV_X1 U3938 ( .A(n6431), .ZN(n5118) );
  INV_X1 U3939 ( .A(n5560), .ZN(n5520) );
  AND2_X1 U3940 ( .A1(n6188), .A2(n6187), .ZN(n6248) );
  NOR2_X2 U3941 ( .A1(n4873), .A2(n6187), .ZN(n6325) );
  AOI22_X1 U3942 ( .A1(n4774), .A2(n6338), .B1(n4773), .B2(n6290), .ZN(n6540)
         );
  INV_X1 U3943 ( .A(n4917), .ZN(n6364) );
  AND2_X1 U3944 ( .A1(n4955), .A2(n4954), .ZN(n5003) );
  NOR2_X1 U3945 ( .A1(n6740), .A2(n4610), .ZN(n6347) );
  NOR2_X1 U3946 ( .A1(n6722), .A2(n4610), .ZN(n6353) );
  AND2_X1 U3947 ( .A1(DATAI_3_), .A2(n4664), .ZN(n6365) );
  NOR2_X1 U3948 ( .A1(n6572), .A2(n4610), .ZN(n6372) );
  NOR2_X1 U3949 ( .A1(n4756), .A2(n4610), .ZN(n6379) );
  NOR2_X1 U3950 ( .A1(n4697), .A2(n4610), .ZN(n6384) );
  AND2_X1 U3951 ( .A1(DATAI_7_), .A2(n4664), .ZN(n6393) );
  INV_X1 U3952 ( .A(n4901), .ZN(n6332) );
  INV_X1 U3953 ( .A(n5177), .ZN(n6352) );
  INV_X1 U3954 ( .A(n6353), .ZN(n5530) );
  INV_X1 U3955 ( .A(n4904), .ZN(n6358) );
  INV_X1 U3956 ( .A(n6359), .ZN(n5534) );
  INV_X1 U3957 ( .A(n4896), .ZN(n6371) );
  INV_X1 U3958 ( .A(n6372), .ZN(n5543) );
  INV_X1 U3959 ( .A(n6536), .ZN(n6378) );
  NAND2_X1 U3960 ( .A1(n4826), .A2(n6217), .ZN(n4849) );
  INV_X1 U3961 ( .A(n6384), .ZN(n5551) );
  NAND2_X1 U3962 ( .A1(n4826), .A2(n6254), .ZN(n4856) );
  INV_X1 U3963 ( .A(n6436), .ZN(n6434) );
  INV_X1 U3964 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6525) );
  NAND2_X1 U3965 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n5204), .ZN(n6431) );
  INV_X1 U3966 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6451) );
  NAND2_X1 U3967 ( .A1(n3159), .A2(n3156), .ZN(U2796) );
  AOI21_X1 U3968 ( .B1(n5565), .B2(n3146), .A(n3145), .ZN(n3159) );
  INV_X1 U3969 ( .A(n3157), .ZN(n3156) );
  AND2_X1 U3970 ( .A1(n5217), .A2(REIP_REG_30__SCAN_IN), .ZN(n3146) );
  NOR2_X1 U3971 ( .A1(n4378), .A2(n4377), .ZN(n4379) );
  INV_X1 U3972 ( .A(n3172), .ZN(n3171) );
  OAI21_X1 U3973 ( .B1(n5320), .B2(n6026), .A(n4186), .ZN(n3172) );
  NOR2_X1 U3974 ( .A1(n4198), .A2(n4197), .ZN(n4199) );
  INV_X1 U3975 ( .A(n4196), .ZN(n4197) );
  AND2_X1 U3976 ( .A1(n5113), .A2(n3201), .ZN(n5302) );
  AND2_X1 U3977 ( .A1(n4275), .A2(n3167), .ZN(n3123) );
  AND3_X1 U3978 ( .A1(n4820), .A2(n3101), .A3(n3195), .ZN(n4765) );
  OR3_X1 U3980 ( .A1(n5294), .A2(n3163), .A3(n5469), .ZN(n3124) );
  NAND2_X1 U3981 ( .A1(n5113), .A2(n5112), .ZN(n5111) );
  NAND2_X1 U3982 ( .A1(n5689), .A2(n3193), .ZN(n3125) );
  INV_X1 U3983 ( .A(n3169), .ZN(n5432) );
  AND2_X1 U3984 ( .A1(n3619), .A2(n3187), .ZN(n3126) );
  AND2_X1 U3985 ( .A1(n5290), .A2(n3197), .ZN(n5274) );
  NAND2_X1 U3986 ( .A1(n5290), .A2(n5292), .ZN(n5277) );
  NAND2_X1 U3987 ( .A1(n5689), .A2(n3624), .ZN(n5703) );
  NAND2_X1 U3988 ( .A1(n5339), .A2(n5338), .ZN(n4188) );
  AND2_X1 U3989 ( .A1(n4760), .A2(n5879), .ZN(n3127) );
  NOR2_X1 U3990 ( .A1(n4354), .A2(n4355), .ZN(n3128) );
  AND2_X1 U3991 ( .A1(n3193), .A2(n3627), .ZN(n3129) );
  OR2_X1 U3992 ( .A1(n3408), .A2(n3409), .ZN(n3130) );
  NOR2_X1 U3993 ( .A1(n5704), .A2(n5981), .ZN(n3131) );
  INV_X1 U3994 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3143) );
  AND2_X1 U3995 ( .A1(n5704), .A2(n5507), .ZN(n3132) );
  AND2_X1 U3996 ( .A1(n3150), .A2(n4257), .ZN(n3133) );
  NOR2_X1 U3997 ( .A1(n5294), .A2(n5295), .ZN(n5280) );
  NOR2_X2 U3998 ( .A1(n3293), .A2(n6522), .ZN(n3877) );
  NOR2_X1 U3999 ( .A1(n4695), .A2(n4696), .ZN(n4819) );
  NAND2_X1 U4000 ( .A1(n4819), .A2(n4820), .ZN(n4758) );
  NAND2_X1 U4001 ( .A1(n3181), .A2(n3185), .ZN(n5500) );
  NAND2_X1 U4002 ( .A1(n5988), .A2(n3615), .ZN(n5980) );
  NAND2_X1 U4003 ( .A1(n4387), .A2(n3332), .ZN(n4413) );
  AND2_X1 U4004 ( .A1(n3570), .A2(n3595), .ZN(n3134) );
  AND2_X1 U4005 ( .A1(n4099), .A2(n4098), .ZN(n3135) );
  INV_X1 U4006 ( .A(n3202), .ZN(n3201) );
  OR2_X1 U4007 ( .A1(n5307), .A2(n3203), .ZN(n3202) );
  AND2_X1 U4008 ( .A1(n3205), .A2(n3204), .ZN(n3136) );
  NAND2_X1 U4009 ( .A1(n5704), .A2(n5427), .ZN(n3137) );
  OR2_X1 U4010 ( .A1(n5294), .A2(n3163), .ZN(n3138) );
  NOR2_X1 U4011 ( .A1(n5704), .A2(n3214), .ZN(n3139) );
  AND2_X1 U4012 ( .A1(n4748), .A2(n4747), .ZN(n4655) );
  AND2_X1 U4013 ( .A1(n5036), .A2(n4290), .ZN(n4931) );
  OAI21_X1 U4014 ( .B1(n4623), .B2(n3472), .A(n3471), .ZN(n6038) );
  AOI21_X1 U4015 ( .B1(n4560), .B2(n4559), .A(n3495), .ZN(n6037) );
  NAND2_X1 U4016 ( .A1(n3736), .A2(n3735), .ZN(n4742) );
  AND2_X1 U4017 ( .A1(n5704), .A2(n5105), .ZN(n3140) );
  AND2_X1 U4018 ( .A1(n3161), .A2(n3160), .ZN(n3141) );
  INV_X1 U4019 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6823) );
  INV_X2 U4020 ( .A(n5727), .ZN(n4228) );
  XNOR2_X1 U4021 ( .A(n4261), .B(n4527), .ZN(n4556) );
  INV_X2 U4022 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6522) );
  INV_X1 U4023 ( .A(n6026), .ZN(n4663) );
  NAND2_X1 U4024 ( .A1(n4170), .A2(n6335), .ZN(n6026) );
  AND2_X1 U4025 ( .A1(REIP_REG_18__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .ZN(
        n3142) );
  INV_X1 U4026 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4495) );
  NOR2_X2 U4027 ( .A1(n4548), .A2(n4359), .ZN(n5891) );
  OR2_X1 U4028 ( .A1(n4358), .A2(n5211), .ZN(n4359) );
  NOR3_X4 U4029 ( .A1(n3114), .A2(n5519), .A3(n5518), .ZN(n6142) );
  INV_X1 U4030 ( .A(n6217), .ZN(n5518) );
  NOR2_X2 U4031 ( .A1(n5639), .A2(n6486), .ZN(n5622) );
  NOR2_X2 U4032 ( .A1(n5799), .A2(n6480), .ZN(n5793) );
  NOR2_X2 U4033 ( .A1(n5214), .A2(n6498), .ZN(n5565) );
  NAND2_X1 U4034 ( .A1(n3148), .A2(n3147), .ZN(n3658) );
  AOI22_X1 U4035 ( .A1(n3208), .A2(n3660), .B1(n3653), .B2(n3667), .ZN(n3148)
         );
  NOR2_X2 U4036 ( .A1(n5872), .A2(n4253), .ZN(n5842) );
  AND2_X2 U4037 ( .A1(n4241), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4918) );
  NAND2_X2 U4038 ( .A1(n6518), .A2(n4231), .ZN(n4241) );
  NAND4_X1 U4039 ( .A1(n3701), .A2(n4367), .A3(n3402), .A4(n4368), .ZN(n4549)
         );
  OAI21_X1 U4040 ( .B1(n4548), .B2(EBX_REG_1__SCAN_IN), .A(n3133), .ZN(n3149)
         );
  OR2_X1 U4041 ( .A1(n5282), .A2(n6625), .ZN(n3150) );
  AND2_X2 U4042 ( .A1(n3169), .A2(n3137), .ZN(n5339) );
  NAND2_X1 U4043 ( .A1(n4187), .A2(n3171), .ZN(U2955) );
  NAND2_X1 U4044 ( .A1(n3173), .A2(n3391), .ZN(n4572) );
  NAND2_X1 U4045 ( .A1(n3178), .A2(n3441), .ZN(n3173) );
  NAND2_X1 U4046 ( .A1(n3175), .A2(n3391), .ZN(n3174) );
  INV_X1 U4047 ( .A(n3441), .ZN(n3175) );
  NAND3_X1 U4048 ( .A1(n3178), .A2(n3441), .A3(n3177), .ZN(n3176) );
  NAND2_X1 U4049 ( .A1(n3380), .A2(n3440), .ZN(n3178) );
  NAND2_X1 U4050 ( .A1(n5973), .A2(n3182), .ZN(n3180) );
  NAND2_X1 U4051 ( .A1(n5987), .A2(n3190), .ZN(n3189) );
  NAND2_X2 U4052 ( .A1(n5689), .A2(n3129), .ZN(n5355) );
  NAND2_X2 U4053 ( .A1(n5355), .A2(n3630), .ZN(n5681) );
  NAND2_X1 U4054 ( .A1(n5290), .A2(n3196), .ZN(n5275) );
  INV_X1 U4055 ( .A(n5275), .ZN(n3973) );
  NAND2_X1 U4056 ( .A1(n4079), .A2(n3205), .ZN(n4192) );
  NAND2_X1 U4057 ( .A1(n4079), .A2(n4078), .ZN(n4190) );
  AND2_X2 U4058 ( .A1(n4079), .A2(n3136), .ZN(n4208) );
  NAND2_X1 U4059 ( .A1(n3571), .A2(n3570), .ZN(n3594) );
  INV_X1 U4060 ( .A(n3546), .ZN(n3548) );
  NAND3_X1 U4061 ( .A1(n3464), .A2(n3465), .A3(n4689), .ZN(n3546) );
  NAND2_X2 U4062 ( .A1(n3464), .A2(n3465), .ZN(n3525) );
  AND2_X1 U4063 ( .A1(n4462), .A2(n4357), .ZN(n5221) );
  NAND2_X1 U4064 ( .A1(n3467), .A2(n3466), .ZN(n3468) );
  OR2_X1 U4065 ( .A1(n4214), .A2(n4168), .ZN(n4169) );
  INV_X1 U4066 ( .A(n5220), .ZN(n4450) );
  NAND2_X1 U4067 ( .A1(n4177), .A2(n4169), .ZN(n4364) );
  INV_X1 U4068 ( .A(n4364), .ZN(n4171) );
  NAND2_X1 U4069 ( .A1(n3525), .A2(n3468), .ZN(n4623) );
  NAND2_X1 U4070 ( .A1(n4171), .A2(n4663), .ZN(n4172) );
  NAND2_X1 U4071 ( .A1(n3114), .A2(n6116), .ZN(n6334) );
  INV_X1 U4072 ( .A(n4498), .ZN(n3369) );
  NOR2_X1 U4073 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4622), .ZN(n4664) );
  OR3_X1 U4074 ( .A1(n4178), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3207) );
  AND2_X1 U4075 ( .A1(n3645), .A2(n3333), .ZN(n3208) );
  OR2_X1 U4076 ( .A1(n3607), .A2(n3611), .ZN(n3209) );
  NAND2_X1 U4077 ( .A1(n3584), .A2(n3583), .ZN(n3595) );
  NOR2_X1 U4078 ( .A1(n3343), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3210)
         );
  INV_X1 U4079 ( .A(n4174), .ZN(n3752) );
  INV_X1 U4080 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5763) );
  INV_X1 U4081 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3693) );
  INV_X1 U4082 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3691) );
  OR2_X1 U4083 ( .A1(n4445), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3211)
         );
  AND3_X1 U4084 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .A3(
        REIP_REG_22__SCAN_IN), .ZN(n3212) );
  NAND2_X1 U4085 ( .A1(n4417), .A2(n3350), .ZN(n4414) );
  AND4_X1 U4086 ( .A1(n5486), .A2(n5462), .A3(n5347), .A4(n6702), .ZN(n3214)
         );
  AND3_X1 U4087 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .A3(
        REIP_REG_7__SCAN_IN), .ZN(n3215) );
  NAND2_X1 U4088 ( .A1(n5704), .A2(n4443), .ZN(n3631) );
  INV_X1 U4089 ( .A(n6452), .ZN(n4805) );
  OR2_X1 U4090 ( .A1(n4529), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3216)
         );
  INV_X1 U4091 ( .A(n5316), .ZN(n5924) );
  NAND2_X1 U4092 ( .A1(n5927), .A2(n3349), .ZN(n5316) );
  AND2_X1 U4093 ( .A1(n3360), .A2(n3359), .ZN(n3217) );
  INV_X1 U4094 ( .A(n3367), .ZN(n3368) );
  AND2_X1 U4095 ( .A1(n4213), .A2(n4212), .ZN(n3218) );
  OR2_X1 U4096 ( .A1(n3682), .A2(n3664), .ZN(n3666) );
  INV_X1 U4097 ( .A(n4414), .ZN(n3291) );
  INV_X1 U4098 ( .A(n3488), .ZN(n3455) );
  OR2_X1 U4099 ( .A1(n3421), .A2(n3420), .ZN(n3606) );
  OR2_X1 U4100 ( .A1(n3453), .A2(n3452), .ZN(n3488) );
  INV_X1 U4101 ( .A(n3403), .ZN(n3517) );
  NOR2_X1 U4102 ( .A1(n4414), .A2(n3333), .ZN(n3364) );
  INV_X1 U4103 ( .A(n5235), .ZN(n4078) );
  OR2_X1 U4104 ( .A1(n3682), .A2(n3562), .ZN(n3560) );
  NAND2_X1 U4105 ( .A1(n3537), .A2(n3536), .ZN(n3547) );
  AND2_X1 U4106 ( .A1(n3351), .A2(n4367), .ZN(n4422) );
  AOI22_X1 U4107 ( .A1(n4122), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3278), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3248) );
  NAND2_X1 U4108 ( .A1(n4143), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3321) );
  NAND2_X1 U4109 ( .A1(n3349), .A2(n3293), .ZN(n3367) );
  AND2_X1 U4110 ( .A1(n4080), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4100)
         );
  INV_X1 U4111 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3692) );
  OAI21_X1 U4112 ( .B1(n4136), .B2(n4823), .A(n3759), .ZN(n3760) );
  OR2_X1 U4113 ( .A1(n5704), .A2(n3629), .ZN(n3630) );
  AOI22_X1 U4114 ( .A1(n3269), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3275) );
  AOI22_X1 U4115 ( .A1(n3105), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3415), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3259) );
  OR2_X1 U4116 ( .A1(n5564), .A2(n3750), .ZN(n4167) );
  NOR2_X1 U4117 ( .A1(n3752), .A2(n3691), .ZN(n3753) );
  NAND2_X1 U4118 ( .A1(n3684), .A2(n3683), .ZN(n3685) );
  NAND2_X1 U4119 ( .A1(n5221), .A2(n5891), .ZN(n4360) );
  NOR2_X1 U4120 ( .A1(n4038), .A2(n3694), .ZN(n4058) );
  INV_X1 U4121 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5874) );
  INV_X1 U4122 ( .A(n5859), .ZN(n5881) );
  INV_X1 U4123 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U4124 ( .A1(n4188), .A2(n4200), .ZN(n4205) );
  NAND2_X1 U4125 ( .A1(n5365), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5345) );
  AND2_X1 U4126 ( .A1(n4314), .A2(n4313), .ZN(n5285) );
  AND2_X1 U4127 ( .A1(n5503), .A2(n4436), .ZN(n5104) );
  OR2_X1 U4128 ( .A1(n5760), .A2(n6438), .ZN(n5727) );
  OR2_X1 U4129 ( .A1(n3114), .A2(n4625), .ZN(n4628) );
  INV_X1 U4130 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6151) );
  AND2_X1 U4131 ( .A1(n3387), .A2(n6330), .ZN(n4629) );
  INV_X1 U4132 ( .A(n5167), .ZN(n4735) );
  AOI21_X1 U4133 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6183), .A(n4610), .ZN(
        n6342) );
  NOR2_X1 U4134 ( .A1(n4219), .A2(n6434), .ZN(n4220) );
  AND2_X1 U4135 ( .A1(n4058), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4080)
         );
  XNOR2_X1 U4136 ( .A(n4183), .B(n5210), .ZN(n4234) );
  AND2_X1 U4137 ( .A1(n4234), .A2(n4232), .ZN(n5886) );
  AND2_X1 U4138 ( .A1(n5927), .A2(n3701), .ZN(n5923) );
  INV_X1 U4139 ( .A(n5965), .ZN(n4808) );
  INV_X1 U4140 ( .A(n5163), .ZN(n5969) );
  NAND2_X1 U4141 ( .A1(n3926), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3940)
         );
  NAND2_X1 U4142 ( .A1(n3898), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3912)
         );
  NOR2_X1 U4143 ( .A1(n6823), .A2(n6822), .ZN(n3726) );
  NOR3_X1 U4144 ( .A1(n4188), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(n5419), 
        .ZN(n4206) );
  OR2_X1 U4145 ( .A1(n5457), .A2(n4438), .ZN(n5442) );
  NOR2_X1 U4146 ( .A1(n3628), .A2(n5726), .ZN(n5485) );
  INV_X1 U4147 ( .A(n6103), .ZN(n6090) );
  INV_X1 U4148 ( .A(n5029), .ZN(n6106) );
  AND2_X1 U4149 ( .A1(n3483), .A2(n3494), .ZN(n4560) );
  INV_X1 U4150 ( .A(n4884), .ZN(n6187) );
  INV_X1 U4151 ( .A(n6335), .ZN(n6340) );
  INV_X1 U4152 ( .A(n6329), .ZN(n6295) );
  AND2_X1 U4153 ( .A1(n4825), .A2(n6187), .ZN(n6254) );
  NAND2_X1 U4154 ( .A1(n4781), .A2(n4780), .ZN(n6543) );
  INV_X1 U4155 ( .A(n6533), .ZN(n6369) );
  INV_X1 U4156 ( .A(n6375), .ZN(n6388) );
  INV_X1 U4157 ( .A(n4912), .ZN(n6391) );
  AND2_X1 U4158 ( .A1(n4885), .A2(n6187), .ZN(n5167) );
  NOR2_X1 U4159 ( .A1(n4705), .A2(n4610), .ZN(n6359) );
  INV_X1 U4160 ( .A(n4907), .ZN(n6383) );
  INV_X1 U4161 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6426) );
  INV_X1 U4162 ( .A(n6532), .ZN(n6495) );
  INV_X1 U4163 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6523) );
  NAND2_X1 U4164 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5842), .ZN(n5841) );
  INV_X1 U4165 ( .A(n5886), .ZN(n5902) );
  OR2_X1 U4166 ( .A1(n4234), .A2(n4233), .ZN(n5903) );
  INV_X1 U4167 ( .A(n5923), .ZN(n5301) );
  INV_X1 U4168 ( .A(n5963), .ZN(n6520) );
  OR2_X1 U4169 ( .A1(n4743), .A2(n4618), .ZN(n6025) );
  AND2_X1 U4170 ( .A1(n4446), .A2(n3211), .ZN(n4447) );
  OR2_X1 U4171 ( .A1(n4426), .A2(n4410), .ZN(n6103) );
  INV_X1 U4172 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U4173 ( .A1(n6426), .A2(n6817), .ZN(n5760) );
  AND2_X1 U4174 ( .A1(n4620), .A2(n4619), .ZN(n4665) );
  AND2_X1 U4175 ( .A1(n5048), .A2(n5047), .ZN(n5082) );
  NAND2_X1 U4176 ( .A1(n5049), .A2(n6187), .ZN(n5560) );
  OR2_X1 U4177 ( .A1(n3114), .A2(n6114), .ZN(n6180) );
  AOI21_X1 U4178 ( .B1(n6340), .B2(n6190), .A(n6186), .ZN(n6216) );
  NAND2_X1 U4179 ( .A1(n6255), .A2(n6217), .ZN(n6289) );
  NAND2_X1 U4180 ( .A1(n6255), .A2(n6254), .ZN(n6329) );
  INV_X1 U4181 ( .A(n6365), .ZN(n5536) );
  INV_X1 U4182 ( .A(n6393), .ZN(n5555) );
  OR2_X1 U4183 ( .A1(n6334), .A2(n5518), .ZN(n6533) );
  OR2_X1 U4184 ( .A1(n6334), .A2(n4949), .ZN(n6375) );
  AND2_X1 U4185 ( .A1(n4711), .A2(n4710), .ZN(n4740) );
  INV_X1 U4186 ( .A(n6347), .ZN(n5526) );
  INV_X1 U4187 ( .A(n6379), .ZN(n6539) );
  INV_X1 U4188 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6817) );
  INV_X1 U4189 ( .A(n6505), .ZN(n6447) );
  INV_X1 U4190 ( .A(n6496), .ZN(n6501) );
  OAI21_X1 U4191 ( .B1(n5413), .B2(n5773), .A(n3218), .ZN(U2958) );
  AND2_X2 U4192 ( .A1(n4581), .A2(n4510), .ZN(n3269) );
  AOI22_X1 U4193 ( .A1(n3269), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3223) );
  AOI22_X1 U4194 ( .A1(n3285), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3278), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3222) );
  AND2_X2 U4195 ( .A1(n4504), .A2(n4606), .ZN(n3872) );
  AOI22_X1 U4196 ( .A1(n3279), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3872), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3221) );
  AOI22_X1 U4197 ( .A1(n3415), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3220) );
  AND2_X2 U4198 ( .A1(n4582), .A2(n4505), .ZN(n3792) );
  AOI22_X1 U4199 ( .A1(n3792), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3229) );
  AND2_X2 U4200 ( .A1(n3144), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3225)
         );
  AND2_X2 U4201 ( .A1(n3225), .A2(n4581), .ZN(n3263) );
  AOI22_X1 U4202 ( .A1(n3263), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3228) );
  AND2_X2 U4203 ( .A1(n4582), .A2(n4510), .ZN(n3443) );
  AOI22_X1 U4204 ( .A1(n3120), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3105), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3227) );
  AND2_X2 U4205 ( .A1(n3225), .A2(n3224), .ZN(n3855) );
  AND2_X2 U4206 ( .A1(n4505), .A2(n4606), .ZN(n3410) );
  AOI22_X1 U4207 ( .A1(n3855), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3102), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3226) );
  AND4_X2 U4208 ( .A1(n3229), .A2(n3228), .A3(n3227), .A4(n3226), .ZN(n3230)
         );
  AOI22_X1 U4209 ( .A1(n3278), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3872), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3235) );
  AOI22_X1 U4210 ( .A1(n3285), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3234) );
  AOI22_X1 U4211 ( .A1(n3104), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3854), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3233) );
  AOI22_X1 U4212 ( .A1(n3269), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3106), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3232) );
  AND4_X2 U4213 ( .A1(n3235), .A2(n3234), .A3(n3233), .A4(n3232), .ZN(n3241)
         );
  AOI22_X1 U4214 ( .A1(n3270), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3239) );
  AOI22_X1 U4215 ( .A1(n4143), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3279), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3238) );
  AOI22_X1 U4216 ( .A1(n3855), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3792), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3237) );
  AOI22_X1 U4217 ( .A1(n3263), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3236) );
  AOI22_X1 U4218 ( .A1(n3269), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3245) );
  AOI22_X1 U4219 ( .A1(n3106), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3415), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3244) );
  AOI22_X1 U4220 ( .A1(n3270), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3243) );
  AOI22_X1 U4221 ( .A1(n3854), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3242) );
  NAND4_X1 U4222 ( .A1(n3245), .A2(n3244), .A3(n3243), .A4(n3242), .ZN(n3251)
         );
  AOI22_X1 U4223 ( .A1(n3792), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3249) );
  BUF_X2 U4224 ( .A(n3263), .Z(n4122) );
  AOI22_X1 U4225 ( .A1(n3855), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3872), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3247) );
  AOI22_X1 U4226 ( .A1(n3279), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3246) );
  NAND4_X1 U4227 ( .A1(n3249), .A2(n3248), .A3(n3247), .A4(n3246), .ZN(n3250)
         );
  AOI22_X1 U4228 ( .A1(n3792), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        INSTQUEUE_REG_8__6__SCAN_IN), .B2(n4143), .ZN(n3255) );
  AOI22_X1 U4229 ( .A1(n3263), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3278), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3254) );
  AOI22_X1 U4230 ( .A1(n3279), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3102), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3253) );
  AOI22_X1 U4231 ( .A1(n3855), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3872), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3252) );
  AOI22_X1 U4232 ( .A1(n3270), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3258) );
  AOI22_X1 U4233 ( .A1(n3269), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3112), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3257) );
  AOI22_X1 U4234 ( .A1(n3854), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3256) );
  OAI21_X1 U4235 ( .B1(n3357), .B2(n3701), .A(n3367), .ZN(n3262) );
  NAND2_X1 U4236 ( .A1(n3262), .A2(n3330), .ZN(n3345) );
  INV_X1 U4237 ( .A(n3345), .ZN(n3292) );
  AOI22_X1 U4238 ( .A1(n3106), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3267) );
  AOI22_X1 U4239 ( .A1(n3278), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3872), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3266) );
  AOI22_X1 U4240 ( .A1(n3279), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3265) );
  AOI22_X1 U4241 ( .A1(n3855), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3792), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3274) );
  AOI22_X1 U4242 ( .A1(n3285), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3273) );
  AOI22_X1 U4243 ( .A1(n3415), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3272) );
  NAND2_X2 U4244 ( .A1(n3277), .A2(n3276), .ZN(n3294) );
  AOI22_X1 U4245 ( .A1(n3792), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3284) );
  AOI22_X1 U4246 ( .A1(n3263), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3278), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3283) );
  AOI22_X1 U4247 ( .A1(n3855), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3872), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3282) );
  AOI21_X1 U4248 ( .B1(n3279), .B2(INSTQUEUE_REG_3__3__SCAN_IN), .A(n3280), 
        .ZN(n3281) );
  AOI22_X1 U4249 ( .A1(n3269), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3112), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3289) );
  AOI22_X1 U4250 ( .A1(n3106), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3288) );
  AOI22_X1 U4251 ( .A1(n3270), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3287) );
  AOI22_X1 U4252 ( .A1(n3120), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3286) );
  NAND2_X2 U4253 ( .A1(n3213), .A2(n3290), .ZN(n3350) );
  NAND2_X1 U4254 ( .A1(n3292), .A2(n3291), .ZN(n3687) );
  INV_X1 U4255 ( .A(n3687), .ZN(n3336) );
  MUX2_X1 U4256 ( .A(n3294), .B(n3706), .S(n3338), .Z(n3298) );
  INV_X1 U4257 ( .A(n3330), .ZN(n4368) );
  NAND2_X1 U4258 ( .A1(n3330), .A2(n3293), .ZN(n3295) );
  NAND2_X1 U4259 ( .A1(n3295), .A2(n3294), .ZN(n3297) );
  AOI22_X1 U4260 ( .A1(n3269), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3302) );
  AOI22_X1 U4261 ( .A1(n3855), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3285), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3301) );
  AOI22_X1 U4262 ( .A1(n3415), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3300) );
  AOI22_X1 U4263 ( .A1(n3263), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3279), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3299) );
  NAND4_X1 U4264 ( .A1(n3302), .A2(n3301), .A3(n3300), .A4(n3299), .ZN(n3308)
         );
  AOI22_X1 U4265 ( .A1(n3106), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3306) );
  AOI22_X1 U4266 ( .A1(n3854), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3305) );
  AOI22_X1 U4267 ( .A1(n3792), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3304) );
  AOI22_X1 U4268 ( .A1(n3278), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3872), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3303) );
  NAND4_X1 U4269 ( .A1(n3306), .A2(n3305), .A3(n3304), .A4(n3303), .ZN(n3307)
         );
  NAND2_X1 U4270 ( .A1(n3115), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3313) );
  NAND2_X1 U4271 ( .A1(n3269), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3312) );
  NAND2_X1 U4272 ( .A1(n3270), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3311)
         );
  NAND2_X1 U4273 ( .A1(n3309), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3310) );
  NAND2_X1 U4274 ( .A1(n3263), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3317)
         );
  NAND2_X1 U4275 ( .A1(n3285), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3316) );
  NAND2_X1 U4276 ( .A1(n3106), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3315) );
  NAND2_X1 U4277 ( .A1(n3278), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3314)
         );
  NAND2_X1 U4278 ( .A1(n3854), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3320)
         );
  NAND2_X1 U4279 ( .A1(n3792), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3319) );
  NAND2_X1 U4280 ( .A1(n3271), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3318) );
  NAND2_X1 U4281 ( .A1(n3855), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3325) );
  NAND2_X1 U4282 ( .A1(n3279), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3324) );
  NAND2_X1 U4283 ( .A1(n3104), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3323)
         );
  NAND2_X1 U4284 ( .A1(n3872), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3322)
         );
  NAND4_X4 U4285 ( .A1(n3329), .A2(n3328), .A3(n3327), .A4(n3326), .ZN(n3332)
         );
  NAND2_X1 U4286 ( .A1(n3373), .A2(n3108), .ZN(n3360) );
  AND2_X2 U4287 ( .A1(n3331), .A2(n3330), .ZN(n4394) );
  NAND2_X1 U4288 ( .A1(n3357), .A2(n4256), .ZN(n4421) );
  XNOR2_X1 U4289 ( .A(n6451), .B(STATE_REG_1__SCAN_IN), .ZN(n4237) );
  OAI21_X1 U4290 ( .B1(n3370), .B2(n3333), .A(n4413), .ZN(n3334) );
  NOR2_X1 U4291 ( .A1(n3353), .A2(n3334), .ZN(n3335) );
  NAND3_X1 U4292 ( .A1(n3336), .A2(n3360), .A3(n3335), .ZN(n3337) );
  NAND2_X1 U4293 ( .A1(n3337), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3363) );
  NAND2_X1 U4294 ( .A1(n3677), .A2(n3339), .ZN(n3362) );
  INV_X1 U4295 ( .A(n3690), .ZN(n3341) );
  INV_X1 U4296 ( .A(n3696), .ZN(n3340) );
  MUX2_X1 U4297 ( .A(n3341), .B(n3340), .S(n6183), .Z(n3343) );
  INV_X1 U4298 ( .A(n3343), .ZN(n3342) );
  AND2_X1 U4299 ( .A1(n3362), .A2(n3342), .ZN(n3344) );
  NAND2_X1 U4300 ( .A1(n3339), .A2(n3338), .ZN(n3346) );
  NAND2_X1 U4301 ( .A1(n3346), .A2(n3350), .ZN(n3347) );
  NOR2_X1 U4302 ( .A1(n5760), .A2(n6525), .ZN(n6437) );
  INV_X1 U4303 ( .A(n3350), .ZN(n3348) );
  NAND2_X1 U4304 ( .A1(n3348), .A2(n3365), .ZN(n4257) );
  OAI211_X1 U4305 ( .C1(n3339), .C2(n4480), .A(n6437), .B(n4257), .ZN(n3352)
         );
  NAND2_X1 U4306 ( .A1(n3349), .A2(n3338), .ZN(n3688) );
  NOR2_X1 U4307 ( .A1(n3688), .A2(n3293), .ZN(n3351) );
  INV_X1 U4308 ( .A(n3353), .ZN(n3354) );
  OAI22_X1 U4309 ( .A1(n3357), .A2(n4413), .B1(n4387), .B2(n4417), .ZN(n3358)
         );
  INV_X1 U4310 ( .A(n3358), .ZN(n3359) );
  NAND2_X1 U4311 ( .A1(n3361), .A2(n3217), .ZN(n3409) );
  NAND2_X1 U4312 ( .A1(n3408), .A2(n3409), .ZN(n3407) );
  INV_X1 U4313 ( .A(n3407), .ZN(n3380) );
  NAND2_X1 U4314 ( .A1(n3363), .A2(n3362), .ZN(n3385) );
  NAND2_X1 U4315 ( .A1(n3385), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3379) );
  XNOR2_X1 U4316 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4952) );
  OAI22_X1 U4317 ( .A1(n3696), .A2(n4952), .B1(n3690), .B2(n6151), .ZN(n3382)
         );
  INV_X1 U4318 ( .A(n3382), .ZN(n3378) );
  NAND2_X1 U4319 ( .A1(n4386), .A2(n3365), .ZN(n4219) );
  NAND3_X1 U4320 ( .A1(n5203), .A2(n3366), .A3(n4367), .ZN(n4498) );
  NAND2_X1 U4321 ( .A1(n3369), .A2(n3368), .ZN(n4406) );
  OAI21_X1 U4322 ( .B1(n4219), .B2(n3370), .A(n4406), .ZN(n3371) );
  NAND2_X1 U4323 ( .A1(n3357), .A2(n4387), .ZN(n3372) );
  NOR2_X2 U4324 ( .A1(n3373), .A2(n3372), .ZN(n5195) );
  AND2_X1 U4325 ( .A1(n3374), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3375) );
  NOR2_X2 U4326 ( .A1(n3377), .A2(n3376), .ZN(n3381) );
  NAND3_X1 U4327 ( .A1(n3379), .A2(n3378), .A3(n3381), .ZN(n3440) );
  INV_X1 U4328 ( .A(n3381), .ZN(n3384) );
  OR2_X1 U4329 ( .A1(n3382), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3383)
         );
  NAND2_X1 U4330 ( .A1(n3385), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3390) );
  NAND2_X1 U4331 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3386) );
  NAND2_X1 U4332 ( .A1(n3386), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3387) );
  NOR2_X1 U4333 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6151), .ZN(n6339)
         );
  NAND2_X1 U4334 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6339), .ZN(n6330) );
  OAI22_X1 U4335 ( .A1(n3696), .A2(n4629), .B1(n3690), .B2(n4866), .ZN(n3388)
         );
  INV_X1 U4336 ( .A(n3388), .ZN(n3389) );
  AOI22_X1 U4337 ( .A1(n3269), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3395) );
  INV_X1 U4338 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n6780) );
  AOI22_X1 U4339 ( .A1(n3422), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4340 ( .A1(n3889), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3393) );
  AOI22_X1 U4341 ( .A1(n3119), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3392) );
  NAND4_X1 U4342 ( .A1(n3395), .A2(n3394), .A3(n3393), .A4(n3392), .ZN(n3401)
         );
  AOI22_X1 U4343 ( .A1(n4087), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3399) );
  AOI22_X1 U4344 ( .A1(n4041), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3398) );
  AOI22_X1 U4345 ( .A1(n3855), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3397) );
  AOI22_X1 U4346 ( .A1(n4148), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3396) );
  NAND4_X1 U4347 ( .A1(n3399), .A2(n3398), .A3(n3397), .A4(n3396), .ZN(n3400)
         );
  INV_X1 U4348 ( .A(n3504), .ZN(n3404) );
  AOI22_X1 U4349 ( .A1(n3677), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3404), 
        .B2(n3403), .ZN(n3405) );
  INV_X1 U4350 ( .A(n3607), .ZN(n3434) );
  AOI22_X1 U4351 ( .A1(n4151), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3414) );
  AOI22_X1 U4352 ( .A1(n4041), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3413) );
  AOI22_X1 U4353 ( .A1(n4149), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3412) );
  AOI22_X1 U4354 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n3975), .B1(n4148), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3411) );
  NAND4_X1 U4355 ( .A1(n3414), .A2(n3413), .A3(n3412), .A4(n3411), .ZN(n3421)
         );
  AOI22_X1 U4356 ( .A1(n4142), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3419) );
  AOI22_X1 U4357 ( .A1(n3415), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3418) );
  AOI22_X1 U4358 ( .A1(n3119), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3417) );
  AOI22_X1 U4359 ( .A1(n3422), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3416) );
  NAND4_X1 U4360 ( .A1(n3419), .A2(n3418), .A3(n3417), .A4(n3416), .ZN(n3420)
         );
  AOI22_X1 U4361 ( .A1(n3854), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3426) );
  AOI22_X1 U4362 ( .A1(n3422), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3425) );
  AOI22_X1 U4363 ( .A1(n4041), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3424) );
  AOI22_X1 U4364 ( .A1(n3121), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3423) );
  NAND4_X1 U4365 ( .A1(n3426), .A2(n3425), .A3(n3424), .A4(n3423), .ZN(n3432)
         );
  AOI22_X1 U4366 ( .A1(n4149), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3430) );
  AOI22_X1 U4367 ( .A1(n4142), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3429) );
  AOI22_X1 U4368 ( .A1(n4151), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3428) );
  AOI22_X1 U4369 ( .A1(n4148), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3427) );
  NAND4_X1 U4370 ( .A1(n3430), .A2(n3429), .A3(n3428), .A4(n3427), .ZN(n3431)
         );
  XNOR2_X1 U4371 ( .A(n3611), .B(n3489), .ZN(n3433) );
  NAND2_X1 U4372 ( .A1(n3434), .A2(n3433), .ZN(n3474) );
  NAND2_X1 U4373 ( .A1(n3677), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3438) );
  NAND2_X1 U4374 ( .A1(n4387), .A2(n3489), .ZN(n3435) );
  OAI211_X1 U4375 ( .C1(n3611), .C2(n3338), .A(STATE2_REG_0__SCAN_IN), .B(
        n3435), .ZN(n3436) );
  INV_X1 U4376 ( .A(n3436), .ZN(n3437) );
  NAND2_X1 U4377 ( .A1(n3438), .A2(n3437), .ZN(n3473) );
  NAND2_X1 U4378 ( .A1(n3439), .A2(n3473), .ZN(n3477) );
  INV_X1 U4379 ( .A(n3485), .ZN(n3459) );
  NAND2_X1 U4380 ( .A1(n3441), .A2(n3440), .ZN(n3442) );
  XNOR2_X2 U4381 ( .A(n3442), .B(n3407), .ZN(n4496) );
  AOI22_X1 U4382 ( .A1(n4142), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3447) );
  AOI22_X1 U4383 ( .A1(n3422), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3446) );
  AOI22_X1 U4384 ( .A1(n3889), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3445) );
  AOI22_X1 U4385 ( .A1(n3120), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3444) );
  NAND4_X1 U4386 ( .A1(n3447), .A2(n3446), .A3(n3445), .A4(n3444), .ZN(n3453)
         );
  AOI22_X1 U4387 ( .A1(n4087), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4388 ( .A1(n4041), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3450) );
  INV_X1 U4389 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n6826) );
  AOI22_X1 U4390 ( .A1(n3855), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4391 ( .A1(n4148), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3448) );
  NAND4_X1 U4392 ( .A1(n3451), .A2(n3450), .A3(n3449), .A4(n3448), .ZN(n3452)
         );
  NAND2_X1 U4393 ( .A1(n3677), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3457) );
  OR2_X1 U4394 ( .A1(n3504), .A2(n3455), .ZN(n3456) );
  OAI211_X1 U4395 ( .C1(n3607), .C2(n3606), .A(n3457), .B(n3456), .ZN(n3461)
         );
  NAND2_X1 U4396 ( .A1(n3460), .A2(n3461), .ZN(n3458) );
  NAND2_X1 U4397 ( .A1(n3459), .A2(n3458), .ZN(n3463) );
  INV_X1 U4398 ( .A(n3461), .ZN(n3484) );
  NAND2_X1 U4399 ( .A1(n3486), .A2(n3484), .ZN(n3462) );
  AND2_X2 U4400 ( .A1(n3463), .A2(n3462), .ZN(n3465) );
  INV_X1 U4401 ( .A(n3464), .ZN(n3467) );
  INV_X1 U4402 ( .A(n3465), .ZN(n3466) );
  INV_X1 U4403 ( .A(n3644), .ZN(n3472) );
  NAND2_X1 U4404 ( .A1(n3489), .A2(n3488), .ZN(n3518) );
  XNOR2_X1 U4405 ( .A(n3518), .B(n3517), .ZN(n3470) );
  INV_X1 U4406 ( .A(n3110), .ZN(n6524) );
  NAND2_X1 U4407 ( .A1(n4387), .A2(n3350), .ZN(n3478) );
  INV_X1 U4408 ( .A(n3478), .ZN(n3469) );
  AOI21_X1 U4409 ( .B1(n3470), .B2(n6524), .A(n3469), .ZN(n3471) );
  NAND2_X1 U4410 ( .A1(n6038), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3496)
         );
  INV_X1 U4411 ( .A(n3473), .ZN(n3475) );
  NAND2_X1 U4412 ( .A1(n3475), .A2(n3474), .ZN(n3476) );
  OAI21_X1 U4413 ( .B1(n3110), .B2(n3489), .A(n3478), .ZN(n3479) );
  INV_X1 U4414 ( .A(n3479), .ZN(n3480) );
  NAND2_X1 U4415 ( .A1(n4513), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3481)
         );
  INV_X1 U4416 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6625) );
  NAND2_X1 U4417 ( .A1(n3481), .A2(n6625), .ZN(n3483) );
  AND2_X1 U4418 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3482) );
  NAND2_X1 U4419 ( .A1(n4513), .A2(n3482), .ZN(n3494) );
  XNOR2_X1 U4420 ( .A(n3485), .B(n3484), .ZN(n3487) );
  XNOR2_X1 U4421 ( .A(n3487), .B(n3486), .ZN(n4624) );
  NAND2_X1 U4422 ( .A1(n4624), .A2(n3644), .ZN(n3493) );
  OAI21_X1 U4423 ( .B1(n3489), .B2(n3488), .A(n3518), .ZN(n3490) );
  OAI211_X1 U4424 ( .C1(n3490), .C2(n3110), .A(n3291), .B(n3333), .ZN(n3491)
         );
  INV_X1 U4425 ( .A(n3491), .ZN(n3492) );
  NAND2_X1 U4426 ( .A1(n3493), .A2(n3492), .ZN(n4559) );
  INV_X1 U4427 ( .A(n3494), .ZN(n3495) );
  NAND2_X1 U4428 ( .A1(n3496), .A2(n6037), .ZN(n3499) );
  INV_X1 U4429 ( .A(n6038), .ZN(n3497) );
  INV_X1 U4430 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U4431 ( .A1(n3497), .A2(n6107), .ZN(n3498) );
  AND2_X1 U4432 ( .A1(n3499), .A2(n3498), .ZN(n6029) );
  NAND2_X1 U4433 ( .A1(n3385), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3503) );
  NAND3_X1 U4434 ( .A1(n6412), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6263) );
  INV_X1 U4435 ( .A(n6263), .ZN(n6261) );
  NAND2_X1 U4436 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6261), .ZN(n6257) );
  NAND2_X1 U4437 ( .A1(n6412), .A2(n6257), .ZN(n3500) );
  NAND3_X1 U4438 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4706) );
  INV_X1 U4439 ( .A(n4706), .ZN(n4830) );
  NAND2_X1 U4440 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4830), .ZN(n4861) );
  NAND2_X1 U4441 ( .A1(n3500), .A2(n4861), .ZN(n4951) );
  OAI22_X1 U4442 ( .A1(n3696), .A2(n4951), .B1(n3690), .B2(n6412), .ZN(n3501)
         );
  INV_X1 U4443 ( .A(n3501), .ZN(n3502) );
  NAND2_X1 U4444 ( .A1(n4578), .A2(n6525), .ZN(n3516) );
  INV_X1 U4445 ( .A(n3682), .ZN(n3656) );
  AOI22_X1 U4446 ( .A1(n4142), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3422), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3508) );
  AOI22_X1 U4447 ( .A1(n3116), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3507) );
  AOI22_X1 U4448 ( .A1(n3120), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3506) );
  AOI22_X1 U4449 ( .A1(n4149), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3505) );
  NAND4_X1 U4450 ( .A1(n3508), .A2(n3507), .A3(n3506), .A4(n3505), .ZN(n3514)
         );
  AOI22_X1 U4451 ( .A1(n4151), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3512) );
  AOI22_X1 U4452 ( .A1(n3121), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3511) );
  AOI22_X1 U4453 ( .A1(n4041), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3510) );
  AOI22_X1 U4454 ( .A1(n4148), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3509) );
  NAND4_X1 U4455 ( .A1(n3512), .A2(n3511), .A3(n3510), .A4(n3509), .ZN(n3513)
         );
  AOI22_X1 U4456 ( .A1(n3656), .A2(n3538), .B1(n3677), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3515) );
  NAND2_X1 U4457 ( .A1(n3725), .A2(n3644), .ZN(n3522) );
  NAND2_X1 U4458 ( .A1(n3518), .A2(n3517), .ZN(n3539) );
  INV_X1 U4459 ( .A(n3538), .ZN(n3519) );
  XNOR2_X1 U4460 ( .A(n3539), .B(n3519), .ZN(n3520) );
  NAND2_X1 U4461 ( .A1(n3520), .A2(n6524), .ZN(n3521) );
  INV_X1 U4462 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6711) );
  XNOR2_X1 U4463 ( .A(n3523), .B(n6711), .ZN(n6027) );
  NAND2_X1 U4464 ( .A1(n6029), .A2(n6027), .ZN(n6028) );
  NAND2_X1 U4465 ( .A1(n3523), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3524)
         );
  NAND2_X1 U4466 ( .A1(n6028), .A2(n3524), .ZN(n6019) );
  AOI22_X1 U4467 ( .A1(n4142), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3529) );
  AOI22_X1 U4468 ( .A1(n3422), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3528) );
  AOI22_X1 U4469 ( .A1(n3889), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3527) );
  AOI22_X1 U4470 ( .A1(n3854), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3526) );
  NAND4_X1 U4471 ( .A1(n3529), .A2(n3528), .A3(n3527), .A4(n3526), .ZN(n3535)
         );
  AOI22_X1 U4472 ( .A1(n4087), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3533) );
  AOI22_X1 U4473 ( .A1(n4041), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3532) );
  AOI22_X1 U4474 ( .A1(n4149), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3531) );
  INV_X1 U4475 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n6820) );
  AOI22_X1 U4476 ( .A1(n4148), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3530) );
  NAND4_X1 U4477 ( .A1(n3533), .A2(n3532), .A3(n3531), .A4(n3530), .ZN(n3534)
         );
  NAND2_X1 U4478 ( .A1(n3677), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3536) );
  XNOR2_X1 U4479 ( .A(n3546), .B(n3547), .ZN(n3737) );
  NAND2_X1 U4480 ( .A1(n3737), .A2(n3644), .ZN(n3542) );
  NAND2_X1 U4481 ( .A1(n3539), .A2(n3538), .ZN(n3588) );
  XNOR2_X1 U4482 ( .A(n3588), .B(n3585), .ZN(n3540) );
  NAND2_X1 U4483 ( .A1(n3540), .A2(n6524), .ZN(n3541) );
  NAND2_X1 U4484 ( .A1(n3542), .A2(n3541), .ZN(n3544) );
  INV_X1 U4485 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3543) );
  XNOR2_X1 U4486 ( .A(n3544), .B(n3543), .ZN(n6018) );
  NAND2_X1 U4487 ( .A1(n6019), .A2(n6018), .ZN(n6017) );
  NAND2_X1 U4488 ( .A1(n3544), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3545)
         );
  NAND2_X1 U4489 ( .A1(n6017), .A2(n3545), .ZN(n4673) );
  AOI22_X1 U4490 ( .A1(n3120), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3552) );
  AOI22_X1 U4491 ( .A1(n4041), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3551) );
  AOI22_X1 U4492 ( .A1(n4149), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3550) );
  AOI22_X1 U4493 ( .A1(n4151), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3549) );
  NAND4_X1 U4494 ( .A1(n3552), .A2(n3551), .A3(n3550), .A4(n3549), .ZN(n3558)
         );
  AOI22_X1 U4495 ( .A1(n4142), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3556) );
  AOI22_X1 U4496 ( .A1(n3121), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3555) );
  AOI22_X1 U4497 ( .A1(n3116), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4498 ( .A1(n3422), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3553) );
  NAND4_X1 U4499 ( .A1(n3556), .A2(n3555), .A3(n3554), .A4(n3553), .ZN(n3557)
         );
  NOR2_X1 U4500 ( .A1(n3558), .A2(n3557), .ZN(n3562) );
  NAND2_X1 U4501 ( .A1(n3677), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3559) );
  NAND2_X1 U4502 ( .A1(n3731), .A2(n3644), .ZN(n3566) );
  OR2_X1 U4503 ( .A1(n3588), .A2(n3561), .ZN(n3563) );
  INV_X1 U4504 ( .A(n3562), .ZN(n3586) );
  XNOR2_X1 U4505 ( .A(n3563), .B(n3586), .ZN(n3564) );
  NAND2_X1 U4506 ( .A1(n3564), .A2(n6524), .ZN(n3565) );
  NAND2_X1 U4507 ( .A1(n3566), .A2(n3565), .ZN(n3567) );
  INV_X1 U4508 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6580) );
  XNOR2_X1 U4509 ( .A(n3567), .B(n6580), .ZN(n4672) );
  NAND2_X1 U4510 ( .A1(n4673), .A2(n4672), .ZN(n4671) );
  NAND2_X1 U4511 ( .A1(n3567), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3568)
         );
  NAND2_X1 U4512 ( .A1(n4671), .A2(n3568), .ZN(n6005) );
  INV_X1 U4513 ( .A(n3569), .ZN(n3571) );
  AOI22_X1 U4514 ( .A1(n4142), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3575) );
  AOI22_X1 U4515 ( .A1(n3422), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3574) );
  AOI22_X1 U4516 ( .A1(n3889), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3573) );
  INV_X1 U4517 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n6563) );
  AOI22_X1 U4518 ( .A1(n3119), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3572) );
  NAND4_X1 U4519 ( .A1(n3575), .A2(n3574), .A3(n3573), .A4(n3572), .ZN(n3581)
         );
  AOI22_X1 U4520 ( .A1(n4087), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3579) );
  AOI22_X1 U4521 ( .A1(n4041), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3578) );
  AOI22_X1 U4522 ( .A1(n4149), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3577) );
  AOI22_X1 U4523 ( .A1(n4148), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3576) );
  NAND4_X1 U4524 ( .A1(n3579), .A2(n3578), .A3(n3577), .A4(n3576), .ZN(n3580)
         );
  INV_X1 U4525 ( .A(n3599), .ZN(n3582) );
  NAND2_X1 U4526 ( .A1(n3677), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3583) );
  XNOR2_X2 U4527 ( .A(n3594), .B(n3595), .ZN(n3756) );
  NAND2_X1 U4528 ( .A1(n3756), .A2(n3644), .ZN(n3591) );
  NAND2_X1 U4529 ( .A1(n3586), .A2(n3585), .ZN(n3587) );
  OR2_X1 U4530 ( .A1(n3588), .A2(n3587), .ZN(n3598) );
  XNOR2_X1 U4531 ( .A(n3598), .B(n3599), .ZN(n3589) );
  NAND2_X1 U4532 ( .A1(n3589), .A2(n6524), .ZN(n3590) );
  NAND2_X1 U4533 ( .A1(n3591), .A2(n3590), .ZN(n3592) );
  INV_X1 U4534 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6654) );
  XNOR2_X1 U4535 ( .A(n3592), .B(n6654), .ZN(n6004) );
  NAND2_X1 U4536 ( .A1(n6005), .A2(n6004), .ZN(n6003) );
  NAND2_X1 U4537 ( .A1(n3592), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3593)
         );
  NAND2_X1 U4538 ( .A1(n6003), .A2(n3593), .ZN(n5996) );
  NAND2_X1 U4539 ( .A1(n3677), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3596) );
  OAI21_X1 U4540 ( .B1(n3682), .B2(n3611), .A(n3596), .ZN(n3597) );
  NAND2_X1 U4541 ( .A1(n3757), .A2(n3644), .ZN(n3603) );
  INV_X1 U4542 ( .A(n3598), .ZN(n3600) );
  NAND2_X1 U4543 ( .A1(n3600), .A2(n3599), .ZN(n3612) );
  XNOR2_X1 U4544 ( .A(n3612), .B(n3606), .ZN(n3601) );
  NAND2_X1 U4545 ( .A1(n3601), .A2(n6524), .ZN(n3602) );
  NAND2_X1 U4546 ( .A1(n3603), .A2(n3602), .ZN(n3604) );
  INV_X1 U4547 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6072) );
  XNOR2_X1 U4548 ( .A(n3604), .B(n6072), .ZN(n5995) );
  NAND2_X1 U4549 ( .A1(n5996), .A2(n5995), .ZN(n5998) );
  NAND2_X1 U4550 ( .A1(n3604), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3605)
         );
  NAND2_X1 U4551 ( .A1(n5998), .A2(n3605), .ZN(n5987) );
  NAND2_X1 U4552 ( .A1(n3644), .A2(n3606), .ZN(n3608) );
  NOR2_X1 U4553 ( .A1(n3608), .A2(n3607), .ZN(n3609) );
  OR3_X1 U4554 ( .A1(n3612), .A2(n3611), .A3(n3110), .ZN(n3613) );
  INV_X1 U4555 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6767) );
  XNOR2_X1 U4556 ( .A(n3614), .B(n6767), .ZN(n5989) );
  NAND2_X1 U4557 ( .A1(n3614), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3615)
         );
  INV_X1 U4558 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U4559 ( .A1(n5704), .A2(n5981), .ZN(n3616) );
  INV_X1 U4560 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3617) );
  NAND2_X1 U4561 ( .A1(n5704), .A2(n3617), .ZN(n5020) );
  AND2_X1 U4562 ( .A1(n5704), .A2(n6052), .ZN(n3620) );
  OR2_X1 U4563 ( .A1(n5704), .A2(n3617), .ZN(n5972) );
  INV_X1 U4564 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5105) );
  NOR2_X1 U4565 ( .A1(n5704), .A2(n5105), .ZN(n5091) );
  XNOR2_X1 U4566 ( .A(n5704), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5501)
         );
  AND2_X1 U4567 ( .A1(n5704), .A2(n5753), .ZN(n3622) );
  OR2_X1 U4568 ( .A1(n5704), .A2(n5753), .ZN(n3621) );
  INV_X1 U4569 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6564) );
  NOR2_X1 U4570 ( .A1(n5704), .A2(n6564), .ZN(n3623) );
  OR2_X2 U4571 ( .A1(n5390), .A2(n3623), .ZN(n5689) );
  NAND2_X1 U4572 ( .A1(n5704), .A2(n6564), .ZN(n3624) );
  INV_X1 U4573 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6579) );
  NAND2_X1 U4574 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3626) );
  NAND2_X1 U4575 ( .A1(n5704), .A2(n3626), .ZN(n3627) );
  INV_X1 U4576 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6717) );
  INV_X1 U4577 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3628) );
  AND3_X1 U4578 ( .A1(n6717), .A2(n3628), .A3(n6579), .ZN(n3629) );
  NOR2_X1 U4579 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5486) );
  NOR2_X1 U4580 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5462) );
  INV_X1 U4581 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5347) );
  INV_X1 U4582 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6702) );
  AND2_X1 U4583 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5463) );
  AND2_X1 U4584 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5487) );
  AND2_X1 U4585 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4437) );
  NAND3_X1 U4586 ( .A1(n5463), .A2(n5487), .A3(n4437), .ZN(n4443) );
  XOR2_X1 U4587 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(n5704), .Z(n5433) );
  INV_X1 U4588 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5427) );
  INV_X1 U4589 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5426) );
  NOR2_X1 U4590 ( .A1(n5693), .A2(n5426), .ZN(n5338) );
  NAND2_X1 U4591 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5405) );
  NOR2_X2 U4592 ( .A1(n4188), .A2(n5405), .ZN(n4380) );
  NOR2_X1 U4593 ( .A1(n5704), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5337)
         );
  NOR2_X1 U4594 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U4595 ( .A1(n5337), .A2(n5406), .ZN(n4178) );
  AOI21_X1 U4596 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n4380), .A(n4382), 
        .ZN(n3633) );
  XNOR2_X1 U4597 ( .A(n3633), .B(n5400), .ZN(n5404) );
  XNOR2_X1 U4598 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3646) );
  NAND2_X1 U4599 ( .A1(n3649), .A2(n3646), .ZN(n3635) );
  NAND2_X1 U4600 ( .A1(n6151), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3634) );
  NAND2_X1 U4601 ( .A1(n3635), .A2(n3634), .ZN(n3663) );
  XNOR2_X1 U4602 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3661) );
  NAND2_X1 U4603 ( .A1(n3663), .A2(n3661), .ZN(n3637) );
  NAND2_X1 U4604 ( .A1(n4866), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3636) );
  XNOR2_X1 U4605 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3673) );
  NAND2_X1 U4606 ( .A1(n3672), .A2(n3673), .ZN(n3639) );
  NAND2_X1 U4607 ( .A1(n6412), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3638) );
  NAND2_X1 U4608 ( .A1(n3639), .A2(n3638), .ZN(n3643) );
  NAND2_X1 U4609 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n5763), .ZN(n3641) );
  OR2_X1 U4610 ( .A1(n3682), .A2(n3374), .ZN(n3645) );
  INV_X1 U4611 ( .A(n3646), .ZN(n3647) );
  XNOR2_X1 U4612 ( .A(n3647), .B(n3649), .ZN(n4223) );
  NAND2_X1 U4613 ( .A1(n4223), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3660) );
  AND2_X1 U4614 ( .A1(n3374), .A2(n3333), .ZN(n3648) );
  NOR2_X1 U4615 ( .A1(n3108), .A2(n3648), .ZN(n3667) );
  INV_X1 U4616 ( .A(n3649), .ZN(n3651) );
  NAND2_X1 U4617 ( .A1(n3144), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3650) );
  NAND2_X1 U4618 ( .A1(n3651), .A2(n3650), .ZN(n3655) );
  OAI21_X1 U4619 ( .B1(n3357), .B2(n3655), .A(n3652), .ZN(n3653) );
  INV_X1 U4620 ( .A(n4223), .ZN(n3654) );
  INV_X1 U4621 ( .A(n3655), .ZN(n3657) );
  OAI211_X1 U4622 ( .C1(n3208), .C2(n3660), .A(n3659), .B(n3658), .ZN(n3671)
         );
  INV_X1 U4623 ( .A(n3677), .ZN(n3665) );
  INV_X1 U4624 ( .A(n3661), .ZN(n3662) );
  XNOR2_X1 U4625 ( .A(n3663), .B(n3662), .ZN(n4222) );
  INV_X1 U4626 ( .A(n4222), .ZN(n3664) );
  OAI211_X1 U4627 ( .C1(n3665), .C2(n4222), .A(n3666), .B(n3667), .ZN(n3670)
         );
  INV_X1 U4628 ( .A(n3666), .ZN(n3669) );
  INV_X1 U4629 ( .A(n3667), .ZN(n3668) );
  AOI22_X1 U4630 ( .A1(n3671), .A2(n3670), .B1(n3669), .B2(n3668), .ZN(n3675)
         );
  XOR2_X1 U4631 ( .A(n3673), .B(n3672), .Z(n4224) );
  NOR2_X1 U4632 ( .A1(n3677), .A2(n4224), .ZN(n3674) );
  OAI22_X1 U4633 ( .A1(n3675), .A2(n3674), .B1(n4224), .B2(n3679), .ZN(n3676)
         );
  OAI21_X1 U4634 ( .B1(n4221), .B2(n3679), .A(n3678), .ZN(n3680) );
  OAI21_X1 U4635 ( .B1(n4226), .B2(n3682), .A(n3681), .ZN(n3686) );
  INV_X1 U4636 ( .A(n4226), .ZN(n3683) );
  AND2_X1 U4637 ( .A1(n4503), .A2(n4387), .ZN(n3689) );
  AND2_X1 U4638 ( .A1(n4398), .A2(n3357), .ZN(n4405) );
  INV_X1 U4639 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5633) );
  INV_X1 U4640 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3992) );
  NAND2_X1 U4641 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3694) );
  INV_X1 U4642 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n3695) );
  XNOR2_X1 U4643 ( .A(n4182), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5564)
         );
  NOR2_X2 U4644 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6335) );
  AND2_X1 U4645 ( .A1(n3696), .A2(n6340), .ZN(n6519) );
  NOR2_X1 U4646 ( .A1(n6519), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3697) );
  NAND2_X1 U4647 ( .A1(n6525), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3699) );
  NAND2_X1 U4648 ( .A1(n6523), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3698) );
  NAND2_X1 U4649 ( .A1(n3699), .A2(n3698), .ZN(n4514) );
  INV_X1 U4650 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4181) );
  NOR2_X1 U4651 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_0__SCAN_IN), .ZN(
        n6446) );
  INV_X1 U4652 ( .A(n6446), .ZN(n6438) );
  NAND2_X1 U4653 ( .A1(n4228), .A2(REIP_REG_30__SCAN_IN), .ZN(n5397) );
  OAI21_X1 U4654 ( .B1(n5393), .B2(n4181), .A(n5397), .ZN(n3700) );
  AOI21_X1 U4655 ( .B1(n5564), .B2(n6022), .A(n3700), .ZN(n4173) );
  INV_X2 U4656 ( .A(n4623), .ZN(n5519) );
  INV_X1 U4657 ( .A(n3877), .ZN(n3708) );
  NOR2_X2 U4658 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6523), .ZN(n4174) );
  NAND2_X1 U4659 ( .A1(n4624), .A2(n3877), .ZN(n3705) );
  NOR2_X1 U4660 ( .A1(n3367), .A2(n6522), .ZN(n3738) );
  INV_X1 U4661 ( .A(EAX_REG_1__SCAN_IN), .ZN(n3702) );
  OAI22_X1 U4662 ( .A1(n4136), .A2(n3702), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6823), .ZN(n3703) );
  AOI21_X1 U4663 ( .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n3738), .A(n3703), 
        .ZN(n3704) );
  NAND2_X1 U4664 ( .A1(n3705), .A2(n3704), .ZN(n4553) );
  AOI21_X1 U4665 ( .B1(n4884), .B2(n3706), .A(n6522), .ZN(n4517) );
  OR2_X1 U4666 ( .A1(n3707), .A2(n3708), .ZN(n3713) );
  INV_X1 U4667 ( .A(EAX_REG_0__SCAN_IN), .ZN(n3710) );
  NAND2_X1 U4668 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n6522), .ZN(n3709)
         );
  OAI21_X1 U4669 ( .B1(n4136), .B2(n3710), .A(n3709), .ZN(n3711) );
  AOI21_X1 U4670 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n3738), .A(n3711), 
        .ZN(n3712) );
  NAND2_X1 U4671 ( .A1(n3713), .A2(n3712), .ZN(n4516) );
  NAND2_X1 U4672 ( .A1(n4517), .A2(n4516), .ZN(n4515) );
  INV_X1 U4673 ( .A(n4516), .ZN(n3714) );
  NAND2_X1 U4674 ( .A1(n6522), .A2(n6523), .ZN(n3750) );
  NAND2_X1 U4675 ( .A1(n3714), .A2(n4141), .ZN(n3715) );
  NAND2_X1 U4676 ( .A1(n4515), .A2(n3715), .ZN(n4552) );
  NAND2_X1 U4677 ( .A1(n4553), .A2(n4552), .ZN(n4555) );
  INV_X1 U4678 ( .A(EAX_REG_2__SCAN_IN), .ZN(n3719) );
  NAND2_X1 U4679 ( .A1(n3738), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3718) );
  AOI21_X1 U4680 ( .B1(n6823), .B2(n6822), .A(n3726), .ZN(n3716) );
  INV_X1 U4681 ( .A(n3716), .ZN(n6046) );
  AOI22_X1 U4682 ( .A1(n6046), .A2(n4141), .B1(PHYADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n4174), .ZN(n3717) );
  OAI211_X1 U4683 ( .C1(n4136), .C2(n3719), .A(n3718), .B(n3717), .ZN(n4702)
         );
  NAND2_X1 U4684 ( .A1(n4703), .A2(n4702), .ZN(n3724) );
  INV_X1 U4685 ( .A(n3720), .ZN(n3722) );
  INV_X1 U4686 ( .A(n4555), .ZN(n3721) );
  NAND2_X1 U4687 ( .A1(n3722), .A2(n3721), .ZN(n3723) );
  NAND2_X1 U4688 ( .A1(n3114), .A2(n3877), .ZN(n3730) );
  INV_X1 U4689 ( .A(EAX_REG_3__SCAN_IN), .ZN(n4700) );
  OAI21_X1 U4690 ( .B1(n3726), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n3743), 
        .ZN(n6035) );
  AOI22_X1 U4691 ( .A1(n4174), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .B1(n4141), 
        .B2(n6035), .ZN(n3727) );
  OAI21_X1 U4692 ( .B1(n4136), .B2(n4700), .A(n3727), .ZN(n3728) );
  AOI21_X1 U4693 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n3738), .A(n3728), 
        .ZN(n3729) );
  NAND2_X1 U4694 ( .A1(n3730), .A2(n3729), .ZN(n4699) );
  INV_X1 U4695 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3733) );
  OAI21_X1 U4696 ( .B1(n3742), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3749), 
        .ZN(n6016) );
  AOI22_X1 U4697 ( .A1(n4174), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .B1(n4141), 
        .B2(n6016), .ZN(n3732) );
  NAND2_X1 U4698 ( .A1(n3737), .A2(n3877), .ZN(n3747) );
  INV_X1 U4699 ( .A(EAX_REG_4__SCAN_IN), .ZN(n3741) );
  NAND2_X1 U4700 ( .A1(n3738), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3740) );
  OAI21_X1 U4701 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n6523), .A(n6522), 
        .ZN(n3739) );
  OAI211_X1 U4702 ( .C1(n4136), .C2(n3741), .A(n3740), .B(n3739), .ZN(n3745)
         );
  AOI21_X1 U4703 ( .B1(n6550), .B2(n3743), .A(n3742), .ZN(n6021) );
  NAND2_X1 U4704 ( .A1(n6021), .A2(n4141), .ZN(n3744) );
  NAND2_X1 U4705 ( .A1(n3745), .A2(n3744), .ZN(n3746) );
  NAND2_X1 U4706 ( .A1(n3747), .A2(n3746), .ZN(n4617) );
  XNOR2_X1 U4707 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .B(n3749), .ZN(n6007) );
  INV_X1 U4708 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3751) );
  OAI22_X1 U4709 ( .A1(n6007), .A2(n3750), .B1(n3751), .B2(n4136), .ZN(n3754)
         );
  NAND2_X1 U4710 ( .A1(n3757), .A2(n3877), .ZN(n3762) );
  INV_X1 U4711 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4823) );
  OAI21_X1 U4712 ( .B1(n3758), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3763), 
        .ZN(n6002) );
  AOI22_X1 U4713 ( .A1(n4174), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .B1(n4141), 
        .B2(n6002), .ZN(n3759) );
  XNOR2_X1 U4714 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3763), .ZN(n5991) );
  INV_X1 U4715 ( .A(n5991), .ZN(n3778) );
  INV_X1 U4716 ( .A(EAX_REG_8__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4717 ( .A1(n3119), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4718 ( .A1(n4151), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4719 ( .A1(n3116), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4720 ( .A1(n4041), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3764) );
  NAND4_X1 U4721 ( .A1(n3767), .A2(n3766), .A3(n3765), .A4(n3764), .ZN(n3773)
         );
  AOI22_X1 U4722 ( .A1(n3422), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3771) );
  AOI22_X1 U4723 ( .A1(n4149), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4724 ( .A1(n4142), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3769) );
  AOI22_X1 U4725 ( .A1(n4148), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3768) );
  NAND4_X1 U4726 ( .A1(n3771), .A2(n3770), .A3(n3769), .A4(n3768), .ZN(n3772)
         );
  OAI21_X1 U4727 ( .B1(n3773), .B2(n3772), .A(n3877), .ZN(n3775) );
  NAND2_X1 U4728 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n4174), .ZN(n3774)
         );
  OAI211_X1 U4729 ( .C1(n3776), .C2(n4136), .A(n3775), .B(n3774), .ZN(n3777)
         );
  AOI21_X1 U4730 ( .B1(n3778), .B2(n4141), .A(n3777), .ZN(n4759) );
  XNOR2_X1 U4731 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3779), .ZN(n5983) );
  AOI22_X1 U4732 ( .A1(n4175), .A2(EAX_REG_9__SCAN_IN), .B1(n4174), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4733 ( .A1(n3116), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4734 ( .A1(n4149), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4735 ( .A1(n3889), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4736 ( .A1(n4148), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3780) );
  NAND4_X1 U4737 ( .A1(n3783), .A2(n3782), .A3(n3781), .A4(n3780), .ZN(n3789)
         );
  AOI22_X1 U4738 ( .A1(n3854), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4739 ( .A1(n3422), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4740 ( .A1(n4041), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4741 ( .A1(n4123), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3784) );
  NAND4_X1 U4742 ( .A1(n3787), .A2(n3786), .A3(n3785), .A4(n3784), .ZN(n3788)
         );
  OAI21_X1 U4743 ( .B1(n3789), .B2(n3788), .A(n3877), .ZN(n3790) );
  OAI211_X1 U4744 ( .C1(n5983), .C2(n3750), .A(n3791), .B(n3790), .ZN(n4768)
         );
  INV_X1 U4745 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5024) );
  AOI22_X1 U4746 ( .A1(n4142), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4747 ( .A1(n4148), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4748 ( .A1(n3116), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4749 ( .A1(n3422), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3793) );
  NAND4_X1 U4750 ( .A1(n3796), .A2(n3795), .A3(n3794), .A4(n3793), .ZN(n3802)
         );
  AOI22_X1 U4751 ( .A1(n3120), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3800) );
  AOI22_X1 U4752 ( .A1(n4041), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3799) );
  AOI22_X1 U4753 ( .A1(n4149), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4754 ( .A1(n3889), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3797) );
  NAND4_X1 U4755 ( .A1(n3800), .A2(n3799), .A3(n3798), .A4(n3797), .ZN(n3801)
         );
  OAI21_X1 U4756 ( .B1(n3802), .B2(n3801), .A(n3877), .ZN(n3803) );
  OAI21_X1 U4757 ( .B1(n5024), .B2(n3752), .A(n3803), .ZN(n3806) );
  XOR2_X1 U4758 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3804), .Z(n5860) );
  NOR2_X1 U4759 ( .A1(n5860), .A2(n3750), .ZN(n3805) );
  AOI211_X1 U4760 ( .C1(n4175), .C2(EAX_REG_10__SCAN_IN), .A(n3806), .B(n3805), 
        .ZN(n4863) );
  NOR2_X2 U4761 ( .A1(n4766), .A2(n4863), .ZN(n4862) );
  AOI21_X1 U4762 ( .B1(n6553), .B2(n3807), .A(n3830), .ZN(n5976) );
  AOI22_X1 U4763 ( .A1(n4175), .A2(EAX_REG_11__SCAN_IN), .B1(n4174), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3819) );
  AOI22_X1 U4764 ( .A1(n4041), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4765 ( .A1(n4149), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4766 ( .A1(n3889), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4767 ( .A1(n3104), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3808) );
  NAND4_X1 U4768 ( .A1(n3811), .A2(n3810), .A3(n3809), .A4(n3808), .ZN(n3817)
         );
  AOI22_X1 U4769 ( .A1(n3119), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3815) );
  AOI22_X1 U4770 ( .A1(n3422), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3814) );
  AOI22_X1 U4771 ( .A1(n4087), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3813) );
  AOI22_X1 U4772 ( .A1(n4123), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3812) );
  NAND4_X1 U4773 ( .A1(n3815), .A2(n3814), .A3(n3813), .A4(n3812), .ZN(n3816)
         );
  OAI21_X1 U4774 ( .B1(n3817), .B2(n3816), .A(n3877), .ZN(n3818) );
  OAI211_X1 U4775 ( .C1(n5976), .C2(n3750), .A(n3819), .B(n3818), .ZN(n4930)
         );
  NAND2_X1 U4776 ( .A1(n4862), .A2(n4930), .ZN(n4928) );
  AOI22_X1 U4777 ( .A1(n3120), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4778 ( .A1(n3889), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4779 ( .A1(n3116), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4780 ( .A1(n4041), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3820) );
  NAND4_X1 U4781 ( .A1(n3823), .A2(n3822), .A3(n3821), .A4(n3820), .ZN(n3829)
         );
  AOI22_X1 U4782 ( .A1(n3422), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4783 ( .A1(n4142), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4784 ( .A1(n4149), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4785 ( .A1(n4151), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3824) );
  NAND4_X1 U4786 ( .A1(n3827), .A2(n3826), .A3(n3825), .A4(n3824), .ZN(n3828)
         );
  OR2_X1 U4787 ( .A1(n3829), .A2(n3828), .ZN(n3834) );
  INV_X1 U4788 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5843) );
  XNOR2_X1 U4789 ( .A(n5843), .B(n3830), .ZN(n5845) );
  OAI21_X1 U4790 ( .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6523), .A(n6522), 
        .ZN(n3832) );
  NAND2_X1 U4791 ( .A1(n4175), .A2(EAX_REG_12__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4792 ( .A1(n5845), .A2(n4141), .B1(n3832), .B2(n3831), .ZN(n3833)
         );
  AOI21_X1 U4793 ( .B1(n3877), .B2(n3834), .A(n3833), .ZN(n5017) );
  NOR2_X2 U4794 ( .A1(n4928), .A2(n5017), .ZN(n3849) );
  XOR2_X1 U4795 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(n3835), .Z(n5712) );
  INV_X1 U4796 ( .A(EAX_REG_13__SCAN_IN), .ZN(n3836) );
  OAI22_X1 U4797 ( .A1(n4136), .A2(n3836), .B1(n3752), .B2(n3693), .ZN(n3837)
         );
  AOI21_X1 U4798 ( .B1(n5712), .B2(n4141), .A(n3837), .ZN(n3850) );
  XNOR2_X1 U4799 ( .A(n3849), .B(n3850), .ZN(n5083) );
  AOI22_X1 U4800 ( .A1(n4142), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4801 ( .A1(n3422), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4802 ( .A1(n3889), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4803 ( .A1(n3120), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3838) );
  NAND4_X1 U4804 ( .A1(n3841), .A2(n3840), .A3(n3839), .A4(n3838), .ZN(n3847)
         );
  AOI22_X1 U4805 ( .A1(n4087), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4806 ( .A1(n4041), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4807 ( .A1(n4149), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3843) );
  AOI22_X1 U4808 ( .A1(n4148), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3842) );
  NAND4_X1 U4809 ( .A1(n3845), .A2(n3844), .A3(n3843), .A4(n3842), .ZN(n3846)
         );
  OR2_X1 U4810 ( .A1(n3847), .A2(n3846), .ZN(n3848) );
  AND2_X1 U4811 ( .A1(n3877), .A2(n3848), .ZN(n5084) );
  NAND2_X1 U4812 ( .A1(n5083), .A2(n5084), .ZN(n5085) );
  INV_X1 U4813 ( .A(n3850), .ZN(n3851) );
  NAND2_X1 U4814 ( .A1(n3849), .A2(n3851), .ZN(n3852) );
  XOR2_X1 U4815 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3853), .Z(n5824) );
  AOI22_X1 U4816 ( .A1(n4175), .A2(EAX_REG_14__SCAN_IN), .B1(n4174), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3867) );
  AOI22_X1 U4817 ( .A1(n3854), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4818 ( .A1(n4151), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4819 ( .A1(n3855), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4820 ( .A1(n3116), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3856) );
  NAND4_X1 U4821 ( .A1(n3859), .A2(n3858), .A3(n3857), .A4(n3856), .ZN(n3865)
         );
  AOI22_X1 U4822 ( .A1(n3269), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4823 ( .A1(n3422), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4824 ( .A1(n4148), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4825 ( .A1(n4041), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3860) );
  NAND4_X1 U4826 ( .A1(n3863), .A2(n3862), .A3(n3861), .A4(n3860), .ZN(n3864)
         );
  OAI21_X1 U4827 ( .B1(n3865), .B2(n3864), .A(n3877), .ZN(n3866) );
  OAI211_X1 U4828 ( .C1(n5824), .C2(n3750), .A(n3867), .B(n3866), .ZN(n5112)
         );
  INV_X1 U4829 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5392) );
  AOI22_X1 U4830 ( .A1(INSTQUEUE_REG_4__7__SCAN_IN), .A2(n4149), .B1(n3422), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4831 ( .A1(n4142), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4832 ( .A1(n3119), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3869) );
  AOI22_X1 U4833 ( .A1(n3121), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3868) );
  NAND4_X1 U4834 ( .A1(n3871), .A2(n3870), .A3(n3869), .A4(n3868), .ZN(n3879)
         );
  AOI22_X1 U4835 ( .A1(n4041), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4836 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n3116), .B1(n3109), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4837 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4123), .B1(n4148), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4838 ( .A1(n4151), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3873) );
  NAND4_X1 U4839 ( .A1(n3876), .A2(n3875), .A3(n3874), .A4(n3873), .ZN(n3878)
         );
  OAI21_X1 U4840 ( .B1(n3879), .B2(n3878), .A(n3877), .ZN(n3880) );
  OAI21_X1 U4841 ( .B1(n5392), .B2(n3752), .A(n3880), .ZN(n3883) );
  XOR2_X1 U4842 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3881), .Z(n5815) );
  NOR2_X1 U4843 ( .A1(n5815), .A2(n3750), .ZN(n3882) );
  AOI211_X1 U4844 ( .C1(n4175), .C2(EAX_REG_15__SCAN_IN), .A(n3883), .B(n3882), 
        .ZN(n5307) );
  XNOR2_X1 U4845 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3884), .ZN(n5805)
         );
  AOI22_X1 U4846 ( .A1(n4175), .A2(EAX_REG_16__SCAN_IN), .B1(n4174), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4847 ( .A1(n4149), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3422), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4848 ( .A1(n4041), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4849 ( .A1(n4151), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4850 ( .A1(n3279), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3885) );
  NAND4_X1 U4851 ( .A1(n3888), .A2(n3887), .A3(n3886), .A4(n3885), .ZN(n3895)
         );
  AOI22_X1 U4852 ( .A1(n3120), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4853 ( .A1(n3889), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4854 ( .A1(n3121), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4855 ( .A1(n4123), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3890) );
  NAND4_X1 U4856 ( .A1(n3893), .A2(n3892), .A3(n3891), .A4(n3890), .ZN(n3894)
         );
  OAI21_X1 U4857 ( .B1(n3895), .B2(n3894), .A(n4138), .ZN(n3896) );
  OAI211_X1 U4858 ( .C1(n5805), .C2(n3750), .A(n3897), .B(n3896), .ZN(n5303)
         );
  OAI21_X1 U4859 ( .B1(n3898), .B2(PHYADDRPOINTER_REG_17__SCAN_IN), .A(n3912), 
        .ZN(n5797) );
  AOI22_X1 U4860 ( .A1(n4175), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6522), .ZN(n3910) );
  AOI22_X1 U4861 ( .A1(n4041), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3902) );
  AOI22_X1 U4862 ( .A1(n3422), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4863 ( .A1(n4149), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4864 ( .A1(n4151), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3899) );
  NAND4_X1 U4865 ( .A1(n3902), .A2(n3901), .A3(n3900), .A4(n3899), .ZN(n3908)
         );
  AOI22_X1 U4866 ( .A1(n3119), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4867 ( .A1(n3889), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4868 ( .A1(n3109), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4869 ( .A1(n3279), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3903) );
  NAND4_X1 U4870 ( .A1(n3906), .A2(n3905), .A3(n3904), .A4(n3903), .ZN(n3907)
         );
  OAI21_X1 U4871 ( .B1(n3908), .B2(n3907), .A(n4138), .ZN(n3909) );
  NAND3_X1 U4872 ( .A1(n3750), .A2(n3910), .A3(n3909), .ZN(n3911) );
  OAI21_X1 U4873 ( .B1(n3750), .B2(n5797), .A(n3911), .ZN(n5299) );
  XNOR2_X1 U4874 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n3912), .ZN(n5789)
         );
  AOI22_X1 U4875 ( .A1(n4087), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4876 ( .A1(n4041), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4877 ( .A1(n4149), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4878 ( .A1(n3279), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3913) );
  NAND4_X1 U4879 ( .A1(n3916), .A2(n3915), .A3(n3914), .A4(n3913), .ZN(n3922)
         );
  AOI22_X1 U4880 ( .A1(n4142), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4881 ( .A1(n3106), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3919) );
  AOI22_X1 U4882 ( .A1(n3889), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4883 ( .A1(n3120), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3917) );
  NAND4_X1 U4884 ( .A1(n3920), .A2(n3919), .A3(n3918), .A4(n3917), .ZN(n3921)
         );
  OR2_X1 U4885 ( .A1(n3922), .A2(n3921), .ZN(n3923) );
  AOI22_X1 U4886 ( .A1(n4138), .A2(n3923), .B1(n4175), .B2(EAX_REG_18__SCAN_IN), .ZN(n3925) );
  OAI21_X1 U4887 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6523), .A(n6522), 
        .ZN(n3924) );
  AOI22_X1 U4888 ( .A1(n4141), .A2(n5789), .B1(n3925), .B2(n3924), .ZN(n5292)
         );
  OAI21_X1 U4889 ( .B1(n3926), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n3940), 
        .ZN(n5688) );
  AOI22_X1 U4890 ( .A1(n4175), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6522), .ZN(n3938) );
  AOI22_X1 U4891 ( .A1(n4142), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4892 ( .A1(n3116), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4893 ( .A1(n3119), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4894 ( .A1(n3422), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3927) );
  NAND4_X1 U4895 ( .A1(n3930), .A2(n3929), .A3(n3928), .A4(n3927), .ZN(n3936)
         );
  AOI22_X1 U4896 ( .A1(n4041), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4897 ( .A1(n4149), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4898 ( .A1(n4151), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4899 ( .A1(n3279), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3931) );
  NAND4_X1 U4900 ( .A1(n3934), .A2(n3933), .A3(n3932), .A4(n3931), .ZN(n3935)
         );
  OAI21_X1 U4901 ( .B1(n3936), .B2(n3935), .A(n4138), .ZN(n3937) );
  NAND3_X1 U4902 ( .A1(n3750), .A2(n3938), .A3(n3937), .ZN(n3939) );
  OAI21_X1 U4903 ( .B1(n3750), .B2(n5688), .A(n3939), .ZN(n5278) );
  XNOR2_X1 U4904 ( .A(n3940), .B(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5385)
         );
  AOI22_X1 U4905 ( .A1(n4142), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4906 ( .A1(n3422), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4907 ( .A1(n3889), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4908 ( .A1(n3119), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3941) );
  NAND4_X1 U4909 ( .A1(n3944), .A2(n3943), .A3(n3942), .A4(n3941), .ZN(n3950)
         );
  AOI22_X1 U4910 ( .A1(n4087), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4911 ( .A1(n4122), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4912 ( .A1(n4149), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4913 ( .A1(n3279), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3945) );
  NAND4_X1 U4914 ( .A1(n3948), .A2(n3947), .A3(n3946), .A4(n3945), .ZN(n3949)
         );
  OR2_X1 U4915 ( .A1(n3950), .A2(n3949), .ZN(n3954) );
  INV_X1 U4916 ( .A(EAX_REG_20__SCAN_IN), .ZN(n3952) );
  OAI21_X1 U4917 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6523), .A(n6522), 
        .ZN(n3951) );
  OAI21_X1 U4918 ( .B1(n4136), .B2(n3952), .A(n3951), .ZN(n3953) );
  AOI21_X1 U4919 ( .B1(n4138), .B2(n3954), .A(n3953), .ZN(n3955) );
  AOI21_X1 U4920 ( .B1(n5385), .B2(n4141), .A(n3955), .ZN(n5276) );
  AND2_X1 U4921 ( .A1(n3956), .A2(n5373), .ZN(n3957) );
  NOR2_X1 U4922 ( .A1(n3974), .A2(n3957), .ZN(n5627) );
  NAND2_X1 U4923 ( .A1(n5627), .A2(n4141), .ZN(n3971) );
  AOI22_X1 U4924 ( .A1(n4175), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6522), .ZN(n3969) );
  AOI22_X1 U4925 ( .A1(n4142), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4926 ( .A1(n3106), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4927 ( .A1(n4041), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4928 ( .A1(n3121), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3958) );
  NAND4_X1 U4929 ( .A1(n3961), .A2(n3960), .A3(n3959), .A4(n3958), .ZN(n3967)
         );
  AOI22_X1 U4930 ( .A1(n4149), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U4931 ( .A1(n3854), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U4932 ( .A1(n4151), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4933 ( .A1(n3279), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3962) );
  NAND4_X1 U4934 ( .A1(n3965), .A2(n3964), .A3(n3963), .A4(n3962), .ZN(n3966)
         );
  OAI21_X1 U4935 ( .B1(n3967), .B2(n3966), .A(n4138), .ZN(n3968) );
  NAND3_X1 U4936 ( .A1(n3750), .A2(n3969), .A3(n3968), .ZN(n3970) );
  NAND2_X1 U4937 ( .A1(n3971), .A2(n3970), .ZN(n5371) );
  NAND2_X1 U4938 ( .A1(n3973), .A2(n3972), .ZN(n5260) );
  INV_X1 U4939 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5367) );
  XNOR2_X1 U4940 ( .A(n3974), .B(n5367), .ZN(n5617) );
  NAND2_X1 U4941 ( .A1(n5617), .A2(n4141), .ZN(n3991) );
  AOI22_X1 U4942 ( .A1(n4149), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4943 ( .A1(n4142), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4944 ( .A1(n4123), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4945 ( .A1(n3889), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3976) );
  NAND4_X1 U4946 ( .A1(n3979), .A2(n3978), .A3(n3977), .A4(n3976), .ZN(n3986)
         );
  AOI22_X1 U4947 ( .A1(n3119), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3106), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U4948 ( .A1(n4151), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U4949 ( .A1(n3116), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4950 ( .A1(n4041), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3981) );
  NAND4_X1 U4951 ( .A1(n3984), .A2(n3983), .A3(n3982), .A4(n3981), .ZN(n3985)
         );
  OAI21_X1 U4952 ( .B1(n3986), .B2(n3985), .A(n4138), .ZN(n3989) );
  OAI21_X1 U4953 ( .B1(n5367), .B2(STATE2_REG_2__SCAN_IN), .A(n3750), .ZN(
        n3987) );
  AOI21_X1 U4954 ( .B1(n4175), .B2(EAX_REG_22__SCAN_IN), .A(n3987), .ZN(n3988)
         );
  NAND2_X1 U4955 ( .A1(n3989), .A2(n3988), .ZN(n3990) );
  NAND2_X1 U4956 ( .A1(n3991), .A2(n3990), .ZN(n5259) );
  NAND2_X1 U4957 ( .A1(n3993), .A2(n3992), .ZN(n3994) );
  NAND2_X1 U4958 ( .A1(n4038), .A2(n3994), .ZN(n5609) );
  INV_X1 U4959 ( .A(n5609), .ZN(n4020) );
  AOI22_X1 U4960 ( .A1(n3854), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4961 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4122), .B1(n3121), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U4962 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n4087), .B1(n3109), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U4963 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n4149), .B1(n3975), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3995) );
  NAND4_X1 U4964 ( .A1(n3998), .A2(n3997), .A3(n3996), .A4(n3995), .ZN(n4004)
         );
  AOI22_X1 U4965 ( .A1(n4142), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3422), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U4966 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n4123), .B1(n4151), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U4967 ( .A1(n3116), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4968 ( .A1(n4148), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3999) );
  NAND4_X1 U4969 ( .A1(n4002), .A2(n4001), .A3(n4000), .A4(n3999), .ZN(n4003)
         );
  NOR2_X1 U4970 ( .A1(n4004), .A2(n4003), .ZN(n4021) );
  AOI22_X1 U4971 ( .A1(n4142), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3422), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4972 ( .A1(n4122), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U4973 ( .A1(n3116), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U4974 ( .A1(n4123), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3279), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4005) );
  NAND4_X1 U4975 ( .A1(n4008), .A2(n4007), .A3(n4006), .A4(n4005), .ZN(n4014)
         );
  AOI22_X1 U4976 ( .A1(n3119), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4977 ( .A1(n4149), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4978 ( .A1(n4087), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U4979 ( .A1(n3104), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4009) );
  NAND4_X1 U4980 ( .A1(n4012), .A2(n4011), .A3(n4010), .A4(n4009), .ZN(n4013)
         );
  NOR2_X1 U4981 ( .A1(n4014), .A2(n4013), .ZN(n4022) );
  XOR2_X1 U4982 ( .A(n4021), .B(n4022), .Z(n4018) );
  INV_X1 U4983 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4016) );
  AOI21_X1 U4984 ( .B1(n6522), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n4141), 
        .ZN(n4015) );
  OAI21_X1 U4985 ( .B1(n4136), .B2(n4016), .A(n4015), .ZN(n4017) );
  AOI21_X1 U4986 ( .B1(n4138), .B2(n4018), .A(n4017), .ZN(n4019) );
  AOI21_X1 U4987 ( .B1(n4020), .B2(n4141), .A(n4019), .ZN(n5357) );
  XNOR2_X1 U4988 ( .A(n4038), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5600)
         );
  INV_X1 U4989 ( .A(n5600), .ZN(n4037) );
  NOR2_X1 U4990 ( .A1(n4022), .A2(n4021), .ZN(n4062) );
  AOI22_X1 U4991 ( .A1(n4087), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U4992 ( .A1(n4122), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U4993 ( .A1(n4149), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U4994 ( .A1(n3279), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4023) );
  NAND4_X1 U4995 ( .A1(n4026), .A2(n4025), .A3(n4024), .A4(n4023), .ZN(n4032)
         );
  AOI22_X1 U4996 ( .A1(n4142), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U4997 ( .A1(n3422), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U4998 ( .A1(n3889), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U4999 ( .A1(n3120), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4027) );
  NAND4_X1 U5000 ( .A1(n4030), .A2(n4029), .A3(n4028), .A4(n4027), .ZN(n4031)
         );
  OR2_X1 U5001 ( .A1(n4032), .A2(n4031), .ZN(n4061) );
  INV_X1 U5002 ( .A(n4138), .ZN(n4163) );
  AOI21_X1 U5003 ( .B1(n4062), .B2(n4061), .A(n4163), .ZN(n4033) );
  OAI21_X1 U5004 ( .B1(n4062), .B2(n4061), .A(n4033), .ZN(n4035) );
  AOI22_X1 U5005 ( .A1(n4175), .A2(EAX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n4174), .ZN(n4034) );
  NAND2_X1 U5006 ( .A1(n4035), .A2(n4034), .ZN(n4036) );
  AOI21_X1 U5007 ( .B1(n4037), .B2(n4141), .A(n4036), .ZN(n5255) );
  INV_X1 U5008 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5350) );
  NOR2_X1 U5009 ( .A1(n4038), .A2(n5350), .ZN(n4039) );
  NOR2_X1 U5010 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n4039), .ZN(n4040)
         );
  OR2_X1 U5011 ( .A1(n4058), .A2(n4040), .ZN(n5674) );
  AOI22_X1 U5012 ( .A1(n4087), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U5013 ( .A1(n4041), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U5014 ( .A1(n4149), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U5015 ( .A1(n3279), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4042) );
  NAND4_X1 U5016 ( .A1(n4045), .A2(n4044), .A3(n4043), .A4(n4042), .ZN(n4051)
         );
  AOI22_X1 U5017 ( .A1(n4142), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4049) );
  AOI22_X1 U5018 ( .A1(n3422), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4048) );
  AOI22_X1 U5019 ( .A1(n3889), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U5020 ( .A1(n3854), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4046) );
  NAND4_X1 U5021 ( .A1(n4049), .A2(n4048), .A3(n4047), .A4(n4046), .ZN(n4050)
         );
  OR2_X1 U5022 ( .A1(n4051), .A2(n4050), .ZN(n4060) );
  NAND2_X1 U5023 ( .A1(n4061), .A2(n4062), .ZN(n4052) );
  XNOR2_X1 U5024 ( .A(n4060), .B(n4052), .ZN(n4053) );
  AOI21_X1 U5025 ( .B1(n4138), .B2(n4053), .A(n4141), .ZN(n4055) );
  AOI22_X1 U5026 ( .A1(n4175), .A2(EAX_REG_25__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6522), .ZN(n4054) );
  NAND2_X1 U5027 ( .A1(n4055), .A2(n4054), .ZN(n4056) );
  OAI21_X1 U5028 ( .B1(n5674), .B2(n3750), .A(n4056), .ZN(n5246) );
  NOR2_X1 U5029 ( .A1(n5255), .A2(n5246), .ZN(n4057) );
  NAND2_X1 U5030 ( .A1(n5243), .A2(n4057), .ZN(n5233) );
  NOR2_X1 U5031 ( .A1(n4058), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4059)
         );
  OR2_X1 U5032 ( .A1(n4080), .A2(n4059), .ZN(n5591) );
  NAND3_X1 U5033 ( .A1(n4062), .A2(n4061), .A3(n4060), .ZN(n4082) );
  AOI22_X1 U5034 ( .A1(n3120), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4066) );
  AOI22_X1 U5035 ( .A1(n4041), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3422), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U5036 ( .A1(n3889), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U5037 ( .A1(n4142), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4063) );
  NAND4_X1 U5038 ( .A1(n4066), .A2(n4065), .A3(n4064), .A4(n4063), .ZN(n4072)
         );
  AOI22_X1 U5039 ( .A1(n4151), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4070) );
  AOI22_X1 U5040 ( .A1(n3109), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4148), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U5041 ( .A1(n3121), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4068) );
  AOI22_X1 U5042 ( .A1(n4149), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4067) );
  NAND4_X1 U5043 ( .A1(n4070), .A2(n4069), .A3(n4068), .A4(n4067), .ZN(n4071)
         );
  NOR2_X1 U5044 ( .A1(n4072), .A2(n4071), .ZN(n4081) );
  XNOR2_X1 U5045 ( .A(n4082), .B(n4081), .ZN(n4076) );
  INV_X1 U5046 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4073) );
  OAI21_X1 U5047 ( .B1(n4073), .B2(STATE2_REG_2__SCAN_IN), .A(n3750), .ZN(
        n4074) );
  AOI21_X1 U5048 ( .B1(n4175), .B2(EAX_REG_26__SCAN_IN), .A(n4074), .ZN(n4075)
         );
  OAI21_X1 U5049 ( .B1(n4076), .B2(n4163), .A(n4075), .ZN(n4077) );
  OAI21_X1 U5050 ( .B1(n5591), .B2(n3750), .A(n4077), .ZN(n5235) );
  INV_X1 U5051 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4194) );
  XNOR2_X1 U5052 ( .A(n4080), .B(n4194), .ZN(n5579) );
  NAND2_X1 U5053 ( .A1(n5579), .A2(n4141), .ZN(n4099) );
  OR2_X1 U5054 ( .A1(n4082), .A2(n4081), .ZN(n4102) );
  AOI22_X1 U5055 ( .A1(n4142), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3422), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4086) );
  AOI22_X1 U5056 ( .A1(n3116), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4085) );
  AOI22_X1 U5057 ( .A1(n3119), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U5058 ( .A1(n3279), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4083) );
  NAND4_X1 U5059 ( .A1(n4086), .A2(n4085), .A3(n4084), .A4(n4083), .ZN(n4093)
         );
  AOI22_X1 U5060 ( .A1(n4151), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4091) );
  AOI22_X1 U5061 ( .A1(n4122), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4090) );
  AOI22_X1 U5062 ( .A1(n4087), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U5063 ( .A1(n4149), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4088) );
  NAND4_X1 U5064 ( .A1(n4091), .A2(n4090), .A3(n4089), .A4(n4088), .ZN(n4092)
         );
  NOR2_X1 U5065 ( .A1(n4093), .A2(n4092), .ZN(n4103) );
  XOR2_X1 U5066 ( .A(n4102), .B(n4103), .Z(n4094) );
  NAND2_X1 U5067 ( .A1(n4094), .A2(n4138), .ZN(n4097) );
  OAI21_X1 U5068 ( .B1(n4194), .B2(STATE2_REG_2__SCAN_IN), .A(n3750), .ZN(
        n4095) );
  AOI21_X1 U5069 ( .B1(n4175), .B2(EAX_REG_27__SCAN_IN), .A(n4095), .ZN(n4096)
         );
  NAND2_X1 U5070 ( .A1(n4097), .A2(n4096), .ZN(n4098) );
  OR2_X1 U5071 ( .A1(n4100), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4101)
         );
  NAND2_X1 U5072 ( .A1(n4119), .A2(n4101), .ZN(n5570) );
  NOR2_X1 U5073 ( .A1(n4103), .A2(n4102), .ZN(n4121) );
  AOI22_X1 U5074 ( .A1(n4087), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U5075 ( .A1(n4122), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4106) );
  AOI22_X1 U5076 ( .A1(n4149), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4105) );
  AOI22_X1 U5077 ( .A1(n3279), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3975), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4104) );
  NAND4_X1 U5078 ( .A1(n4107), .A2(n4106), .A3(n4105), .A4(n4104), .ZN(n4113)
         );
  AOI22_X1 U5079 ( .A1(n4142), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4111) );
  AOI22_X1 U5080 ( .A1(n3422), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4110) );
  AOI22_X1 U5081 ( .A1(n3889), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U5082 ( .A1(n3120), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4108) );
  NAND4_X1 U5083 ( .A1(n4111), .A2(n4110), .A3(n4109), .A4(n4108), .ZN(n4112)
         );
  OR2_X1 U5084 ( .A1(n4113), .A2(n4112), .ZN(n4120) );
  XNOR2_X1 U5085 ( .A(n4121), .B(n4120), .ZN(n4117) );
  INV_X1 U5086 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4114) );
  OAI21_X1 U5087 ( .B1(n4114), .B2(STATE2_REG_2__SCAN_IN), .A(n3750), .ZN(
        n4115) );
  AOI21_X1 U5088 ( .B1(n4175), .B2(EAX_REG_28__SCAN_IN), .A(n4115), .ZN(n4116)
         );
  OAI21_X1 U5089 ( .B1(n4117), .B2(n4163), .A(n4116), .ZN(n4118) );
  OAI21_X1 U5090 ( .B1(n5570), .B2(n3750), .A(n4118), .ZN(n4209) );
  XNOR2_X1 U5091 ( .A(n4119), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4451)
         );
  NAND2_X1 U5092 ( .A1(n4121), .A2(n4120), .ZN(n4158) );
  AOI22_X1 U5093 ( .A1(n4142), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4127) );
  AOI22_X1 U5094 ( .A1(n4122), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3889), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4126) );
  AOI22_X1 U5095 ( .A1(n4149), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U5096 ( .A1(n3279), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4124) );
  NAND4_X1 U5097 ( .A1(n4127), .A2(n4126), .A3(n4125), .A4(n4124), .ZN(n4133)
         );
  AOI22_X1 U5098 ( .A1(n3119), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U5099 ( .A1(n3422), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4130) );
  AOI22_X1 U5100 ( .A1(n3116), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4129) );
  AOI22_X1 U5101 ( .A1(n3109), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4128) );
  NAND4_X1 U5102 ( .A1(n4131), .A2(n4130), .A3(n4129), .A4(n4128), .ZN(n4132)
         );
  NOR2_X1 U5103 ( .A1(n4133), .A2(n4132), .ZN(n4159) );
  XOR2_X1 U5104 ( .A(n4158), .B(n4159), .Z(n4139) );
  INV_X1 U5105 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4135) );
  AOI21_X1 U5106 ( .B1(n6522), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n4141), 
        .ZN(n4134) );
  OAI21_X1 U5107 ( .B1(n4136), .B2(n4135), .A(n4134), .ZN(n4137) );
  AOI21_X1 U5108 ( .B1(n4139), .B2(n4138), .A(n4137), .ZN(n4140) );
  AOI21_X1 U5109 ( .B1(n4451), .B2(n4141), .A(n4140), .ZN(n4215) );
  AND2_X2 U5110 ( .A1(n4208), .A2(n4215), .ZN(n4214) );
  AOI22_X1 U5111 ( .A1(n3854), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4147) );
  AOI22_X1 U5112 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n3889), .B1(n4087), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4146) );
  AOI22_X1 U5113 ( .A1(n3121), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4123), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4145) );
  AOI22_X1 U5114 ( .A1(n3103), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3980), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4144) );
  NAND4_X1 U5115 ( .A1(n4147), .A2(n4146), .A3(n4145), .A4(n4144), .ZN(n4157)
         );
  AOI22_X1 U5116 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n4041), .B1(n3106), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4155) );
  AOI22_X1 U5117 ( .A1(n3116), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U5118 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(n4149), .B1(n4148), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4153) );
  AOI22_X1 U5119 ( .A1(n4151), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4152) );
  NAND4_X1 U5120 ( .A1(n4155), .A2(n4154), .A3(n4153), .A4(n4152), .ZN(n4156)
         );
  NOR2_X1 U5121 ( .A1(n4157), .A2(n4156), .ZN(n4161) );
  NOR2_X1 U5122 ( .A1(n4159), .A2(n4158), .ZN(n4160) );
  XOR2_X1 U5123 ( .A(n4161), .B(n4160), .Z(n4164) );
  AOI22_X1 U5124 ( .A1(n4175), .A2(EAX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6522), .ZN(n4162) );
  OAI21_X1 U5125 ( .B1(n4164), .B2(n4163), .A(n4162), .ZN(n4165) );
  NAND2_X1 U5126 ( .A1(n4165), .A2(n3750), .ZN(n4166) );
  NAND2_X1 U5127 ( .A1(n4167), .A2(n4166), .ZN(n4168) );
  NAND2_X1 U5128 ( .A1(n4214), .A2(n4168), .ZN(n4177) );
  NAND3_X1 U5129 ( .A1(n6525), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6444) );
  INV_X1 U5130 ( .A(n6444), .ZN(n4170) );
  OAI211_X1 U5131 ( .C1(n5404), .C2(n5773), .A(n4173), .B(n4172), .ZN(U2956)
         );
  AOI22_X1 U5132 ( .A1(n4175), .A2(EAX_REG_31__SCAN_IN), .B1(n4174), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4176) );
  XNOR2_X2 U5133 ( .A(n4177), .B(n4176), .ZN(n5320) );
  AND2_X1 U5134 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4468) );
  AOI21_X1 U5135 ( .B1(n4380), .B2(n4468), .A(n4179), .ZN(n4180) );
  NAND2_X1 U5136 ( .A1(n4459), .A2(n6040), .ZN(n4187) );
  INV_X1 U5137 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5210) );
  NAND2_X1 U5138 ( .A1(n4234), .A2(n6022), .ZN(n4184) );
  NAND2_X1 U5139 ( .A1(n4228), .A2(REIP_REG_31__SCAN_IN), .ZN(n4469) );
  OAI211_X1 U5140 ( .C1(n5210), .C2(n5393), .A(n4184), .B(n4469), .ZN(n4185)
         );
  INV_X1 U5141 ( .A(n4185), .ZN(n4186) );
  NAND2_X1 U5142 ( .A1(n5432), .A2(n5337), .ZN(n4201) );
  NAND2_X1 U5143 ( .A1(n4188), .A2(n4201), .ZN(n4189) );
  XNOR2_X1 U5144 ( .A(n4189), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5422)
         );
  INV_X1 U5145 ( .A(n4190), .ZN(n4191) );
  NOR2_X1 U5146 ( .A1(n5584), .A2(n6026), .ZN(n4198) );
  NAND2_X1 U5147 ( .A1(n4228), .A2(REIP_REG_27__SCAN_IN), .ZN(n5415) );
  OAI21_X1 U5148 ( .B1(n5393), .B2(n4194), .A(n5415), .ZN(n4195) );
  OAI21_X1 U5149 ( .B1(n5422), .B2(n5773), .A(n4199), .ZN(U2959) );
  INV_X1 U5150 ( .A(n5405), .ZN(n4200) );
  INV_X1 U5151 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6630) );
  NOR2_X1 U5152 ( .A1(n6630), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4202)
         );
  MUX2_X1 U5153 ( .A(n5406), .B(n4202), .S(n4201), .Z(n4203) );
  INV_X1 U5154 ( .A(n4203), .ZN(n4204) );
  NAND2_X1 U5155 ( .A1(n4205), .A2(n4204), .ZN(n4207) );
  INV_X1 U5156 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5419) );
  NAND2_X1 U5157 ( .A1(n5653), .A2(n5700), .ZN(n4213) );
  INV_X1 U5158 ( .A(REIP_REG_28__SCAN_IN), .ZN(n4210) );
  NOR2_X1 U5159 ( .A1(n5727), .A2(n4210), .ZN(n5407) );
  NOR2_X1 U5160 ( .A1(n5570), .A2(n6045), .ZN(n4211) );
  AOI211_X1 U5161 ( .C1(PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n6036), .A(n5407), 
        .B(n4211), .ZN(n4212) );
  INV_X1 U5162 ( .A(n4214), .ZN(n4218) );
  OR2_X1 U5163 ( .A1(n4216), .A2(n4215), .ZN(n4217) );
  NAND2_X1 U5164 ( .A1(n4218), .A2(n4217), .ZN(n5220) );
  NAND4_X1 U5165 ( .A1(n4224), .A2(n4223), .A3(n4222), .A4(n4221), .ZN(n4225)
         );
  NAND2_X1 U5166 ( .A1(n4226), .A2(n4225), .ZN(n5194) );
  INV_X1 U5167 ( .A(n5194), .ZN(n4227) );
  NAND2_X1 U5168 ( .A1(n5195), .A2(n4227), .ZN(n5201) );
  NAND2_X1 U5169 ( .A1(n6426), .A2(n6522), .ZN(n6521) );
  NOR3_X1 U5170 ( .A1(n6817), .A2(n6525), .A3(n6521), .ZN(n6427) );
  NOR3_X1 U5171 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n6438), .A3(n6426), .ZN(
        n4229) );
  OR2_X1 U5172 ( .A1(n4229), .A2(n4228), .ZN(n4230) );
  NOR2_X1 U5173 ( .A1(n6427), .A2(n4230), .ZN(n4231) );
  NAND2_X1 U5174 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n4241), .ZN(n4233) );
  INV_X1 U5175 ( .A(n4233), .ZN(n4232) );
  INV_X1 U5176 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6486) );
  NAND2_X1 U5177 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n4235) );
  INV_X1 U5178 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6726) );
  INV_X1 U5179 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6651) );
  NOR2_X1 U5180 ( .A1(n6726), .A2(n6651), .ZN(n6832) );
  NAND2_X1 U5181 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .ZN(
        n4254) );
  NAND3_X1 U5182 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .ZN(n4253) );
  INV_X1 U5183 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6467) );
  INV_X1 U5184 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6765) );
  NAND3_X1 U5185 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n4972) );
  NOR4_X1 U5186 ( .A1(n4971), .A2(n6467), .A3(n6765), .A4(n4972), .ZN(n5882)
         );
  NAND4_X1 U5187 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_6__SCAN_IN), .A4(n5882), .ZN(n5858) );
  NOR2_X1 U5188 ( .A1(n4253), .A2(n5858), .ZN(n5852) );
  NAND2_X1 U5189 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5852), .ZN(n5832) );
  NOR2_X1 U5190 ( .A1(n4254), .A2(n5832), .ZN(n5810) );
  NAND3_X1 U5191 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6832), .A3(n5810), .ZN(
        n5643) );
  NOR3_X1 U5192 ( .A1(n6486), .A2(n4235), .A3(n5643), .ZN(n5615) );
  NAND4_X1 U5193 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5615), .ZN(n5596) );
  NAND3_X1 U5194 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4255) );
  NAND2_X1 U5195 ( .A1(n6523), .A2(n4918), .ZN(n4240) );
  INV_X1 U5196 ( .A(STATE_REG_0__SCAN_IN), .ZN(n4236) );
  NAND2_X1 U5197 ( .A1(n4237), .A2(n4236), .ZN(n6452) );
  AOI21_X1 U5198 ( .B1(n3374), .B2(n6452), .A(READY_N), .ZN(n4238) );
  NAND2_X1 U5199 ( .A1(n3365), .A2(n4238), .ZN(n4239) );
  NAND2_X1 U5200 ( .A1(n4241), .A2(n5208), .ZN(n5859) );
  OAI21_X1 U5201 ( .B1(n5596), .B2(n4255), .A(n5859), .ZN(n5586) );
  INV_X1 U5202 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6655) );
  NOR2_X1 U5203 ( .A1(n4210), .A2(n6655), .ZN(n4242) );
  OR2_X1 U5204 ( .A1(n5208), .A2(n4242), .ZN(n4243) );
  AND2_X1 U5205 ( .A1(n5586), .A2(n4243), .ZN(n5571) );
  INV_X1 U5206 ( .A(n5571), .ZN(n5206) );
  AOI22_X1 U5207 ( .A1(n4451), .A2(n5892), .B1(REIP_REG_29__SCAN_IN), .B2(
        n5206), .ZN(n4249) );
  NOR2_X1 U5208 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4358) );
  NAND2_X1 U5209 ( .A1(n4805), .A2(n4358), .ZN(n6423) );
  INV_X1 U5210 ( .A(n6423), .ZN(n4244) );
  OR2_X1 U5211 ( .A1(n3110), .A2(n4244), .ZN(n5212) );
  NOR2_X1 U5212 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4358), .ZN(n4245) );
  NAND2_X1 U5213 ( .A1(n3365), .A2(n4245), .ZN(n4246) );
  NAND2_X1 U5214 ( .A1(n5212), .A2(n4246), .ZN(n4247) );
  NOR2_X2 U5215 ( .A1(n4971), .A2(n6817), .ZN(n5893) );
  AOI22_X1 U5216 ( .A1(EBX_REG_29__SCAN_IN), .A2(n5908), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n5893), .ZN(n4248) );
  OAI21_X1 U5217 ( .B1(n5220), .B2(n5902), .A(n4250), .ZN(n4251) );
  INV_X1 U5218 ( .A(n4251), .ZN(n4363) );
  NAND2_X1 U5219 ( .A1(REIP_REG_3__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .ZN(
        n4252) );
  NOR2_X2 U5220 ( .A1(n5009), .A2(n4252), .ZN(n4946) );
  NOR2_X2 U5221 ( .A1(n5841), .A2(n4254), .ZN(n5820) );
  INV_X1 U5222 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6480) );
  NOR2_X2 U5223 ( .A1(n5597), .A2(n4255), .ZN(n5580) );
  NAND3_X1 U5224 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .A3(
        n5580), .ZN(n5214) );
  INV_X1 U5225 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4921) );
  INV_X1 U5226 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4258) );
  OR2_X1 U5227 ( .A1(n4257), .A2(n4258), .ZN(n4260) );
  NAND2_X1 U5228 ( .A1(n5282), .A2(n4258), .ZN(n4259) );
  NAND2_X1 U5229 ( .A1(n4260), .A2(n4259), .ZN(n4527) );
  INV_X1 U5230 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4262) );
  NAND2_X1 U5231 ( .A1(n4341), .A2(n4262), .ZN(n4265) );
  NAND2_X1 U5232 ( .A1(n4557), .A2(n4262), .ZN(n4263) );
  OAI211_X1 U5233 ( .C1(n5282), .C2(n6107), .A(n4263), .B(n4257), .ZN(n4264)
         );
  AND2_X1 U5234 ( .A1(n4265), .A2(n4264), .ZN(n4747) );
  INV_X1 U5235 ( .A(n4341), .ZN(n4293) );
  MUX2_X1 U5236 ( .A(n4293), .B(n4461), .S(EBX_REG_4__SCAN_IN), .Z(n4267) );
  OR2_X1 U5237 ( .A1(n4529), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4266)
         );
  NAND2_X1 U5238 ( .A1(n4267), .A2(n4266), .ZN(n4657) );
  INV_X1 U5239 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4974) );
  NAND2_X1 U5240 ( .A1(n4352), .A2(n4974), .ZN(n4270) );
  OAI21_X1 U5241 ( .B1(n5282), .B2(n6711), .A(n4346), .ZN(n4268) );
  OAI21_X1 U5242 ( .B1(EBX_REG_3__SCAN_IN), .B2(n4548), .A(n4268), .ZN(n4269)
         );
  AND2_X1 U5243 ( .A1(n4270), .A2(n4269), .ZN(n4656) );
  NOR2_X1 U5244 ( .A1(n4657), .A2(n4656), .ZN(n4271) );
  INV_X1 U5245 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4744) );
  NAND2_X1 U5246 ( .A1(n4352), .A2(n4744), .ZN(n4274) );
  NAND2_X1 U5247 ( .A1(n4346), .A2(n6580), .ZN(n4272) );
  OAI211_X1 U5248 ( .C1(n4548), .C2(EBX_REG_5__SCAN_IN), .A(n4272), .B(n4461), 
        .ZN(n4273) );
  AND2_X1 U5249 ( .A1(n4274), .A2(n4273), .ZN(n4680) );
  INV_X1 U5250 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U5251 ( .A1(n4341), .A2(n5896), .ZN(n4278) );
  NAND2_X1 U5252 ( .A1(n4557), .A2(n5896), .ZN(n4276) );
  OAI211_X1 U5253 ( .C1(n5282), .C2(n6654), .A(n4276), .B(n4346), .ZN(n4277)
         );
  NAND2_X1 U5254 ( .A1(n4278), .A2(n4277), .ZN(n4752) );
  MUX2_X1 U5255 ( .A(n4341), .B(n5282), .S(EBX_REG_8__SCAN_IN), .Z(n4280) );
  NOR2_X1 U5256 ( .A1(n4529), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4279)
         );
  NOR2_X1 U5257 ( .A1(n4280), .A2(n4279), .ZN(n4760) );
  INV_X1 U5258 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5926) );
  NAND2_X1 U5259 ( .A1(n4352), .A2(n5926), .ZN(n4283) );
  NAND2_X1 U5260 ( .A1(n4257), .A2(n6072), .ZN(n4281) );
  OAI211_X1 U5261 ( .C1(n4548), .C2(EBX_REG_7__SCAN_IN), .A(n4281), .B(n4461), 
        .ZN(n4282) );
  NAND2_X1 U5262 ( .A1(n4283), .A2(n4282), .ZN(n5879) );
  INV_X1 U5263 ( .A(n4529), .ZN(n4284) );
  NAND2_X1 U5264 ( .A1(n3617), .A2(n4284), .ZN(n4286) );
  MUX2_X1 U5265 ( .A(n4293), .B(n4461), .S(EBX_REG_10__SCAN_IN), .Z(n4285) );
  NAND2_X1 U5266 ( .A1(n4286), .A2(n4285), .ZN(n5038) );
  INV_X1 U5267 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U5268 ( .A1(n4352), .A2(n5867), .ZN(n4289) );
  NAND2_X1 U5269 ( .A1(n4346), .A2(n5981), .ZN(n4287) );
  OAI211_X1 U5270 ( .C1(n4548), .C2(EBX_REG_9__SCAN_IN), .A(n4287), .B(n4461), 
        .ZN(n4288) );
  NOR2_X1 U5271 ( .A1(n5038), .A2(n5034), .ZN(n4290) );
  NAND2_X1 U5272 ( .A1(n4346), .A2(n6052), .ZN(n4291) );
  OAI211_X1 U5273 ( .C1(n4548), .C2(EBX_REG_11__SCAN_IN), .A(n4291), .B(n4461), 
        .ZN(n4292) );
  OAI21_X1 U5274 ( .B1(n4349), .B2(EBX_REG_11__SCAN_IN), .A(n4292), .ZN(n4932)
         );
  NAND2_X1 U5275 ( .A1(n4931), .A2(n4932), .ZN(n5097) );
  MUX2_X1 U5276 ( .A(n4293), .B(n4461), .S(EBX_REG_12__SCAN_IN), .Z(n4294) );
  NAND2_X1 U5277 ( .A1(n3216), .A2(n4294), .ZN(n5096) );
  INV_X1 U5278 ( .A(EBX_REG_13__SCAN_IN), .ZN(n4295) );
  NAND2_X1 U5279 ( .A1(n4352), .A2(n4295), .ZN(n4298) );
  OAI21_X1 U5280 ( .B1(n5282), .B2(n5507), .A(n4257), .ZN(n4296) );
  OAI21_X1 U5281 ( .B1(EBX_REG_13__SCAN_IN), .B2(n4548), .A(n4296), .ZN(n4297)
         );
  AND2_X1 U5282 ( .A1(n4298), .A2(n4297), .ZN(n5087) );
  INV_X1 U5283 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6658) );
  NAND2_X1 U5284 ( .A1(n4341), .A2(n6658), .ZN(n4301) );
  INV_X1 U5285 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U5286 ( .A1(n4557), .A2(n6658), .ZN(n4299) );
  OAI211_X1 U5287 ( .C1(n5282), .C2(n5753), .A(n4299), .B(n4346), .ZN(n4300)
         );
  NAND2_X1 U5288 ( .A1(n4301), .A2(n4300), .ZN(n5115) );
  NAND2_X1 U5289 ( .A1(n4346), .A2(n6564), .ZN(n4302) );
  OAI211_X1 U5290 ( .C1(n4548), .C2(EBX_REG_15__SCAN_IN), .A(n4302), .B(n4461), 
        .ZN(n4303) );
  OAI21_X1 U5291 ( .B1(n4349), .B2(EBX_REG_15__SCAN_IN), .A(n4303), .ZN(n5309)
         );
  INV_X1 U5292 ( .A(EBX_REG_16__SCAN_IN), .ZN(n4304) );
  NAND2_X1 U5293 ( .A1(n4341), .A2(n4304), .ZN(n4307) );
  NAND2_X1 U5294 ( .A1(n4557), .A2(n4304), .ZN(n4305) );
  OAI211_X1 U5295 ( .C1(n5282), .C2(n6579), .A(n4305), .B(n4346), .ZN(n4306)
         );
  NAND2_X1 U5296 ( .A1(n4307), .A2(n4306), .ZN(n5305) );
  INV_X1 U5297 ( .A(EBX_REG_17__SCAN_IN), .ZN(n4308) );
  NAND2_X1 U5298 ( .A1(n4352), .A2(n4308), .ZN(n4311) );
  OAI21_X1 U5299 ( .B1(n5282), .B2(n6717), .A(n4257), .ZN(n4309) );
  OAI21_X1 U5300 ( .B1(EBX_REG_17__SCAN_IN), .B2(n4548), .A(n4309), .ZN(n4310)
         );
  INV_X1 U5301 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5287) );
  NAND2_X1 U5302 ( .A1(n4341), .A2(n5287), .ZN(n4314) );
  INV_X1 U5303 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5722) );
  NAND2_X1 U5304 ( .A1(n4557), .A2(n5287), .ZN(n4312) );
  OAI211_X1 U5305 ( .C1(n5282), .C2(n5722), .A(n4312), .B(n4346), .ZN(n4313)
         );
  OR2_X1 U5306 ( .A1(n4529), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4317)
         );
  INV_X1 U5307 ( .A(EBX_REG_20__SCAN_IN), .ZN(n4315) );
  NAND2_X1 U5308 ( .A1(n4557), .A2(n4315), .ZN(n4316) );
  AND2_X1 U5309 ( .A1(n4317), .A2(n4316), .ZN(n5272) );
  OR2_X1 U5310 ( .A1(n4529), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4318)
         );
  INV_X1 U5311 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U5312 ( .A1(n4557), .A2(n5293), .ZN(n5281) );
  NAND2_X1 U5313 ( .A1(n4318), .A2(n5281), .ZN(n5270) );
  NAND2_X1 U5314 ( .A1(n5282), .A2(EBX_REG_20__SCAN_IN), .ZN(n4320) );
  NAND2_X1 U5315 ( .A1(n5270), .A2(n4461), .ZN(n4319) );
  OAI211_X1 U5316 ( .C1(n5272), .C2(n5270), .A(n4320), .B(n4319), .ZN(n4321)
         );
  INV_X1 U5317 ( .A(n4321), .ZN(n4322) );
  INV_X1 U5318 ( .A(EBX_REG_21__SCAN_IN), .ZN(n6566) );
  NAND2_X1 U5319 ( .A1(n4341), .A2(n6566), .ZN(n4326) );
  INV_X1 U5320 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4324) );
  NAND2_X1 U5321 ( .A1(n4557), .A2(n6566), .ZN(n4323) );
  OAI211_X1 U5322 ( .C1(n5282), .C2(n4324), .A(n4323), .B(n4346), .ZN(n4325)
         );
  NAND2_X1 U5323 ( .A1(n4326), .A2(n4325), .ZN(n5469) );
  INV_X1 U5324 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5267) );
  NAND2_X1 U5325 ( .A1(n4352), .A2(n5267), .ZN(n4329) );
  INV_X1 U5326 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5364) );
  NAND2_X1 U5327 ( .A1(n4257), .A2(n5364), .ZN(n4327) );
  OAI211_X1 U5328 ( .C1(n4548), .C2(EBX_REG_22__SCAN_IN), .A(n4327), .B(n4461), 
        .ZN(n4328) );
  AND2_X1 U5329 ( .A1(n4329), .A2(n4328), .ZN(n5265) );
  INV_X1 U5330 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5649) );
  NAND2_X1 U5331 ( .A1(n4341), .A2(n5649), .ZN(n4332) );
  NAND2_X1 U5332 ( .A1(n4557), .A2(n5649), .ZN(n4330) );
  OAI211_X1 U5333 ( .C1(n5282), .C2(n6702), .A(n4330), .B(n4346), .ZN(n4331)
         );
  AND2_X1 U5334 ( .A1(n4332), .A2(n4331), .ZN(n5447) );
  NAND2_X1 U5335 ( .A1(n4346), .A2(n5347), .ZN(n4333) );
  OAI211_X1 U5336 ( .C1(EBX_REG_24__SCAN_IN), .C2(n4548), .A(n4333), .B(n4461), 
        .ZN(n4334) );
  OAI21_X1 U5337 ( .B1(n4349), .B2(EBX_REG_24__SCAN_IN), .A(n4334), .ZN(n5256)
         );
  INV_X1 U5338 ( .A(EBX_REG_25__SCAN_IN), .ZN(n6607) );
  NAND2_X1 U5339 ( .A1(n4352), .A2(n6607), .ZN(n4337) );
  NAND2_X1 U5340 ( .A1(n4257), .A2(n5427), .ZN(n4335) );
  OAI211_X1 U5341 ( .C1(n4548), .C2(EBX_REG_25__SCAN_IN), .A(n4335), .B(n4461), 
        .ZN(n4336) );
  AND2_X1 U5342 ( .A1(n4337), .A2(n4336), .ZN(n5249) );
  INV_X1 U5343 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5240) );
  NAND2_X1 U5344 ( .A1(n4352), .A2(n5240), .ZN(n4340) );
  NAND2_X1 U5345 ( .A1(n4346), .A2(n5426), .ZN(n4338) );
  OAI211_X1 U5346 ( .C1(n4548), .C2(EBX_REG_26__SCAN_IN), .A(n4338), .B(n4461), 
        .ZN(n4339) );
  AND2_X1 U5347 ( .A1(n4340), .A2(n4339), .ZN(n5237) );
  INV_X1 U5348 ( .A(EBX_REG_27__SCAN_IN), .ZN(n4342) );
  NAND2_X1 U5349 ( .A1(n4341), .A2(n4342), .ZN(n4345) );
  NAND2_X1 U5350 ( .A1(n4557), .A2(n4342), .ZN(n4343) );
  OAI211_X1 U5351 ( .C1(n5282), .C2(n5419), .A(n4343), .B(n4346), .ZN(n4344)
         );
  AND2_X1 U5352 ( .A1(n4345), .A2(n4344), .ZN(n5228) );
  NAND2_X1 U5353 ( .A1(n4346), .A2(n6630), .ZN(n4347) );
  OAI211_X1 U5354 ( .C1(n4548), .C2(EBX_REG_28__SCAN_IN), .A(n4347), .B(n4461), 
        .ZN(n4348) );
  OAI21_X1 U5355 ( .B1(n4349), .B2(EBX_REG_28__SCAN_IN), .A(n4348), .ZN(n5224)
         );
  NAND2_X1 U5356 ( .A1(n5229), .A2(n5224), .ZN(n4354) );
  OR2_X1 U5357 ( .A1(n4529), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4351)
         );
  INV_X1 U5358 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5223) );
  NAND2_X1 U5359 ( .A1(n4557), .A2(n5223), .ZN(n4350) );
  NAND2_X1 U5360 ( .A1(n4351), .A2(n4350), .ZN(n4356) );
  NAND2_X1 U5361 ( .A1(n4352), .A2(n5223), .ZN(n4355) );
  NOR2_X1 U5362 ( .A1(n4353), .A2(n3128), .ZN(n4462) );
  OAI211_X1 U5363 ( .C1(n5282), .C2(n4356), .A(n4354), .B(n4355), .ZN(n4357)
         );
  NAND2_X1 U5364 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4918), .ZN(n5211) );
  OAI21_X1 U5365 ( .B1(n5214), .B2(REIP_REG_29__SCAN_IN), .A(n4360), .ZN(n4361) );
  INV_X1 U5366 ( .A(n4361), .ZN(n4362) );
  NAND2_X1 U5367 ( .A1(n4363), .A2(n4362), .ZN(U2798) );
  AND2_X1 U5368 ( .A1(n4398), .A2(n3108), .ZN(n4579) );
  NAND2_X1 U5369 ( .A1(n5204), .A2(n4579), .ZN(n4366) );
  AND2_X1 U5370 ( .A1(n5195), .A2(n3374), .ZN(n4571) );
  NOR2_X1 U5371 ( .A1(READY_N), .A2(n5194), .ZN(n4392) );
  NAND2_X1 U5372 ( .A1(n4571), .A2(n4392), .ZN(n4365) );
  NAND2_X1 U5373 ( .A1(n4366), .A2(n4365), .ZN(n4485) );
  NOR2_X1 U5374 ( .A1(n4549), .A2(n3107), .ZN(n4369) );
  INV_X1 U5375 ( .A(READY_N), .ZN(n4388) );
  NAND2_X1 U5376 ( .A1(n3332), .A2(n4388), .ZN(n4370) );
  NAND2_X1 U5377 ( .A1(n3339), .A2(n3349), .ZN(n4372) );
  NAND2_X2 U5378 ( .A1(n5317), .A2(n4372), .ZN(n5652) );
  AND2_X1 U5379 ( .A1(n3366), .A2(n3349), .ZN(n4374) );
  AOI22_X1 U5380 ( .A1(n5932), .A2(DATAI_14_), .B1(n5931), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n4375) );
  INV_X1 U5381 ( .A(n4375), .ZN(n4378) );
  AND2_X1 U5382 ( .A1(n5317), .A2(n3368), .ZN(n5928) );
  INV_X1 U5383 ( .A(n5928), .ZN(n5669) );
  INV_X1 U5384 ( .A(DATAI_30_), .ZN(n4376) );
  NOR2_X1 U5385 ( .A1(n5669), .A2(n4376), .ZN(n4377) );
  OAI21_X1 U5386 ( .B1(n4364), .B2(n5652), .A(n4379), .ZN(U2861) );
  INV_X1 U5387 ( .A(n4380), .ZN(n4385) );
  NAND3_X1 U5388 ( .A1(n4385), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n4381), .ZN(n4384) );
  INV_X1 U5389 ( .A(n4382), .ZN(n4383) );
  OAI211_X1 U5390 ( .C1(n4385), .C2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n4384), .B(n4383), .ZN(n4449) );
  AOI21_X1 U5391 ( .B1(n4386), .B2(n4388), .A(n4387), .ZN(n4389) );
  NAND2_X1 U5392 ( .A1(n5204), .A2(n4389), .ZN(n4391) );
  OR2_X1 U5393 ( .A1(n3110), .A2(n4805), .ZN(n4390) );
  AOI21_X1 U5394 ( .B1(n4391), .B2(n4390), .A(n3368), .ZN(n4403) );
  NOR2_X1 U5395 ( .A1(n4503), .A2(n3374), .ZN(n4424) );
  AOI21_X1 U5396 ( .B1(n5204), .B2(n4417), .A(n4424), .ZN(n4402) );
  NAND2_X1 U5397 ( .A1(n3332), .A2(n6452), .ZN(n4393) );
  NAND3_X1 U5398 ( .A1(n4393), .A2(n4392), .A3(n3294), .ZN(n4401) );
  INV_X1 U5399 ( .A(n4394), .ZN(n4395) );
  NAND2_X1 U5400 ( .A1(n4395), .A2(n3365), .ZN(n4397) );
  INV_X1 U5401 ( .A(n3339), .ZN(n4396) );
  MUX2_X1 U5402 ( .A(n4397), .B(n3110), .S(n4396), .Z(n4419) );
  NAND2_X1 U5403 ( .A1(n4398), .A2(n4419), .ZN(n4400) );
  INV_X1 U5404 ( .A(n5195), .ZN(n4399) );
  NAND2_X1 U5405 ( .A1(n4400), .A2(n4399), .ZN(n4490) );
  OAI211_X1 U5406 ( .C1(n4403), .C2(n4402), .A(n4401), .B(n4490), .ZN(n4404)
         );
  OR2_X1 U5407 ( .A1(n4579), .A2(n4405), .ZN(n5193) );
  NAND2_X1 U5408 ( .A1(n4386), .A2(n4557), .ZN(n4407) );
  OR2_X1 U5409 ( .A1(n4571), .A2(n4408), .ZN(n4409) );
  NOR2_X1 U5410 ( .A1(n5193), .A2(n4409), .ZN(n4410) );
  NAND2_X1 U5411 ( .A1(n4449), .A2(n6090), .ZN(n4448) );
  NAND2_X1 U5412 ( .A1(n4386), .A2(n6524), .ZN(n6424) );
  OAI21_X1 U5413 ( .B1(n4406), .B2(n3338), .A(n6424), .ZN(n4411) );
  INV_X1 U5414 ( .A(n4411), .ZN(n4412) );
  NAND2_X1 U5415 ( .A1(n5195), .A2(n3332), .ZN(n4599) );
  NAND2_X1 U5416 ( .A1(n3345), .A2(n5282), .ZN(n4416) );
  NOR2_X1 U5417 ( .A1(n4413), .A2(n3294), .ZN(n4488) );
  OAI21_X1 U5418 ( .B1(n4488), .B2(n4529), .A(n4414), .ZN(n4415) );
  OAI211_X1 U5419 ( .C1(n3368), .C2(n4417), .A(n4416), .B(n4415), .ZN(n4418)
         );
  INV_X1 U5420 ( .A(n4418), .ZN(n4420) );
  NAND3_X1 U5421 ( .A1(n3217), .A2(n4420), .A3(n4419), .ZN(n4497) );
  INV_X1 U5422 ( .A(n4422), .ZN(n4597) );
  OAI21_X1 U5423 ( .B1(n4421), .B2(n3365), .A(n4597), .ZN(n4423) );
  NOR2_X1 U5424 ( .A1(n4497), .A2(n4423), .ZN(n4425) );
  OR2_X1 U5425 ( .A1(n4426), .A2(n4425), .ZN(n4436) );
  NAND2_X1 U5426 ( .A1(n4425), .A2(n4424), .ZN(n5196) );
  NAND2_X1 U5427 ( .A1(n5727), .A2(n4426), .ZN(n4525) );
  NAND2_X1 U5428 ( .A1(n6095), .A2(n4436), .ZN(n5505) );
  NAND2_X1 U5429 ( .A1(n4435), .A2(n5505), .ZN(n4530) );
  NAND2_X1 U5430 ( .A1(n4525), .A2(n4530), .ZN(n4675) );
  INV_X1 U5431 ( .A(n4675), .ZN(n4427) );
  AND2_X1 U5432 ( .A1(n6095), .A2(n4427), .ZN(n5480) );
  NAND2_X1 U5433 ( .A1(n5104), .A2(n5480), .ZN(n4429) );
  NAND3_X1 U5434 ( .A1(n5487), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4428) );
  NAND2_X1 U5435 ( .A1(n4429), .A2(n4428), .ZN(n4433) );
  NAND2_X1 U5436 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5028) );
  NAND2_X1 U5437 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6819) );
  NAND2_X1 U5438 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6081) );
  NOR2_X1 U5439 ( .A1(n6819), .A2(n6081), .ZN(n5027) );
  NOR2_X1 U5440 ( .A1(n6072), .A2(n6767), .ZN(n6061) );
  NAND4_X1 U5441 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n5027), .A4(n6061), .ZN(n4431)
         );
  NOR2_X1 U5442 ( .A1(n5028), .A2(n4431), .ZN(n5103) );
  NAND2_X1 U5443 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6824) );
  INV_X1 U5444 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U5445 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5506) );
  NOR2_X1 U5446 ( .A1(n5507), .A2(n5506), .ZN(n5754) );
  NAND2_X1 U5447 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5754), .ZN(n5740) );
  NOR2_X1 U5448 ( .A1(n6824), .A2(n5740), .ZN(n5478) );
  AND2_X1 U5449 ( .A1(n5103), .A2(n5478), .ZN(n4430) );
  OR2_X1 U5450 ( .A1(n5104), .A2(n4430), .ZN(n5479) );
  NAND2_X1 U5451 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U5452 ( .A1(n6107), .A2(n6097), .ZN(n6096) );
  INV_X1 U5453 ( .A(n6096), .ZN(n4678) );
  AND2_X1 U5454 ( .A1(n5478), .A2(n5102), .ZN(n5481) );
  OR2_X1 U5455 ( .A1(n5480), .A2(n5481), .ZN(n4432) );
  NAND2_X1 U5456 ( .A1(n5104), .A2(n6095), .ZN(n5493) );
  INV_X1 U5457 ( .A(n5463), .ZN(n5454) );
  NAND2_X1 U5458 ( .A1(n5493), .A2(n5454), .ZN(n4434) );
  NAND2_X1 U5459 ( .A1(n5460), .A2(n4434), .ZN(n5457) );
  INV_X1 U5460 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4435) );
  AOI21_X1 U5461 ( .B1(n5029), .B2(n6095), .A(n4437), .ZN(n4438) );
  NAND2_X1 U5462 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5424) );
  AND2_X1 U5463 ( .A1(n5493), .A2(n5424), .ZN(n4439) );
  NOR2_X1 U5464 ( .A1(n5442), .A2(n4439), .ZN(n5417) );
  NAND2_X1 U5465 ( .A1(n5493), .A2(n5405), .ZN(n4440) );
  AND2_X1 U5466 ( .A1(n5417), .A2(n4440), .ZN(n4467) );
  INV_X1 U5467 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4441) );
  NAND2_X1 U5468 ( .A1(n4228), .A2(REIP_REG_29__SCAN_IN), .ZN(n4453) );
  OAI21_X1 U5469 ( .B1(n4467), .B2(n4441), .A(n4453), .ZN(n4442) );
  AOI21_X1 U5470 ( .B1(n5221), .B2(n6099), .A(n4442), .ZN(n4446) );
  INV_X1 U5471 ( .A(n5102), .ZN(n5748) );
  NAND2_X1 U5472 ( .A1(n5103), .A2(n6106), .ZN(n5484) );
  NAND2_X1 U5473 ( .A1(n5748), .A2(n5484), .ZN(n5752) );
  NAND3_X1 U5474 ( .A1(n5478), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5752), .ZN(n5726) );
  INV_X1 U5475 ( .A(n4443), .ZN(n4444) );
  NAND2_X1 U5476 ( .A1(n5485), .A2(n4444), .ZN(n5436) );
  NOR2_X1 U5477 ( .A1(n5414), .A2(n5405), .ZN(n5401) );
  INV_X1 U5478 ( .A(n5401), .ZN(n4445) );
  NAND2_X1 U5479 ( .A1(n4448), .A2(n4447), .ZN(U2989) );
  NAND2_X1 U5480 ( .A1(n4449), .A2(n6040), .ZN(n4458) );
  NAND2_X1 U5481 ( .A1(n4450), .A2(n5700), .ZN(n4457) );
  INV_X1 U5482 ( .A(n4451), .ZN(n4454) );
  NAND2_X1 U5483 ( .A1(n6036), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4452)
         );
  OAI211_X1 U5484 ( .C1(n4454), .C2(n6045), .A(n4453), .B(n4452), .ZN(n4455)
         );
  INV_X1 U5485 ( .A(n4455), .ZN(n4456) );
  NAND3_X1 U5486 ( .A1(n4458), .A2(n4457), .A3(n4456), .ZN(U2957) );
  NAND2_X1 U5487 ( .A1(n4459), .A2(n6090), .ZN(n4475) );
  AND2_X1 U5488 ( .A1(n4548), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4460)
         );
  AOI21_X1 U5489 ( .B1(n4529), .B2(EBX_REG_30__SCAN_IN), .A(n4460), .ZN(n5179)
         );
  INV_X1 U5490 ( .A(n5179), .ZN(n5181) );
  NAND2_X1 U5491 ( .A1(n5182), .A2(n4461), .ZN(n5184) );
  OAI22_X1 U5492 ( .A1(n4529), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4548), .ZN(n4463) );
  XNOR2_X1 U5493 ( .A(n4464), .B(n4463), .ZN(n5219) );
  INV_X1 U5494 ( .A(n5219), .ZN(n4473) );
  INV_X1 U5495 ( .A(n4468), .ZN(n4465) );
  NAND2_X1 U5496 ( .A1(n5493), .A2(n4465), .ZN(n4466) );
  AND2_X1 U5497 ( .A1(n4467), .A2(n4466), .ZN(n5398) );
  INV_X1 U5498 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4471) );
  NAND3_X1 U5499 ( .A1(n5401), .A2(n4468), .A3(n4471), .ZN(n4470) );
  OAI211_X1 U5500 ( .C1(n5398), .C2(n4471), .A(n4470), .B(n4469), .ZN(n4472)
         );
  AOI21_X1 U5501 ( .B1(n4473), .B2(n6099), .A(n4472), .ZN(n4474) );
  NAND2_X1 U5502 ( .A1(n4475), .A2(n4474), .ZN(U2987) );
  NAND2_X1 U5503 ( .A1(n6335), .A2(n6426), .ZN(n5768) );
  INV_X1 U5504 ( .A(n5768), .ZN(n4478) );
  AOI21_X1 U5505 ( .B1(n4476), .B2(MEMORYFETCH_REG_SCAN_IN), .A(n4478), .ZN(
        n4477) );
  NAND2_X1 U5506 ( .A1(n4482), .A2(n4477), .ZN(U2788) );
  NAND2_X1 U5507 ( .A1(n4413), .A2(n3110), .ZN(n5205) );
  OAI21_X1 U5508 ( .B1(n4478), .B2(READREQUEST_REG_SCAN_IN), .A(n6518), .ZN(
        n4479) );
  OAI21_X1 U5509 ( .B1(n6518), .B2(n5205), .A(n4479), .ZN(U3474) );
  INV_X1 U5510 ( .A(DATAI_15_), .ZN(n4484) );
  INV_X1 U5511 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4483) );
  AND2_X1 U5512 ( .A1(n3110), .A2(READY_N), .ZN(n4481) );
  INV_X1 U5513 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6704) );
  OAI222_X1 U5514 ( .A1(n4484), .A2(n4536), .B1(n4483), .B2(n4547), .C1(n5163), 
        .C2(n6704), .ZN(U2954) );
  INV_X1 U5515 ( .A(n4485), .ZN(n4494) );
  OR2_X1 U5516 ( .A1(n4599), .A2(n6452), .ZN(n4487) );
  OAI21_X1 U5517 ( .B1(n4805), .B2(n4557), .A(n4386), .ZN(n4486) );
  AOI21_X1 U5518 ( .B1(n4487), .B2(n4486), .A(READY_N), .ZN(n4492) );
  INV_X1 U5519 ( .A(n4488), .ZN(n4489) );
  NAND2_X1 U5520 ( .A1(n4490), .A2(n4489), .ZN(n4491) );
  AOI21_X1 U5521 ( .B1(n5204), .B2(n4492), .A(n4491), .ZN(n4493) );
  NAND3_X1 U5522 ( .A1(n4494), .A2(n4493), .A3(n4551), .ZN(n6399) );
  NAND2_X1 U5523 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4807) );
  NOR2_X1 U5524 ( .A1(n6525), .A2(n4807), .ZN(n6443) );
  AOI22_X1 U5525 ( .A1(n6399), .A2(n6436), .B1(FLUSH_REG_SCAN_IN), .B2(n6443), 
        .ZN(n5761) );
  NAND2_X1 U5526 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6525), .ZN(n4621) );
  NAND2_X1 U5527 ( .A1(n5761), .A2(n4621), .ZN(n5764) );
  OAI21_X1 U5528 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6431), .A(n5764), 
        .ZN(n4523) );
  INV_X1 U5529 ( .A(n4523), .ZN(n4512) );
  AOI22_X1 U5530 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4471), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6625), .ZN(n5119) );
  NOR2_X1 U5531 ( .A1(n6426), .A2(n4435), .ZN(n4509) );
  INV_X1 U5532 ( .A(n4496), .ZN(n4877) );
  INV_X1 U5533 ( .A(n4497), .ZN(n4502) );
  INV_X1 U5534 ( .A(n4386), .ZN(n4499) );
  NAND3_X1 U5535 ( .A1(n4499), .A2(n4498), .A3(n4421), .ZN(n4500) );
  NOR2_X1 U5536 ( .A1(n4571), .A2(n4500), .ZN(n4501) );
  NAND2_X1 U5537 ( .A1(n4502), .A2(n4501), .ZN(n4595) );
  NAND2_X1 U5538 ( .A1(n4877), .A2(n4595), .ZN(n4508) );
  INV_X1 U5539 ( .A(n4503), .ZN(n4521) );
  INV_X1 U5540 ( .A(n4504), .ZN(n5120) );
  INV_X1 U5541 ( .A(n4505), .ZN(n4506) );
  NAND3_X1 U5542 ( .A1(n4521), .A2(n5120), .A3(n4506), .ZN(n4507) );
  OAI211_X1 U5543 ( .C1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n4599), .A(n4508), .B(n4507), .ZN(n6403) );
  INV_X1 U5544 ( .A(n5760), .ZN(n5123) );
  AOI222_X1 U5545 ( .A1(n5118), .A2(n4510), .B1(n5119), .B2(n4509), .C1(n6403), 
        .C2(n5123), .ZN(n4511) );
  INV_X1 U5546 ( .A(n5764), .ZN(n5124) );
  OAI22_X1 U5547 ( .A1(n4512), .A2(n4495), .B1(n4511), .B2(n5124), .ZN(U3460)
         );
  XNOR2_X1 U5548 ( .A(n4513), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4535)
         );
  OAI21_X1 U5549 ( .B1(n6036), .B2(n4514), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4520) );
  OAI21_X1 U5550 ( .B1(n4517), .B2(n4516), .A(n4515), .ZN(n4941) );
  INV_X1 U5551 ( .A(n4941), .ZN(n4518) );
  AOI22_X1 U5552 ( .A1(n4518), .A2(n5700), .B1(n4228), .B2(REIP_REG_0__SCAN_IN), .ZN(n4519) );
  OAI211_X1 U5553 ( .C1(n4535), .C2(n5773), .A(n4520), .B(n4519), .ZN(U2986)
         );
  INV_X1 U5554 ( .A(n4599), .ZN(n4803) );
  NAND2_X1 U5555 ( .A1(n4803), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6401) );
  INV_X1 U5556 ( .A(n3707), .ZN(n6337) );
  AOI22_X1 U5557 ( .A1(n6337), .A2(n4595), .B1(n4521), .B2(n3144), .ZN(n6402)
         );
  OAI22_X1 U5558 ( .A1(n6402), .A2(n5760), .B1(n6426), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4522) );
  OAI22_X1 U5559 ( .A1(n4523), .A2(n4522), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5764), .ZN(n4524) );
  OAI21_X1 U5560 ( .B1(n6401), .B2(n5760), .A(n4524), .ZN(U3461) );
  INV_X1 U5561 ( .A(n5503), .ZN(n4526) );
  INV_X1 U5562 ( .A(n4525), .ZN(n5031) );
  OAI21_X1 U5563 ( .B1(n4526), .B2(n5031), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4534) );
  INV_X1 U5564 ( .A(n4527), .ZN(n4528) );
  OAI21_X1 U5565 ( .B1(n4529), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4528), 
        .ZN(n4936) );
  INV_X1 U5566 ( .A(n4936), .ZN(n4532) );
  INV_X1 U5567 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6575) );
  OAI21_X1 U5568 ( .B1(n5727), .B2(n6575), .A(n4530), .ZN(n4531) );
  AOI21_X1 U5569 ( .B1(n6099), .B2(n4532), .A(n4531), .ZN(n4533) );
  OAI211_X1 U5570 ( .C1(n4535), .C2(n6103), .A(n4534), .B(n4533), .ZN(U3018)
         );
  INV_X1 U5571 ( .A(LWORD_REG_6__SCAN_IN), .ZN(n6737) );
  NAND2_X1 U5572 ( .A1(n5966), .A2(DATAI_6_), .ZN(n5155) );
  NAND2_X1 U5573 ( .A1(n5969), .A2(EAX_REG_6__SCAN_IN), .ZN(n4537) );
  OAI211_X1 U5574 ( .C1(n4547), .C2(n6737), .A(n5155), .B(n4537), .ZN(U2945)
         );
  INV_X1 U5575 ( .A(LWORD_REG_2__SCAN_IN), .ZN(n6628) );
  NAND2_X1 U5576 ( .A1(n5966), .A2(DATAI_2_), .ZN(n5159) );
  NAND2_X1 U5577 ( .A1(n5969), .A2(EAX_REG_2__SCAN_IN), .ZN(n4538) );
  OAI211_X1 U5578 ( .C1(n4547), .C2(n6628), .A(n5159), .B(n4538), .ZN(U2941)
         );
  INV_X1 U5579 ( .A(LWORD_REG_13__SCAN_IN), .ZN(n5944) );
  NAND2_X1 U5580 ( .A1(n5966), .A2(DATAI_13_), .ZN(n4544) );
  NAND2_X1 U5581 ( .A1(n5969), .A2(EAX_REG_13__SCAN_IN), .ZN(n4539) );
  OAI211_X1 U5582 ( .C1(n4547), .C2(n5944), .A(n4544), .B(n4539), .ZN(U2952)
         );
  INV_X1 U5583 ( .A(LWORD_REG_11__SCAN_IN), .ZN(n6640) );
  NAND2_X1 U5584 ( .A1(n5966), .A2(DATAI_11_), .ZN(n5152) );
  NAND2_X1 U5585 ( .A1(n5969), .A2(EAX_REG_11__SCAN_IN), .ZN(n4540) );
  OAI211_X1 U5586 ( .C1(n4547), .C2(n6640), .A(n5152), .B(n4540), .ZN(U2950)
         );
  INV_X1 U5587 ( .A(LWORD_REG_4__SCAN_IN), .ZN(n5956) );
  NAND2_X1 U5588 ( .A1(n5966), .A2(DATAI_4_), .ZN(n5157) );
  NAND2_X1 U5589 ( .A1(n5969), .A2(EAX_REG_4__SCAN_IN), .ZN(n4541) );
  OAI211_X1 U5590 ( .C1(n4547), .C2(n5956), .A(n5157), .B(n4541), .ZN(U2943)
         );
  INV_X1 U5591 ( .A(UWORD_REG_8__SCAN_IN), .ZN(n6614) );
  NAND2_X1 U5592 ( .A1(n5966), .A2(DATAI_8_), .ZN(n5139) );
  NAND2_X1 U5593 ( .A1(n5969), .A2(EAX_REG_24__SCAN_IN), .ZN(n4542) );
  OAI211_X1 U5594 ( .C1(n4547), .C2(n6614), .A(n5139), .B(n4542), .ZN(U2932)
         );
  INV_X1 U5595 ( .A(UWORD_REG_13__SCAN_IN), .ZN(n6592) );
  NAND2_X1 U5596 ( .A1(n5969), .A2(EAX_REG_29__SCAN_IN), .ZN(n4543) );
  OAI211_X1 U5597 ( .C1(n4547), .C2(n6592), .A(n4544), .B(n4543), .ZN(U2937)
         );
  INV_X1 U5598 ( .A(UWORD_REG_7__SCAN_IN), .ZN(n6545) );
  NAND2_X1 U5599 ( .A1(n5966), .A2(DATAI_7_), .ZN(n5147) );
  NAND2_X1 U5600 ( .A1(n5969), .A2(EAX_REG_23__SCAN_IN), .ZN(n4545) );
  OAI211_X1 U5601 ( .C1(n4547), .C2(n6545), .A(n5147), .B(n4545), .ZN(U2931)
         );
  INV_X1 U5602 ( .A(UWORD_REG_12__SCAN_IN), .ZN(n6677) );
  NAND2_X1 U5603 ( .A1(n5966), .A2(DATAI_12_), .ZN(n5141) );
  NAND2_X1 U5604 ( .A1(n5969), .A2(EAX_REG_28__SCAN_IN), .ZN(n4546) );
  OAI211_X1 U5605 ( .C1(n4547), .C2(n6677), .A(n5141), .B(n4546), .ZN(U2936)
         );
  OR2_X1 U5606 ( .A1(n4549), .A2(n4548), .ZN(n4550) );
  AOI21_X4 U5607 ( .B1(n4551), .B2(n4550), .A(n6434), .ZN(n5927) );
  OR2_X1 U5608 ( .A1(n4553), .A2(n4552), .ZN(n4554) );
  NAND2_X1 U5609 ( .A1(n4555), .A2(n4554), .ZN(n4927) );
  XNOR2_X1 U5610 ( .A(n4556), .B(n4557), .ZN(n4567) );
  INV_X1 U5611 ( .A(n5927), .ZN(n5313) );
  AOI22_X1 U5612 ( .A1(n5923), .A2(n4567), .B1(n5313), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4558) );
  OAI21_X1 U5613 ( .B1(n5316), .B2(n4927), .A(n4558), .ZN(U2858) );
  XNOR2_X1 U5614 ( .A(n4559), .B(n4560), .ZN(n4570) );
  INV_X1 U5615 ( .A(n6026), .ZN(n5700) );
  INV_X1 U5616 ( .A(n4927), .ZN(n4563) );
  AND2_X1 U5617 ( .A1(n4228), .A2(REIP_REG_1__SCAN_IN), .ZN(n4566) );
  AOI21_X1 U5618 ( .B1(n6036), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4566), 
        .ZN(n4561) );
  OAI21_X1 U5619 ( .B1(n6045), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4561), 
        .ZN(n4562) );
  AOI21_X1 U5620 ( .B1(n5700), .B2(n4563), .A(n4562), .ZN(n4564) );
  OAI21_X1 U5621 ( .B1(n4570), .B2(n5773), .A(n4564), .ZN(U2985) );
  INV_X1 U5622 ( .A(n5493), .ZN(n5032) );
  AOI21_X1 U5623 ( .B1(n5503), .B2(n4435), .A(n5032), .ZN(n4565) );
  AOI22_X1 U5624 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4675), .B1(n4565), 
        .B2(n6625), .ZN(n4569) );
  AOI21_X1 U5625 ( .B1(n6099), .B2(n4567), .A(n4566), .ZN(n4568) );
  OAI211_X1 U5626 ( .C1(n4570), .C2(n6103), .A(n4569), .B(n4568), .ZN(U3017)
         );
  OAI222_X1 U5627 ( .A1(n4936), .A2(n5301), .B1(n4258), .B2(n5927), .C1(n4941), 
        .C2(n5316), .ZN(U2859) );
  INV_X1 U5628 ( .A(n4571), .ZN(n5759) );
  INV_X1 U5629 ( .A(n6182), .ZN(n6218) );
  OR2_X1 U5630 ( .A1(n4572), .A2(n6218), .ZN(n4573) );
  XNOR2_X1 U5631 ( .A(n4573), .B(n5763), .ZN(n5758) );
  OAI22_X1 U5632 ( .A1(n6399), .A2(n5763), .B1(n5759), .B2(n5758), .ZN(n4576)
         );
  INV_X1 U5633 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6708) );
  NAND2_X1 U5634 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6708), .ZN(n4577) );
  INV_X1 U5635 ( .A(n4577), .ZN(n4574) );
  AND2_X1 U5636 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n4574), .ZN(n4575)
         );
  AOI21_X1 U5637 ( .B1(n4576), .B2(n6426), .A(n4575), .ZN(n4609) );
  OAI21_X1 U5638 ( .B1(n6399), .B2(STATE2_REG_1__SCAN_IN), .A(n4577), .ZN(
        n4607) );
  NAND2_X1 U5639 ( .A1(n3113), .A2(n4595), .ZN(n4593) );
  INV_X1 U5640 ( .A(n4579), .ZN(n4580) );
  NAND2_X1 U5641 ( .A1(n5196), .A2(n4580), .ZN(n4602) );
  INV_X1 U5642 ( .A(n4581), .ZN(n4587) );
  MUX2_X1 U5643 ( .A(n4587), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4504), 
        .Z(n4584) );
  INV_X1 U5644 ( .A(n4582), .ZN(n4583) );
  NAND2_X1 U5645 ( .A1(n4584), .A2(n4583), .ZN(n4591) );
  XNOR2_X1 U5646 ( .A(n4585), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4589)
         );
  OAI21_X1 U5647 ( .B1(n4504), .B2(n4586), .A(n4587), .ZN(n4588) );
  NOR2_X1 U5648 ( .A1(n4588), .A2(n3116), .ZN(n5511) );
  OAI22_X1 U5649 ( .A1(n4599), .A2(n4589), .B1(n5511), .B2(n4597), .ZN(n4590)
         );
  AOI21_X1 U5650 ( .B1(n4602), .B2(n4591), .A(n4590), .ZN(n4592) );
  NAND2_X1 U5651 ( .A1(n4593), .A2(n4592), .ZN(n6398) );
  INV_X1 U5652 ( .A(n4595), .ZN(n4596) );
  OR2_X1 U5653 ( .A1(n3122), .A2(n4596), .ZN(n4604) );
  XNOR2_X1 U5654 ( .A(n4504), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4601)
         );
  XNOR2_X1 U5655 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4598) );
  OAI22_X1 U5656 ( .A1(n4599), .A2(n4598), .B1(n4597), .B2(n4601), .ZN(n4600)
         );
  AOI21_X1 U5657 ( .B1(n4602), .B2(n4601), .A(n4600), .ZN(n4603) );
  NAND2_X1 U5658 ( .A1(n4604), .A2(n4603), .ZN(n6400) );
  AND3_X1 U5659 ( .A1(n6398), .A2(n6426), .A3(n6400), .ZN(n4605) );
  AOI22_X1 U5660 ( .A1(n4607), .A2(n4606), .B1(n4605), .B2(n6399), .ZN(n4608)
         );
  AND2_X1 U5661 ( .A1(n4609), .A2(n4608), .ZN(n6420) );
  AOI21_X1 U5662 ( .B1(n4609), .B2(n4505), .A(n6420), .ZN(n4612) );
  OAI21_X1 U5663 ( .B1(n4612), .B2(FLUSH_REG_SCAN_IN), .A(n6443), .ZN(n4611)
         );
  INV_X1 U5664 ( .A(n4664), .ZN(n4610) );
  NAND2_X1 U5665 ( .A1(n4611), .A2(n4610), .ZN(n6112) );
  NOR2_X1 U5666 ( .A1(n4612), .A2(n4807), .ZN(n6428) );
  NAND2_X1 U5667 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6817), .ZN(n4687) );
  INV_X1 U5668 ( .A(n4687), .ZN(n4613) );
  OAI22_X1 U5669 ( .A1(n4884), .A2(n6340), .B1(n3707), .B2(n4613), .ZN(n4614)
         );
  OAI21_X1 U5670 ( .B1(n6428), .B2(n4614), .A(n6112), .ZN(n4615) );
  OAI21_X1 U5671 ( .B1(n6112), .B2(n6183), .A(n4615), .ZN(U3465) );
  INV_X1 U5672 ( .A(DATAI_1_), .ZN(n6722) );
  OAI222_X1 U5673 ( .A1(n4927), .A2(n5652), .B1(n5089), .B2(n6722), .C1(n5317), 
        .C2(n3702), .ZN(U2890) );
  AND2_X1 U5674 ( .A1(n4616), .A2(n4617), .ZN(n4743) );
  NOR2_X1 U5675 ( .A1(n4616), .A2(n4617), .ZN(n4618) );
  INV_X1 U5676 ( .A(DATAI_4_), .ZN(n6572) );
  OAI222_X1 U5677 ( .A1(n6025), .A2(n5652), .B1(n5089), .B2(n6572), .C1(n5317), 
        .C2(n3741), .ZN(U2887) );
  INV_X1 U5678 ( .A(DATAI_0_), .ZN(n6740) );
  OAI222_X1 U5679 ( .A1(n4941), .A2(n5652), .B1(n5089), .B2(n6740), .C1(n5317), 
        .C2(n3710), .ZN(U2891) );
  OR2_X1 U5680 ( .A1(n3113), .A2(n6340), .ZN(n6150) );
  NAND2_X1 U5681 ( .A1(n3122), .A2(n4496), .ZN(n6297) );
  OR2_X1 U5682 ( .A1(n6150), .A2(n6297), .ZN(n4620) );
  AND2_X1 U5683 ( .A1(n4629), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6290) );
  AND2_X1 U5684 ( .A1(n4951), .A2(n4952), .ZN(n6148) );
  NAND2_X1 U5685 ( .A1(n6290), .A2(n6148), .ZN(n4619) );
  NAND2_X1 U5686 ( .A1(n4661), .A2(n3338), .ZN(n4896) );
  NAND3_X1 U5687 ( .A1(n6412), .A2(n4866), .A3(n6151), .ZN(n5051) );
  NOR2_X1 U5688 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5051), .ZN(n4652)
         );
  NAND2_X1 U5689 ( .A1(n6116), .A2(n6154), .ZN(n4625) );
  NAND2_X1 U5690 ( .A1(n5049), .A2(n4884), .ZN(n5078) );
  NAND2_X1 U5691 ( .A1(n4663), .A2(DATAI_20_), .ZN(n6376) );
  NAND2_X1 U5692 ( .A1(n4663), .A2(DATAI_28_), .ZN(n6318) );
  INV_X1 U5693 ( .A(n4689), .ZN(n4626) );
  OAI22_X1 U5694 ( .A1(n5078), .A2(n6376), .B1(n6318), .B2(n4856), .ZN(n4627)
         );
  AOI21_X1 U5695 ( .B1(n6371), .B2(n4652), .A(n4627), .ZN(n4634) );
  AND2_X1 U5696 ( .A1(n6335), .A2(n6523), .ZN(n6157) );
  AOI21_X1 U5697 ( .B1(n4628), .B2(n6335), .A(n6157), .ZN(n5050) );
  OAI22_X1 U5698 ( .A1(n4856), .A2(n6157), .B1(n3113), .B2(n6297), .ZN(n4632)
         );
  INV_X1 U5699 ( .A(n4652), .ZN(n4670) );
  OAI21_X1 U5700 ( .B1(n6148), .B2(n6522), .A(n4664), .ZN(n6152) );
  AOI21_X1 U5701 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n4670), .A(n6152), .ZN(
        n4631) );
  INV_X1 U5702 ( .A(n4629), .ZN(n4630) );
  NAND2_X1 U5703 ( .A1(n4630), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6300) );
  OAI211_X1 U5704 ( .C1(n5050), .C2(n4632), .A(n4631), .B(n6300), .ZN(n4662)
         );
  NAND2_X1 U5705 ( .A1(n4662), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4633) );
  OAI211_X1 U5706 ( .C1(n5543), .C2(n4665), .A(n4634), .B(n4633), .ZN(U3024)
         );
  NAND2_X1 U5707 ( .A1(n4661), .A2(n3332), .ZN(n5177) );
  NAND2_X1 U5708 ( .A1(n5700), .A2(DATAI_17_), .ZN(n6356) );
  NAND2_X1 U5709 ( .A1(n4663), .A2(DATAI_25_), .ZN(n6308) );
  OAI22_X1 U5710 ( .A1(n5078), .A2(n6356), .B1(n6308), .B2(n4856), .ZN(n4635)
         );
  AOI21_X1 U5711 ( .B1(n6352), .B2(n4652), .A(n4635), .ZN(n4637) );
  NAND2_X1 U5712 ( .A1(n4662), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4636) );
  OAI211_X1 U5713 ( .C1(n5530), .C2(n4665), .A(n4637), .B(n4636), .ZN(U3021)
         );
  INV_X1 U5714 ( .A(DATAI_2_), .ZN(n4705) );
  NAND2_X1 U5715 ( .A1(n4661), .A2(n3294), .ZN(n4904) );
  NAND2_X1 U5716 ( .A1(n4663), .A2(DATAI_18_), .ZN(n6237) );
  NAND2_X1 U5717 ( .A1(n4663), .A2(DATAI_26_), .ZN(n6362) );
  OAI22_X1 U5718 ( .A1(n5078), .A2(n6237), .B1(n6362), .B2(n4856), .ZN(n4638)
         );
  AOI21_X1 U5719 ( .B1(n6358), .B2(n4652), .A(n4638), .ZN(n4640) );
  NAND2_X1 U5720 ( .A1(n4662), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4639) );
  OAI211_X1 U5721 ( .C1(n5534), .C2(n4665), .A(n4640), .B(n4639), .ZN(U3022)
         );
  NAND2_X1 U5722 ( .A1(n4661), .A2(n3365), .ZN(n4901) );
  NAND2_X1 U5723 ( .A1(n5700), .A2(DATAI_16_), .ZN(n6231) );
  NAND2_X1 U5724 ( .A1(n5700), .A2(DATAI_24_), .ZN(n6350) );
  OAI22_X1 U5725 ( .A1(n5078), .A2(n6231), .B1(n6350), .B2(n4856), .ZN(n4641)
         );
  AOI21_X1 U5726 ( .B1(n6332), .B2(n4652), .A(n4641), .ZN(n4643) );
  NAND2_X1 U5727 ( .A1(n4662), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4642) );
  OAI211_X1 U5728 ( .C1(n5526), .C2(n4665), .A(n4643), .B(n4642), .ZN(U3020)
         );
  INV_X1 U5729 ( .A(DATAI_6_), .ZN(n4697) );
  NAND2_X1 U5730 ( .A1(n4661), .A2(n3293), .ZN(n4907) );
  NAND2_X1 U5731 ( .A1(n4663), .A2(DATAI_22_), .ZN(n6283) );
  NAND2_X1 U5732 ( .A1(n4663), .A2(DATAI_30_), .ZN(n6387) );
  OAI22_X1 U5733 ( .A1(n5078), .A2(n6283), .B1(n6387), .B2(n4856), .ZN(n4644)
         );
  AOI21_X1 U5734 ( .B1(n6383), .B2(n4652), .A(n4644), .ZN(n4646) );
  NAND2_X1 U5735 ( .A1(n4662), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4645) );
  OAI211_X1 U5736 ( .C1(n5551), .C2(n4665), .A(n4646), .B(n4645), .ZN(U3026)
         );
  INV_X1 U5737 ( .A(DATAI_5_), .ZN(n4756) );
  NAND2_X1 U5738 ( .A1(n4661), .A2(n3333), .ZN(n6536) );
  NAND2_X1 U5739 ( .A1(n4663), .A2(DATAI_21_), .ZN(n6534) );
  NAND2_X1 U5740 ( .A1(n4663), .A2(DATAI_29_), .ZN(n6537) );
  OAI22_X1 U5741 ( .A1(n5078), .A2(n6534), .B1(n6537), .B2(n4856), .ZN(n4647)
         );
  AOI21_X1 U5742 ( .B1(n6378), .B2(n4652), .A(n4647), .ZN(n4649) );
  NAND2_X1 U5743 ( .A1(n4662), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4648) );
  OAI211_X1 U5744 ( .C1(n6539), .C2(n4665), .A(n4649), .B(n4648), .ZN(U3025)
         );
  INV_X1 U5745 ( .A(n4662), .ZN(n4654) );
  INV_X1 U5746 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n6772) );
  NAND2_X1 U5747 ( .A1(n4661), .A2(n3350), .ZN(n4917) );
  NAND2_X1 U5748 ( .A1(n4663), .A2(DATAI_19_), .ZN(n6368) );
  NOR2_X1 U5749 ( .A1(n5078), .A2(n6368), .ZN(n4651) );
  NAND2_X1 U5750 ( .A1(n4663), .A2(DATAI_27_), .ZN(n6314) );
  OAI22_X1 U5751 ( .A1(n4856), .A2(n6314), .B1(n4665), .B2(n5536), .ZN(n4650)
         );
  AOI211_X1 U5752 ( .C1(n6364), .C2(n4652), .A(n4651), .B(n4650), .ZN(n4653)
         );
  OAI21_X1 U5753 ( .B1(n4654), .B2(n6772), .A(n4653), .ZN(U3023) );
  INV_X1 U5754 ( .A(n4656), .ZN(n4741) );
  NAND2_X1 U5755 ( .A1(n4655), .A2(n4741), .ZN(n4658) );
  NAND2_X1 U5756 ( .A1(n4658), .A2(n4657), .ZN(n4659) );
  AND2_X1 U5757 ( .A1(n4659), .A2(n4681), .ZN(n6082) );
  INV_X1 U5758 ( .A(n6082), .ZN(n4660) );
  INV_X1 U5759 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6743) );
  OAI222_X1 U5760 ( .A1(n4660), .A2(n5301), .B1(n5927), .B2(n6743), .C1(n6025), 
        .C2(n5316), .ZN(U2855) );
  NAND2_X1 U5761 ( .A1(n4661), .A2(n3349), .ZN(n4912) );
  NAND2_X1 U5762 ( .A1(n4662), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4669) );
  INV_X1 U5763 ( .A(n5078), .ZN(n4667) );
  NAND2_X1 U5764 ( .A1(n4663), .A2(DATAI_23_), .ZN(n6253) );
  INV_X1 U5765 ( .A(n6253), .ZN(n6389) );
  NAND2_X1 U5766 ( .A1(n4663), .A2(DATAI_31_), .ZN(n6397) );
  OAI22_X1 U5767 ( .A1(n4856), .A2(n6397), .B1(n4665), .B2(n5555), .ZN(n4666)
         );
  AOI21_X1 U5768 ( .B1(n4667), .B2(n6389), .A(n4666), .ZN(n4668) );
  OAI211_X1 U5769 ( .C1(n4670), .C2(n4912), .A(n4669), .B(n4668), .ZN(U3027)
         );
  OAI21_X1 U5770 ( .B1(n4673), .B2(n4672), .A(n4671), .ZN(n6011) );
  NOR3_X1 U5771 ( .A1(n4678), .A2(n6081), .A3(n6580), .ZN(n6077) );
  INV_X1 U5772 ( .A(n5028), .ZN(n4674) );
  OR2_X1 U5773 ( .A1(n5104), .A2(n4674), .ZN(n4677) );
  NAND2_X1 U5774 ( .A1(n6095), .A2(n4675), .ZN(n4676) );
  OAI21_X1 U5775 ( .B1(n5032), .B2(n6077), .A(n6104), .ZN(n6074) );
  OR2_X1 U5776 ( .A1(n6081), .A2(n4678), .ZN(n4679) );
  OAI21_X1 U5777 ( .B1(n6095), .B2(n4679), .A(n6580), .ZN(n4685) );
  NAND2_X1 U5778 ( .A1(n4681), .A2(n4680), .ZN(n4682) );
  NAND2_X1 U5779 ( .A1(n4753), .A2(n4682), .ZN(n5915) );
  OAI22_X1 U5780 ( .A1(n5733), .A2(n5915), .B1(n5727), .B2(n6467), .ZN(n4684)
         );
  NOR4_X1 U5781 ( .A1(n5029), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n5028), 
        .A4(n6081), .ZN(n4683) );
  AOI211_X1 U5782 ( .C1(n6074), .C2(n4685), .A(n4684), .B(n4683), .ZN(n4686)
         );
  OAI21_X1 U5783 ( .B1(n6103), .B2(n6011), .A(n4686), .ZN(U3013) );
  INV_X1 U5784 ( .A(n3113), .ZN(n6298) );
  NAND2_X1 U5785 ( .A1(n6112), .A2(n4687), .ZN(n5191) );
  NAND2_X1 U5786 ( .A1(n6112), .A2(n6335), .ZN(n5187) );
  INV_X1 U5787 ( .A(n5187), .ZN(n4692) );
  NAND2_X1 U5788 ( .A1(n4885), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4876) );
  NAND2_X1 U5789 ( .A1(n3114), .A2(n6523), .ZN(n4690) );
  NAND2_X1 U5790 ( .A1(n4825), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6333) );
  INV_X1 U5791 ( .A(n6333), .ZN(n6117) );
  NAND2_X1 U5792 ( .A1(n6255), .A2(n6117), .ZN(n6256) );
  NAND4_X1 U5793 ( .A1(n4876), .A2(n6334), .A3(n4690), .A4(n6256), .ZN(n4691)
         );
  INV_X1 U5794 ( .A(n6112), .ZN(n5189) );
  AOI22_X1 U5795 ( .A1(n4692), .A2(n4691), .B1(n5189), .B2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4693) );
  OAI21_X1 U5796 ( .B1(n6298), .B2(n5191), .A(n4693), .ZN(U3462) );
  XNOR2_X1 U5797 ( .A(n6116), .B(n6333), .ZN(n4694) );
  OAI222_X1 U5798 ( .A1(n5191), .A2(n3122), .B1(n6112), .B2(n4866), .C1(n5187), 
        .C2(n4694), .ZN(U3463) );
  XNOR2_X1 U5799 ( .A(n4696), .B(n4695), .ZN(n6010) );
  OAI222_X1 U5800 ( .A1(n5652), .A2(n6010), .B1(n5317), .B2(n3751), .C1(n4697), 
        .C2(n5089), .ZN(U2885) );
  XNOR2_X1 U5801 ( .A(n4698), .B(n4699), .ZN(n6031) );
  INV_X1 U5802 ( .A(DATAI_3_), .ZN(n4701) );
  OAI222_X1 U5803 ( .A1(n6031), .A2(n5652), .B1(n4701), .B2(n5089), .C1(n5317), 
        .C2(n4700), .ZN(U2888) );
  NOR2_X1 U5804 ( .A1(n4703), .A2(n4702), .ZN(n4704) );
  NOR2_X1 U5805 ( .A1(n4698), .A2(n4704), .ZN(n6042) );
  INV_X1 U5806 ( .A(n6042), .ZN(n4751) );
  OAI222_X1 U5807 ( .A1(n4751), .A2(n5652), .B1(n5089), .B2(n4705), .C1(n5317), 
        .C2(n3719), .ZN(U2889) );
  NOR2_X1 U5808 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4706), .ZN(n4737)
         );
  INV_X1 U5809 ( .A(n4737), .ZN(n4727) );
  OR2_X1 U5810 ( .A1(n3122), .A2(n4496), .ZN(n6259) );
  AOI21_X1 U5811 ( .B1(n6259), .B2(n6157), .A(n6290), .ZN(n6222) );
  OAI21_X1 U5812 ( .B1(n6817), .B2(n4737), .A(n6222), .ZN(n4708) );
  NAND2_X1 U5813 ( .A1(n6259), .A2(n6335), .ZN(n6223) );
  INV_X1 U5814 ( .A(n4849), .ZN(n4858) );
  AOI211_X1 U5815 ( .C1(n6223), .C2(n6150), .A(n4858), .B(n5167), .ZN(n4707)
         );
  NOR2_X1 U5816 ( .A1(n4708), .A2(n4707), .ZN(n4709) );
  INV_X1 U5817 ( .A(n4952), .ZN(n5514) );
  NAND2_X1 U5818 ( .A1(n5514), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4772) );
  AOI21_X1 U5819 ( .B1(n4772), .B2(STATE2_REG_2__SCAN_IN), .A(n4610), .ZN(
        n4777) );
  NAND2_X1 U5820 ( .A1(n4709), .A2(n4777), .ZN(n4734) );
  NAND2_X1 U5821 ( .A1(n4734), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4714)
         );
  INV_X1 U5822 ( .A(n6314), .ZN(n6363) );
  NAND2_X1 U5823 ( .A1(n3113), .A2(n6335), .ZN(n6293) );
  OR2_X1 U5824 ( .A1(n6259), .A2(n6293), .ZN(n4711) );
  OR2_X1 U5825 ( .A1(n6300), .A2(n4772), .ZN(n4710) );
  OAI22_X1 U5826 ( .A1(n4849), .A2(n6368), .B1(n4740), .B2(n5536), .ZN(n4712)
         );
  AOI21_X1 U5827 ( .B1(n6363), .B2(n5167), .A(n4712), .ZN(n4713) );
  OAI211_X1 U5828 ( .C1(n4727), .C2(n4917), .A(n4714), .B(n4713), .ZN(U3135)
         );
  NAND2_X1 U5829 ( .A1(n4734), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4717)
         );
  OAI22_X1 U5830 ( .A1(n4735), .A2(n6362), .B1(n6237), .B2(n4849), .ZN(n4715)
         );
  AOI21_X1 U5831 ( .B1(n6358), .B2(n4737), .A(n4715), .ZN(n4716) );
  OAI211_X1 U5832 ( .C1(n4740), .C2(n5534), .A(n4717), .B(n4716), .ZN(U3134)
         );
  NAND2_X1 U5833 ( .A1(n4734), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4720)
         );
  OAI22_X1 U5834 ( .A1(n4735), .A2(n6308), .B1(n6356), .B2(n4849), .ZN(n4718)
         );
  AOI21_X1 U5835 ( .B1(n6352), .B2(n4737), .A(n4718), .ZN(n4719) );
  OAI211_X1 U5836 ( .C1(n4740), .C2(n5530), .A(n4720), .B(n4719), .ZN(U3133)
         );
  NAND2_X1 U5837 ( .A1(n4734), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4723)
         );
  OAI22_X1 U5838 ( .A1(n4735), .A2(n6350), .B1(n6231), .B2(n4849), .ZN(n4721)
         );
  AOI21_X1 U5839 ( .B1(n6332), .B2(n4737), .A(n4721), .ZN(n4722) );
  OAI211_X1 U5840 ( .C1(n4740), .C2(n5526), .A(n4723), .B(n4722), .ZN(U3132)
         );
  NAND2_X1 U5841 ( .A1(n4734), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4726)
         );
  INV_X1 U5842 ( .A(n6397), .ZN(n6249) );
  OAI22_X1 U5843 ( .A1(n4849), .A2(n6253), .B1(n4740), .B2(n5555), .ZN(n4724)
         );
  AOI21_X1 U5844 ( .B1(n6249), .B2(n5167), .A(n4724), .ZN(n4725) );
  OAI211_X1 U5845 ( .C1(n4727), .C2(n4912), .A(n4726), .B(n4725), .ZN(U3139)
         );
  NAND2_X1 U5846 ( .A1(n4734), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4730)
         );
  OAI22_X1 U5847 ( .A1(n4735), .A2(n6387), .B1(n6283), .B2(n4849), .ZN(n4728)
         );
  AOI21_X1 U5848 ( .B1(n6383), .B2(n4737), .A(n4728), .ZN(n4729) );
  OAI211_X1 U5849 ( .C1(n4740), .C2(n5551), .A(n4730), .B(n4729), .ZN(U3138)
         );
  NAND2_X1 U5850 ( .A1(n4734), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4733)
         );
  OAI22_X1 U5851 ( .A1(n4735), .A2(n6537), .B1(n6534), .B2(n4849), .ZN(n4731)
         );
  AOI21_X1 U5852 ( .B1(n6378), .B2(n4737), .A(n4731), .ZN(n4732) );
  OAI211_X1 U5853 ( .C1(n4740), .C2(n6539), .A(n4733), .B(n4732), .ZN(U3137)
         );
  NAND2_X1 U5854 ( .A1(n4734), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4739)
         );
  OAI22_X1 U5855 ( .A1(n4735), .A2(n6318), .B1(n6376), .B2(n4849), .ZN(n4736)
         );
  AOI21_X1 U5856 ( .B1(n6371), .B2(n4737), .A(n4736), .ZN(n4738) );
  OAI211_X1 U5857 ( .C1(n4740), .C2(n5543), .A(n4739), .B(n4738), .ZN(U3136)
         );
  XNOR2_X1 U5858 ( .A(n4655), .B(n4741), .ZN(n6087) );
  OAI222_X1 U5859 ( .A1(n5316), .A2(n6031), .B1(n4974), .B2(n5927), .C1(n5301), 
        .C2(n6087), .ZN(U2856) );
  XOR2_X1 U5860 ( .A(n4742), .B(n4743), .Z(n6013) );
  OAI22_X1 U5861 ( .A1(n5301), .A2(n5915), .B1(n4744), .B2(n5927), .ZN(n4745)
         );
  AOI21_X1 U5862 ( .B1(n6013), .B2(n5924), .A(n4745), .ZN(n4746) );
  INV_X1 U5863 ( .A(n4746), .ZN(U2854) );
  NOR2_X1 U5864 ( .A1(n4748), .A2(n4747), .ZN(n4749) );
  OR2_X1 U5865 ( .A1(n4655), .A2(n4749), .ZN(n5007) );
  INV_X1 U5866 ( .A(n5007), .ZN(n6098) );
  AOI22_X1 U5867 ( .A1(n5923), .A2(n6098), .B1(n5313), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4750) );
  OAI21_X1 U5868 ( .B1(n4751), .B2(n5316), .A(n4750), .ZN(U2857) );
  NAND2_X1 U5869 ( .A1(n4753), .A2(n4752), .ZN(n4754) );
  AND2_X1 U5870 ( .A1(n5880), .A2(n4754), .ZN(n6073) );
  AOI22_X1 U5871 ( .A1(n5923), .A2(n6073), .B1(n5313), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4755) );
  OAI21_X1 U5872 ( .B1(n6010), .B2(n5316), .A(n4755), .ZN(U2853) );
  INV_X1 U5873 ( .A(n6013), .ZN(n4757) );
  OAI222_X1 U5874 ( .A1(n5652), .A2(n4757), .B1(n5317), .B2(n3733), .C1(n4756), 
        .C2(n5089), .ZN(U2886) );
  XNOR2_X1 U5875 ( .A(n4758), .B(n4759), .ZN(n5994) );
  INV_X1 U5876 ( .A(n5880), .ZN(n4761) );
  AOI21_X1 U5877 ( .B1(n4761), .B2(n5879), .A(n4760), .ZN(n4762) );
  NOR2_X1 U5878 ( .A1(n4762), .A2(n5036), .ZN(n6060) );
  AOI22_X1 U5879 ( .A1(n5923), .A2(n6060), .B1(n5313), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n4763) );
  OAI21_X1 U5880 ( .B1(n5316), .B2(n5994), .A(n4763), .ZN(U2851) );
  INV_X1 U5881 ( .A(DATAI_8_), .ZN(n4764) );
  OAI222_X1 U5882 ( .A1(n5994), .A2(n5652), .B1(n5089), .B2(n4764), .C1(n5317), 
        .C2(n3776), .ZN(U2883) );
  OAI21_X1 U5883 ( .B1(n4765), .B2(n4768), .A(n4767), .ZN(n5986) );
  XNOR2_X1 U5884 ( .A(n5036), .B(n5034), .ZN(n6054) );
  AOI22_X1 U5885 ( .A1(n5923), .A2(n6054), .B1(n5313), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n4769) );
  OAI21_X1 U5886 ( .B1(n5986), .B2(n5316), .A(n4769), .ZN(U2850) );
  AOI22_X1 U5887 ( .A1(n5335), .A2(DATAI_9_), .B1(n5931), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n4770) );
  OAI21_X1 U5888 ( .B1(n5986), .B2(n5652), .A(n4770), .ZN(U2882) );
  NOR2_X1 U5889 ( .A1(n4873), .A2(n4884), .ZN(n5174) );
  OAI21_X1 U5890 ( .B1(n5174), .B2(n6369), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4771) );
  NAND2_X1 U5891 ( .A1(n4771), .A2(n6335), .ZN(n4776) );
  INV_X1 U5892 ( .A(n4776), .ZN(n4774) );
  NAND2_X1 U5893 ( .A1(n3122), .A2(n4877), .ZN(n6119) );
  INV_X1 U5894 ( .A(n6119), .ZN(n5516) );
  AND2_X1 U5895 ( .A1(n5516), .A2(n3113), .ZN(n6338) );
  INV_X1 U5896 ( .A(n4772), .ZN(n4773) );
  NAND3_X1 U5897 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6339), .A3(n6183), .ZN(n6535) );
  INV_X1 U5898 ( .A(n6535), .ZN(n4800) );
  INV_X1 U5899 ( .A(n5174), .ZN(n6538) );
  OAI22_X1 U5900 ( .A1(n6538), .A2(n6362), .B1(n6237), .B2(n6533), .ZN(n4775)
         );
  AOI21_X1 U5901 ( .B1(n6358), .B2(n4800), .A(n4775), .ZN(n4783) );
  OR2_X1 U5902 ( .A1(n4776), .A2(n6338), .ZN(n4781) );
  INV_X1 U5903 ( .A(n4777), .ZN(n4778) );
  AOI21_X1 U5904 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6535), .A(n4778), .ZN(
        n4779) );
  AND2_X1 U5905 ( .A1(n6300), .A2(n4779), .ZN(n4780) );
  NAND2_X1 U5906 ( .A1(n6543), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4782)
         );
  OAI211_X1 U5907 ( .C1(n6540), .C2(n5534), .A(n4783), .B(n4782), .ZN(U3102)
         );
  OAI22_X1 U5908 ( .A1(n6538), .A2(n6397), .B1(n6253), .B2(n6533), .ZN(n4784)
         );
  AOI21_X1 U5909 ( .B1(n6391), .B2(n4800), .A(n4784), .ZN(n4786) );
  NAND2_X1 U5910 ( .A1(n6543), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4785)
         );
  OAI211_X1 U5911 ( .C1(n6540), .C2(n5555), .A(n4786), .B(n4785), .ZN(U3107)
         );
  OAI22_X1 U5912 ( .A1(n6538), .A2(n6308), .B1(n6356), .B2(n6533), .ZN(n4787)
         );
  AOI21_X1 U5913 ( .B1(n6352), .B2(n4800), .A(n4787), .ZN(n4789) );
  NAND2_X1 U5914 ( .A1(n6543), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4788)
         );
  OAI211_X1 U5915 ( .C1(n6540), .C2(n5530), .A(n4789), .B(n4788), .ZN(U3101)
         );
  OAI22_X1 U5916 ( .A1(n6538), .A2(n6314), .B1(n6368), .B2(n6533), .ZN(n4790)
         );
  AOI21_X1 U5917 ( .B1(n6364), .B2(n4800), .A(n4790), .ZN(n4792) );
  NAND2_X1 U5918 ( .A1(n6543), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4791)
         );
  OAI211_X1 U5919 ( .C1(n6540), .C2(n5536), .A(n4792), .B(n4791), .ZN(U3103)
         );
  OAI22_X1 U5920 ( .A1(n6538), .A2(n6318), .B1(n6376), .B2(n6533), .ZN(n4793)
         );
  AOI21_X1 U5921 ( .B1(n6371), .B2(n4800), .A(n4793), .ZN(n4795) );
  NAND2_X1 U5922 ( .A1(n6543), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4794)
         );
  OAI211_X1 U5923 ( .C1(n6540), .C2(n5543), .A(n4795), .B(n4794), .ZN(U3104)
         );
  OAI22_X1 U5924 ( .A1(n6538), .A2(n6350), .B1(n6231), .B2(n6533), .ZN(n4796)
         );
  AOI21_X1 U5925 ( .B1(n6332), .B2(n4800), .A(n4796), .ZN(n4798) );
  NAND2_X1 U5926 ( .A1(n6543), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4797)
         );
  OAI211_X1 U5927 ( .C1(n6540), .C2(n5526), .A(n4798), .B(n4797), .ZN(U3100)
         );
  OAI22_X1 U5928 ( .A1(n6538), .A2(n6387), .B1(n6283), .B2(n6533), .ZN(n4799)
         );
  AOI21_X1 U5929 ( .B1(n6383), .B2(n4800), .A(n4799), .ZN(n4802) );
  NAND2_X1 U5930 ( .A1(n6543), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4801)
         );
  OAI211_X1 U5931 ( .C1(n6540), .C2(n5551), .A(n4802), .B(n4801), .ZN(U3106)
         );
  INV_X1 U5932 ( .A(EAX_REG_22__SCAN_IN), .ZN(n6559) );
  NAND3_X1 U5933 ( .A1(n5204), .A2(n6436), .A3(n4803), .ZN(n4804) );
  NAND2_X1 U5934 ( .A1(n4808), .A2(n3365), .ZN(n5935) );
  NOR2_X1 U5935 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4807), .ZN(n5963) );
  AOI22_X1 U5936 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n5960), .B1(n5962), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4809) );
  OAI21_X1 U5937 ( .B1(n6559), .B2(n5935), .A(n4809), .ZN(U2901) );
  INV_X1 U5938 ( .A(EAX_REG_18__SCAN_IN), .ZN(n5160) );
  AOI22_X1 U5939 ( .A1(n5963), .A2(UWORD_REG_2__SCAN_IN), .B1(n5962), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4810) );
  OAI21_X1 U5940 ( .B1(n5160), .B2(n5935), .A(n4810), .ZN(U2905) );
  INV_X1 U5941 ( .A(EAX_REG_19__SCAN_IN), .ZN(n5130) );
  AOI22_X1 U5942 ( .A1(n5963), .A2(UWORD_REG_3__SCAN_IN), .B1(n5962), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4811) );
  OAI21_X1 U5943 ( .B1(n5130), .B2(n5935), .A(n4811), .ZN(U2904) );
  AOI22_X1 U5944 ( .A1(n5963), .A2(UWORD_REG_4__SCAN_IN), .B1(n5962), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4812) );
  OAI21_X1 U5945 ( .B1(n3952), .B2(n5935), .A(n4812), .ZN(U2903) );
  INV_X1 U5946 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6622) );
  AOI22_X1 U5947 ( .A1(n5960), .A2(UWORD_REG_5__SCAN_IN), .B1(n5962), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4813) );
  OAI21_X1 U5948 ( .B1(n6622), .B2(n5935), .A(n4813), .ZN(U2902) );
  INV_X1 U5949 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6707) );
  AOI22_X1 U5950 ( .A1(n5960), .A2(UWORD_REG_14__SCAN_IN), .B1(n5962), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4814) );
  OAI21_X1 U5951 ( .B1(n6707), .B2(n5935), .A(n4814), .ZN(U2893) );
  INV_X1 U5952 ( .A(EAX_REG_16__SCAN_IN), .ZN(n5164) );
  AOI22_X1 U5953 ( .A1(n5960), .A2(UWORD_REG_0__SCAN_IN), .B1(n5962), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4815) );
  OAI21_X1 U5954 ( .B1(n5164), .B2(n5935), .A(n4815), .ZN(U2907) );
  INV_X1 U5955 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6751) );
  AOI22_X1 U5956 ( .A1(n5960), .A2(UWORD_REG_10__SCAN_IN), .B1(n5962), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4816) );
  OAI21_X1 U5957 ( .B1(n6751), .B2(n5935), .A(n4816), .ZN(U2897) );
  INV_X1 U5958 ( .A(EAX_REG_27__SCAN_IN), .ZN(n5153) );
  AOI22_X1 U5959 ( .A1(n5960), .A2(UWORD_REG_11__SCAN_IN), .B1(n5962), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4817) );
  OAI21_X1 U5960 ( .B1(n5153), .B2(n5935), .A(n4817), .ZN(U2896) );
  INV_X1 U5961 ( .A(EAX_REG_17__SCAN_IN), .ZN(n5128) );
  AOI22_X1 U5962 ( .A1(n5960), .A2(UWORD_REG_1__SCAN_IN), .B1(n5962), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4818) );
  OAI21_X1 U5963 ( .B1(n5128), .B2(n5935), .A(n4818), .ZN(U2906) );
  INV_X1 U5964 ( .A(DATAI_7_), .ZN(n4822) );
  XOR2_X1 U5965 ( .A(n4819), .B(n4820), .Z(n5999) );
  INV_X1 U5966 ( .A(n5999), .ZN(n4821) );
  OAI222_X1 U5967 ( .A1(n4823), .A2(n5317), .B1(n4822), .B2(n5089), .C1(n5652), 
        .C2(n4821), .ZN(U2884) );
  AND2_X1 U5968 ( .A1(n3113), .A2(n6337), .ZN(n4879) );
  INV_X1 U5969 ( .A(n6259), .ZN(n6219) );
  INV_X1 U5970 ( .A(n4861), .ZN(n4851) );
  AOI21_X1 U5971 ( .B1(n4879), .B2(n6219), .A(n4851), .ZN(n4827) );
  INV_X1 U5972 ( .A(n4827), .ZN(n4824) );
  AOI22_X1 U5973 ( .A1(n4824), .A2(n6335), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4830), .ZN(n4855) );
  AOI21_X1 U5974 ( .B1(n4826), .B2(n4825), .A(n6026), .ZN(n4828) );
  OAI21_X1 U5975 ( .B1(n4828), .B2(n6157), .A(n4827), .ZN(n4829) );
  OAI211_X1 U5976 ( .C1(n6335), .C2(n4830), .A(n6342), .B(n4829), .ZN(n4854)
         );
  NAND2_X1 U5977 ( .A1(n4854), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4833)
         );
  OAI22_X1 U5978 ( .A1(n6308), .A2(n4849), .B1(n4856), .B2(n6356), .ZN(n4831)
         );
  AOI21_X1 U5979 ( .B1(n6352), .B2(n4851), .A(n4831), .ZN(n4832) );
  OAI211_X1 U5980 ( .C1(n4855), .C2(n5530), .A(n4833), .B(n4832), .ZN(U3141)
         );
  NAND2_X1 U5981 ( .A1(n4854), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4836)
         );
  OAI22_X1 U5982 ( .A1(n6362), .A2(n4849), .B1(n4856), .B2(n6237), .ZN(n4834)
         );
  AOI21_X1 U5983 ( .B1(n6358), .B2(n4851), .A(n4834), .ZN(n4835) );
  OAI211_X1 U5984 ( .C1(n4855), .C2(n5534), .A(n4836), .B(n4835), .ZN(U3142)
         );
  NAND2_X1 U5985 ( .A1(n4854), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4839)
         );
  OAI22_X1 U5986 ( .A1(n6350), .A2(n4849), .B1(n4856), .B2(n6231), .ZN(n4837)
         );
  AOI21_X1 U5987 ( .B1(n6332), .B2(n4851), .A(n4837), .ZN(n4838) );
  OAI211_X1 U5988 ( .C1(n4855), .C2(n5526), .A(n4839), .B(n4838), .ZN(U3140)
         );
  NAND2_X1 U5989 ( .A1(n4854), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4842)
         );
  OAI22_X1 U5990 ( .A1(n6387), .A2(n4849), .B1(n4856), .B2(n6283), .ZN(n4840)
         );
  AOI21_X1 U5991 ( .B1(n6383), .B2(n4851), .A(n4840), .ZN(n4841) );
  OAI211_X1 U5992 ( .C1(n4855), .C2(n5551), .A(n4842), .B(n4841), .ZN(U3146)
         );
  NAND2_X1 U5993 ( .A1(n4854), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4845)
         );
  OAI22_X1 U5994 ( .A1(n4856), .A2(n6253), .B1(n4855), .B2(n5555), .ZN(n4843)
         );
  AOI21_X1 U5995 ( .B1(n6249), .B2(n4858), .A(n4843), .ZN(n4844) );
  OAI211_X1 U5996 ( .C1(n4912), .C2(n4861), .A(n4845), .B(n4844), .ZN(U3147)
         );
  NAND2_X1 U5997 ( .A1(n4854), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4848)
         );
  OAI22_X1 U5998 ( .A1(n6318), .A2(n4849), .B1(n4856), .B2(n6376), .ZN(n4846)
         );
  AOI21_X1 U5999 ( .B1(n6371), .B2(n4851), .A(n4846), .ZN(n4847) );
  OAI211_X1 U6000 ( .C1(n4855), .C2(n5543), .A(n4848), .B(n4847), .ZN(U3144)
         );
  NAND2_X1 U6001 ( .A1(n4854), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4853)
         );
  OAI22_X1 U6002 ( .A1(n6537), .A2(n4849), .B1(n4856), .B2(n6534), .ZN(n4850)
         );
  AOI21_X1 U6003 ( .B1(n6378), .B2(n4851), .A(n4850), .ZN(n4852) );
  OAI211_X1 U6004 ( .C1(n4855), .C2(n6539), .A(n4853), .B(n4852), .ZN(U3145)
         );
  NAND2_X1 U6005 ( .A1(n4854), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4860)
         );
  OAI22_X1 U6006 ( .A1(n4856), .A2(n6368), .B1(n4855), .B2(n5536), .ZN(n4857)
         );
  AOI21_X1 U6007 ( .B1(n6363), .B2(n4858), .A(n4857), .ZN(n4859) );
  OAI211_X1 U6008 ( .C1(n4917), .C2(n4861), .A(n4860), .B(n4859), .ZN(U3143)
         );
  AOI21_X1 U6009 ( .B1(n4767), .B2(n4863), .A(n4862), .ZN(n5921) );
  INV_X1 U6010 ( .A(n5921), .ZN(n4865) );
  AOI22_X1 U6011 ( .A1(n5335), .A2(DATAI_10_), .B1(n5931), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n4864) );
  OAI21_X1 U6012 ( .B1(n4865), .B2(n5652), .A(n4864), .ZN(U2881) );
  NAND3_X1 U6013 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4866), .A3(n6151), .ZN(n6294) );
  NOR2_X1 U6014 ( .A1(n6183), .A2(n6294), .ZN(n4867) );
  INV_X1 U6015 ( .A(n4867), .ZN(n5178) );
  OAI21_X1 U6016 ( .B1(n4873), .B2(n6523), .A(n6335), .ZN(n4872) );
  INV_X1 U6017 ( .A(n6297), .ZN(n4868) );
  AOI21_X1 U6018 ( .B1(n4879), .B2(n4868), .A(n4867), .ZN(n4871) );
  INV_X1 U6019 ( .A(n4871), .ZN(n4870) );
  NAND2_X1 U6020 ( .A1(n6340), .A2(n6294), .ZN(n4869) );
  OAI211_X1 U6021 ( .C1(n4872), .C2(n4870), .A(n6342), .B(n4869), .ZN(n5173)
         );
  OAI22_X1 U6022 ( .A1(n4872), .A2(n4871), .B1(n6522), .B2(n6294), .ZN(n5172)
         );
  AOI22_X1 U6023 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n5173), .B1(n6359), 
        .B2(n5172), .ZN(n4875) );
  INV_X1 U6024 ( .A(n6362), .ZN(n6234) );
  INV_X1 U6025 ( .A(n6237), .ZN(n6357) );
  AOI22_X1 U6026 ( .A1(n6325), .A2(n6234), .B1(n5174), .B2(n6357), .ZN(n4874)
         );
  OAI211_X1 U6027 ( .C1(n5178), .C2(n4904), .A(n4875), .B(n4874), .ZN(U3094)
         );
  NAND3_X1 U6028 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6151), .ZN(n4950) );
  NOR2_X1 U6029 ( .A1(n6183), .A2(n4950), .ZN(n4878) );
  INV_X1 U6030 ( .A(n4878), .ZN(n5171) );
  NAND2_X1 U6031 ( .A1(n6335), .A2(n4876), .ZN(n4882) );
  NOR2_X1 U6032 ( .A1(n3122), .A2(n4877), .ZN(n6155) );
  AOI21_X1 U6033 ( .B1(n4879), .B2(n6155), .A(n4878), .ZN(n4883) );
  INV_X1 U6034 ( .A(n4883), .ZN(n4881) );
  NAND2_X1 U6035 ( .A1(n6340), .A2(n4950), .ZN(n4880) );
  OAI211_X1 U6036 ( .C1(n4882), .C2(n4881), .A(n6342), .B(n4880), .ZN(n5166)
         );
  OAI22_X1 U6037 ( .A1(n4883), .A2(n4882), .B1(n6522), .B2(n4950), .ZN(n5165)
         );
  AOI22_X1 U6038 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n5166), .B1(n6384), 
        .B2(n5165), .ZN(n4887) );
  INV_X1 U6039 ( .A(n6387), .ZN(n6280) );
  AND2_X1 U6040 ( .A1(n4885), .A2(n4884), .ZN(n5168) );
  INV_X1 U6041 ( .A(n6283), .ZN(n6382) );
  AOI22_X1 U6042 ( .A1(n6280), .A2(n5168), .B1(n5167), .B2(n6382), .ZN(n4886)
         );
  OAI211_X1 U6043 ( .C1(n4907), .C2(n5171), .A(n4887), .B(n4886), .ZN(U3130)
         );
  AOI22_X1 U6044 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n5166), .B1(n6347), 
        .B2(n5165), .ZN(n4889) );
  INV_X1 U6045 ( .A(n6350), .ZN(n6228) );
  INV_X1 U6046 ( .A(n6231), .ZN(n6331) );
  AOI22_X1 U6047 ( .A1(n6228), .A2(n5168), .B1(n5167), .B2(n6331), .ZN(n4888)
         );
  OAI211_X1 U6048 ( .C1(n4901), .C2(n5171), .A(n4889), .B(n4888), .ZN(U3124)
         );
  AOI22_X1 U6049 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n5166), .B1(n6372), 
        .B2(n5165), .ZN(n4891) );
  INV_X1 U6050 ( .A(n6318), .ZN(n6370) );
  INV_X1 U6051 ( .A(n6376), .ZN(n6315) );
  AOI22_X1 U6052 ( .A1(n6370), .A2(n5168), .B1(n5167), .B2(n6315), .ZN(n4890)
         );
  OAI211_X1 U6053 ( .C1(n4896), .C2(n5171), .A(n4891), .B(n4890), .ZN(U3128)
         );
  AOI22_X1 U6054 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n5166), .B1(n6365), 
        .B2(n5165), .ZN(n4893) );
  INV_X1 U6055 ( .A(n6368), .ZN(n6311) );
  AOI22_X1 U6056 ( .A1(n6363), .A2(n5168), .B1(n5167), .B2(n6311), .ZN(n4892)
         );
  OAI211_X1 U6057 ( .C1(n4917), .C2(n5171), .A(n4893), .B(n4892), .ZN(U3127)
         );
  AOI22_X1 U6058 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5173), .B1(n6372), 
        .B2(n5172), .ZN(n4895) );
  AOI22_X1 U6059 ( .A1(n6325), .A2(n6370), .B1(n5174), .B2(n6315), .ZN(n4894)
         );
  OAI211_X1 U6060 ( .C1(n5178), .C2(n4896), .A(n4895), .B(n4894), .ZN(U3096)
         );
  AOI22_X1 U6061 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n5166), .B1(n6379), 
        .B2(n5165), .ZN(n4898) );
  INV_X1 U6062 ( .A(n6537), .ZN(n6276) );
  INV_X1 U6063 ( .A(n6534), .ZN(n6377) );
  AOI22_X1 U6064 ( .A1(n6276), .A2(n5168), .B1(n5167), .B2(n6377), .ZN(n4897)
         );
  OAI211_X1 U6065 ( .C1(n6536), .C2(n5171), .A(n4898), .B(n4897), .ZN(U3129)
         );
  AOI22_X1 U6066 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5173), .B1(n6347), 
        .B2(n5172), .ZN(n4900) );
  AOI22_X1 U6067 ( .A1(n6228), .A2(n6325), .B1(n5174), .B2(n6331), .ZN(n4899)
         );
  OAI211_X1 U6068 ( .C1(n5178), .C2(n4901), .A(n4900), .B(n4899), .ZN(U3092)
         );
  AOI22_X1 U6069 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n5166), .B1(n6359), 
        .B2(n5165), .ZN(n4903) );
  AOI22_X1 U6070 ( .A1(n6234), .A2(n5168), .B1(n5167), .B2(n6357), .ZN(n4902)
         );
  OAI211_X1 U6071 ( .C1(n4904), .C2(n5171), .A(n4903), .B(n4902), .ZN(U3126)
         );
  AOI22_X1 U6072 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n5173), .B1(n6384), 
        .B2(n5172), .ZN(n4906) );
  AOI22_X1 U6073 ( .A1(n6325), .A2(n6280), .B1(n5174), .B2(n6382), .ZN(n4905)
         );
  OAI211_X1 U6074 ( .C1(n5178), .C2(n4907), .A(n4906), .B(n4905), .ZN(U3098)
         );
  AOI22_X1 U6075 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n5166), .B1(n6393), 
        .B2(n5165), .ZN(n4909) );
  AOI22_X1 U6076 ( .A1(n6249), .A2(n5168), .B1(n5167), .B2(n6389), .ZN(n4908)
         );
  OAI211_X1 U6077 ( .C1(n4912), .C2(n5171), .A(n4909), .B(n4908), .ZN(U3131)
         );
  AOI22_X1 U6078 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5173), .B1(n6393), 
        .B2(n5172), .ZN(n4911) );
  AOI22_X1 U6079 ( .A1(n6325), .A2(n6249), .B1(n5174), .B2(n6389), .ZN(n4910)
         );
  OAI211_X1 U6080 ( .C1(n5178), .C2(n4912), .A(n4911), .B(n4910), .ZN(U3099)
         );
  AOI22_X1 U6081 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n5173), .B1(n6379), 
        .B2(n5172), .ZN(n4914) );
  AOI22_X1 U6082 ( .A1(n6325), .A2(n6276), .B1(n5174), .B2(n6377), .ZN(n4913)
         );
  OAI211_X1 U6083 ( .C1(n5178), .C2(n6536), .A(n4914), .B(n4913), .ZN(U3097)
         );
  AOI22_X1 U6084 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n5173), .B1(n6365), 
        .B2(n5172), .ZN(n4916) );
  AOI22_X1 U6085 ( .A1(n6325), .A2(n6363), .B1(n5174), .B2(n6311), .ZN(n4915)
         );
  OAI211_X1 U6086 ( .C1(n5178), .C2(n4917), .A(n4916), .B(n4915), .ZN(U3095)
         );
  AOI21_X1 U6087 ( .B1(n3108), .B2(n4918), .A(n5886), .ZN(n5004) );
  INV_X1 U6088 ( .A(n4918), .ZN(n4919) );
  OR2_X1 U6089 ( .A1(n4413), .A2(n4919), .ZN(n4935) );
  NOR2_X1 U6090 ( .A1(n5208), .A2(REIP_REG_1__SCAN_IN), .ZN(n4970) );
  AOI21_X1 U6091 ( .B1(n5893), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4970), 
        .ZN(n4920) );
  OAI21_X1 U6092 ( .B1(n5897), .B2(n4921), .A(n4920), .ZN(n4922) );
  AOI21_X1 U6093 ( .B1(n5891), .B2(n4556), .A(n4922), .ZN(n4923) );
  OAI21_X1 U6094 ( .B1(n4496), .B2(n4935), .A(n4923), .ZN(n4925) );
  NOR2_X1 U6095 ( .A1(n5903), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4924)
         );
  AOI211_X1 U6096 ( .C1(n4971), .C2(REIP_REG_1__SCAN_IN), .A(n4925), .B(n4924), 
        .ZN(n4926) );
  OAI21_X1 U6097 ( .B1(n5004), .B2(n4927), .A(n4926), .ZN(U2826) );
  OAI21_X1 U6098 ( .B1(n4862), .B2(n4930), .A(n4929), .ZN(n5979) );
  OR2_X1 U6099 ( .A1(n4931), .A2(n4932), .ZN(n4933) );
  AND2_X1 U6100 ( .A1(n5097), .A2(n4933), .ZN(n6048) );
  AOI22_X1 U6101 ( .A1(n5923), .A2(n6048), .B1(n5313), .B2(EBX_REG_11__SCAN_IN), .ZN(n4934) );
  OAI21_X1 U6102 ( .B1(n5979), .B2(n5316), .A(n4934), .ZN(U2848) );
  INV_X1 U6103 ( .A(n4935), .ZN(n5014) );
  OAI22_X1 U6104 ( .A1(n5897), .A2(n4258), .B1(n4936), .B2(n5916), .ZN(n4938)
         );
  NOR2_X1 U6105 ( .A1(n5881), .A2(n6575), .ZN(n4937) );
  AOI211_X1 U6106 ( .C1(n6337), .C2(n5014), .A(n4938), .B(n4937), .ZN(n4940)
         );
  OAI21_X1 U6107 ( .B1(n5892), .B2(n5893), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4939) );
  OAI211_X1 U6108 ( .C1(n5004), .C2(n4941), .A(n4940), .B(n4939), .ZN(U2827)
         );
  OAI21_X1 U6109 ( .B1(n4971), .B2(n4972), .A(n5859), .ZN(n4979) );
  NOR2_X1 U6110 ( .A1(n4979), .A2(n6765), .ZN(n4945) );
  INV_X1 U6111 ( .A(n5758), .ZN(n4942) );
  AOI22_X1 U6112 ( .A1(n4942), .A2(n5014), .B1(n5893), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4943) );
  INV_X1 U6113 ( .A(n5907), .ZN(n5894) );
  OAI211_X1 U6114 ( .C1(n5897), .C2(n6743), .A(n4943), .B(n5894), .ZN(n4944)
         );
  AOI211_X1 U6115 ( .C1(n5892), .C2(n6021), .A(n4945), .B(n4944), .ZN(n4948)
         );
  AOI22_X1 U6116 ( .A1(n4946), .A2(n6765), .B1(n6082), .B2(n5891), .ZN(n4947)
         );
  OAI211_X1 U6117 ( .C1(n5004), .C2(n6025), .A(n4948), .B(n4947), .ZN(U2823)
         );
  INV_X1 U6118 ( .A(n6254), .ZN(n4949) );
  NOR2_X1 U6119 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4950), .ZN(n5001)
         );
  NAND2_X1 U6120 ( .A1(n6364), .A2(n5001), .ZN(n4964) );
  INV_X1 U6121 ( .A(n6155), .ZN(n6185) );
  OR2_X1 U6122 ( .A1(n6185), .A2(n6293), .ZN(n4955) );
  INV_X1 U6123 ( .A(n4951), .ZN(n4953) );
  NAND2_X1 U6124 ( .A1(n4953), .A2(n4952), .ZN(n6291) );
  OR2_X1 U6125 ( .A1(n6300), .A2(n6291), .ZN(n4954) );
  INV_X1 U6126 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4961) );
  AOI21_X1 U6127 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6291), .A(n4610), .ZN(
        n6302) );
  INV_X1 U6128 ( .A(n5001), .ZN(n4959) );
  INV_X1 U6129 ( .A(n5168), .ZN(n4956) );
  AOI21_X1 U6130 ( .B1(n4956), .B2(n6375), .A(n6523), .ZN(n4957) );
  AOI211_X1 U6131 ( .C1(n6155), .C2(n6182), .A(n4957), .B(n6340), .ZN(n4958)
         );
  AOI211_X1 U6132 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4959), .A(n4958), .B(
        n6290), .ZN(n4960) );
  NAND2_X1 U6133 ( .A1(n6302), .A2(n4960), .ZN(n4998) );
  INV_X1 U6134 ( .A(n4998), .ZN(n4965) );
  OAI22_X1 U6135 ( .A1(n5003), .A2(n5536), .B1(n4961), .B2(n4965), .ZN(n4962)
         );
  AOI21_X1 U6136 ( .B1(n5168), .B2(n6311), .A(n4962), .ZN(n4963) );
  OAI211_X1 U6137 ( .C1(n6375), .C2(n6314), .A(n4964), .B(n4963), .ZN(U3119)
         );
  NAND2_X1 U6138 ( .A1(n6391), .A2(n5001), .ZN(n4969) );
  INV_X1 U6139 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4966) );
  OAI22_X1 U6140 ( .A1(n5003), .A2(n5555), .B1(n4966), .B2(n4965), .ZN(n4967)
         );
  AOI21_X1 U6141 ( .B1(n5168), .B2(n6389), .A(n4967), .ZN(n4968) );
  OAI211_X1 U6142 ( .C1(n6375), .C2(n6397), .A(n4969), .B(n4968), .ZN(U3123)
         );
  INV_X1 U6143 ( .A(EAX_REG_11__SCAN_IN), .ZN(n5947) );
  INV_X1 U6144 ( .A(DATAI_11_), .ZN(n6690) );
  OAI222_X1 U6145 ( .A1(n5652), .A2(n5979), .B1(n5317), .B2(n5947), .C1(n6690), 
        .C2(n5089), .ZN(U2880) );
  INV_X1 U6146 ( .A(n6035), .ZN(n4981) );
  INV_X1 U6147 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6464) );
  INV_X1 U6148 ( .A(REIP_REG_2__SCAN_IN), .ZN(n5010) );
  NOR3_X1 U6149 ( .A1(n4971), .A2(n4970), .A3(n5010), .ZN(n5008) );
  NAND3_X1 U6150 ( .A1(n5008), .A2(n5207), .A3(n4972), .ZN(n4978) );
  NOR2_X1 U6151 ( .A1(n6087), .A2(n5916), .ZN(n4976) );
  INV_X1 U6152 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4973) );
  OAI22_X1 U6153 ( .A1(n5897), .A2(n4974), .B1(n4973), .B2(n5904), .ZN(n4975)
         );
  AOI211_X1 U6154 ( .C1(n3113), .C2(n5014), .A(n4976), .B(n4975), .ZN(n4977)
         );
  OAI211_X1 U6155 ( .C1(n6464), .C2(n4979), .A(n4978), .B(n4977), .ZN(n4980)
         );
  AOI21_X1 U6156 ( .B1(n5892), .B2(n4981), .A(n4980), .ZN(n4982) );
  OAI21_X1 U6157 ( .B1(n5004), .B2(n6031), .A(n4982), .ZN(U2824) );
  AOI22_X1 U6158 ( .A1(n5168), .A2(n6377), .B1(INSTQUEUE_REG_12__5__SCAN_IN), 
        .B2(n4998), .ZN(n4983) );
  OAI21_X1 U6159 ( .B1(n6537), .B2(n6375), .A(n4983), .ZN(n4984) );
  AOI21_X1 U6160 ( .B1(n6378), .B2(n5001), .A(n4984), .ZN(n4985) );
  OAI21_X1 U6161 ( .B1(n6539), .B2(n5003), .A(n4985), .ZN(U3121) );
  AOI22_X1 U6162 ( .A1(n5168), .A2(n6331), .B1(INSTQUEUE_REG_12__0__SCAN_IN), 
        .B2(n4998), .ZN(n4986) );
  OAI21_X1 U6163 ( .B1(n6350), .B2(n6375), .A(n4986), .ZN(n4987) );
  AOI21_X1 U6164 ( .B1(n6332), .B2(n5001), .A(n4987), .ZN(n4988) );
  OAI21_X1 U6165 ( .B1(n5526), .B2(n5003), .A(n4988), .ZN(U3116) );
  INV_X1 U6166 ( .A(n6356), .ZN(n6305) );
  AOI22_X1 U6167 ( .A1(n5168), .A2(n6305), .B1(INSTQUEUE_REG_12__1__SCAN_IN), 
        .B2(n4998), .ZN(n4989) );
  OAI21_X1 U6168 ( .B1(n6308), .B2(n6375), .A(n4989), .ZN(n4990) );
  AOI21_X1 U6169 ( .B1(n6352), .B2(n5001), .A(n4990), .ZN(n4991) );
  OAI21_X1 U6170 ( .B1(n5530), .B2(n5003), .A(n4991), .ZN(U3117) );
  AOI22_X1 U6171 ( .A1(n5168), .A2(n6315), .B1(INSTQUEUE_REG_12__4__SCAN_IN), 
        .B2(n4998), .ZN(n4992) );
  OAI21_X1 U6172 ( .B1(n6318), .B2(n6375), .A(n4992), .ZN(n4993) );
  AOI21_X1 U6173 ( .B1(n6371), .B2(n5001), .A(n4993), .ZN(n4994) );
  OAI21_X1 U6174 ( .B1(n5543), .B2(n5003), .A(n4994), .ZN(U3120) );
  AOI22_X1 U6175 ( .A1(n5168), .A2(n6382), .B1(INSTQUEUE_REG_12__6__SCAN_IN), 
        .B2(n4998), .ZN(n4995) );
  OAI21_X1 U6176 ( .B1(n6387), .B2(n6375), .A(n4995), .ZN(n4996) );
  AOI21_X1 U6177 ( .B1(n6383), .B2(n5001), .A(n4996), .ZN(n4997) );
  OAI21_X1 U6178 ( .B1(n5551), .B2(n5003), .A(n4997), .ZN(U3122) );
  AOI22_X1 U6179 ( .A1(n5168), .A2(n6357), .B1(INSTQUEUE_REG_12__2__SCAN_IN), 
        .B2(n4998), .ZN(n4999) );
  OAI21_X1 U6180 ( .B1(n6362), .B2(n6375), .A(n4999), .ZN(n5000) );
  AOI21_X1 U6181 ( .B1(n6358), .B2(n5001), .A(n5000), .ZN(n5002) );
  OAI21_X1 U6182 ( .B1(n5534), .B2(n5003), .A(n5002), .ZN(U3118) );
  INV_X1 U6183 ( .A(n5004), .ZN(n5912) );
  NAND2_X1 U6184 ( .A1(n5912), .A2(n6042), .ZN(n5016) );
  INV_X1 U6185 ( .A(n3122), .ZN(n5013) );
  NOR2_X1 U6186 ( .A1(n5904), .A2(n6822), .ZN(n5005) );
  AOI21_X1 U6187 ( .B1(n5908), .B2(EBX_REG_2__SCAN_IN), .A(n5005), .ZN(n5006)
         );
  OAI21_X1 U6188 ( .B1(n5007), .B2(n5916), .A(n5006), .ZN(n5012) );
  AOI21_X1 U6189 ( .B1(n5010), .B2(n5009), .A(n5008), .ZN(n5011) );
  AOI211_X1 U6190 ( .C1(n5014), .C2(n5013), .A(n5012), .B(n5011), .ZN(n5015)
         );
  OAI211_X1 U6191 ( .C1(n6046), .C2(n5903), .A(n5016), .B(n5015), .ZN(U2825)
         );
  AOI21_X1 U6192 ( .B1(n4929), .B2(n5017), .A(n3849), .ZN(n5918) );
  INV_X1 U6193 ( .A(n5918), .ZN(n5019) );
  AOI22_X1 U6194 ( .A1(n5335), .A2(DATAI_12_), .B1(n5931), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n5018) );
  OAI21_X1 U6195 ( .B1(n5019), .B2(n5652), .A(n5018), .ZN(U2879) );
  NAND2_X1 U6196 ( .A1(n5972), .A2(n5020), .ZN(n5022) );
  XOR2_X1 U6197 ( .A(n5022), .B(n5021), .Z(n5043) );
  NAND2_X1 U6198 ( .A1(n6022), .A2(n5860), .ZN(n5023) );
  NAND2_X1 U6199 ( .A1(n4228), .A2(REIP_REG_10__SCAN_IN), .ZN(n5039) );
  OAI211_X1 U6200 ( .C1(n5393), .C2(n5024), .A(n5023), .B(n5039), .ZN(n5025)
         );
  AOI21_X1 U6201 ( .B1(n5921), .B2(n4663), .A(n5025), .ZN(n5026) );
  OAI21_X1 U6202 ( .B1(n5043), .B2(n5773), .A(n5026), .ZN(U2976) );
  INV_X1 U6203 ( .A(n5027), .ZN(n5030) );
  OAI21_X1 U6204 ( .B1(n5029), .B2(n5028), .A(n6095), .ZN(n6076) );
  NAND2_X1 U6205 ( .A1(n6096), .A2(n6076), .ZN(n6094) );
  NOR2_X1 U6206 ( .A1(n5030), .A2(n6094), .ZN(n6068) );
  NAND2_X1 U6207 ( .A1(n6061), .A2(n6068), .ZN(n6059) );
  AOI21_X1 U6208 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6059), .ZN(n5033) );
  OAI21_X1 U6209 ( .B1(n6096), .B2(n6095), .A(n6104), .ZN(n6091) );
  OAI22_X1 U6210 ( .A1(n5031), .A2(n5493), .B1(n5030), .B2(n6091), .ZN(n6071)
         );
  OAI21_X1 U6211 ( .B1(n5032), .B2(n6061), .A(n6071), .ZN(n6056) );
  AOI222_X1 U6212 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n5033), .B1(
        INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6056), .C1(n5033), .C2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5042) );
  INV_X1 U6213 ( .A(n5034), .ZN(n5035) );
  NAND2_X1 U6214 ( .A1(n5036), .A2(n5035), .ZN(n5037) );
  AOI21_X1 U6215 ( .B1(n5038), .B2(n5037), .A(n4931), .ZN(n5920) );
  INV_X1 U6216 ( .A(n5039), .ZN(n5040) );
  AOI21_X1 U6217 ( .B1(n6099), .B2(n5920), .A(n5040), .ZN(n5041) );
  OAI211_X1 U6218 ( .C1(n5043), .C2(n6103), .A(n5042), .B(n5041), .ZN(U3008)
         );
  OR2_X1 U6219 ( .A1(n3707), .A2(n3113), .ZN(n6120) );
  OR2_X1 U6220 ( .A1(n6120), .A2(n6297), .ZN(n5045) );
  NOR2_X1 U6221 ( .A1(n6183), .A2(n5051), .ZN(n5080) );
  INV_X1 U6222 ( .A(n5080), .ZN(n5044) );
  AND2_X1 U6223 ( .A1(n5045), .A2(n5044), .ZN(n5053) );
  OR2_X1 U6224 ( .A1(n5050), .A2(n5053), .ZN(n5048) );
  INV_X1 U6225 ( .A(n5051), .ZN(n5046) );
  NAND2_X1 U6226 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5046), .ZN(n5047) );
  INV_X1 U6227 ( .A(n5050), .ZN(n5052) );
  AOI22_X1 U6228 ( .A1(n5053), .A2(n5052), .B1(n5051), .B2(n6340), .ZN(n5054)
         );
  NAND2_X1 U6229 ( .A1(n6342), .A2(n5054), .ZN(n5076) );
  AOI22_X1 U6230 ( .A1(n5520), .A2(n6315), .B1(INSTQUEUE_REG_1__4__SCAN_IN), 
        .B2(n5076), .ZN(n5055) );
  OAI21_X1 U6231 ( .B1(n6318), .B2(n5078), .A(n5055), .ZN(n5056) );
  AOI21_X1 U6232 ( .B1(n6371), .B2(n5080), .A(n5056), .ZN(n5057) );
  OAI21_X1 U6233 ( .B1(n5543), .B2(n5082), .A(n5057), .ZN(U3032) );
  AOI22_X1 U6234 ( .A1(n5520), .A2(n6305), .B1(INSTQUEUE_REG_1__1__SCAN_IN), 
        .B2(n5076), .ZN(n5058) );
  OAI21_X1 U6235 ( .B1(n6308), .B2(n5078), .A(n5058), .ZN(n5059) );
  AOI21_X1 U6236 ( .B1(n6352), .B2(n5080), .A(n5059), .ZN(n5060) );
  OAI21_X1 U6237 ( .B1(n5530), .B2(n5082), .A(n5060), .ZN(U3029) );
  AOI22_X1 U6238 ( .A1(n5520), .A2(n6382), .B1(INSTQUEUE_REG_1__6__SCAN_IN), 
        .B2(n5076), .ZN(n5061) );
  OAI21_X1 U6239 ( .B1(n6387), .B2(n5078), .A(n5061), .ZN(n5062) );
  AOI21_X1 U6240 ( .B1(n6383), .B2(n5080), .A(n5062), .ZN(n5063) );
  OAI21_X1 U6241 ( .B1(n5551), .B2(n5082), .A(n5063), .ZN(U3034) );
  AOI22_X1 U6242 ( .A1(n5520), .A2(n6377), .B1(INSTQUEUE_REG_1__5__SCAN_IN), 
        .B2(n5076), .ZN(n5064) );
  OAI21_X1 U6243 ( .B1(n6537), .B2(n5078), .A(n5064), .ZN(n5065) );
  AOI21_X1 U6244 ( .B1(n6378), .B2(n5080), .A(n5065), .ZN(n5066) );
  OAI21_X1 U6245 ( .B1(n6539), .B2(n5082), .A(n5066), .ZN(U3033) );
  AOI22_X1 U6246 ( .A1(n5520), .A2(n6357), .B1(INSTQUEUE_REG_1__2__SCAN_IN), 
        .B2(n5076), .ZN(n5067) );
  OAI21_X1 U6247 ( .B1(n6362), .B2(n5078), .A(n5067), .ZN(n5068) );
  AOI21_X1 U6248 ( .B1(n6358), .B2(n5080), .A(n5068), .ZN(n5069) );
  OAI21_X1 U6249 ( .B1(n5534), .B2(n5082), .A(n5069), .ZN(U3030) );
  AOI22_X1 U6250 ( .A1(n5520), .A2(n6331), .B1(INSTQUEUE_REG_1__0__SCAN_IN), 
        .B2(n5076), .ZN(n5070) );
  OAI21_X1 U6251 ( .B1(n6350), .B2(n5078), .A(n5070), .ZN(n5071) );
  AOI21_X1 U6252 ( .B1(n6332), .B2(n5080), .A(n5071), .ZN(n5072) );
  OAI21_X1 U6253 ( .B1(n5526), .B2(n5082), .A(n5072), .ZN(U3028) );
  AOI22_X1 U6254 ( .A1(n5520), .A2(n6311), .B1(INSTQUEUE_REG_1__3__SCAN_IN), 
        .B2(n5076), .ZN(n5073) );
  OAI21_X1 U6255 ( .B1(n6314), .B2(n5078), .A(n5073), .ZN(n5074) );
  AOI21_X1 U6256 ( .B1(n6364), .B2(n5080), .A(n5074), .ZN(n5075) );
  OAI21_X1 U6257 ( .B1(n5082), .B2(n5536), .A(n5075), .ZN(U3031) );
  AOI22_X1 U6258 ( .A1(n5520), .A2(n6389), .B1(INSTQUEUE_REG_1__7__SCAN_IN), 
        .B2(n5076), .ZN(n5077) );
  OAI21_X1 U6259 ( .B1(n6397), .B2(n5078), .A(n5077), .ZN(n5079) );
  AOI21_X1 U6260 ( .B1(n6391), .B2(n5080), .A(n5079), .ZN(n5081) );
  OAI21_X1 U6261 ( .B1(n5082), .B2(n5555), .A(n5081), .ZN(U3035) );
  OR2_X1 U6262 ( .A1(n5084), .A2(n5083), .ZN(n5086) );
  NAND2_X1 U6263 ( .A1(n5086), .A2(n5085), .ZN(n5833) );
  NAND2_X1 U6264 ( .A1(n5099), .A2(n5087), .ZN(n5088) );
  NAND2_X1 U6265 ( .A1(n5114), .A2(n5088), .ZN(n5837) );
  OAI222_X1 U6266 ( .A1(n5833), .A2(n5316), .B1(n5927), .B2(n4295), .C1(n5837), 
        .C2(n5301), .ZN(U2846) );
  INV_X1 U6267 ( .A(DATAI_13_), .ZN(n6785) );
  OAI222_X1 U6268 ( .A1(n5833), .A2(n5652), .B1(n5089), .B2(n6785), .C1(n5317), 
        .C2(n3836), .ZN(U2878) );
  NOR2_X1 U6269 ( .A1(n5091), .A2(n3140), .ZN(n5092) );
  XNOR2_X1 U6270 ( .A(n5090), .B(n5092), .ZN(n5110) );
  NAND2_X1 U6271 ( .A1(n6022), .A2(n5845), .ZN(n5093) );
  NAND2_X1 U6272 ( .A1(n4228), .A2(REIP_REG_12__SCAN_IN), .ZN(n5100) );
  OAI211_X1 U6273 ( .C1(n5393), .C2(n5843), .A(n5093), .B(n5100), .ZN(n5094)
         );
  AOI21_X1 U6274 ( .B1(n5918), .B2(n5700), .A(n5094), .ZN(n5095) );
  OAI21_X1 U6275 ( .B1(n5110), .B2(n5773), .A(n5095), .ZN(U2974) );
  NAND2_X1 U6276 ( .A1(n5097), .A2(n5096), .ZN(n5098) );
  AND2_X1 U6277 ( .A1(n5099), .A2(n5098), .ZN(n5917) );
  INV_X1 U6278 ( .A(n5100), .ZN(n5101) );
  AOI21_X1 U6279 ( .B1(n6099), .B2(n5917), .A(n5101), .ZN(n5109) );
  INV_X1 U6280 ( .A(n5506), .ZN(n5502) );
  AOI21_X1 U6281 ( .B1(n6095), .B2(n5484), .A(n5502), .ZN(n5107) );
  OAI22_X1 U6282 ( .A1(n5104), .A2(n5103), .B1(n5480), .B2(n5102), .ZN(n6047)
         );
  INV_X1 U6283 ( .A(n5752), .ZN(n6053) );
  INV_X1 U6284 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6052) );
  OAI21_X1 U6285 ( .B1(n6053), .B2(n6052), .A(n5105), .ZN(n5106) );
  OAI21_X1 U6286 ( .B1(n5107), .B2(n6047), .A(n5106), .ZN(n5108) );
  OAI211_X1 U6287 ( .C1(n5110), .C2(n6103), .A(n5109), .B(n5108), .ZN(U3006)
         );
  OAI21_X1 U6288 ( .B1(n5113), .B2(n5112), .A(n5111), .ZN(n5831) );
  AOI21_X1 U6289 ( .B1(n5115), .B2(n5114), .A(n5310), .ZN(n5823) );
  AOI22_X1 U6290 ( .A1(n5923), .A2(n5823), .B1(n5313), .B2(EBX_REG_14__SCAN_IN), .ZN(n5116) );
  OAI21_X1 U6291 ( .B1(n5831), .B2(n5316), .A(n5116), .ZN(U2845) );
  AOI22_X1 U6292 ( .A1(n5335), .A2(DATAI_14_), .B1(n5931), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5117) );
  OAI21_X1 U6293 ( .B1(n5831), .B2(n5652), .A(n5117), .ZN(U2877) );
  AOI21_X1 U6294 ( .B1(n5120), .B2(n5118), .A(n5124), .ZN(n5126) );
  NOR3_X1 U6295 ( .A1(n6426), .A2(n4435), .A3(n5119), .ZN(n5122) );
  NOR3_X1 U6296 ( .A1(n5120), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n6431), 
        .ZN(n5121) );
  AOI211_X1 U6297 ( .C1(n6400), .C2(n5123), .A(n5122), .B(n5121), .ZN(n5125)
         );
  OAI22_X1 U6298 ( .A1(n5126), .A2(n3143), .B1(n5125), .B2(n5124), .ZN(U3459)
         );
  NAND2_X1 U6299 ( .A1(n5966), .A2(DATAI_1_), .ZN(n5135) );
  NAND2_X1 U6300 ( .A1(n5968), .A2(UWORD_REG_1__SCAN_IN), .ZN(n5127) );
  OAI211_X1 U6301 ( .C1(n5128), .C2(n5163), .A(n5135), .B(n5127), .ZN(U2925)
         );
  NAND2_X1 U6302 ( .A1(n5966), .A2(DATAI_3_), .ZN(n5149) );
  NAND2_X1 U6303 ( .A1(n5968), .A2(UWORD_REG_3__SCAN_IN), .ZN(n5129) );
  OAI211_X1 U6304 ( .C1(n5130), .C2(n5163), .A(n5149), .B(n5129), .ZN(U2927)
         );
  NAND2_X1 U6305 ( .A1(n5966), .A2(DATAI_5_), .ZN(n5137) );
  NAND2_X1 U6306 ( .A1(n5968), .A2(UWORD_REG_5__SCAN_IN), .ZN(n5131) );
  OAI211_X1 U6307 ( .C1(n6622), .C2(n5163), .A(n5137), .B(n5131), .ZN(U2929)
         );
  NAND2_X1 U6308 ( .A1(n5966), .A2(DATAI_10_), .ZN(n5145) );
  NAND2_X1 U6309 ( .A1(n5968), .A2(UWORD_REG_10__SCAN_IN), .ZN(n5132) );
  OAI211_X1 U6310 ( .C1(n6751), .C2(n5163), .A(n5145), .B(n5132), .ZN(U2934)
         );
  NAND2_X1 U6311 ( .A1(n5966), .A2(DATAI_14_), .ZN(n5143) );
  NAND2_X1 U6312 ( .A1(n5968), .A2(UWORD_REG_14__SCAN_IN), .ZN(n5133) );
  OAI211_X1 U6313 ( .C1(n6707), .C2(n5163), .A(n5143), .B(n5133), .ZN(U2938)
         );
  NAND2_X1 U6314 ( .A1(n5968), .A2(LWORD_REG_1__SCAN_IN), .ZN(n5134) );
  OAI211_X1 U6315 ( .C1(n3702), .C2(n5163), .A(n5135), .B(n5134), .ZN(U2940)
         );
  NAND2_X1 U6316 ( .A1(n5968), .A2(LWORD_REG_5__SCAN_IN), .ZN(n5136) );
  OAI211_X1 U6317 ( .C1(n3733), .C2(n5163), .A(n5137), .B(n5136), .ZN(U2944)
         );
  NAND2_X1 U6318 ( .A1(n5968), .A2(LWORD_REG_8__SCAN_IN), .ZN(n5138) );
  OAI211_X1 U6319 ( .C1(n3776), .C2(n5163), .A(n5139), .B(n5138), .ZN(U2947)
         );
  INV_X1 U6320 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U6321 ( .A1(n5968), .A2(LWORD_REG_12__SCAN_IN), .ZN(n5140) );
  OAI211_X1 U6322 ( .C1(n5946), .C2(n5163), .A(n5141), .B(n5140), .ZN(U2951)
         );
  INV_X1 U6323 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6686) );
  NAND2_X1 U6324 ( .A1(n5968), .A2(LWORD_REG_14__SCAN_IN), .ZN(n5142) );
  OAI211_X1 U6325 ( .C1(n6686), .C2(n5163), .A(n5143), .B(n5142), .ZN(U2953)
         );
  INV_X1 U6326 ( .A(EAX_REG_10__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U6327 ( .A1(n5968), .A2(LWORD_REG_10__SCAN_IN), .ZN(n5144) );
  OAI211_X1 U6328 ( .C1(n5949), .C2(n5163), .A(n5145), .B(n5144), .ZN(U2949)
         );
  NAND2_X1 U6329 ( .A1(n5968), .A2(LWORD_REG_7__SCAN_IN), .ZN(n5146) );
  OAI211_X1 U6330 ( .C1(n4823), .C2(n5163), .A(n5147), .B(n5146), .ZN(U2946)
         );
  NAND2_X1 U6331 ( .A1(n5968), .A2(LWORD_REG_3__SCAN_IN), .ZN(n5148) );
  OAI211_X1 U6332 ( .C1(n4700), .C2(n5163), .A(n5149), .B(n5148), .ZN(U2942)
         );
  NAND2_X1 U6333 ( .A1(n5966), .A2(DATAI_0_), .ZN(n5162) );
  NAND2_X1 U6334 ( .A1(n5968), .A2(LWORD_REG_0__SCAN_IN), .ZN(n5150) );
  OAI211_X1 U6335 ( .C1(n3710), .C2(n5163), .A(n5162), .B(n5150), .ZN(U2939)
         );
  NAND2_X1 U6336 ( .A1(n5968), .A2(UWORD_REG_11__SCAN_IN), .ZN(n5151) );
  OAI211_X1 U6337 ( .C1(n5153), .C2(n5163), .A(n5152), .B(n5151), .ZN(U2935)
         );
  NAND2_X1 U6338 ( .A1(n5968), .A2(UWORD_REG_6__SCAN_IN), .ZN(n5154) );
  OAI211_X1 U6339 ( .C1(n6559), .C2(n5163), .A(n5155), .B(n5154), .ZN(U2930)
         );
  NAND2_X1 U6340 ( .A1(n5968), .A2(UWORD_REG_4__SCAN_IN), .ZN(n5156) );
  OAI211_X1 U6341 ( .C1(n3952), .C2(n5163), .A(n5157), .B(n5156), .ZN(U2928)
         );
  NAND2_X1 U6342 ( .A1(n5968), .A2(UWORD_REG_2__SCAN_IN), .ZN(n5158) );
  OAI211_X1 U6343 ( .C1(n5160), .C2(n5163), .A(n5159), .B(n5158), .ZN(U2926)
         );
  NAND2_X1 U6344 ( .A1(n5968), .A2(UWORD_REG_0__SCAN_IN), .ZN(n5161) );
  OAI211_X1 U6345 ( .C1(n5164), .C2(n5163), .A(n5162), .B(n5161), .ZN(U2924)
         );
  AOI22_X1 U6346 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n5166), .B1(n6353), 
        .B2(n5165), .ZN(n5170) );
  INV_X1 U6347 ( .A(n6308), .ZN(n6351) );
  AOI22_X1 U6348 ( .A1(n6351), .A2(n5168), .B1(n5167), .B2(n6305), .ZN(n5169)
         );
  OAI211_X1 U6349 ( .C1(n5177), .C2(n5171), .A(n5170), .B(n5169), .ZN(U3125)
         );
  AOI22_X1 U6350 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n5173), .B1(n6353), 
        .B2(n5172), .ZN(n5176) );
  AOI22_X1 U6351 ( .A1(n6325), .A2(n6351), .B1(n5174), .B2(n6305), .ZN(n5175)
         );
  OAI211_X1 U6352 ( .C1(n5178), .C2(n5177), .A(n5176), .B(n5175), .ZN(U3093)
         );
  INV_X1 U6353 ( .A(n4354), .ZN(n5180) );
  AOI21_X1 U6354 ( .B1(n5182), .B2(n5180), .A(n5179), .ZN(n5185) );
  AOI21_X1 U6355 ( .B1(n4354), .B2(n5282), .A(n5181), .ZN(n5183) );
  AOI22_X1 U6356 ( .A1(n5185), .A2(n5184), .B1(n5183), .B2(n5182), .ZN(n5566)
         );
  AOI22_X1 U6357 ( .A1(n5566), .A2(n5923), .B1(EBX_REG_30__SCAN_IN), .B2(n5313), .ZN(n5186) );
  OAI21_X1 U6358 ( .B1(n4364), .B2(n5316), .A(n5186), .ZN(U2829) );
  AOI211_X1 U6359 ( .C1(n6523), .C2(n6154), .A(n6117), .B(n5187), .ZN(n5188)
         );
  AOI21_X1 U6360 ( .B1(n5189), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n5188), 
        .ZN(n5190) );
  OAI21_X1 U6361 ( .B1(n4496), .B2(n5191), .A(n5190), .ZN(U3464) );
  INV_X1 U6362 ( .A(n4219), .ZN(n5192) );
  NOR2_X1 U6363 ( .A1(n5193), .A2(n5192), .ZN(n5200) );
  NAND2_X1 U6364 ( .A1(n5195), .A2(n5194), .ZN(n5199) );
  INV_X1 U6365 ( .A(n5196), .ZN(n5197) );
  NAND2_X1 U6366 ( .A1(n5204), .A2(n5197), .ZN(n5198) );
  OAI211_X1 U6367 ( .C1(n5204), .C2(n5200), .A(n5199), .B(n5198), .ZN(n6418)
         );
  NAND2_X1 U6368 ( .A1(n5201), .A2(n4219), .ZN(n5202) );
  OAI21_X1 U6369 ( .B1(n5204), .B2(n3108), .A(n5202), .ZN(n5766) );
  AOI21_X1 U6370 ( .B1(n5205), .B2(n6452), .A(READY_N), .ZN(n6527) );
  NOR2_X1 U6371 ( .A1(n5766), .A2(n6527), .ZN(n6414) );
  OR2_X1 U6372 ( .A1(n6414), .A2(n6434), .ZN(n5772) );
  MUX2_X1 U6373 ( .A(n6418), .B(MORE_REG_SCAN_IN), .S(n5772), .Z(U3471) );
  INV_X1 U6374 ( .A(REIP_REG_31__SCAN_IN), .ZN(n5217) );
  INV_X1 U6375 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6498) );
  AOI21_X1 U6376 ( .B1(n5207), .B2(n6498), .A(n5206), .ZN(n5562) );
  OAI21_X1 U6377 ( .B1(REIP_REG_30__SCAN_IN), .B2(n5208), .A(n5562), .ZN(n5209) );
  INV_X1 U6378 ( .A(n5209), .ZN(n5216) );
  OAI22_X1 U6379 ( .A1(n5212), .A2(n5211), .B1(n5210), .B2(n5904), .ZN(n5213)
         );
  INV_X1 U6380 ( .A(n5213), .ZN(n5215) );
  INV_X1 U6381 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5218) );
  OAI22_X1 U6382 ( .A1(n5219), .A2(n5301), .B1(n5927), .B2(n5218), .ZN(U2828)
         );
  INV_X1 U6383 ( .A(n5221), .ZN(n5222) );
  OAI222_X1 U6384 ( .A1(n5220), .A2(n5316), .B1(n5223), .B2(n5927), .C1(n5301), 
        .C2(n5222), .ZN(U2830) );
  OR2_X1 U6385 ( .A1(n5229), .A2(n5224), .ZN(n5225) );
  NAND2_X1 U6386 ( .A1(n4354), .A2(n5225), .ZN(n5576) );
  INV_X1 U6387 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5569) );
  OAI22_X1 U6388 ( .A1(n5576), .A2(n5301), .B1(n5569), .B2(n5927), .ZN(n5226)
         );
  AOI21_X1 U6389 ( .B1(n5653), .B2(n5924), .A(n5226), .ZN(n5227) );
  INV_X1 U6390 ( .A(n5227), .ZN(U2831) );
  INV_X1 U6391 ( .A(n5228), .ZN(n5231) );
  INV_X1 U6392 ( .A(n5238), .ZN(n5230) );
  AOI21_X1 U6393 ( .B1(n5231), .B2(n5230), .A(n5229), .ZN(n5581) );
  AOI22_X1 U6394 ( .A1(n5581), .A2(n5923), .B1(EBX_REG_27__SCAN_IN), .B2(n5313), .ZN(n5232) );
  OAI21_X1 U6395 ( .B1(n5584), .B2(n5316), .A(n5232), .ZN(U2832) );
  NAND2_X1 U6397 ( .A1(n5234), .A2(n5235), .ZN(n5236) );
  AND2_X1 U6398 ( .A1(n4190), .A2(n5236), .ZN(n5656) );
  AND2_X1 U6399 ( .A1(n5252), .A2(n5237), .ZN(n5239) );
  OR2_X1 U6400 ( .A1(n5239), .A2(n5238), .ZN(n5585) );
  OAI22_X1 U6401 ( .A1(n5585), .A2(n5301), .B1(n5240), .B2(n5927), .ZN(n5241)
         );
  AOI21_X1 U6402 ( .B1(n5656), .B2(n5924), .A(n5241), .ZN(n5242) );
  INV_X1 U6403 ( .A(n5242), .ZN(U2833) );
  INV_X1 U6405 ( .A(n5255), .ZN(n5245) );
  AND2_X1 U6406 ( .A1(n5244), .A2(n5245), .ZN(n5248) );
  INV_X1 U6407 ( .A(n5246), .ZN(n5247) );
  OAI21_X1 U6408 ( .B1(n5248), .B2(n5247), .A(n5234), .ZN(n5679) );
  NAND2_X1 U6409 ( .A1(n5250), .A2(n5249), .ZN(n5251) );
  NAND2_X1 U6410 ( .A1(n5252), .A2(n5251), .ZN(n5592) );
  OAI22_X1 U6411 ( .A1(n5592), .A2(n5301), .B1(n6607), .B2(n5927), .ZN(n5253)
         );
  INV_X1 U6412 ( .A(n5253), .ZN(n5254) );
  OAI21_X1 U6413 ( .B1(n5679), .B2(n5316), .A(n5254), .ZN(U2834) );
  XNOR2_X1 U6414 ( .A(n5244), .B(n5255), .ZN(n5659) );
  INV_X1 U6415 ( .A(n5659), .ZN(n5258) );
  XOR2_X1 U6416 ( .A(n5256), .B(n5449), .Z(n5602) );
  AOI22_X1 U6417 ( .A1(n5602), .A2(n5923), .B1(EBX_REG_24__SCAN_IN), .B2(n5313), .ZN(n5257) );
  OAI21_X1 U6418 ( .B1(n5258), .B2(n5316), .A(n5257), .ZN(U2835) );
  INV_X1 U6419 ( .A(n5259), .ZN(n5264) );
  INV_X1 U6420 ( .A(n5261), .ZN(n5263) );
  INV_X1 U6421 ( .A(n5262), .ZN(n5358) );
  AND2_X1 U6422 ( .A1(n3124), .A2(n5265), .ZN(n5266) );
  OR2_X1 U6423 ( .A1(n5266), .A2(n5448), .ZN(n5619) );
  OAI22_X1 U6424 ( .A1(n5619), .A2(n5301), .B1(n5267), .B2(n5927), .ZN(n5268)
         );
  INV_X1 U6425 ( .A(n5268), .ZN(n5269) );
  OAI21_X1 U6426 ( .B1(n5625), .B2(n5316), .A(n5269), .ZN(U2837) );
  INV_X1 U6427 ( .A(n5270), .ZN(n5284) );
  MUX2_X1 U6428 ( .A(n5282), .B(n5284), .S(n5271), .Z(n5273) );
  XNOR2_X1 U6429 ( .A(n5273), .B(n5272), .ZN(n5635) );
  OAI21_X1 U6430 ( .B1(n5274), .B2(n5276), .A(n5275), .ZN(n5634) );
  OAI222_X1 U6431 ( .A1(n5635), .A2(n5301), .B1(n5927), .B2(n4315), .C1(n5634), 
        .C2(n5316), .ZN(U2839) );
  AND2_X1 U6432 ( .A1(n5277), .A2(n5278), .ZN(n5279) );
  OR2_X1 U6433 ( .A1(n5279), .A2(n5274), .ZN(n5684) );
  INV_X1 U6434 ( .A(n5281), .ZN(n5283) );
  MUX2_X1 U6435 ( .A(n5284), .B(n5283), .S(n5282), .Z(n5289) );
  NAND2_X1 U6436 ( .A1(n5280), .A2(n5289), .ZN(n5288) );
  XNOR2_X1 U6437 ( .A(n5288), .B(n5285), .ZN(n5716) );
  INV_X1 U6438 ( .A(n5716), .ZN(n5286) );
  OAI222_X1 U6439 ( .A1(n5684), .A2(n5316), .B1(n5287), .B2(n5927), .C1(n5301), 
        .C2(n5286), .ZN(U2840) );
  OAI21_X1 U6440 ( .B1(n5280), .B2(n5289), .A(n5288), .ZN(n5724) );
  OAI21_X1 U6441 ( .B1(n5291), .B2(n5292), .A(n5277), .ZN(n5796) );
  OAI222_X1 U6442 ( .A1(n5724), .A2(n5301), .B1(n5316), .B2(n5796), .C1(n5293), 
        .C2(n5927), .ZN(U2841) );
  INV_X1 U6443 ( .A(n5294), .ZN(n5304) );
  INV_X1 U6444 ( .A(n5295), .ZN(n5297) );
  INV_X1 U6445 ( .A(n5280), .ZN(n5296) );
  OAI21_X1 U6446 ( .B1(n5304), .B2(n5297), .A(n5296), .ZN(n5804) );
  AOI21_X1 U6447 ( .B1(n5298), .B2(n5299), .A(n5291), .ZN(n5930) );
  INV_X1 U6448 ( .A(n5930), .ZN(n5300) );
  OAI222_X1 U6449 ( .A1(n5301), .A2(n5804), .B1(n5927), .B2(n4308), .C1(n5316), 
        .C2(n5300), .ZN(U2842) );
  OAI21_X1 U6450 ( .B1(n5302), .B2(n5303), .A(n5298), .ZN(n5814) );
  AOI21_X1 U6451 ( .B1(n5305), .B2(n5312), .A(n5304), .ZN(n5809) );
  AOI22_X1 U6452 ( .A1(n5809), .A2(n5923), .B1(EBX_REG_16__SCAN_IN), .B2(n5313), .ZN(n5306) );
  OAI21_X1 U6453 ( .B1(n5814), .B2(n5316), .A(n5306), .ZN(U2843) );
  AOI21_X1 U6454 ( .B1(n5111), .B2(n5307), .A(n5302), .ZN(n5308) );
  INV_X1 U6455 ( .A(n5308), .ZN(n5822) );
  OR2_X1 U6456 ( .A1(n5310), .A2(n5309), .ZN(n5311) );
  NAND2_X1 U6457 ( .A1(n5312), .A2(n5311), .ZN(n5818) );
  INV_X1 U6458 ( .A(n5818), .ZN(n5314) );
  AOI22_X1 U6459 ( .A1(n5923), .A2(n5314), .B1(n5313), .B2(EBX_REG_15__SCAN_IN), .ZN(n5315) );
  OAI21_X1 U6460 ( .B1(n5822), .B2(n5316), .A(n5315), .ZN(U2844) );
  NAND2_X1 U6461 ( .A1(n5317), .A2(n3701), .ZN(n5319) );
  AOI22_X1 U6462 ( .A1(n5928), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n5931), .ZN(n5318) );
  OAI21_X1 U6463 ( .B1(n5320), .B2(n5319), .A(n5318), .ZN(U2860) );
  AOI22_X1 U6464 ( .A1(n5932), .A2(DATAI_13_), .B1(n5931), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U6465 ( .A1(n5928), .A2(DATAI_29_), .ZN(n5321) );
  OAI211_X1 U6466 ( .C1(n5220), .C2(n5652), .A(n5322), .B(n5321), .ZN(U2862)
         );
  AOI22_X1 U6467 ( .A1(n5932), .A2(DATAI_11_), .B1(n5931), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5324) );
  NAND2_X1 U6468 ( .A1(n5928), .A2(DATAI_27_), .ZN(n5323) );
  OAI211_X1 U6469 ( .C1(n5584), .C2(n5652), .A(n5324), .B(n5323), .ZN(U2864)
         );
  AOI22_X1 U6470 ( .A1(n5932), .A2(DATAI_9_), .B1(n5931), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5326) );
  NAND2_X1 U6471 ( .A1(n5928), .A2(DATAI_25_), .ZN(n5325) );
  OAI211_X1 U6472 ( .C1(n5679), .C2(n5652), .A(n5326), .B(n5325), .ZN(U2866)
         );
  AOI22_X1 U6473 ( .A1(n5932), .A2(DATAI_6_), .B1(n5931), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5328) );
  NAND2_X1 U6474 ( .A1(n5928), .A2(DATAI_22_), .ZN(n5327) );
  OAI211_X1 U6475 ( .C1(n5625), .C2(n5652), .A(n5328), .B(n5327), .ZN(U2869)
         );
  AOI22_X1 U6476 ( .A1(n5932), .A2(DATAI_4_), .B1(n5931), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5330) );
  NAND2_X1 U6477 ( .A1(n5928), .A2(DATAI_20_), .ZN(n5329) );
  OAI211_X1 U6478 ( .C1(n5634), .C2(n5652), .A(n5330), .B(n5329), .ZN(U2871)
         );
  AOI22_X1 U6479 ( .A1(n5932), .A2(DATAI_2_), .B1(n5931), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U6480 ( .A1(n5928), .A2(DATAI_18_), .ZN(n5331) );
  OAI211_X1 U6481 ( .C1(n5796), .C2(n5652), .A(n5332), .B(n5331), .ZN(U2873)
         );
  AOI22_X1 U6482 ( .A1(n5932), .A2(DATAI_0_), .B1(n5931), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U6483 ( .A1(n5928), .A2(DATAI_16_), .ZN(n5333) );
  OAI211_X1 U6484 ( .C1(n5814), .C2(n5652), .A(n5334), .B(n5333), .ZN(U2875)
         );
  AOI22_X1 U6485 ( .A1(n5335), .A2(DATAI_15_), .B1(n5931), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5336) );
  OAI21_X1 U6486 ( .B1(n5822), .B2(n5652), .A(n5336), .ZN(U2876) );
  NOR2_X1 U6487 ( .A1(n5338), .A2(n5337), .ZN(n5340) );
  XOR2_X1 U6488 ( .A(n5340), .B(n5339), .Z(n5431) );
  NAND2_X1 U6489 ( .A1(n4228), .A2(REIP_REG_26__SCAN_IN), .ZN(n5423) );
  NAND2_X1 U6490 ( .A1(n6036), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5341)
         );
  OAI211_X1 U6491 ( .C1(n5591), .C2(n6045), .A(n5423), .B(n5341), .ZN(n5342)
         );
  AOI21_X1 U6492 ( .B1(n5656), .B2(n4663), .A(n5342), .ZN(n5343) );
  OAI21_X1 U6493 ( .B1(n5431), .B2(n5773), .A(n5343), .ZN(U2960) );
  XNOR2_X1 U6494 ( .A(n5704), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5680)
         );
  NAND2_X1 U6495 ( .A1(n5681), .A2(n5680), .ZN(n5683) );
  OAI21_X1 U6496 ( .B1(n5704), .B2(n5722), .A(n5683), .ZN(n5384) );
  INV_X1 U6497 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5344) );
  NOR2_X1 U6498 ( .A1(n5704), .A2(n5344), .ZN(n5382) );
  NAND2_X1 U6499 ( .A1(n5704), .A2(n5344), .ZN(n5380) );
  XNOR2_X1 U6500 ( .A(n5704), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5375)
         );
  NAND2_X1 U6501 ( .A1(n5376), .A2(n5375), .ZN(n5353) );
  OAI21_X1 U6502 ( .B1(n5693), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5353), 
        .ZN(n5365) );
  MUX2_X1 U6503 ( .A(n5364), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .S(n5704), 
        .Z(n5346) );
  OAI211_X1 U6504 ( .C1(n5365), .C2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5346), .B(n5345), .ZN(n5348) );
  XNOR2_X1 U6505 ( .A(n5348), .B(n5347), .ZN(n5446) );
  NAND2_X1 U6506 ( .A1(n6022), .A2(n5600), .ZN(n5349) );
  NAND2_X1 U6507 ( .A1(n4228), .A2(REIP_REG_24__SCAN_IN), .ZN(n5440) );
  OAI211_X1 U6508 ( .C1(n5350), .C2(n5393), .A(n5349), .B(n5440), .ZN(n5351)
         );
  AOI21_X1 U6509 ( .B1(n5659), .B2(n5700), .A(n5351), .ZN(n5352) );
  OAI21_X1 U6510 ( .B1(n5446), .B2(n5773), .A(n5352), .ZN(U2962) );
  NAND2_X1 U6511 ( .A1(n5693), .A2(n5364), .ZN(n5363) );
  NAND3_X1 U6512 ( .A1(n5704), .A2(n5463), .A3(n5487), .ZN(n5354) );
  OAI22_X1 U6513 ( .A1(n5353), .A2(n5363), .B1(n5355), .B2(n5354), .ZN(n5356)
         );
  XNOR2_X1 U6514 ( .A(n5356), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5459)
         );
  INV_X1 U6515 ( .A(n5357), .ZN(n5359) );
  AOI21_X1 U6516 ( .B1(n5359), .B2(n5358), .A(n5244), .ZN(n5662) );
  NAND2_X1 U6517 ( .A1(n4228), .A2(REIP_REG_23__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U6518 ( .A1(n6036), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5360)
         );
  OAI211_X1 U6519 ( .C1(n6045), .C2(n5609), .A(n5452), .B(n5360), .ZN(n5361)
         );
  AOI21_X1 U6520 ( .B1(n5662), .B2(n4663), .A(n5361), .ZN(n5362) );
  OAI21_X1 U6521 ( .B1(n5459), .B2(n5773), .A(n5362), .ZN(U2963) );
  OAI21_X1 U6522 ( .B1(n5693), .B2(n5364), .A(n5363), .ZN(n5366) );
  XOR2_X1 U6523 ( .A(n5366), .B(n5365), .Z(n5467) );
  NAND2_X1 U6524 ( .A1(n4228), .A2(REIP_REG_22__SCAN_IN), .ZN(n5461) );
  OAI21_X1 U6525 ( .B1(n5393), .B2(n5367), .A(n5461), .ZN(n5369) );
  NOR2_X1 U6526 ( .A1(n5625), .A2(n6026), .ZN(n5368) );
  AOI211_X1 U6527 ( .C1(n6022), .C2(n5617), .A(n5369), .B(n5368), .ZN(n5370)
         );
  OAI21_X1 U6528 ( .B1(n5467), .B2(n5773), .A(n5370), .ZN(U2964) );
  NAND2_X1 U6529 ( .A1(n5275), .A2(n5371), .ZN(n5372) );
  AND2_X1 U6530 ( .A1(n5261), .A2(n5372), .ZN(n5665) );
  INV_X1 U6531 ( .A(n5665), .ZN(n5379) );
  NAND2_X1 U6532 ( .A1(n4228), .A2(REIP_REG_21__SCAN_IN), .ZN(n5471) );
  OAI21_X1 U6533 ( .B1(n5393), .B2(n5373), .A(n5471), .ZN(n5374) );
  AOI21_X1 U6534 ( .B1(n6022), .B2(n5627), .A(n5374), .ZN(n5378) );
  OAI21_X1 U6535 ( .B1(n5376), .B2(n5375), .A(n5353), .ZN(n5468) );
  NAND2_X1 U6536 ( .A1(n5468), .A2(n6040), .ZN(n5377) );
  OAI211_X1 U6537 ( .C1(n5379), .C2(n6026), .A(n5378), .B(n5377), .ZN(U2965)
         );
  INV_X1 U6538 ( .A(n5380), .ZN(n5381) );
  NOR2_X1 U6539 ( .A1(n5382), .A2(n5381), .ZN(n5383) );
  XNOR2_X1 U6540 ( .A(n5384), .B(n5383), .ZN(n5492) );
  INV_X1 U6541 ( .A(n5634), .ZN(n5388) );
  INV_X1 U6542 ( .A(n5385), .ZN(n5632) );
  AOI22_X1 U6543 ( .A1(n6036), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .B1(n4228), 
        .B2(REIP_REG_20__SCAN_IN), .ZN(n5386) );
  OAI21_X1 U6544 ( .B1(n5632), .B2(n6045), .A(n5386), .ZN(n5387) );
  AOI21_X1 U6545 ( .B1(n5388), .B2(n4663), .A(n5387), .ZN(n5389) );
  OAI21_X1 U6546 ( .B1(n5492), .B2(n5773), .A(n5389), .ZN(U2966) );
  XNOR2_X1 U6547 ( .A(n5704), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5391)
         );
  XNOR2_X1 U6548 ( .A(n5390), .B(n5391), .ZN(n5499) );
  NAND2_X1 U6549 ( .A1(n4228), .A2(REIP_REG_15__SCAN_IN), .ZN(n5494) );
  OAI21_X1 U6550 ( .B1(n5393), .B2(n5392), .A(n5494), .ZN(n5395) );
  NOR2_X1 U6551 ( .A1(n5822), .A2(n6026), .ZN(n5394) );
  AOI211_X1 U6552 ( .C1(n5815), .C2(n6022), .A(n5395), .B(n5394), .ZN(n5396)
         );
  OAI21_X1 U6553 ( .B1(n5499), .B2(n5773), .A(n5396), .ZN(U2971) );
  INV_X1 U6554 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5400) );
  OAI21_X1 U6555 ( .B1(n5398), .B2(n5400), .A(n5397), .ZN(n5399) );
  AOI21_X1 U6556 ( .B1(n5566), .B2(n6099), .A(n5399), .ZN(n5403) );
  NAND3_X1 U6557 ( .A1(n5401), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5400), .ZN(n5402) );
  OAI211_X1 U6558 ( .C1(n5404), .C2(n6103), .A(n5403), .B(n5402), .ZN(U2988)
         );
  INV_X1 U6559 ( .A(n5417), .ZN(n5411) );
  NOR3_X1 U6560 ( .A1(n5414), .A2(n5406), .A3(n4200), .ZN(n5410) );
  INV_X1 U6561 ( .A(n5407), .ZN(n5408) );
  OAI21_X1 U6562 ( .B1(n5576), .B2(n5733), .A(n5408), .ZN(n5409) );
  AOI211_X1 U6563 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n5411), .A(n5410), .B(n5409), .ZN(n5412) );
  OAI21_X1 U6564 ( .B1(n5413), .B2(n6103), .A(n5412), .ZN(U2990) );
  INV_X1 U6565 ( .A(n5414), .ZN(n5420) );
  NAND2_X1 U6566 ( .A1(n5581), .A2(n6099), .ZN(n5416) );
  OAI211_X1 U6567 ( .C1(n5417), .C2(n5419), .A(n5416), .B(n5415), .ZN(n5418)
         );
  AOI21_X1 U6568 ( .B1(n5420), .B2(n5419), .A(n5418), .ZN(n5421) );
  OAI21_X1 U6569 ( .B1(n5422), .B2(n6103), .A(n5421), .ZN(U2991) );
  OAI21_X1 U6570 ( .B1(n5585), .B2(n5733), .A(n5423), .ZN(n5429) );
  INV_X1 U6571 ( .A(n5424), .ZN(n5425) );
  AOI211_X1 U6572 ( .C1(n5427), .C2(n5426), .A(n5425), .B(n5436), .ZN(n5428)
         );
  AOI211_X1 U6573 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n5442), .A(n5429), .B(n5428), .ZN(n5430) );
  OAI21_X1 U6574 ( .B1(n5431), .B2(n6103), .A(n5430), .ZN(U2992) );
  AOI21_X1 U6575 ( .B1(n5434), .B2(n5433), .A(n5432), .ZN(n5673) );
  NAND2_X1 U6576 ( .A1(n4228), .A2(REIP_REG_25__SCAN_IN), .ZN(n5435) );
  OAI21_X1 U6577 ( .B1(n5592), .B2(n5733), .A(n5435), .ZN(n5438) );
  NOR2_X1 U6578 ( .A1(n5436), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5437)
         );
  AOI211_X1 U6579 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n5442), .A(n5438), .B(n5437), .ZN(n5439) );
  OAI21_X1 U6580 ( .B1(n5673), .B2(n6103), .A(n5439), .ZN(U2993) );
  INV_X1 U6581 ( .A(n5440), .ZN(n5441) );
  AOI21_X1 U6582 ( .B1(n5602), .B2(n6099), .A(n5441), .ZN(n5445) );
  NAND2_X1 U6583 ( .A1(n5485), .A2(n5487), .ZN(n5477) );
  NOR3_X1 U6584 ( .A1(n5477), .A2(n6702), .A3(n5454), .ZN(n5443) );
  OAI21_X1 U6585 ( .B1(n5443), .B2(INSTADDRPOINTER_REG_24__SCAN_IN), .A(n5442), 
        .ZN(n5444) );
  OAI211_X1 U6586 ( .C1(n5446), .C2(n6103), .A(n5445), .B(n5444), .ZN(U2994)
         );
  INV_X1 U6587 ( .A(n5447), .ZN(n5451) );
  INV_X1 U6588 ( .A(n5448), .ZN(n5450) );
  AOI21_X1 U6589 ( .B1(n5451), .B2(n5450), .A(n5449), .ZN(n5647) );
  INV_X1 U6590 ( .A(n5647), .ZN(n5453) );
  OAI21_X1 U6591 ( .B1(n5453), .B2(n5733), .A(n5452), .ZN(n5456) );
  NOR3_X1 U6592 ( .A1(n5477), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n5454), 
        .ZN(n5455) );
  AOI211_X1 U6593 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5457), .A(n5456), .B(n5455), .ZN(n5458) );
  OAI21_X1 U6594 ( .B1(n5459), .B2(n6103), .A(n5458), .ZN(U2995) );
  INV_X1 U6595 ( .A(n5460), .ZN(n5474) );
  OAI21_X1 U6596 ( .B1(n5619), .B2(n5733), .A(n5461), .ZN(n5465) );
  NOR3_X1 U6597 ( .A1(n5477), .A2(n5463), .A3(n5462), .ZN(n5464) );
  AOI211_X1 U6598 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5474), .A(n5465), .B(n5464), .ZN(n5466) );
  OAI21_X1 U6599 ( .B1(n5467), .B2(n6103), .A(n5466), .ZN(U2996) );
  NAND2_X1 U6600 ( .A1(n5468), .A2(n6090), .ZN(n5476) );
  NAND2_X1 U6601 ( .A1(n3138), .A2(n5469), .ZN(n5470) );
  AND2_X1 U6602 ( .A1(n3124), .A2(n5470), .ZN(n5650) );
  INV_X1 U6603 ( .A(n5650), .ZN(n5472) );
  OAI21_X1 U6604 ( .B1(n5472), .B2(n5733), .A(n5471), .ZN(n5473) );
  AOI21_X1 U6605 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5474), .A(n5473), 
        .ZN(n5475) );
  OAI211_X1 U6606 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5477), .A(n5476), .B(n5475), .ZN(U2997) );
  NAND2_X1 U6607 ( .A1(n5478), .A2(n6717), .ZN(n5739) );
  INV_X1 U6608 ( .A(n5479), .ZN(n5483) );
  AOI21_X1 U6609 ( .B1(n5481), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5480), 
        .ZN(n5482) );
  NOR2_X1 U6610 ( .A1(n5483), .A2(n5482), .ZN(n5734) );
  OAI21_X1 U6611 ( .B1(n5484), .B2(n5739), .A(n5734), .ZN(n5729) );
  AOI21_X1 U6612 ( .B1(n3628), .B2(n5493), .A(n5729), .ZN(n5723) );
  INV_X1 U6613 ( .A(n5723), .ZN(n5490) );
  INV_X1 U6614 ( .A(n5485), .ZN(n5717) );
  NOR3_X1 U6615 ( .A1(n5717), .A2(n5487), .A3(n5486), .ZN(n5489) );
  OAI22_X1 U6616 ( .A1(n5635), .A2(n5733), .B1(n6486), .B2(n5727), .ZN(n5488)
         );
  AOI211_X1 U6617 ( .C1(n5490), .C2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5489), .B(n5488), .ZN(n5491) );
  OAI21_X1 U6618 ( .B1(n5492), .B2(n6103), .A(n5491), .ZN(U2998) );
  NOR2_X1 U6619 ( .A1(n6053), .A2(n5740), .ZN(n5497) );
  AOI21_X1 U6620 ( .B1(n5493), .B2(n5740), .A(n6047), .ZN(n5745) );
  NOR2_X1 U6621 ( .A1(n5745), .A2(n6564), .ZN(n5496) );
  OAI21_X1 U6622 ( .B1(n5733), .B2(n5818), .A(n5494), .ZN(n5495) );
  AOI211_X1 U6623 ( .C1(n5497), .C2(n6564), .A(n5496), .B(n5495), .ZN(n5498)
         );
  OAI21_X1 U6624 ( .B1(n5499), .B2(n6103), .A(n5498), .ZN(U3003) );
  XNOR2_X1 U6625 ( .A(n5500), .B(n5501), .ZN(n5713) );
  NAND2_X1 U6626 ( .A1(n5502), .A2(n5507), .ZN(n5749) );
  NOR2_X1 U6627 ( .A1(n5754), .A2(n5503), .ZN(n5504) );
  AOI211_X1 U6628 ( .C1(n5506), .C2(n5505), .A(n5504), .B(n6047), .ZN(n5746)
         );
  OAI22_X1 U6629 ( .A1(n6053), .A2(n5749), .B1(n5746), .B2(n5507), .ZN(n5509)
         );
  OAI22_X1 U6630 ( .A1(n5733), .A2(n5837), .B1(n5727), .B2(n6476), .ZN(n5508)
         );
  AOI211_X1 U6631 ( .C1(n5713), .C2(n6090), .A(n5509), .B(n5508), .ZN(n5510)
         );
  INV_X1 U6632 ( .A(n5510), .ZN(U3005) );
  INV_X1 U6633 ( .A(n6398), .ZN(n5512) );
  OAI22_X1 U6634 ( .A1(n5512), .A2(n5760), .B1(n5511), .B2(n6431), .ZN(n5513)
         );
  MUX2_X1 U6635 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5513), .S(n5764), 
        .Z(U3456) );
  INV_X1 U6636 ( .A(n6150), .ZN(n5517) );
  NAND2_X1 U6637 ( .A1(n5514), .A2(n6412), .ZN(n6221) );
  INV_X1 U6638 ( .A(n6221), .ZN(n5515) );
  AOI22_X1 U6639 ( .A1(n5517), .A2(n5516), .B1(n6290), .B2(n5515), .ZN(n5556)
         );
  NAND2_X1 U6640 ( .A1(n6339), .A2(n6412), .ZN(n6125) );
  NOR2_X1 U6641 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6125), .ZN(n5552)
         );
  NOR2_X1 U6642 ( .A1(n5520), .A2(n6142), .ZN(n5521) );
  OAI22_X1 U6643 ( .A1(n6157), .A2(n5521), .B1(n3113), .B2(n6119), .ZN(n5522)
         );
  AOI21_X1 U6644 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6221), .A(n4610), .ZN(
        n6226) );
  OAI221_X1 U6645 ( .B1(n5552), .B2(n6817), .C1(n5552), .C2(n5522), .A(n6226), 
        .ZN(n5547) );
  AOI22_X1 U6646 ( .A1(n6142), .A2(n6331), .B1(INSTQUEUE_REG_2__0__SCAN_IN), 
        .B2(n5547), .ZN(n5523) );
  OAI21_X1 U6647 ( .B1(n6350), .B2(n5560), .A(n5523), .ZN(n5524) );
  AOI21_X1 U6648 ( .B1(n6332), .B2(n5552), .A(n5524), .ZN(n5525) );
  OAI21_X1 U6649 ( .B1(n5526), .B2(n5556), .A(n5525), .ZN(U3036) );
  AOI22_X1 U6650 ( .A1(n6142), .A2(n6305), .B1(INSTQUEUE_REG_2__1__SCAN_IN), 
        .B2(n5547), .ZN(n5527) );
  OAI21_X1 U6651 ( .B1(n6308), .B2(n5560), .A(n5527), .ZN(n5528) );
  AOI21_X1 U6652 ( .B1(n6352), .B2(n5552), .A(n5528), .ZN(n5529) );
  OAI21_X1 U6653 ( .B1(n5530), .B2(n5556), .A(n5529), .ZN(U3037) );
  AOI22_X1 U6654 ( .A1(n6142), .A2(n6357), .B1(INSTQUEUE_REG_2__2__SCAN_IN), 
        .B2(n5547), .ZN(n5531) );
  OAI21_X1 U6655 ( .B1(n6362), .B2(n5560), .A(n5531), .ZN(n5532) );
  AOI21_X1 U6656 ( .B1(n6358), .B2(n5552), .A(n5532), .ZN(n5533) );
  OAI21_X1 U6657 ( .B1(n5534), .B2(n5556), .A(n5533), .ZN(U3038) );
  NAND2_X1 U6658 ( .A1(n6364), .A2(n5552), .ZN(n5539) );
  INV_X1 U6659 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5535) );
  INV_X1 U6660 ( .A(n5547), .ZN(n5553) );
  OAI22_X1 U6661 ( .A1(n5556), .A2(n5536), .B1(n5535), .B2(n5553), .ZN(n5537)
         );
  AOI21_X1 U6662 ( .B1(n6142), .B2(n6311), .A(n5537), .ZN(n5538) );
  OAI211_X1 U6663 ( .C1(n5560), .C2(n6314), .A(n5539), .B(n5538), .ZN(U3039)
         );
  AOI22_X1 U6664 ( .A1(n6142), .A2(n6315), .B1(INSTQUEUE_REG_2__4__SCAN_IN), 
        .B2(n5547), .ZN(n5540) );
  OAI21_X1 U6665 ( .B1(n6318), .B2(n5560), .A(n5540), .ZN(n5541) );
  AOI21_X1 U6666 ( .B1(n6371), .B2(n5552), .A(n5541), .ZN(n5542) );
  OAI21_X1 U6667 ( .B1(n5543), .B2(n5556), .A(n5542), .ZN(U3040) );
  AOI22_X1 U6668 ( .A1(n6142), .A2(n6377), .B1(INSTQUEUE_REG_2__5__SCAN_IN), 
        .B2(n5547), .ZN(n5544) );
  OAI21_X1 U6669 ( .B1(n6537), .B2(n5560), .A(n5544), .ZN(n5545) );
  AOI21_X1 U6670 ( .B1(n6378), .B2(n5552), .A(n5545), .ZN(n5546) );
  OAI21_X1 U6671 ( .B1(n6539), .B2(n5556), .A(n5546), .ZN(U3041) );
  AOI22_X1 U6672 ( .A1(n6142), .A2(n6382), .B1(INSTQUEUE_REG_2__6__SCAN_IN), 
        .B2(n5547), .ZN(n5548) );
  OAI21_X1 U6673 ( .B1(n6387), .B2(n5560), .A(n5548), .ZN(n5549) );
  AOI21_X1 U6674 ( .B1(n6383), .B2(n5552), .A(n5549), .ZN(n5550) );
  OAI21_X1 U6675 ( .B1(n5551), .B2(n5556), .A(n5550), .ZN(U3042) );
  NAND2_X1 U6676 ( .A1(n6391), .A2(n5552), .ZN(n5559) );
  INV_X1 U6677 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5554) );
  OAI22_X1 U6678 ( .A1(n5556), .A2(n5555), .B1(n5554), .B2(n5553), .ZN(n5557)
         );
  AOI21_X1 U6679 ( .B1(n6142), .B2(n6389), .A(n5557), .ZN(n5558) );
  OAI211_X1 U6680 ( .C1(n5560), .C2(n6397), .A(n5559), .B(n5558), .ZN(U3043)
         );
  AND2_X1 U6681 ( .A1(n5962), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U6682 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6500) );
  AOI22_X1 U6683 ( .A1(EBX_REG_30__SCAN_IN), .A2(n5908), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n5893), .ZN(n5561) );
  OAI21_X1 U6684 ( .B1(n5562), .B2(n6500), .A(n5561), .ZN(n5563) );
  AOI21_X1 U6685 ( .B1(n5564), .B2(n5892), .A(n5563), .ZN(n5568) );
  AOI22_X1 U6686 ( .A1(n5566), .A2(n5891), .B1(n5565), .B2(n6500), .ZN(n5567)
         );
  OAI211_X1 U6687 ( .C1(n4364), .C2(n5902), .A(n5568), .B(n5567), .ZN(U2797)
         );
  OAI22_X1 U6688 ( .A1(n5569), .A2(n5897), .B1(n4114), .B2(n5904), .ZN(n5573)
         );
  OAI22_X1 U6689 ( .A1(n5571), .A2(n4210), .B1(n5570), .B2(n5903), .ZN(n5572)
         );
  AOI211_X1 U6690 ( .C1(n5653), .C2(n5886), .A(n5573), .B(n5572), .ZN(n5575)
         );
  NAND3_X1 U6691 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5580), .A3(n4210), .ZN(
        n5574) );
  OAI211_X1 U6692 ( .C1(n5916), .C2(n5576), .A(n5575), .B(n5574), .ZN(U2799)
         );
  AOI22_X1 U6693 ( .A1(EBX_REG_27__SCAN_IN), .A2(n5908), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n5893), .ZN(n5577) );
  OAI21_X1 U6694 ( .B1(n6655), .B2(n5586), .A(n5577), .ZN(n5578) );
  AOI21_X1 U6695 ( .B1(n5579), .B2(n5892), .A(n5578), .ZN(n5583) );
  AOI22_X1 U6696 ( .A1(n5891), .A2(n5581), .B1(n5580), .B2(n6655), .ZN(n5582)
         );
  OAI211_X1 U6697 ( .C1(n5584), .C2(n5902), .A(n5583), .B(n5582), .ZN(U2800)
         );
  AOI22_X1 U6698 ( .A1(EBX_REG_26__SCAN_IN), .A2(n5908), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n5893), .ZN(n5590) );
  INV_X1 U6699 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6627) );
  NOR2_X1 U6700 ( .A1(n6627), .A2(n5597), .ZN(n5595) );
  AOI21_X1 U6701 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5595), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5587) );
  OAI22_X1 U6702 ( .A1(n5587), .A2(n5586), .B1(n5585), .B2(n5916), .ZN(n5588)
         );
  AOI21_X1 U6703 ( .B1(n5656), .B2(n5886), .A(n5588), .ZN(n5589) );
  OAI211_X1 U6704 ( .C1(n5591), .C2(n5903), .A(n5590), .B(n5589), .ZN(U2801)
         );
  INV_X1 U6705 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6491) );
  INV_X1 U6706 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6720) );
  OAI22_X1 U6707 ( .A1(n6607), .A2(n5897), .B1(n6720), .B2(n5904), .ZN(n5594)
         );
  OAI22_X1 U6708 ( .A1(n5674), .A2(n5903), .B1(n5916), .B2(n5592), .ZN(n5593)
         );
  AOI211_X1 U6709 ( .C1(n5595), .C2(n6491), .A(n5594), .B(n5593), .ZN(n5599)
         );
  NAND2_X1 U6710 ( .A1(n5859), .A2(n5596), .ZN(n5613) );
  INV_X1 U6711 ( .A(n5613), .ZN(n5601) );
  NOR2_X1 U6712 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5597), .ZN(n5603) );
  OAI21_X1 U6713 ( .B1(n5601), .B2(n5603), .A(REIP_REG_25__SCAN_IN), .ZN(n5598) );
  OAI211_X1 U6714 ( .C1(n5679), .C2(n5902), .A(n5599), .B(n5598), .ZN(U2802)
         );
  AOI22_X1 U6715 ( .A1(EBX_REG_24__SCAN_IN), .A2(n5908), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n5893), .ZN(n5607) );
  AOI22_X1 U6716 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5601), .B1(n5600), .B2(
        n5892), .ZN(n5606) );
  AOI22_X1 U6717 ( .A1(n5602), .A2(n5891), .B1(n5659), .B2(n5886), .ZN(n5605)
         );
  INV_X1 U6718 ( .A(n5603), .ZN(n5604) );
  NAND4_X1 U6719 ( .A1(n5607), .A2(n5606), .A3(n5605), .A4(n5604), .ZN(U2803)
         );
  INV_X1 U6720 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6489) );
  INV_X1 U6721 ( .A(REIP_REG_21__SCAN_IN), .ZN(n5616) );
  NOR2_X1 U6722 ( .A1(n6489), .A2(n5616), .ZN(n5608) );
  AOI21_X1 U6723 ( .B1(n5622), .B2(n5608), .A(REIP_REG_23__SCAN_IN), .ZN(n5614) );
  OAI22_X1 U6724 ( .A1(n5649), .A2(n5897), .B1(n5609), .B2(n5903), .ZN(n5610)
         );
  AOI21_X1 U6725 ( .B1(PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n5893), .A(n5610), 
        .ZN(n5612) );
  AOI22_X1 U6726 ( .A1(n5662), .A2(n5886), .B1(n5647), .B2(n5891), .ZN(n5611)
         );
  OAI211_X1 U6727 ( .C1(n5614), .C2(n5613), .A(n5612), .B(n5611), .ZN(U2804)
         );
  NOR2_X1 U6728 ( .A1(n5881), .A2(n5615), .ZN(n5626) );
  INV_X1 U6729 ( .A(n5626), .ZN(n5640) );
  NAND2_X1 U6730 ( .A1(n5622), .A2(n5616), .ZN(n5628) );
  AOI21_X1 U6731 ( .B1(n5640), .B2(n5628), .A(n6489), .ZN(n5621) );
  AOI22_X1 U6732 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n5893), .B1(n5617), 
        .B2(n5892), .ZN(n5618) );
  OAI21_X1 U6733 ( .B1(n5619), .B2(n5916), .A(n5618), .ZN(n5620) );
  AOI211_X1 U6734 ( .C1(n5908), .C2(EBX_REG_22__SCAN_IN), .A(n5621), .B(n5620), 
        .ZN(n5624) );
  NAND3_X1 U6735 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5622), .A3(n6489), .ZN(
        n5623) );
  OAI211_X1 U6736 ( .C1(n5902), .C2(n5625), .A(n5624), .B(n5623), .ZN(U2805)
         );
  AOI22_X1 U6737 ( .A1(EBX_REG_21__SCAN_IN), .A2(n5908), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n5893), .ZN(n5631) );
  AOI22_X1 U6738 ( .A1(n5627), .A2(n5892), .B1(REIP_REG_21__SCAN_IN), .B2(
        n5626), .ZN(n5630) );
  AOI22_X1 U6739 ( .A1(n5665), .A2(n5886), .B1(n5650), .B2(n5891), .ZN(n5629)
         );
  NAND4_X1 U6740 ( .A1(n5631), .A2(n5630), .A3(n5629), .A4(n5628), .ZN(U2806)
         );
  OAI22_X1 U6741 ( .A1(n5633), .A2(n5904), .B1(n5632), .B2(n5903), .ZN(n5637)
         );
  OAI22_X1 U6742 ( .A1(n5635), .A2(n5916), .B1(n5902), .B2(n5634), .ZN(n5636)
         );
  AOI211_X1 U6743 ( .C1(EBX_REG_20__SCAN_IN), .C2(n5908), .A(n5637), .B(n5636), 
        .ZN(n5638) );
  OAI221_X1 U6744 ( .B1(n5640), .B2(n6486), .C1(n5640), .C2(n5639), .A(n5638), 
        .ZN(U2807) );
  AOI22_X1 U6745 ( .A1(EBX_REG_19__SCAN_IN), .A2(n5908), .B1(n5891), .B2(n5716), .ZN(n5641) );
  OAI21_X1 U6746 ( .B1(n5688), .B2(n5903), .A(n5641), .ZN(n5642) );
  AOI211_X1 U6747 ( .C1(n5893), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5907), 
        .B(n5642), .ZN(n5646) );
  AND2_X1 U6748 ( .A1(n5859), .A2(n5643), .ZN(n5801) );
  INV_X1 U6749 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6483) );
  XNOR2_X1 U6750 ( .A(REIP_REG_19__SCAN_IN), .B(n6483), .ZN(n5644) );
  AOI22_X1 U6751 ( .A1(REIP_REG_19__SCAN_IN), .A2(n5801), .B1(n5793), .B2(
        n5644), .ZN(n5645) );
  OAI211_X1 U6752 ( .C1(n5902), .C2(n5684), .A(n5646), .B(n5645), .ZN(U2808)
         );
  AOI22_X1 U6753 ( .A1(n5662), .A2(n5924), .B1(n5923), .B2(n5647), .ZN(n5648)
         );
  OAI21_X1 U6754 ( .B1(n5927), .B2(n5649), .A(n5648), .ZN(U2836) );
  AOI22_X1 U6755 ( .A1(n5665), .A2(n5924), .B1(n5923), .B2(n5650), .ZN(n5651)
         );
  OAI21_X1 U6756 ( .B1(n5927), .B2(n6566), .A(n5651), .ZN(U2838) );
  INV_X1 U6757 ( .A(n5652), .ZN(n5929) );
  AOI22_X1 U6758 ( .A1(n5653), .A2(n5929), .B1(n5928), .B2(DATAI_28_), .ZN(
        n5655) );
  AOI22_X1 U6759 ( .A1(n5932), .A2(DATAI_12_), .B1(n5931), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U6760 ( .A1(n5655), .A2(n5654), .ZN(U2863) );
  AOI22_X1 U6761 ( .A1(n5656), .A2(n5929), .B1(n5928), .B2(DATAI_26_), .ZN(
        n5658) );
  AOI22_X1 U6762 ( .A1(n5932), .A2(DATAI_10_), .B1(n5931), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U6763 ( .A1(n5658), .A2(n5657), .ZN(U2865) );
  AOI22_X1 U6764 ( .A1(n5659), .A2(n5929), .B1(DATAI_24_), .B2(n5928), .ZN(
        n5661) );
  AOI22_X1 U6765 ( .A1(n5932), .A2(DATAI_8_), .B1(n5931), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5660) );
  NAND2_X1 U6766 ( .A1(n5661), .A2(n5660), .ZN(U2867) );
  AOI22_X1 U6767 ( .A1(n5662), .A2(n5929), .B1(n5928), .B2(DATAI_23_), .ZN(
        n5664) );
  AOI22_X1 U6768 ( .A1(n5932), .A2(DATAI_7_), .B1(n5931), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U6769 ( .A1(n5664), .A2(n5663), .ZN(U2868) );
  AOI22_X1 U6770 ( .A1(n5665), .A2(n5929), .B1(n5928), .B2(DATAI_21_), .ZN(
        n5667) );
  AOI22_X1 U6771 ( .A1(n5932), .A2(DATAI_5_), .B1(n5931), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5666) );
  NAND2_X1 U6772 ( .A1(n5667), .A2(n5666), .ZN(U2870) );
  INV_X1 U6773 ( .A(DATAI_19_), .ZN(n5668) );
  OAI22_X1 U6774 ( .A1(n5684), .A2(n5652), .B1(n5669), .B2(n5668), .ZN(n5670)
         );
  INV_X1 U6775 ( .A(n5670), .ZN(n5672) );
  AOI22_X1 U6776 ( .A1(n5932), .A2(DATAI_3_), .B1(n5931), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U6777 ( .A1(n5672), .A2(n5671), .ZN(U2872) );
  AOI22_X1 U6778 ( .A1(n4228), .A2(REIP_REG_25__SCAN_IN), .B1(n6036), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5678) );
  INV_X1 U6779 ( .A(n5673), .ZN(n5676) );
  INV_X1 U6780 ( .A(n5674), .ZN(n5675) );
  AOI22_X1 U6781 ( .A1(n5676), .A2(n6040), .B1(n6022), .B2(n5675), .ZN(n5677)
         );
  OAI211_X1 U6782 ( .C1(n6026), .C2(n5679), .A(n5678), .B(n5677), .ZN(U2961)
         );
  AOI22_X1 U6783 ( .A1(n4228), .A2(REIP_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6036), .ZN(n5687) );
  OR2_X1 U6784 ( .A1(n5681), .A2(n5680), .ZN(n5682) );
  NAND2_X1 U6785 ( .A1(n5683), .A2(n5682), .ZN(n5718) );
  OAI22_X1 U6786 ( .A1(n5684), .A2(n6026), .B1(n5773), .B2(n5718), .ZN(n5685)
         );
  INV_X1 U6787 ( .A(n5685), .ZN(n5686) );
  OAI211_X1 U6788 ( .C1(n5688), .C2(n6045), .A(n5687), .B(n5686), .ZN(U2967)
         );
  AOI22_X1 U6789 ( .A1(n4228), .A2(REIP_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6036), .ZN(n5692) );
  NOR3_X1 U6790 ( .A1(n3125), .A2(n5693), .A3(n6717), .ZN(n5698) );
  NAND2_X1 U6791 ( .A1(n5693), .A2(n6579), .ZN(n5695) );
  NOR3_X1 U6792 ( .A1(n5689), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5695), 
        .ZN(n5696) );
  NOR2_X1 U6793 ( .A1(n5698), .A2(n5696), .ZN(n5690) );
  XNOR2_X1 U6794 ( .A(n5690), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5725)
         );
  AOI22_X1 U6795 ( .A1(n5789), .A2(n6022), .B1(n6040), .B2(n5725), .ZN(n5691)
         );
  OAI211_X1 U6796 ( .C1(n6026), .C2(n5796), .A(n5692), .B(n5691), .ZN(U2968)
         );
  AOI22_X1 U6797 ( .A1(n4228), .A2(REIP_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6036), .ZN(n5702) );
  AOI21_X1 U6798 ( .B1(n5693), .B2(n6717), .A(n3125), .ZN(n5694) );
  AOI21_X1 U6799 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5695), .A(n5694), 
        .ZN(n5699) );
  INV_X1 U6800 ( .A(n5696), .ZN(n5697) );
  OAI21_X1 U6801 ( .B1(n5699), .B2(n5698), .A(n5697), .ZN(n5736) );
  AOI22_X1 U6802 ( .A1(n5700), .A2(n5930), .B1(n6040), .B2(n5736), .ZN(n5701)
         );
  OAI211_X1 U6803 ( .C1(n5797), .C2(n6045), .A(n5702), .B(n5701), .ZN(U2969)
         );
  AOI22_X1 U6804 ( .A1(n4228), .A2(REIP_REG_16__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n6036), .ZN(n5707) );
  XNOR2_X1 U6805 ( .A(n5704), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5705)
         );
  XNOR2_X1 U6806 ( .A(n5703), .B(n5705), .ZN(n5742) );
  AOI22_X1 U6807 ( .A1(n5742), .A2(n6040), .B1(n6022), .B2(n5805), .ZN(n5706)
         );
  OAI211_X1 U6808 ( .C1(n6026), .C2(n5814), .A(n5707), .B(n5706), .ZN(U2970)
         );
  AOI22_X1 U6809 ( .A1(n4228), .A2(REIP_REG_14__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n6036), .ZN(n5711) );
  XNOR2_X1 U6810 ( .A(n5704), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5709)
         );
  XNOR2_X1 U6811 ( .A(n5708), .B(n5709), .ZN(n5751) );
  AOI22_X1 U6812 ( .A1(n5751), .A2(n6040), .B1(n6022), .B2(n5824), .ZN(n5710)
         );
  OAI211_X1 U6813 ( .C1(n6026), .C2(n5831), .A(n5711), .B(n5710), .ZN(U2972)
         );
  AOI22_X1 U6814 ( .A1(n4228), .A2(REIP_REG_13__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n6036), .ZN(n5715) );
  INV_X1 U6815 ( .A(n5712), .ZN(n5834) );
  AOI22_X1 U6816 ( .A1(n5713), .A2(n6040), .B1(n6022), .B2(n5834), .ZN(n5714)
         );
  OAI211_X1 U6817 ( .C1(n6026), .C2(n5833), .A(n5715), .B(n5714), .ZN(U2973)
         );
  AOI22_X1 U6818 ( .A1(n5716), .A2(n6099), .B1(n4228), .B2(
        REIP_REG_19__SCAN_IN), .ZN(n5721) );
  OAI22_X1 U6819 ( .A1(n5718), .A2(n6103), .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5717), .ZN(n5719) );
  INV_X1 U6820 ( .A(n5719), .ZN(n5720) );
  OAI211_X1 U6821 ( .C1(n5723), .C2(n5722), .A(n5721), .B(n5720), .ZN(U2999)
         );
  INV_X1 U6822 ( .A(n5724), .ZN(n5788) );
  AOI22_X1 U6823 ( .A1(n5725), .A2(n6090), .B1(n6099), .B2(n5788), .ZN(n5732)
         );
  INV_X1 U6824 ( .A(n5726), .ZN(n5730) );
  NOR2_X1 U6825 ( .A1(n5727), .A2(n6483), .ZN(n5728) );
  AOI221_X1 U6826 ( .B1(n5730), .B2(n3628), .C1(n5729), .C2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .A(n5728), .ZN(n5731) );
  NAND2_X1 U6827 ( .A1(n5732), .A2(n5731), .ZN(U3000) );
  OAI22_X1 U6828 ( .A1(n5734), .A2(n6717), .B1(n5733), .B2(n5804), .ZN(n5735)
         );
  AOI21_X1 U6829 ( .B1(n5736), .B2(n6090), .A(n5735), .ZN(n5738) );
  NAND2_X1 U6830 ( .A1(n4228), .A2(REIP_REG_17__SCAN_IN), .ZN(n5737) );
  OAI211_X1 U6831 ( .C1(n6053), .C2(n5739), .A(n5738), .B(n5737), .ZN(U3001)
         );
  AOI22_X1 U6832 ( .A1(n5809), .A2(n6099), .B1(n4228), .B2(
        REIP_REG_16__SCAN_IN), .ZN(n5744) );
  AOI211_X1 U6833 ( .C1(n6564), .C2(n6579), .A(n6053), .B(n5740), .ZN(n5741)
         );
  AOI22_X1 U6834 ( .A1(n5742), .A2(n6090), .B1(n5741), .B2(n6824), .ZN(n5743)
         );
  OAI211_X1 U6835 ( .C1(n5745), .C2(n6579), .A(n5744), .B(n5743), .ZN(U3002)
         );
  AOI22_X1 U6836 ( .A1(n6099), .A2(n5823), .B1(n4228), .B2(
        REIP_REG_14__SCAN_IN), .ZN(n5757) );
  OAI221_X1 U6837 ( .B1(n5749), .B2(n5748), .C1(n5749), .C2(n5747), .A(n5746), 
        .ZN(n5750) );
  AOI22_X1 U6838 ( .A1(n5751), .A2(n6090), .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n5750), .ZN(n5756) );
  NAND3_X1 U6839 ( .A1(n5754), .A2(n5753), .A3(n5752), .ZN(n5755) );
  NAND3_X1 U6840 ( .A1(n5757), .A2(n5756), .A3(n5755), .ZN(U3004) );
  OR4_X1 U6841 ( .A1(n5761), .A2(n5760), .A3(n5759), .A4(n5758), .ZN(n5762) );
  OAI21_X1 U6842 ( .B1(n5764), .B2(n5763), .A(n5762), .ZN(U3455) );
  AOI21_X1 U6843 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6451), .A(n4236), .ZN(n5770) );
  INV_X1 U6844 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5765) );
  INV_X1 U6845 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6448) );
  NOR2_X4 U6846 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6448), .ZN(n6532) );
  AOI21_X1 U6847 ( .B1(n5770), .B2(n5765), .A(n6532), .ZN(U2789) );
  OAI21_X1 U6848 ( .B1(n5766), .B2(n6434), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5767) );
  OAI21_X1 U6849 ( .B1(n5768), .B2(n6525), .A(n5767), .ZN(U2790) );
  INV_X1 U6850 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6548) );
  NOR2_X1 U6851 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n5771) );
  NOR2_X1 U6852 ( .A1(n6532), .A2(n5771), .ZN(n5769) );
  AOI22_X1 U6853 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n6532), .B1(n6548), .B2(
        n5769), .ZN(U2791) );
  NOR2_X1 U6854 ( .A1(n6532), .A2(n5770), .ZN(n6505) );
  OAI21_X1 U6855 ( .B1(BS16_N), .B2(n5771), .A(n6505), .ZN(n6503) );
  OAI21_X1 U6856 ( .B1(n6505), .B2(n6523), .A(n6503), .ZN(U2792) );
  INV_X1 U6857 ( .A(n5772), .ZN(n5774) );
  OAI21_X1 U6858 ( .B1(n5774), .B2(n6708), .A(n5773), .ZN(U2793) );
  NOR4_X1 U6859 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n5778) );
  NOR4_X1 U6860 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(
        DATAWIDTH_REG_13__SCAN_IN), .ZN(n5777) );
  NOR4_X1 U6861 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_27__SCAN_IN), .A3(DATAWIDTH_REG_28__SCAN_IN), .A4(
        DATAWIDTH_REG_29__SCAN_IN), .ZN(n5776) );
  NOR4_X1 U6862 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n5775) );
  NAND4_X1 U6863 ( .A1(n5778), .A2(n5777), .A3(n5776), .A4(n5775), .ZN(n5784)
         );
  NOR4_X1 U6864 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(
        DATAWIDTH_REG_31__SCAN_IN), .A3(DATAWIDTH_REG_17__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n5782) );
  AOI211_X1 U6865 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_5__SCAN_IN), .B(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n5781) );
  NOR4_X1 U6866 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_9__SCAN_IN), .ZN(
        n5780) );
  NOR4_X1 U6867 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_4__SCAN_IN), .ZN(n5779) );
  NAND4_X1 U6868 ( .A1(n5782), .A2(n5781), .A3(n5780), .A4(n5779), .ZN(n5783)
         );
  NOR2_X1 U6869 ( .A1(n5784), .A2(n5783), .ZN(n6513) );
  INV_X1 U6870 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6786) );
  INV_X1 U6871 ( .A(n6513), .ZN(n6515) );
  INV_X1 U6872 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6516) );
  NOR2_X1 U6873 ( .A1(REIP_REG_0__SCAN_IN), .A2(n6515), .ZN(n6517) );
  NOR2_X1 U6874 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .ZN(n6510) );
  NAND2_X1 U6875 ( .A1(n6517), .A2(n6510), .ZN(n5786) );
  OAI221_X1 U6876 ( .B1(n6513), .B2(n6786), .C1(n6515), .C2(n6516), .A(n5786), 
        .ZN(U2794) );
  OAI21_X1 U6877 ( .B1(REIP_REG_1__SCAN_IN), .B2(DATAWIDTH_REG_1__SCAN_IN), 
        .A(n6513), .ZN(n5785) );
  OAI21_X1 U6878 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(n6513), .A(n5785), .ZN(
        n5787) );
  NAND2_X1 U6879 ( .A1(n5787), .A2(n5786), .ZN(U2795) );
  AOI22_X1 U6880 ( .A1(n5789), .A2(n5892), .B1(n5891), .B2(n5788), .ZN(n5790)
         );
  OAI211_X1 U6881 ( .C1(n5904), .C2(n5791), .A(n5790), .B(n5894), .ZN(n5792)
         );
  AOI21_X1 U6882 ( .B1(EBX_REG_18__SCAN_IN), .B2(n5908), .A(n5792), .ZN(n5795)
         );
  AOI22_X1 U6883 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5801), .B1(n5793), .B2(
        n6483), .ZN(n5794) );
  OAI211_X1 U6884 ( .C1(n5902), .C2(n5796), .A(n5795), .B(n5794), .ZN(U2809)
         );
  INV_X1 U6885 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6779) );
  OAI22_X1 U6886 ( .A1(n6779), .A2(n5904), .B1(n5797), .B2(n5903), .ZN(n5798)
         );
  AOI211_X1 U6887 ( .C1(n5908), .C2(EBX_REG_17__SCAN_IN), .A(n5907), .B(n5798), 
        .ZN(n5803) );
  NAND2_X1 U6888 ( .A1(n6480), .A2(n5799), .ZN(n5800) );
  AOI22_X1 U6889 ( .A1(n5886), .A2(n5930), .B1(n5801), .B2(n5800), .ZN(n5802)
         );
  OAI211_X1 U6890 ( .C1(n5916), .C2(n5804), .A(n5803), .B(n5802), .ZN(U2810)
         );
  AOI22_X1 U6891 ( .A1(EBX_REG_16__SCAN_IN), .A2(n5908), .B1(n5805), .B2(n5892), .ZN(n5806) );
  OAI211_X1 U6892 ( .C1(n5904), .C2(n5807), .A(n5806), .B(n5894), .ZN(n5808)
         );
  AOI21_X1 U6893 ( .B1(n5891), .B2(n5809), .A(n5808), .ZN(n5813) );
  NOR2_X1 U6894 ( .A1(n5881), .A2(n5810), .ZN(n5828) );
  AOI21_X1 U6895 ( .B1(n6726), .B2(n6651), .A(n6832), .ZN(n5811) );
  AOI22_X1 U6896 ( .A1(REIP_REG_16__SCAN_IN), .A2(n5828), .B1(n5820), .B2(
        n5811), .ZN(n5812) );
  OAI211_X1 U6897 ( .C1(n5902), .C2(n5814), .A(n5813), .B(n5812), .ZN(U2811)
         );
  AOI21_X1 U6898 ( .B1(n5893), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5907), 
        .ZN(n5817) );
  AOI22_X1 U6899 ( .A1(EBX_REG_15__SCAN_IN), .A2(n5908), .B1(n5815), .B2(n5892), .ZN(n5816) );
  OAI211_X1 U6900 ( .C1(n5916), .C2(n5818), .A(n5817), .B(n5816), .ZN(n5819)
         );
  AOI221_X1 U6901 ( .B1(n5828), .B2(REIP_REG_15__SCAN_IN), .C1(n5820), .C2(
        n6726), .A(n5819), .ZN(n5821) );
  OAI21_X1 U6902 ( .B1(n5902), .B2(n5822), .A(n5821), .ZN(U2812) );
  AOI22_X1 U6903 ( .A1(n5824), .A2(n5892), .B1(n5891), .B2(n5823), .ZN(n5825)
         );
  OAI21_X1 U6904 ( .B1(n6658), .B2(n5897), .A(n5825), .ZN(n5826) );
  AOI211_X1 U6905 ( .C1(n5893), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n5907), 
        .B(n5826), .ZN(n5830) );
  NOR2_X1 U6906 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5841), .ZN(n5827) );
  AOI22_X1 U6907 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5828), .B1(
        REIP_REG_13__SCAN_IN), .B2(n5827), .ZN(n5829) );
  OAI211_X1 U6908 ( .C1(n5902), .C2(n5831), .A(n5830), .B(n5829), .ZN(U2813)
         );
  INV_X1 U6909 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6476) );
  NAND2_X1 U6910 ( .A1(n5859), .A2(n5832), .ZN(n5848) );
  INV_X1 U6911 ( .A(n5833), .ZN(n5839) );
  AOI21_X1 U6912 ( .B1(n5893), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5907), 
        .ZN(n5836) );
  AOI22_X1 U6913 ( .A1(EBX_REG_13__SCAN_IN), .A2(n5908), .B1(n5834), .B2(n5892), .ZN(n5835) );
  OAI211_X1 U6914 ( .C1(n5916), .C2(n5837), .A(n5836), .B(n5835), .ZN(n5838)
         );
  AOI21_X1 U6915 ( .B1(n5886), .B2(n5839), .A(n5838), .ZN(n5840) );
  OAI221_X1 U6916 ( .B1(REIP_REG_13__SCAN_IN), .B2(n5841), .C1(n6476), .C2(
        n5848), .A(n5840), .ZN(U2814) );
  NOR2_X1 U6917 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5842), .ZN(n5849) );
  INV_X1 U6918 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6723) );
  OAI22_X1 U6919 ( .A1(n6723), .A2(n5897), .B1(n5843), .B2(n5904), .ZN(n5844)
         );
  AOI211_X1 U6920 ( .C1(n5892), .C2(n5845), .A(n5907), .B(n5844), .ZN(n5847)
         );
  AOI22_X1 U6921 ( .A1(n5891), .A2(n5917), .B1(n5886), .B2(n5918), .ZN(n5846)
         );
  OAI211_X1 U6922 ( .C1(n5849), .C2(n5848), .A(n5847), .B(n5846), .ZN(U2815)
         );
  INV_X1 U6923 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5850) );
  OAI22_X1 U6924 ( .A1(n5850), .A2(n5897), .B1(n6553), .B2(n5904), .ZN(n5851)
         );
  AOI211_X1 U6925 ( .C1(n5892), .C2(n5976), .A(n5907), .B(n5851), .ZN(n5856)
         );
  NAND2_X1 U6926 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n5857) );
  NOR3_X1 U6927 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5872), .A3(n5857), .ZN(n5854) );
  INV_X1 U6928 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6473) );
  NOR3_X1 U6929 ( .A1(n5881), .A2(n5852), .A3(n6473), .ZN(n5853) );
  AOI211_X1 U6930 ( .C1(n6048), .C2(n5891), .A(n5854), .B(n5853), .ZN(n5855)
         );
  OAI211_X1 U6931 ( .C1(n5902), .C2(n5979), .A(n5856), .B(n5855), .ZN(U2816)
         );
  OAI21_X1 U6932 ( .B1(REIP_REG_10__SCAN_IN), .B2(REIP_REG_9__SCAN_IN), .A(
        n5857), .ZN(n5865) );
  AND2_X1 U6933 ( .A1(n5859), .A2(n5858), .ZN(n5876) );
  AOI22_X1 U6934 ( .A1(n5891), .A2(n5920), .B1(REIP_REG_10__SCAN_IN), .B2(
        n5876), .ZN(n5864) );
  INV_X1 U6935 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6621) );
  AOI22_X1 U6936 ( .A1(PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n5893), .B1(n5860), 
        .B2(n5892), .ZN(n5861) );
  OAI211_X1 U6937 ( .C1(n5897), .C2(n6621), .A(n5861), .B(n5894), .ZN(n5862)
         );
  AOI21_X1 U6938 ( .B1(n5886), .B2(n5921), .A(n5862), .ZN(n5863) );
  OAI211_X1 U6939 ( .C1(n5872), .C2(n5865), .A(n5864), .B(n5863), .ZN(U2817)
         );
  AOI22_X1 U6940 ( .A1(n5891), .A2(n6054), .B1(REIP_REG_9__SCAN_IN), .B2(n5876), .ZN(n5871) );
  INV_X1 U6941 ( .A(n5986), .ZN(n5869) );
  AOI22_X1 U6942 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n5893), .B1(n5983), 
        .B2(n5892), .ZN(n5866) );
  OAI211_X1 U6943 ( .C1(n5897), .C2(n5867), .A(n5866), .B(n5894), .ZN(n5868)
         );
  AOI21_X1 U6944 ( .B1(n5886), .B2(n5869), .A(n5868), .ZN(n5870) );
  OAI211_X1 U6945 ( .C1(REIP_REG_9__SCAN_IN), .C2(n5872), .A(n5871), .B(n5870), 
        .ZN(U2818) );
  AOI22_X1 U6946 ( .A1(EBX_REG_8__SCAN_IN), .A2(n5908), .B1(n5991), .B2(n5892), 
        .ZN(n5873) );
  OAI211_X1 U6947 ( .C1(n5904), .C2(n5874), .A(n5873), .B(n5894), .ZN(n5875)
         );
  AOI21_X1 U6948 ( .B1(n5891), .B2(n6060), .A(n5875), .ZN(n5878) );
  INV_X1 U6949 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6674) );
  INV_X1 U6950 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6468) );
  NOR2_X1 U6951 ( .A1(n6674), .A2(n6468), .ZN(n5885) );
  OAI221_X1 U6952 ( .B1(REIP_REG_8__SCAN_IN), .B2(n5899), .C1(
        REIP_REG_8__SCAN_IN), .C2(n5885), .A(n5876), .ZN(n5877) );
  OAI211_X1 U6953 ( .C1(n5994), .C2(n5902), .A(n5878), .B(n5877), .ZN(U2819)
         );
  XNOR2_X1 U6954 ( .A(n5880), .B(n5879), .ZN(n6066) );
  NOR2_X1 U6955 ( .A1(n5882), .A2(n5881), .ZN(n5910) );
  AOI22_X1 U6956 ( .A1(n5891), .A2(n6066), .B1(REIP_REG_7__SCAN_IN), .B2(n5910), .ZN(n5890) );
  INV_X1 U6957 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5883) );
  OAI22_X1 U6958 ( .A1(n5883), .A2(n5904), .B1(n6002), .B2(n5903), .ZN(n5884)
         );
  AOI211_X1 U6959 ( .C1(n5908), .C2(EBX_REG_7__SCAN_IN), .A(n5907), .B(n5884), 
        .ZN(n5889) );
  AOI21_X1 U6960 ( .B1(n6674), .B2(n6468), .A(n5885), .ZN(n5887) );
  AOI22_X1 U6961 ( .A1(n5899), .A2(n5887), .B1(n5886), .B2(n5999), .ZN(n5888)
         );
  NAND3_X1 U6962 ( .A1(n5890), .A2(n5889), .A3(n5888), .ZN(U2820) );
  AOI22_X1 U6963 ( .A1(n5891), .A2(n6073), .B1(REIP_REG_6__SCAN_IN), .B2(n5910), .ZN(n5901) );
  AOI22_X1 U6964 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n5893), .B1(n6007), 
        .B2(n5892), .ZN(n5895) );
  OAI211_X1 U6965 ( .C1(n5897), .C2(n5896), .A(n5895), .B(n5894), .ZN(n5898)
         );
  AOI21_X1 U6966 ( .B1(n5899), .B2(n6468), .A(n5898), .ZN(n5900) );
  OAI211_X1 U6967 ( .C1(n5902), .C2(n6010), .A(n5901), .B(n5900), .ZN(U2821)
         );
  INV_X1 U6968 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5905) );
  OAI22_X1 U6969 ( .A1(n5905), .A2(n5904), .B1(n6016), .B2(n5903), .ZN(n5906)
         );
  AOI211_X1 U6970 ( .C1(n5908), .C2(EBX_REG_5__SCAN_IN), .A(n5907), .B(n5906), 
        .ZN(n5914) );
  NAND2_X1 U6971 ( .A1(n6467), .A2(n5909), .ZN(n5911) );
  AOI22_X1 U6972 ( .A1(n5912), .A2(n6013), .B1(n5911), .B2(n5910), .ZN(n5913)
         );
  OAI211_X1 U6973 ( .C1(n5916), .C2(n5915), .A(n5914), .B(n5913), .ZN(U2822)
         );
  AOI22_X1 U6974 ( .A1(n5918), .A2(n5924), .B1(n5923), .B2(n5917), .ZN(n5919)
         );
  OAI21_X1 U6975 ( .B1(n5927), .B2(n6723), .A(n5919), .ZN(U2847) );
  AOI22_X1 U6976 ( .A1(n5921), .A2(n5924), .B1(n5923), .B2(n5920), .ZN(n5922)
         );
  OAI21_X1 U6977 ( .B1(n5927), .B2(n6621), .A(n5922), .ZN(U2849) );
  AOI22_X1 U6978 ( .A1(n5999), .A2(n5924), .B1(n5923), .B2(n6066), .ZN(n5925)
         );
  OAI21_X1 U6979 ( .B1(n5927), .B2(n5926), .A(n5925), .ZN(U2852) );
  AOI22_X1 U6980 ( .A1(n5930), .A2(n5929), .B1(n5928), .B2(DATAI_17_), .ZN(
        n5934) );
  AOI22_X1 U6981 ( .A1(n5932), .A2(DATAI_1_), .B1(n5931), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5933) );
  NAND2_X1 U6982 ( .A1(n5934), .A2(n5933), .ZN(U2874) );
  INV_X1 U6983 ( .A(n5935), .ZN(n5940) );
  AOI22_X1 U6984 ( .A1(n5962), .A2(DATAO_REG_29__SCAN_IN), .B1(n5940), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5936) );
  OAI21_X1 U6985 ( .B1(n6592), .B2(n6520), .A(n5936), .ZN(U2894) );
  AOI22_X1 U6986 ( .A1(n5962), .A2(DATAO_REG_28__SCAN_IN), .B1(n5940), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5937) );
  OAI21_X1 U6987 ( .B1(n6677), .B2(n6520), .A(n5937), .ZN(U2895) );
  INV_X1 U6988 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n6770) );
  AOI22_X1 U6989 ( .A1(n5940), .A2(EAX_REG_25__SCAN_IN), .B1(n5960), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n5938) );
  OAI21_X1 U6990 ( .B1(n6770), .B2(n5957), .A(n5938), .ZN(U2898) );
  AOI22_X1 U6991 ( .A1(n5962), .A2(DATAO_REG_24__SCAN_IN), .B1(n5940), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5939) );
  OAI21_X1 U6992 ( .B1(n6614), .B2(n6520), .A(n5939), .ZN(U2899) );
  AOI22_X1 U6993 ( .A1(n5962), .A2(DATAO_REG_23__SCAN_IN), .B1(n5940), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5941) );
  OAI21_X1 U6994 ( .B1(n6545), .B2(n6520), .A(n5941), .ZN(U2900) );
  AOI22_X1 U6995 ( .A1(n5960), .A2(LWORD_REG_15__SCAN_IN), .B1(n5962), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n5942) );
  OAI21_X1 U6996 ( .B1(n6704), .B2(n5965), .A(n5942), .ZN(U2908) );
  INV_X1 U6997 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n6759) );
  INV_X1 U6998 ( .A(LWORD_REG_14__SCAN_IN), .ZN(n5943) );
  OAI222_X1 U6999 ( .A1(n5957), .A2(n6759), .B1(n5965), .B2(n6686), .C1(n6520), 
        .C2(n5943), .ZN(U2909) );
  INV_X1 U7000 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n6768) );
  OAI222_X1 U7001 ( .A1(n5957), .A2(n6768), .B1(n5965), .B2(n3836), .C1(n6520), 
        .C2(n5944), .ZN(U2910) );
  AOI22_X1 U7002 ( .A1(n5960), .A2(LWORD_REG_12__SCAN_IN), .B1(n5962), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n5945) );
  OAI21_X1 U7003 ( .B1(n5946), .B2(n5965), .A(n5945), .ZN(U2911) );
  INV_X1 U7004 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n6624) );
  OAI222_X1 U7005 ( .A1(n6520), .A2(n6640), .B1(n5965), .B2(n5947), .C1(n6624), 
        .C2(n5957), .ZN(U2912) );
  AOI22_X1 U7006 ( .A1(n5960), .A2(LWORD_REG_10__SCAN_IN), .B1(n5962), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n5948) );
  OAI21_X1 U7007 ( .B1(n5949), .B2(n5965), .A(n5948), .ZN(U2913) );
  INV_X1 U7008 ( .A(EAX_REG_9__SCAN_IN), .ZN(n5951) );
  AOI22_X1 U7009 ( .A1(n5960), .A2(LWORD_REG_9__SCAN_IN), .B1(n5962), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n5950) );
  OAI21_X1 U7010 ( .B1(n5951), .B2(n5965), .A(n5950), .ZN(U2914) );
  AOI22_X1 U7011 ( .A1(n5960), .A2(LWORD_REG_8__SCAN_IN), .B1(n5962), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n5952) );
  OAI21_X1 U7012 ( .B1(n3776), .B2(n5965), .A(n5952), .ZN(U2915) );
  AOI22_X1 U7013 ( .A1(n5960), .A2(LWORD_REG_7__SCAN_IN), .B1(n5962), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n5953) );
  OAI21_X1 U7014 ( .B1(n4823), .B2(n5965), .A(n5953), .ZN(U2916) );
  AOI22_X1 U7015 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n5963), .B1(n5962), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n5954) );
  OAI21_X1 U7016 ( .B1(n3751), .B2(n5965), .A(n5954), .ZN(U2917) );
  INV_X1 U7017 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n6551) );
  INV_X1 U7018 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n5955) );
  OAI222_X1 U7019 ( .A1(n5957), .A2(n6551), .B1(n5965), .B2(n3733), .C1(n6520), 
        .C2(n5955), .ZN(U2918) );
  INV_X1 U7020 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n6589) );
  OAI222_X1 U7021 ( .A1(n5957), .A2(n6589), .B1(n5965), .B2(n3741), .C1(n6520), 
        .C2(n5956), .ZN(U2919) );
  AOI22_X1 U7022 ( .A1(n5960), .A2(LWORD_REG_3__SCAN_IN), .B1(n5962), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n5958) );
  OAI21_X1 U7023 ( .B1(n4700), .B2(n5965), .A(n5958), .ZN(U2920) );
  AOI22_X1 U7024 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n5963), .B1(n5962), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n5959) );
  OAI21_X1 U7025 ( .B1(n3719), .B2(n5965), .A(n5959), .ZN(U2921) );
  AOI22_X1 U7026 ( .A1(n5960), .A2(LWORD_REG_1__SCAN_IN), .B1(n5962), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n5961) );
  OAI21_X1 U7027 ( .B1(n3702), .B2(n5965), .A(n5961), .ZN(U2922) );
  AOI22_X1 U7028 ( .A1(n5963), .A2(LWORD_REG_0__SCAN_IN), .B1(n5962), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n5964) );
  OAI21_X1 U7029 ( .B1(n3710), .B2(n5965), .A(n5964), .ZN(U2923) );
  AOI22_X1 U7030 ( .A1(n5969), .A2(EAX_REG_25__SCAN_IN), .B1(
        UWORD_REG_9__SCAN_IN), .B2(n5968), .ZN(n5967) );
  NAND2_X1 U7031 ( .A1(n5966), .A2(DATAI_9_), .ZN(n5970) );
  NAND2_X1 U7032 ( .A1(n5967), .A2(n5970), .ZN(U2933) );
  AOI22_X1 U7033 ( .A1(n5969), .A2(EAX_REG_9__SCAN_IN), .B1(
        LWORD_REG_9__SCAN_IN), .B2(n5968), .ZN(n5971) );
  NAND2_X1 U7034 ( .A1(n5971), .A2(n5970), .ZN(U2948) );
  AOI22_X1 U7035 ( .A1(n4228), .A2(REIP_REG_11__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n6036), .ZN(n5978) );
  NAND2_X1 U7036 ( .A1(n5973), .A2(n5972), .ZN(n5975) );
  XNOR2_X1 U7037 ( .A(n5704), .B(n6052), .ZN(n5974) );
  XNOR2_X1 U7038 ( .A(n5975), .B(n5974), .ZN(n6049) );
  AOI22_X1 U7039 ( .A1(n5976), .A2(n6022), .B1(n6040), .B2(n6049), .ZN(n5977)
         );
  OAI211_X1 U7040 ( .C1(n6026), .C2(n5979), .A(n5978), .B(n5977), .ZN(U2975)
         );
  AOI22_X1 U7041 ( .A1(n4228), .A2(REIP_REG_9__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n6036), .ZN(n5985) );
  XNOR2_X1 U7042 ( .A(n5704), .B(n5981), .ZN(n5982) );
  XNOR2_X1 U7043 ( .A(n5980), .B(n5982), .ZN(n6055) );
  AOI22_X1 U7044 ( .A1(n6055), .A2(n6040), .B1(n6022), .B2(n5983), .ZN(n5984)
         );
  OAI211_X1 U7045 ( .C1(n6026), .C2(n5986), .A(n5985), .B(n5984), .ZN(U2977)
         );
  AOI22_X1 U7046 ( .A1(n4228), .A2(REIP_REG_8__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n6036), .ZN(n5993) );
  OAI21_X1 U7047 ( .B1(n5987), .B2(n5989), .A(n5988), .ZN(n5990) );
  INV_X1 U7048 ( .A(n5990), .ZN(n6063) );
  AOI22_X1 U7049 ( .A1(n6063), .A2(n6040), .B1(n6022), .B2(n5991), .ZN(n5992)
         );
  OAI211_X1 U7050 ( .C1(n6026), .C2(n5994), .A(n5993), .B(n5992), .ZN(U2978)
         );
  AOI22_X1 U7051 ( .A1(n4228), .A2(REIP_REG_7__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n6036), .ZN(n6001) );
  OR2_X1 U7052 ( .A1(n5996), .A2(n5995), .ZN(n5997) );
  AND2_X1 U7053 ( .A1(n5998), .A2(n5997), .ZN(n6067) );
  AOI22_X1 U7054 ( .A1(n5999), .A2(n5700), .B1(n6040), .B2(n6067), .ZN(n6000)
         );
  OAI211_X1 U7055 ( .C1(n6002), .C2(n6045), .A(n6001), .B(n6000), .ZN(U2979)
         );
  AOI22_X1 U7056 ( .A1(n4228), .A2(REIP_REG_6__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6036), .ZN(n6009) );
  OAI21_X1 U7057 ( .B1(n6005), .B2(n6004), .A(n6003), .ZN(n6006) );
  INV_X1 U7058 ( .A(n6006), .ZN(n6075) );
  AOI22_X1 U7059 ( .A1(n6075), .A2(n6040), .B1(n6022), .B2(n6007), .ZN(n6008)
         );
  OAI211_X1 U7060 ( .C1(n6026), .C2(n6010), .A(n6009), .B(n6008), .ZN(U2980)
         );
  AOI22_X1 U7061 ( .A1(n4228), .A2(REIP_REG_5__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n6036), .ZN(n6015) );
  INV_X1 U7062 ( .A(n6011), .ZN(n6012) );
  AOI22_X1 U7063 ( .A1(n4663), .A2(n6013), .B1(n6012), .B2(n6040), .ZN(n6014)
         );
  OAI211_X1 U7064 ( .C1(n6016), .C2(n6045), .A(n6015), .B(n6014), .ZN(U2981)
         );
  AOI22_X1 U7065 ( .A1(n4228), .A2(REIP_REG_4__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n6036), .ZN(n6024) );
  OAI21_X1 U7066 ( .B1(n6019), .B2(n6018), .A(n6017), .ZN(n6020) );
  INV_X1 U7067 ( .A(n6020), .ZN(n6083) );
  AOI22_X1 U7068 ( .A1(n6083), .A2(n6040), .B1(n6022), .B2(n6021), .ZN(n6023)
         );
  OAI211_X1 U7069 ( .C1(n6026), .C2(n6025), .A(n6024), .B(n6023), .ZN(U2982)
         );
  AOI22_X1 U7070 ( .A1(n4228), .A2(REIP_REG_3__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n6036), .ZN(n6034) );
  OAI21_X1 U7071 ( .B1(n6027), .B2(n6029), .A(n6028), .ZN(n6030) );
  INV_X1 U7072 ( .A(n6030), .ZN(n6089) );
  INV_X1 U7073 ( .A(n6031), .ZN(n6032) );
  AOI22_X1 U7074 ( .A1(n6040), .A2(n6089), .B1(n6032), .B2(n5700), .ZN(n6033)
         );
  OAI211_X1 U7075 ( .C1(n6035), .C2(n6045), .A(n6034), .B(n6033), .ZN(U2983)
         );
  AOI22_X1 U7076 ( .A1(n4228), .A2(REIP_REG_2__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n6036), .ZN(n6044) );
  XNOR2_X1 U7077 ( .A(n6038), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6039)
         );
  XNOR2_X1 U7078 ( .A(n6037), .B(n6039), .ZN(n6102) );
  INV_X1 U7079 ( .A(n6102), .ZN(n6041) );
  AOI22_X1 U7080 ( .A1(n5700), .A2(n6042), .B1(n6041), .B2(n6040), .ZN(n6043)
         );
  OAI211_X1 U7081 ( .C1(n6046), .C2(n6045), .A(n6044), .B(n6043), .ZN(U2984)
         );
  INV_X1 U7082 ( .A(n6047), .ZN(n6051) );
  AOI222_X1 U7083 ( .A1(n6049), .A2(n6090), .B1(n6099), .B2(n6048), .C1(
        REIP_REG_11__SCAN_IN), .C2(n4228), .ZN(n6050) );
  OAI221_X1 U7084 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6053), .C1(
        n6052), .C2(n6051), .A(n6050), .ZN(U3007) );
  AOI22_X1 U7085 ( .A1(n6099), .A2(n6054), .B1(n4228), .B2(REIP_REG_9__SCAN_IN), .ZN(n6058) );
  AOI22_X1 U7086 ( .A1(n6056), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .B1(n6090), 
        .B2(n6055), .ZN(n6057) );
  OAI211_X1 U7087 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6059), .A(n6058), 
        .B(n6057), .ZN(U3009) );
  AOI22_X1 U7088 ( .A1(n6099), .A2(n6060), .B1(n4228), .B2(REIP_REG_8__SCAN_IN), .ZN(n6065) );
  AOI21_X1 U7089 ( .B1(n6072), .B2(n6767), .A(n6061), .ZN(n6062) );
  AOI22_X1 U7090 ( .A1(n6063), .A2(n6090), .B1(n6068), .B2(n6062), .ZN(n6064)
         );
  OAI211_X1 U7091 ( .C1(n6767), .C2(n6071), .A(n6065), .B(n6064), .ZN(U3010)
         );
  AOI22_X1 U7092 ( .A1(n6099), .A2(n6066), .B1(n4228), .B2(REIP_REG_7__SCAN_IN), .ZN(n6070) );
  AOI22_X1 U7093 ( .A1(n6068), .A2(n6072), .B1(n6090), .B2(n6067), .ZN(n6069)
         );
  OAI211_X1 U7094 ( .C1(n6072), .C2(n6071), .A(n6070), .B(n6069), .ZN(U3011)
         );
  AOI22_X1 U7095 ( .A1(n6099), .A2(n6073), .B1(n4228), .B2(REIP_REG_6__SCAN_IN), .ZN(n6080) );
  AOI22_X1 U7096 ( .A1(n6075), .A2(n6090), .B1(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .B2(n6074), .ZN(n6079) );
  NAND3_X1 U7097 ( .A1(n6077), .A2(n6654), .A3(n6076), .ZN(n6078) );
  NAND3_X1 U7098 ( .A1(n6080), .A2(n6079), .A3(n6078), .ZN(U3012) );
  OAI21_X1 U7099 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6081), .ZN(n6086) );
  AOI22_X1 U7100 ( .A1(n6099), .A2(n6082), .B1(n4228), .B2(REIP_REG_4__SCAN_IN), .ZN(n6085) );
  AOI22_X1 U7101 ( .A1(n6091), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .B1(n6090), 
        .B2(n6083), .ZN(n6084) );
  OAI211_X1 U7102 ( .C1(n6094), .C2(n6086), .A(n6085), .B(n6084), .ZN(U3014)
         );
  INV_X1 U7103 ( .A(n6087), .ZN(n6088) );
  AOI22_X1 U7104 ( .A1(n6099), .A2(n6088), .B1(n4228), .B2(REIP_REG_3__SCAN_IN), .ZN(n6093) );
  AOI22_X1 U7105 ( .A1(n6091), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .B1(n6090), 
        .B2(n6089), .ZN(n6092) );
  OAI211_X1 U7106 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n6094), .A(n6093), 
        .B(n6092), .ZN(U3015) );
  INV_X1 U7107 ( .A(n6095), .ZN(n6101) );
  OAI21_X1 U7108 ( .B1(n6097), .B2(n6107), .A(n6096), .ZN(n6100) );
  AOI22_X1 U7109 ( .A1(n6101), .A2(n6100), .B1(n6099), .B2(n6098), .ZN(n6111)
         );
  OAI22_X1 U7110 ( .A1(n6104), .A2(n6107), .B1(n6103), .B2(n6102), .ZN(n6105)
         );
  INV_X1 U7111 ( .A(n6105), .ZN(n6110) );
  NAND2_X1 U7112 ( .A1(n4228), .A2(REIP_REG_2__SCAN_IN), .ZN(n6109) );
  NAND3_X1 U7113 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6107), .A3(n6106), 
        .ZN(n6108) );
  NAND4_X1 U7114 ( .A1(n6111), .A2(n6110), .A3(n6109), .A4(n6108), .ZN(U3016)
         );
  NOR2_X1 U7115 ( .A1(n6113), .A2(n6112), .ZN(U3019) );
  NAND2_X1 U7116 ( .A1(n6116), .A2(n6254), .ZN(n6114) );
  INV_X1 U7117 ( .A(n6330), .ZN(n6115) );
  NAND2_X1 U7118 ( .A1(n6115), .A2(n6412), .ZN(n6121) );
  INV_X1 U7119 ( .A(n6121), .ZN(n6143) );
  AOI22_X1 U7120 ( .A1(n6332), .A2(n6143), .B1(n6228), .B2(n6142), .ZN(n6129)
         );
  NAND2_X1 U7121 ( .A1(n6117), .A2(n6116), .ZN(n6118) );
  OAI21_X1 U7122 ( .B1(n3114), .B2(n6118), .A(n6335), .ZN(n6127) );
  OR2_X1 U7123 ( .A1(n6120), .A2(n6119), .ZN(n6122) );
  NAND2_X1 U7124 ( .A1(n6122), .A2(n6121), .ZN(n6124) );
  NAND2_X1 U7125 ( .A1(n6340), .A2(n6125), .ZN(n6123) );
  OAI211_X1 U7126 ( .C1(n6127), .C2(n6124), .A(n6342), .B(n6123), .ZN(n6145)
         );
  INV_X1 U7127 ( .A(n6124), .ZN(n6126) );
  OAI22_X1 U7128 ( .A1(n6127), .A2(n6126), .B1(n6125), .B2(n6522), .ZN(n6144)
         );
  AOI22_X1 U7129 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6145), .B1(n6347), 
        .B2(n6144), .ZN(n6128) );
  OAI211_X1 U7130 ( .C1(n6231), .C2(n6180), .A(n6129), .B(n6128), .ZN(U3044)
         );
  AOI22_X1 U7131 ( .A1(n6352), .A2(n6143), .B1(n6351), .B2(n6142), .ZN(n6131)
         );
  AOI22_X1 U7132 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6145), .B1(n6353), 
        .B2(n6144), .ZN(n6130) );
  OAI211_X1 U7133 ( .C1(n6356), .C2(n6180), .A(n6131), .B(n6130), .ZN(U3045)
         );
  AOI22_X1 U7134 ( .A1(n6358), .A2(n6143), .B1(n6234), .B2(n6142), .ZN(n6133)
         );
  AOI22_X1 U7135 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6145), .B1(n6359), 
        .B2(n6144), .ZN(n6132) );
  OAI211_X1 U7136 ( .C1(n6237), .C2(n6180), .A(n6133), .B(n6132), .ZN(U3046)
         );
  AOI22_X1 U7137 ( .A1(n6364), .A2(n6143), .B1(n6363), .B2(n6142), .ZN(n6135)
         );
  AOI22_X1 U7138 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6145), .B1(n6365), 
        .B2(n6144), .ZN(n6134) );
  OAI211_X1 U7139 ( .C1(n6368), .C2(n6180), .A(n6135), .B(n6134), .ZN(U3047)
         );
  AOI22_X1 U7140 ( .A1(n6371), .A2(n6143), .B1(n6370), .B2(n6142), .ZN(n6137)
         );
  AOI22_X1 U7141 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6145), .B1(n6372), 
        .B2(n6144), .ZN(n6136) );
  OAI211_X1 U7142 ( .C1(n6376), .C2(n6180), .A(n6137), .B(n6136), .ZN(U3048)
         );
  AOI22_X1 U7143 ( .A1(n6378), .A2(n6143), .B1(n6276), .B2(n6142), .ZN(n6139)
         );
  AOI22_X1 U7144 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6145), .B1(n6379), 
        .B2(n6144), .ZN(n6138) );
  OAI211_X1 U7145 ( .C1(n6534), .C2(n6180), .A(n6139), .B(n6138), .ZN(U3049)
         );
  AOI22_X1 U7146 ( .A1(n6383), .A2(n6143), .B1(n6280), .B2(n6142), .ZN(n6141)
         );
  AOI22_X1 U7147 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6145), .B1(n6384), 
        .B2(n6144), .ZN(n6140) );
  OAI211_X1 U7148 ( .C1(n6283), .C2(n6180), .A(n6141), .B(n6140), .ZN(U3050)
         );
  AOI22_X1 U7149 ( .A1(n6391), .A2(n6143), .B1(n6249), .B2(n6142), .ZN(n6147)
         );
  AOI22_X1 U7150 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6145), .B1(n6393), 
        .B2(n6144), .ZN(n6146) );
  OAI211_X1 U7151 ( .C1(n6253), .C2(n6180), .A(n6147), .B(n6146), .ZN(U3051)
         );
  INV_X1 U7152 ( .A(n6148), .ZN(n6149) );
  OAI22_X1 U7153 ( .A1(n6185), .A2(n6150), .B1(n6300), .B2(n6149), .ZN(n6175)
         );
  NAND3_X1 U7154 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6412), .A3(n6151), .ZN(n6190) );
  NOR2_X1 U7155 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6190), .ZN(n6176)
         );
  AOI22_X1 U7156 ( .A1(n6347), .A2(n6175), .B1(n6332), .B2(n6176), .ZN(n6162)
         );
  INV_X1 U7157 ( .A(n6176), .ZN(n6153) );
  AOI211_X1 U7158 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6153), .A(n6290), .B(
        n6152), .ZN(n6159) );
  AOI21_X1 U7159 ( .B1(n6188), .B2(STATEBS16_REG_SCAN_IN), .A(n6340), .ZN(
        n6181) );
  NAND2_X1 U7160 ( .A1(n6155), .A2(n6218), .ZN(n6156) );
  OAI211_X1 U7161 ( .C1(n6157), .C2(n6180), .A(n6181), .B(n6156), .ZN(n6158)
         );
  NAND2_X1 U7162 ( .A1(n6159), .A2(n6158), .ZN(n6177) );
  INV_X1 U7163 ( .A(n6188), .ZN(n6160) );
  NOR2_X2 U7164 ( .A1(n6160), .A2(n6187), .ZN(n6212) );
  AOI22_X1 U7165 ( .A1(n6177), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n6331), 
        .B2(n6212), .ZN(n6161) );
  OAI211_X1 U7166 ( .C1(n6350), .C2(n6180), .A(n6162), .B(n6161), .ZN(U3052)
         );
  AOI22_X1 U7167 ( .A1(n6353), .A2(n6175), .B1(n6352), .B2(n6176), .ZN(n6164)
         );
  AOI22_X1 U7168 ( .A1(n6177), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n6305), 
        .B2(n6212), .ZN(n6163) );
  OAI211_X1 U7169 ( .C1(n6308), .C2(n6180), .A(n6164), .B(n6163), .ZN(U3053)
         );
  AOI22_X1 U7170 ( .A1(n6359), .A2(n6175), .B1(n6358), .B2(n6176), .ZN(n6166)
         );
  AOI22_X1 U7171 ( .A1(n6177), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n6357), 
        .B2(n6212), .ZN(n6165) );
  OAI211_X1 U7172 ( .C1(n6362), .C2(n6180), .A(n6166), .B(n6165), .ZN(U3054)
         );
  AOI22_X1 U7173 ( .A1(n6364), .A2(n6176), .B1(n6365), .B2(n6175), .ZN(n6168)
         );
  AOI22_X1 U7174 ( .A1(n6177), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n6311), 
        .B2(n6212), .ZN(n6167) );
  OAI211_X1 U7175 ( .C1(n6314), .C2(n6180), .A(n6168), .B(n6167), .ZN(U3055)
         );
  AOI22_X1 U7176 ( .A1(n6372), .A2(n6175), .B1(n6371), .B2(n6176), .ZN(n6170)
         );
  AOI22_X1 U7177 ( .A1(n6177), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n6315), 
        .B2(n6212), .ZN(n6169) );
  OAI211_X1 U7178 ( .C1(n6318), .C2(n6180), .A(n6170), .B(n6169), .ZN(U3056)
         );
  AOI22_X1 U7179 ( .A1(n6379), .A2(n6175), .B1(n6378), .B2(n6176), .ZN(n6172)
         );
  AOI22_X1 U7180 ( .A1(n6177), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n6377), 
        .B2(n6212), .ZN(n6171) );
  OAI211_X1 U7181 ( .C1(n6537), .C2(n6180), .A(n6172), .B(n6171), .ZN(U3057)
         );
  AOI22_X1 U7182 ( .A1(n6384), .A2(n6175), .B1(n6383), .B2(n6176), .ZN(n6174)
         );
  AOI22_X1 U7183 ( .A1(n6177), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n6382), 
        .B2(n6212), .ZN(n6173) );
  OAI211_X1 U7184 ( .C1(n6387), .C2(n6180), .A(n6174), .B(n6173), .ZN(U3058)
         );
  AOI22_X1 U7185 ( .A1(n6391), .A2(n6176), .B1(n6393), .B2(n6175), .ZN(n6179)
         );
  AOI22_X1 U7186 ( .A1(n6177), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n6389), 
        .B2(n6212), .ZN(n6178) );
  OAI211_X1 U7187 ( .C1(n6397), .C2(n6180), .A(n6179), .B(n6178), .ZN(U3059)
         );
  INV_X1 U7188 ( .A(n6181), .ZN(n6192) );
  OR2_X1 U7189 ( .A1(n3707), .A2(n6182), .ZN(n6258) );
  NOR2_X1 U7190 ( .A1(n6183), .A2(n6190), .ZN(n6211) );
  INV_X1 U7191 ( .A(n6211), .ZN(n6184) );
  OAI21_X1 U7192 ( .B1(n6185), .B2(n6258), .A(n6184), .ZN(n6189) );
  OAI21_X1 U7193 ( .B1(n6192), .B2(n6189), .A(n6342), .ZN(n6186) );
  INV_X1 U7194 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n6595) );
  AOI22_X1 U7195 ( .A1(n6332), .A2(n6211), .B1(n6331), .B2(n6248), .ZN(n6194)
         );
  INV_X1 U7196 ( .A(n6189), .ZN(n6191) );
  OAI22_X1 U7197 ( .A1(n6192), .A2(n6191), .B1(n6190), .B2(n6522), .ZN(n6213)
         );
  AOI22_X1 U7198 ( .A1(n6347), .A2(n6213), .B1(n6228), .B2(n6212), .ZN(n6193)
         );
  OAI211_X1 U7199 ( .C1(n6216), .C2(n6595), .A(n6194), .B(n6193), .ZN(U3060)
         );
  INV_X1 U7200 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n6827) );
  AOI22_X1 U7201 ( .A1(n6352), .A2(n6211), .B1(n6305), .B2(n6248), .ZN(n6196)
         );
  AOI22_X1 U7202 ( .A1(n6353), .A2(n6213), .B1(n6351), .B2(n6212), .ZN(n6195)
         );
  OAI211_X1 U7203 ( .C1(n6216), .C2(n6827), .A(n6196), .B(n6195), .ZN(U3061)
         );
  INV_X1 U7204 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n6199) );
  AOI22_X1 U7205 ( .A1(n6358), .A2(n6211), .B1(n6357), .B2(n6248), .ZN(n6198)
         );
  AOI22_X1 U7206 ( .A1(n6359), .A2(n6213), .B1(n6234), .B2(n6212), .ZN(n6197)
         );
  OAI211_X1 U7207 ( .C1(n6216), .C2(n6199), .A(n6198), .B(n6197), .ZN(U3062)
         );
  INV_X1 U7208 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n6202) );
  AOI22_X1 U7209 ( .A1(n6364), .A2(n6211), .B1(n6311), .B2(n6248), .ZN(n6201)
         );
  AOI22_X1 U7210 ( .A1(n6213), .A2(n6365), .B1(n6363), .B2(n6212), .ZN(n6200)
         );
  OAI211_X1 U7211 ( .C1(n6216), .C2(n6202), .A(n6201), .B(n6200), .ZN(U3063)
         );
  INV_X1 U7212 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n6205) );
  AOI22_X1 U7213 ( .A1(n6371), .A2(n6211), .B1(n6315), .B2(n6248), .ZN(n6204)
         );
  AOI22_X1 U7214 ( .A1(n6372), .A2(n6213), .B1(n6370), .B2(n6212), .ZN(n6203)
         );
  OAI211_X1 U7215 ( .C1(n6216), .C2(n6205), .A(n6204), .B(n6203), .ZN(U3064)
         );
  INV_X1 U7216 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n6660) );
  AOI22_X1 U7217 ( .A1(n6378), .A2(n6211), .B1(n6377), .B2(n6248), .ZN(n6207)
         );
  AOI22_X1 U7218 ( .A1(n6379), .A2(n6213), .B1(n6276), .B2(n6212), .ZN(n6206)
         );
  OAI211_X1 U7219 ( .C1(n6216), .C2(n6660), .A(n6207), .B(n6206), .ZN(U3065)
         );
  INV_X1 U7220 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6210) );
  AOI22_X1 U7221 ( .A1(n6383), .A2(n6211), .B1(n6382), .B2(n6248), .ZN(n6209)
         );
  AOI22_X1 U7222 ( .A1(n6384), .A2(n6213), .B1(n6280), .B2(n6212), .ZN(n6208)
         );
  OAI211_X1 U7223 ( .C1(n6216), .C2(n6210), .A(n6209), .B(n6208), .ZN(U3066)
         );
  INV_X1 U7224 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n6611) );
  AOI22_X1 U7225 ( .A1(n6391), .A2(n6211), .B1(n6389), .B2(n6248), .ZN(n6215)
         );
  AOI22_X1 U7226 ( .A1(n6213), .A2(n6393), .B1(n6249), .B2(n6212), .ZN(n6214)
         );
  OAI211_X1 U7227 ( .C1(n6216), .C2(n6611), .A(n6215), .B(n6214), .ZN(U3067)
         );
  NAND3_X1 U7228 ( .A1(n6219), .A2(n6218), .A3(n6335), .ZN(n6220) );
  OAI21_X1 U7229 ( .B1(n6300), .B2(n6221), .A(n6220), .ZN(n6246) );
  NOR2_X1 U7230 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6263), .ZN(n6247)
         );
  AOI22_X1 U7231 ( .A1(n6347), .A2(n6246), .B1(n6332), .B2(n6247), .ZN(n6230)
         );
  OAI21_X1 U7232 ( .B1(n6817), .B2(n6247), .A(n6222), .ZN(n6225) );
  INV_X1 U7233 ( .A(n6289), .ZN(n6279) );
  AOI211_X1 U7234 ( .C1(n6293), .C2(n6223), .A(n6279), .B(n6248), .ZN(n6224)
         );
  NOR2_X1 U7235 ( .A1(n6225), .A2(n6224), .ZN(n6227) );
  NAND2_X1 U7236 ( .A1(n6227), .A2(n6226), .ZN(n6250) );
  AOI22_X1 U7237 ( .A1(n6250), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6228), 
        .B2(n6248), .ZN(n6229) );
  OAI211_X1 U7238 ( .C1(n6231), .C2(n6289), .A(n6230), .B(n6229), .ZN(U3068)
         );
  AOI22_X1 U7239 ( .A1(n6353), .A2(n6246), .B1(n6352), .B2(n6247), .ZN(n6233)
         );
  AOI22_X1 U7240 ( .A1(n6250), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6351), 
        .B2(n6248), .ZN(n6232) );
  OAI211_X1 U7241 ( .C1(n6356), .C2(n6289), .A(n6233), .B(n6232), .ZN(U3069)
         );
  AOI22_X1 U7242 ( .A1(n6359), .A2(n6246), .B1(n6358), .B2(n6247), .ZN(n6236)
         );
  AOI22_X1 U7243 ( .A1(n6250), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6234), 
        .B2(n6248), .ZN(n6235) );
  OAI211_X1 U7244 ( .C1(n6237), .C2(n6289), .A(n6236), .B(n6235), .ZN(U3070)
         );
  AOI22_X1 U7245 ( .A1(n6364), .A2(n6247), .B1(n6365), .B2(n6246), .ZN(n6239)
         );
  AOI22_X1 U7246 ( .A1(n6250), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6363), 
        .B2(n6248), .ZN(n6238) );
  OAI211_X1 U7247 ( .C1(n6368), .C2(n6289), .A(n6239), .B(n6238), .ZN(U3071)
         );
  AOI22_X1 U7248 ( .A1(n6372), .A2(n6246), .B1(n6371), .B2(n6247), .ZN(n6241)
         );
  AOI22_X1 U7249 ( .A1(n6250), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6370), 
        .B2(n6248), .ZN(n6240) );
  OAI211_X1 U7250 ( .C1(n6376), .C2(n6289), .A(n6241), .B(n6240), .ZN(U3072)
         );
  AOI22_X1 U7251 ( .A1(n6379), .A2(n6246), .B1(n6378), .B2(n6247), .ZN(n6243)
         );
  AOI22_X1 U7252 ( .A1(n6250), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6276), 
        .B2(n6248), .ZN(n6242) );
  OAI211_X1 U7253 ( .C1(n6534), .C2(n6289), .A(n6243), .B(n6242), .ZN(U3073)
         );
  AOI22_X1 U7254 ( .A1(n6384), .A2(n6246), .B1(n6383), .B2(n6247), .ZN(n6245)
         );
  AOI22_X1 U7255 ( .A1(n6250), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6280), 
        .B2(n6248), .ZN(n6244) );
  OAI211_X1 U7256 ( .C1(n6283), .C2(n6289), .A(n6245), .B(n6244), .ZN(U3074)
         );
  AOI22_X1 U7257 ( .A1(n6391), .A2(n6247), .B1(n6393), .B2(n6246), .ZN(n6252)
         );
  AOI22_X1 U7258 ( .A1(n6250), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6249), 
        .B2(n6248), .ZN(n6251) );
  OAI211_X1 U7259 ( .C1(n6253), .C2(n6289), .A(n6252), .B(n6251), .ZN(U3075)
         );
  INV_X1 U7260 ( .A(n6257), .ZN(n6284) );
  AOI22_X1 U7261 ( .A1(n6332), .A2(n6284), .B1(n6331), .B2(n6295), .ZN(n6267)
         );
  NAND2_X1 U7262 ( .A1(n6256), .A2(n6335), .ZN(n6265) );
  OAI21_X1 U7263 ( .B1(n6259), .B2(n6258), .A(n6257), .ZN(n6262) );
  OR2_X1 U7264 ( .A1(n6265), .A2(n6262), .ZN(n6260) );
  OAI211_X1 U7265 ( .C1(n6335), .C2(n6261), .A(n6342), .B(n6260), .ZN(n6286)
         );
  INV_X1 U7266 ( .A(n6262), .ZN(n6264) );
  OAI22_X1 U7267 ( .A1(n6265), .A2(n6264), .B1(n6263), .B2(n6522), .ZN(n6285)
         );
  AOI22_X1 U7268 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6286), .B1(n6347), 
        .B2(n6285), .ZN(n6266) );
  OAI211_X1 U7269 ( .C1(n6350), .C2(n6289), .A(n6267), .B(n6266), .ZN(U3076)
         );
  AOI22_X1 U7270 ( .A1(n6352), .A2(n6284), .B1(n6305), .B2(n6295), .ZN(n6269)
         );
  AOI22_X1 U7271 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6286), .B1(n6353), 
        .B2(n6285), .ZN(n6268) );
  OAI211_X1 U7272 ( .C1(n6308), .C2(n6289), .A(n6269), .B(n6268), .ZN(U3077)
         );
  AOI22_X1 U7273 ( .A1(n6358), .A2(n6284), .B1(n6357), .B2(n6295), .ZN(n6271)
         );
  AOI22_X1 U7274 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6286), .B1(n6359), 
        .B2(n6285), .ZN(n6270) );
  OAI211_X1 U7275 ( .C1(n6362), .C2(n6289), .A(n6271), .B(n6270), .ZN(U3078)
         );
  AOI22_X1 U7276 ( .A1(n6364), .A2(n6284), .B1(n6363), .B2(n6279), .ZN(n6273)
         );
  AOI22_X1 U7277 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6286), .B1(n6365), 
        .B2(n6285), .ZN(n6272) );
  OAI211_X1 U7278 ( .C1(n6368), .C2(n6329), .A(n6273), .B(n6272), .ZN(U3079)
         );
  AOI22_X1 U7279 ( .A1(n6371), .A2(n6284), .B1(n6315), .B2(n6295), .ZN(n6275)
         );
  AOI22_X1 U7280 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6286), .B1(n6372), 
        .B2(n6285), .ZN(n6274) );
  OAI211_X1 U7281 ( .C1(n6318), .C2(n6289), .A(n6275), .B(n6274), .ZN(U3080)
         );
  AOI22_X1 U7282 ( .A1(n6378), .A2(n6284), .B1(n6276), .B2(n6279), .ZN(n6278)
         );
  AOI22_X1 U7283 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6286), .B1(n6379), 
        .B2(n6285), .ZN(n6277) );
  OAI211_X1 U7284 ( .C1(n6534), .C2(n6329), .A(n6278), .B(n6277), .ZN(U3081)
         );
  AOI22_X1 U7285 ( .A1(n6383), .A2(n6284), .B1(n6280), .B2(n6279), .ZN(n6282)
         );
  AOI22_X1 U7286 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6286), .B1(n6384), 
        .B2(n6285), .ZN(n6281) );
  OAI211_X1 U7287 ( .C1(n6283), .C2(n6329), .A(n6282), .B(n6281), .ZN(U3082)
         );
  AOI22_X1 U7288 ( .A1(n6391), .A2(n6284), .B1(n6389), .B2(n6295), .ZN(n6288)
         );
  AOI22_X1 U7289 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6286), .B1(n6393), 
        .B2(n6285), .ZN(n6287) );
  OAI211_X1 U7290 ( .C1(n6397), .C2(n6289), .A(n6288), .B(n6287), .ZN(U3083)
         );
  INV_X1 U7291 ( .A(n6290), .ZN(n6292) );
  OAI22_X1 U7292 ( .A1(n6293), .A2(n6297), .B1(n6292), .B2(n6291), .ZN(n6323)
         );
  NOR2_X1 U7293 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6294), .ZN(n6324)
         );
  AOI22_X1 U7294 ( .A1(n6347), .A2(n6323), .B1(n6332), .B2(n6324), .ZN(n6304)
         );
  OR2_X1 U7295 ( .A1(n6817), .A2(n6324), .ZN(n6301) );
  OAI21_X1 U7296 ( .B1(n6325), .B2(n6295), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6296) );
  OAI211_X1 U7297 ( .C1(n6298), .C2(n6297), .A(n6296), .B(n6335), .ZN(n6299)
         );
  NAND4_X1 U7298 ( .A1(n6302), .A2(n6301), .A3(n6300), .A4(n6299), .ZN(n6326)
         );
  AOI22_X1 U7299 ( .A1(n6326), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6325), 
        .B2(n6331), .ZN(n6303) );
  OAI211_X1 U7300 ( .C1(n6350), .C2(n6329), .A(n6304), .B(n6303), .ZN(U3084)
         );
  AOI22_X1 U7301 ( .A1(n6353), .A2(n6323), .B1(n6352), .B2(n6324), .ZN(n6307)
         );
  AOI22_X1 U7302 ( .A1(n6326), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6325), 
        .B2(n6305), .ZN(n6306) );
  OAI211_X1 U7303 ( .C1(n6308), .C2(n6329), .A(n6307), .B(n6306), .ZN(U3085)
         );
  AOI22_X1 U7304 ( .A1(n6359), .A2(n6323), .B1(n6358), .B2(n6324), .ZN(n6310)
         );
  AOI22_X1 U7305 ( .A1(n6326), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6325), 
        .B2(n6357), .ZN(n6309) );
  OAI211_X1 U7306 ( .C1(n6362), .C2(n6329), .A(n6310), .B(n6309), .ZN(U3086)
         );
  AOI22_X1 U7307 ( .A1(n6364), .A2(n6324), .B1(n6365), .B2(n6323), .ZN(n6313)
         );
  AOI22_X1 U7308 ( .A1(n6326), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6325), 
        .B2(n6311), .ZN(n6312) );
  OAI211_X1 U7309 ( .C1(n6314), .C2(n6329), .A(n6313), .B(n6312), .ZN(U3087)
         );
  AOI22_X1 U7310 ( .A1(n6372), .A2(n6323), .B1(n6371), .B2(n6324), .ZN(n6317)
         );
  AOI22_X1 U7311 ( .A1(n6326), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6325), 
        .B2(n6315), .ZN(n6316) );
  OAI211_X1 U7312 ( .C1(n6318), .C2(n6329), .A(n6317), .B(n6316), .ZN(U3088)
         );
  AOI22_X1 U7313 ( .A1(n6379), .A2(n6323), .B1(n6378), .B2(n6324), .ZN(n6320)
         );
  AOI22_X1 U7314 ( .A1(n6326), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6325), 
        .B2(n6377), .ZN(n6319) );
  OAI211_X1 U7315 ( .C1(n6537), .C2(n6329), .A(n6320), .B(n6319), .ZN(U3089)
         );
  AOI22_X1 U7316 ( .A1(n6384), .A2(n6323), .B1(n6383), .B2(n6324), .ZN(n6322)
         );
  AOI22_X1 U7317 ( .A1(n6326), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6325), 
        .B2(n6382), .ZN(n6321) );
  OAI211_X1 U7318 ( .C1(n6387), .C2(n6329), .A(n6322), .B(n6321), .ZN(U3090)
         );
  AOI22_X1 U7319 ( .A1(n6391), .A2(n6324), .B1(n6393), .B2(n6323), .ZN(n6328)
         );
  AOI22_X1 U7320 ( .A1(n6326), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6325), 
        .B2(n6389), .ZN(n6327) );
  OAI211_X1 U7321 ( .C1(n6397), .C2(n6329), .A(n6328), .B(n6327), .ZN(U3091)
         );
  NOR2_X1 U7322 ( .A1(n6412), .A2(n6330), .ZN(n6390) );
  AOI22_X1 U7323 ( .A1(n6332), .A2(n6390), .B1(n6331), .B2(n6388), .ZN(n6349)
         );
  OR2_X1 U7324 ( .A1(n6334), .A2(n6333), .ZN(n6336) );
  AND2_X1 U7325 ( .A1(n6336), .A2(n6335), .ZN(n6343) );
  AOI21_X1 U7326 ( .B1(n6338), .B2(n6337), .A(n6390), .ZN(n6345) );
  NAND2_X1 U7327 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6339), .ZN(n6344) );
  AOI22_X1 U7328 ( .A1(n6343), .A2(n6345), .B1(n6344), .B2(n6340), .ZN(n6341)
         );
  NAND2_X1 U7329 ( .A1(n6342), .A2(n6341), .ZN(n6394) );
  INV_X1 U7330 ( .A(n6343), .ZN(n6346) );
  OAI22_X1 U7331 ( .A1(n6346), .A2(n6345), .B1(n6344), .B2(n6522), .ZN(n6392)
         );
  AOI22_X1 U7332 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6394), .B1(n6347), 
        .B2(n6392), .ZN(n6348) );
  OAI211_X1 U7333 ( .C1(n6533), .C2(n6350), .A(n6349), .B(n6348), .ZN(U3108)
         );
  AOI22_X1 U7334 ( .A1(n6352), .A2(n6390), .B1(n6351), .B2(n6369), .ZN(n6355)
         );
  AOI22_X1 U7335 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6394), .B1(n6353), 
        .B2(n6392), .ZN(n6354) );
  OAI211_X1 U7336 ( .C1(n6356), .C2(n6375), .A(n6355), .B(n6354), .ZN(U3109)
         );
  AOI22_X1 U7337 ( .A1(n6358), .A2(n6390), .B1(n6357), .B2(n6388), .ZN(n6361)
         );
  AOI22_X1 U7338 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6394), .B1(n6359), 
        .B2(n6392), .ZN(n6360) );
  OAI211_X1 U7339 ( .C1(n6533), .C2(n6362), .A(n6361), .B(n6360), .ZN(U3110)
         );
  AOI22_X1 U7340 ( .A1(n6364), .A2(n6390), .B1(n6363), .B2(n6369), .ZN(n6367)
         );
  AOI22_X1 U7341 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6394), .B1(n6365), 
        .B2(n6392), .ZN(n6366) );
  OAI211_X1 U7342 ( .C1(n6368), .C2(n6375), .A(n6367), .B(n6366), .ZN(U3111)
         );
  AOI22_X1 U7343 ( .A1(n6371), .A2(n6390), .B1(n6370), .B2(n6369), .ZN(n6374)
         );
  AOI22_X1 U7344 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6394), .B1(n6372), 
        .B2(n6392), .ZN(n6373) );
  OAI211_X1 U7345 ( .C1(n6376), .C2(n6375), .A(n6374), .B(n6373), .ZN(U3112)
         );
  AOI22_X1 U7346 ( .A1(n6378), .A2(n6390), .B1(n6377), .B2(n6388), .ZN(n6381)
         );
  AOI22_X1 U7347 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6394), .B1(n6379), 
        .B2(n6392), .ZN(n6380) );
  OAI211_X1 U7348 ( .C1(n6537), .C2(n6533), .A(n6381), .B(n6380), .ZN(U3113)
         );
  AOI22_X1 U7349 ( .A1(n6383), .A2(n6390), .B1(n6382), .B2(n6388), .ZN(n6386)
         );
  AOI22_X1 U7350 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6394), .B1(n6384), 
        .B2(n6392), .ZN(n6385) );
  OAI211_X1 U7351 ( .C1(n6533), .C2(n6387), .A(n6386), .B(n6385), .ZN(U3114)
         );
  AOI22_X1 U7352 ( .A1(n6391), .A2(n6390), .B1(n6389), .B2(n6388), .ZN(n6396)
         );
  AOI22_X1 U7353 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6394), .B1(n6393), 
        .B2(n6392), .ZN(n6395) );
  OAI211_X1 U7354 ( .C1(n6533), .C2(n6397), .A(n6396), .B(n6395), .ZN(U3115)
         );
  AND2_X1 U7355 ( .A1(n6399), .A2(n6398), .ZN(n6413) );
  INV_X1 U7356 ( .A(n6399), .ZN(n6406) );
  NAND2_X1 U7357 ( .A1(n6399), .A2(n6400), .ZN(n6410) );
  AND3_X1 U7358 ( .A1(n6402), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6401), 
        .ZN(n6404) );
  NAND2_X1 U7359 ( .A1(n6404), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6408) );
  INV_X1 U7360 ( .A(n6403), .ZN(n6405) );
  OAI22_X1 U7361 ( .A1(n6406), .A2(n6405), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6404), .ZN(n6407) );
  NAND2_X1 U7362 ( .A1(n6408), .A2(n6407), .ZN(n6409) );
  AOI222_X1 U7363 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6410), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6409), .C1(n6410), .C2(n6409), 
        .ZN(n6411) );
  AOI222_X1 U7364 ( .A1(n6413), .A2(n6412), .B1(n6413), .B2(n6411), .C1(n6412), 
        .C2(n6411), .ZN(n6416) );
  OAI21_X1 U7365 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6414), 
        .ZN(n6415) );
  OAI21_X1 U7366 ( .B1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n6416), .A(n6415), 
        .ZN(n6422) );
  NOR2_X1 U7367 ( .A1(n6418), .A2(n6417), .ZN(n6419) );
  NAND2_X1 U7368 ( .A1(n6420), .A2(n6419), .ZN(n6421) );
  NOR2_X1 U7369 ( .A1(n6422), .A2(n6421), .ZN(n6435) );
  OAI21_X1 U7370 ( .B1(n6424), .B2(n6423), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n6425) );
  AOI221_X1 U7371 ( .B1(n6426), .B2(n6525), .C1(n4388), .C2(n6525), .A(n6425), 
        .ZN(n6429) );
  OAI221_X1 U7372 ( .B1(n6525), .B2(n6435), .C1(n6525), .C2(n6426), .A(n6429), 
        .ZN(n6507) );
  OAI21_X1 U7373 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4388), .A(n6507), .ZN(
        n6439) );
  AOI221_X1 U7374 ( .B1(n6428), .B2(STATE2_REG_0__SCAN_IN), .C1(n6439), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6427), .ZN(n6433) );
  INV_X1 U7375 ( .A(n6429), .ZN(n6430) );
  OAI211_X1 U7376 ( .C1(n6521), .C2(n6431), .A(n6525), .B(n6430), .ZN(n6432)
         );
  OAI211_X1 U7377 ( .C1(n6435), .C2(n6434), .A(n6433), .B(n6432), .ZN(U3148)
         );
  INV_X1 U7378 ( .A(n6507), .ZN(n6442) );
  AOI21_X1 U7379 ( .B1(n6437), .B2(n4388), .A(n6436), .ZN(n6441) );
  OAI221_X1 U7380 ( .B1(n6446), .B2(n6439), .C1(n6438), .C2(n6523), .A(
        STATE2_REG_1__SCAN_IN), .ZN(n6440) );
  OAI21_X1 U7381 ( .B1(n6442), .B2(n6441), .A(n6440), .ZN(U3149) );
  INV_X1 U7382 ( .A(n6443), .ZN(n6506) );
  OAI211_X1 U7383 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n4388), .A(n6506), .B(
        n6521), .ZN(n6445) );
  OAI21_X1 U7384 ( .B1(n6446), .B2(n6445), .A(n6444), .ZN(U3150) );
  INV_X1 U7385 ( .A(DATAWIDTH_REG_31__SCAN_IN), .ZN(n6680) );
  NOR2_X1 U7386 ( .A1(n6505), .A2(n6680), .ZN(U3151) );
  AND2_X1 U7387 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6447), .ZN(U3152) );
  AND2_X1 U7388 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6447), .ZN(U3153) );
  AND2_X1 U7389 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6447), .ZN(U3154) );
  AND2_X1 U7390 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6447), .ZN(U3155) );
  AND2_X1 U7391 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6447), .ZN(U3156) );
  INV_X1 U7392 ( .A(DATAWIDTH_REG_25__SCAN_IN), .ZN(n6696) );
  NOR2_X1 U7393 ( .A1(n6505), .A2(n6696), .ZN(U3157) );
  AND2_X1 U7394 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6447), .ZN(U3158) );
  AND2_X1 U7395 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6447), .ZN(U3159) );
  INV_X1 U7396 ( .A(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6586) );
  NOR2_X1 U7397 ( .A1(n6505), .A2(n6586), .ZN(U3160) );
  INV_X1 U7398 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n6689) );
  NOR2_X1 U7399 ( .A1(n6505), .A2(n6689), .ZN(U3161) );
  AND2_X1 U7400 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6447), .ZN(U3162) );
  INV_X1 U7401 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n6710) );
  NOR2_X1 U7402 ( .A1(n6505), .A2(n6710), .ZN(U3163) );
  AND2_X1 U7403 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6447), .ZN(U3164) );
  INV_X1 U7404 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n6783) );
  NOR2_X1 U7405 ( .A1(n6505), .A2(n6783), .ZN(U3165) );
  AND2_X1 U7406 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6447), .ZN(U3166) );
  AND2_X1 U7407 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6447), .ZN(U3167) );
  AND2_X1 U7408 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6447), .ZN(U3168) );
  AND2_X1 U7409 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6447), .ZN(U3169) );
  AND2_X1 U7410 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6447), .ZN(U3170) );
  AND2_X1 U7411 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6447), .ZN(U3171) );
  AND2_X1 U7412 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6447), .ZN(U3172) );
  AND2_X1 U7413 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6447), .ZN(U3173) );
  AND2_X1 U7414 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6447), .ZN(U3174) );
  AND2_X1 U7415 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6447), .ZN(U3175) );
  AND2_X1 U7416 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6447), .ZN(U3176) );
  INV_X1 U7417 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6736) );
  NOR2_X1 U7418 ( .A1(n6505), .A2(n6736), .ZN(U3177) );
  AND2_X1 U7419 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6447), .ZN(U3178) );
  AND2_X1 U7420 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6447), .ZN(U3179) );
  AND2_X1 U7421 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6447), .ZN(U3180) );
  NAND2_X1 U7422 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n6458) );
  INV_X1 U7423 ( .A(HOLD), .ZN(n6673) );
  OAI221_X1 U7424 ( .B1(n6673), .B2(n6448), .C1(n6673), .C2(n6451), .A(
        REQUESTPENDING_REG_SCAN_IN), .ZN(n6449) );
  INV_X1 U7425 ( .A(NA_N), .ZN(n6456) );
  AOI221_X1 U7426 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6456), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6460) );
  AOI21_X1 U7427 ( .B1(n6495), .B2(n6449), .A(n6460), .ZN(n6450) );
  OAI21_X1 U7428 ( .B1(STATE_REG_2__SCAN_IN), .B2(n6458), .A(n6450), .ZN(U3181) );
  NOR2_X1 U7429 ( .A1(n6451), .A2(n6673), .ZN(n6454) );
  INV_X1 U7430 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6645) );
  NOR2_X1 U7431 ( .A1(n4236), .A2(n6645), .ZN(n6457) );
  AOI21_X1 U7432 ( .B1(HOLD), .B2(STATE_REG_1__SCAN_IN), .A(n6457), .ZN(n6453)
         );
  OAI211_X1 U7433 ( .C1(n6454), .C2(n6453), .A(n6452), .B(n6458), .ZN(U3182)
         );
  AOI221_X1 U7434 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n4388), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6455) );
  AOI221_X1 U7435 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6455), .C2(HOLD), .A(n4236), .ZN(n6461) );
  AOI21_X1 U7436 ( .B1(n6457), .B2(n6456), .A(STATE_REG_2__SCAN_IN), .ZN(n6459) );
  OAI22_X1 U7437 ( .A1(n6461), .A2(n6460), .B1(n6459), .B2(n6458), .ZN(U3183)
         );
  NAND2_X1 U7438 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6532), .ZN(n6499) );
  NOR2_X2 U7439 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6495), .ZN(n6496) );
  AOI22_X1 U7440 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6496), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6495), .ZN(n6462) );
  OAI21_X1 U7441 ( .B1(n6516), .B2(n6499), .A(n6462), .ZN(U3184) );
  INV_X1 U7442 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n6574) );
  OAI222_X1 U7443 ( .A1(n6499), .A2(n5010), .B1(n6574), .B2(n6532), .C1(n6464), 
        .C2(n6501), .ZN(U3185) );
  AOI22_X1 U7444 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6496), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6495), .ZN(n6463) );
  OAI21_X1 U7445 ( .B1(n6464), .B2(n6499), .A(n6463), .ZN(U3186) );
  AOI22_X1 U7446 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6496), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6495), .ZN(n6465) );
  OAI21_X1 U7447 ( .B1(n6765), .B2(n6499), .A(n6465), .ZN(U3187) );
  AOI22_X1 U7448 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6496), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6495), .ZN(n6466) );
  OAI21_X1 U7449 ( .B1(n6467), .B2(n6499), .A(n6466), .ZN(U3188) );
  INV_X1 U7450 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n6687) );
  OAI222_X1 U7451 ( .A1(n6499), .A2(n6468), .B1(n6687), .B2(n6532), .C1(n6674), 
        .C2(n6501), .ZN(U3189) );
  AOI22_X1 U7452 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6496), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6495), .ZN(n6469) );
  OAI21_X1 U7453 ( .B1(n6674), .B2(n6499), .A(n6469), .ZN(U3190) );
  INV_X1 U7454 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6471) );
  INV_X1 U7455 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n6590) );
  INV_X1 U7456 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6705) );
  OAI222_X1 U7457 ( .A1(n6501), .A2(n6471), .B1(n6590), .B2(n6532), .C1(n6705), 
        .C2(n6499), .ZN(U3191) );
  AOI22_X1 U7458 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6496), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6495), .ZN(n6470) );
  OAI21_X1 U7459 ( .B1(n6471), .B2(n6499), .A(n6470), .ZN(U3192) );
  INV_X1 U7460 ( .A(n6499), .ZN(n6492) );
  AOI22_X1 U7461 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6492), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6495), .ZN(n6472) );
  OAI21_X1 U7462 ( .B1(n6473), .B2(n6501), .A(n6472), .ZN(U3193) );
  INV_X1 U7463 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n6756) );
  INV_X1 U7464 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6745) );
  OAI222_X1 U7465 ( .A1(n6499), .A2(n6473), .B1(n6756), .B2(n6532), .C1(n6745), 
        .C2(n6501), .ZN(U3194) );
  AOI22_X1 U7466 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6496), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6495), .ZN(n6474) );
  OAI21_X1 U7467 ( .B1(n6745), .B2(n6499), .A(n6474), .ZN(U3195) );
  AOI22_X1 U7468 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6496), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6495), .ZN(n6475) );
  OAI21_X1 U7469 ( .B1(n6476), .B2(n6499), .A(n6475), .ZN(U3196) );
  AOI22_X1 U7470 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6492), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6495), .ZN(n6477) );
  OAI21_X1 U7471 ( .B1(n6726), .B2(n6501), .A(n6477), .ZN(U3197) );
  AOI22_X1 U7472 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6496), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6495), .ZN(n6478) );
  OAI21_X1 U7473 ( .B1(n6726), .B2(n6499), .A(n6478), .ZN(U3198) );
  AOI22_X1 U7474 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6492), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6495), .ZN(n6479) );
  OAI21_X1 U7475 ( .B1(n6480), .B2(n6501), .A(n6479), .ZN(U3199) );
  AOI22_X1 U7476 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6492), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6495), .ZN(n6481) );
  OAI21_X1 U7477 ( .B1(n6483), .B2(n6501), .A(n6481), .ZN(U3200) );
  AOI22_X1 U7478 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6496), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6495), .ZN(n6482) );
  OAI21_X1 U7479 ( .B1(n6483), .B2(n6499), .A(n6482), .ZN(U3201) );
  INV_X1 U7480 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6484) );
  INV_X1 U7481 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n6606) );
  OAI222_X1 U7482 ( .A1(n6499), .A2(n6484), .B1(n6606), .B2(n6532), .C1(n6486), 
        .C2(n6501), .ZN(U3202) );
  AOI22_X1 U7483 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6496), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6495), .ZN(n6485) );
  OAI21_X1 U7484 ( .B1(n6486), .B2(n6499), .A(n6485), .ZN(U3203) );
  AOI22_X1 U7485 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6492), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6495), .ZN(n6487) );
  OAI21_X1 U7486 ( .B1(n6489), .B2(n6501), .A(n6487), .ZN(U3204) );
  AOI22_X1 U7487 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6496), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6495), .ZN(n6488) );
  OAI21_X1 U7488 ( .B1(n6489), .B2(n6499), .A(n6488), .ZN(U3205) );
  AOI22_X1 U7489 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6492), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6495), .ZN(n6490) );
  OAI21_X1 U7490 ( .B1(n6627), .B2(n6501), .A(n6490), .ZN(U3206) );
  INV_X1 U7491 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6695) );
  OAI222_X1 U7492 ( .A1(n6501), .A2(n6491), .B1(n6695), .B2(n6532), .C1(n6627), 
        .C2(n6499), .ZN(U3207) );
  INV_X1 U7493 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6692) );
  AOI22_X1 U7494 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6492), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6495), .ZN(n6493) );
  OAI21_X1 U7495 ( .B1(n6692), .B2(n6501), .A(n6493), .ZN(U3208) );
  INV_X1 U7496 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n6757) );
  OAI222_X1 U7497 ( .A1(n6499), .A2(n6692), .B1(n6757), .B2(n6532), .C1(n6655), 
        .C2(n6501), .ZN(U3209) );
  INV_X1 U7498 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6609) );
  OAI222_X1 U7499 ( .A1(n6499), .A2(n6655), .B1(n6609), .B2(n6532), .C1(n4210), 
        .C2(n6501), .ZN(U3210) );
  AOI22_X1 U7500 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6496), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6495), .ZN(n6494) );
  OAI21_X1 U7501 ( .B1(n4210), .B2(n6499), .A(n6494), .ZN(U3211) );
  AOI22_X1 U7502 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6496), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6495), .ZN(n6497) );
  OAI21_X1 U7503 ( .B1(n6498), .B2(n6499), .A(n6497), .ZN(U3212) );
  INV_X1 U7504 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n6657) );
  OAI222_X1 U7505 ( .A1(n6501), .A2(n5217), .B1(n6657), .B2(n6532), .C1(n6500), 
        .C2(n6499), .ZN(U3213) );
  MUX2_X1 U7506 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6532), .Z(U3445) );
  MUX2_X1 U7507 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6532), .Z(U3446) );
  MUX2_X1 U7508 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6532), .Z(U3447) );
  MUX2_X1 U7509 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6532), .Z(U3448) );
  OAI21_X1 U7510 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6505), .A(n6503), .ZN(
        n6502) );
  INV_X1 U7511 ( .A(n6502), .ZN(U3451) );
  INV_X1 U7512 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6504) );
  OAI21_X1 U7513 ( .B1(n6505), .B2(n6504), .A(n6503), .ZN(U3452) );
  OAI221_X1 U7514 ( .B1(n6817), .B2(STATE2_REG_0__SCAN_IN), .C1(n6817), .C2(
        n6507), .A(n6506), .ZN(U3453) );
  INV_X1 U7515 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6508) );
  OAI21_X1 U7516 ( .B1(REIP_REG_0__SCAN_IN), .B2(n6508), .A(n6516), .ZN(n6509)
         );
  OAI22_X1 U7517 ( .A1(n6510), .A2(n6509), .B1(REIP_REG_0__SCAN_IN), .B2(n6516), .ZN(n6512) );
  INV_X1 U7518 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6511) );
  AOI22_X1 U7519 ( .A1(n6513), .A2(n6512), .B1(n6511), .B2(n6515), .ZN(U3468)
         );
  INV_X1 U7520 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6514) );
  AOI22_X1 U7521 ( .A1(n6517), .A2(n6516), .B1(n6515), .B2(n6514), .ZN(U3469)
         );
  INV_X1 U7522 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6753) );
  MUX2_X1 U7523 ( .A(W_R_N_REG_SCAN_IN), .B(n6753), .S(n6532), .Z(U3470) );
  OAI211_X1 U7524 ( .C1(READY_N), .C2(n6520), .A(n6519), .B(n6518), .ZN(n6531)
         );
  INV_X1 U7525 ( .A(n6521), .ZN(n6529) );
  AOI21_X1 U7526 ( .B1(n6524), .B2(n6523), .A(n6522), .ZN(n6526) );
  AOI21_X1 U7527 ( .B1(n6527), .B2(n6526), .A(n6525), .ZN(n6528) );
  OAI21_X1 U7528 ( .B1(n6529), .B2(n6528), .A(n6531), .ZN(n6530) );
  OAI21_X1 U7529 ( .B1(n6531), .B2(n6645), .A(n6530), .ZN(U3472) );
  MUX2_X1 U7530 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6532), .Z(U3473) );
  OAI22_X1 U7531 ( .A1(n6536), .A2(n6535), .B1(n6534), .B2(n6533), .ZN(n6542)
         );
  OAI22_X1 U7532 ( .A1(n6540), .A2(n6539), .B1(n6538), .B2(n6537), .ZN(n6541)
         );
  AOI211_X1 U7533 ( .C1(INSTQUEUE_REG_10__5__SCAN_IN), .C2(n6543), .A(n6542), 
        .B(n6541), .ZN(n6802) );
  INV_X1 U7534 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n6546) );
  AOI22_X1 U7535 ( .A1(n6546), .A2(keyinput40), .B1(keyinput17), .B2(n6545), 
        .ZN(n6544) );
  OAI221_X1 U7536 ( .B1(n6546), .B2(keyinput40), .C1(n6545), .C2(keyinput17), 
        .A(n6544), .ZN(n6557) );
  AOI22_X1 U7537 ( .A1(n6548), .A2(keyinput8), .B1(n4376), .B2(keyinput0), 
        .ZN(n6547) );
  OAI221_X1 U7538 ( .B1(n6548), .B2(keyinput8), .C1(n4376), .C2(keyinput0), 
        .A(n6547), .ZN(n6556) );
  AOI22_X1 U7539 ( .A1(n6551), .A2(keyinput77), .B1(n6550), .B2(keyinput126), 
        .ZN(n6549) );
  OAI221_X1 U7540 ( .B1(n6551), .B2(keyinput77), .C1(n6550), .C2(keyinput126), 
        .A(n6549), .ZN(n6555) );
  NOR4_X1 U7541 ( .A1(n6557), .A2(n6556), .A3(n6555), .A4(n6554), .ZN(n6604)
         );
  AOI22_X1 U7542 ( .A1(n6559), .A2(keyinput84), .B1(n5347), .B2(keyinput50), 
        .ZN(n6558) );
  OAI221_X1 U7543 ( .B1(n6559), .B2(keyinput84), .C1(n5347), .C2(keyinput50), 
        .A(n6558), .ZN(n6570) );
  INV_X1 U7544 ( .A(EAX_REG_31__SCAN_IN), .ZN(n6561) );
  AOI22_X1 U7545 ( .A1(n5293), .A2(keyinput12), .B1(keyinput11), .B2(n6561), 
        .ZN(n6560) );
  OAI221_X1 U7546 ( .B1(n5293), .B2(keyinput12), .C1(n6561), .C2(keyinput11), 
        .A(n6560), .ZN(n6569) );
  AOI22_X1 U7547 ( .A1(n6564), .A2(keyinput62), .B1(n6563), .B2(keyinput89), 
        .ZN(n6562) );
  OAI221_X1 U7548 ( .B1(n6564), .B2(keyinput62), .C1(n6563), .C2(keyinput89), 
        .A(n6562), .ZN(n6568) );
  AOI22_X1 U7549 ( .A1(n6566), .A2(keyinput2), .B1(keyinput24), .B2(n6823), 
        .ZN(n6565) );
  OAI221_X1 U7550 ( .B1(n6566), .B2(keyinput2), .C1(n6823), .C2(keyinput24), 
        .A(n6565), .ZN(n6567) );
  NOR4_X1 U7551 ( .A1(n6570), .A2(n6569), .A3(n6568), .A4(n6567), .ZN(n6603)
         );
  INV_X1 U7552 ( .A(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n6835) );
  AOI22_X1 U7553 ( .A1(n6572), .A2(keyinput37), .B1(n6835), .B2(keyinput97), 
        .ZN(n6571) );
  OAI221_X1 U7554 ( .B1(n6572), .B2(keyinput37), .C1(n6835), .C2(keyinput97), 
        .A(n6571), .ZN(n6584) );
  AOI22_X1 U7555 ( .A1(n6575), .A2(keyinput53), .B1(n6574), .B2(keyinput19), 
        .ZN(n6573) );
  OAI221_X1 U7556 ( .B1(n6575), .B2(keyinput53), .C1(n6574), .C2(keyinput19), 
        .A(n6573), .ZN(n6583) );
  INV_X1 U7557 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n6577) );
  AOI22_X1 U7558 ( .A1(n3776), .A2(keyinput127), .B1(n6577), .B2(keyinput119), 
        .ZN(n6576) );
  OAI221_X1 U7559 ( .B1(n3776), .B2(keyinput127), .C1(n6577), .C2(keyinput119), 
        .A(n6576), .ZN(n6582) );
  AOI22_X1 U7560 ( .A1(n6580), .A2(keyinput59), .B1(keyinput85), .B2(n6579), 
        .ZN(n6578) );
  OAI221_X1 U7561 ( .B1(n6580), .B2(keyinput59), .C1(n6579), .C2(keyinput85), 
        .A(n6578), .ZN(n6581) );
  NOR4_X1 U7562 ( .A1(n6584), .A2(n6583), .A3(n6582), .A4(n6581), .ZN(n6602)
         );
  INV_X1 U7563 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6587) );
  AOI22_X1 U7564 ( .A1(n6587), .A2(keyinput125), .B1(keyinput78), .B2(n6586), 
        .ZN(n6585) );
  OAI221_X1 U7565 ( .B1(n6587), .B2(keyinput125), .C1(n6586), .C2(keyinput78), 
        .A(n6585), .ZN(n6600) );
  AOI22_X1 U7566 ( .A1(n6590), .A2(keyinput63), .B1(keyinput88), .B2(n6589), 
        .ZN(n6588) );
  OAI221_X1 U7567 ( .B1(n6590), .B2(keyinput63), .C1(n6589), .C2(keyinput88), 
        .A(n6588), .ZN(n6599) );
  INV_X1 U7568 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n6593) );
  AOI22_X1 U7569 ( .A1(n6593), .A2(keyinput33), .B1(keyinput14), .B2(n6592), 
        .ZN(n6591) );
  OAI221_X1 U7570 ( .B1(n6593), .B2(keyinput33), .C1(n6592), .C2(keyinput14), 
        .A(n6591), .ZN(n6598) );
  INV_X1 U7571 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6596) );
  AOI22_X1 U7572 ( .A1(n6596), .A2(keyinput118), .B1(n6595), .B2(keyinput48), 
        .ZN(n6594) );
  OAI221_X1 U7573 ( .B1(n6596), .B2(keyinput118), .C1(n6595), .C2(keyinput48), 
        .A(n6594), .ZN(n6597) );
  NOR4_X1 U7574 ( .A1(n6600), .A2(n6599), .A3(n6598), .A4(n6597), .ZN(n6601)
         );
  NAND4_X1 U7575 ( .A1(n6604), .A2(n6603), .A3(n6602), .A4(n6601), .ZN(n6800)
         );
  AOI22_X1 U7576 ( .A1(n6607), .A2(keyinput111), .B1(keyinput101), .B2(n6606), 
        .ZN(n6605) );
  OAI221_X1 U7577 ( .B1(n6607), .B2(keyinput111), .C1(n6606), .C2(keyinput101), 
        .A(n6605), .ZN(n6619) );
  AOI22_X1 U7578 ( .A1(n6609), .A2(keyinput106), .B1(n6820), .B2(keyinput10), 
        .ZN(n6608) );
  OAI221_X1 U7579 ( .B1(n6609), .B2(keyinput106), .C1(n6820), .C2(keyinput10), 
        .A(n6608), .ZN(n6618) );
  INV_X1 U7580 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n6612) );
  AOI22_X1 U7581 ( .A1(n6612), .A2(keyinput79), .B1(keyinput61), .B2(n6611), 
        .ZN(n6610) );
  OAI221_X1 U7582 ( .B1(n6612), .B2(keyinput79), .C1(n6611), .C2(keyinput61), 
        .A(n6610), .ZN(n6617) );
  INV_X1 U7583 ( .A(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n6615) );
  AOI22_X1 U7584 ( .A1(n6615), .A2(keyinput75), .B1(keyinput30), .B2(n6614), 
        .ZN(n6613) );
  OAI221_X1 U7585 ( .B1(n6615), .B2(keyinput75), .C1(n6614), .C2(keyinput30), 
        .A(n6613), .ZN(n6616) );
  NOR4_X1 U7586 ( .A1(n6619), .A2(n6618), .A3(n6617), .A4(n6616), .ZN(n6669)
         );
  AOI22_X1 U7587 ( .A1(n6622), .A2(keyinput38), .B1(n6621), .B2(keyinput56), 
        .ZN(n6620) );
  OAI221_X1 U7588 ( .B1(n6622), .B2(keyinput38), .C1(n6621), .C2(keyinput56), 
        .A(n6620), .ZN(n6635) );
  AOI22_X1 U7589 ( .A1(n6625), .A2(keyinput65), .B1(keyinput104), .B2(n6624), 
        .ZN(n6623) );
  OAI221_X1 U7590 ( .B1(n6625), .B2(keyinput65), .C1(n6624), .C2(keyinput104), 
        .A(n6623), .ZN(n6634) );
  AOI22_X1 U7591 ( .A1(n6628), .A2(keyinput39), .B1(n6627), .B2(keyinput3), 
        .ZN(n6626) );
  OAI221_X1 U7592 ( .B1(n6628), .B2(keyinput39), .C1(n6627), .C2(keyinput3), 
        .A(n6626), .ZN(n6633) );
  INV_X1 U7593 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n6631) );
  AOI22_X1 U7594 ( .A1(n6631), .A2(keyinput55), .B1(keyinput21), .B2(n6630), 
        .ZN(n6629) );
  OAI221_X1 U7595 ( .B1(n6631), .B2(keyinput55), .C1(n6630), .C2(keyinput21), 
        .A(n6629), .ZN(n6632) );
  NOR4_X1 U7596 ( .A1(n6635), .A2(n6634), .A3(n6633), .A4(n6632), .ZN(n6668)
         );
  INV_X1 U7597 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n6840) );
  INV_X1 U7598 ( .A(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n6637) );
  AOI22_X1 U7599 ( .A1(n6840), .A2(keyinput121), .B1(n6637), .B2(keyinput9), 
        .ZN(n6636) );
  OAI221_X1 U7600 ( .B1(n6840), .B2(keyinput121), .C1(n6637), .C2(keyinput9), 
        .A(n6636), .ZN(n6649) );
  INV_X1 U7601 ( .A(UWORD_REG_6__SCAN_IN), .ZN(n6639) );
  AOI22_X1 U7602 ( .A1(n6640), .A2(keyinput95), .B1(n6639), .B2(keyinput36), 
        .ZN(n6638) );
  OAI221_X1 U7603 ( .B1(n6640), .B2(keyinput95), .C1(n6639), .C2(keyinput36), 
        .A(n6638), .ZN(n6648) );
  INV_X1 U7604 ( .A(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n6641) );
  XOR2_X1 U7605 ( .A(n6641), .B(keyinput45), .Z(n6644) );
  XNOR2_X1 U7606 ( .A(INSTQUEUE_REG_9__6__SCAN_IN), .B(keyinput99), .ZN(n6643)
         );
  XNOR2_X1 U7607 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput26), .ZN(
        n6642) );
  NAND3_X1 U7608 ( .A1(n6644), .A2(n6643), .A3(n6642), .ZN(n6647) );
  XNOR2_X1 U7609 ( .A(n6645), .B(keyinput69), .ZN(n6646) );
  NOR4_X1 U7610 ( .A1(n6649), .A2(n6648), .A3(n6647), .A4(n6646), .ZN(n6667)
         );
  INV_X1 U7611 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n6652) );
  AOI22_X1 U7612 ( .A1(n6652), .A2(keyinput41), .B1(keyinput122), .B2(n6651), 
        .ZN(n6650) );
  OAI221_X1 U7613 ( .B1(n6652), .B2(keyinput41), .C1(n6651), .C2(keyinput122), 
        .A(n6650), .ZN(n6665) );
  AOI22_X1 U7614 ( .A1(n6655), .A2(keyinput71), .B1(n6654), .B2(keyinput94), 
        .ZN(n6653) );
  OAI221_X1 U7615 ( .B1(n6655), .B2(keyinput71), .C1(n6654), .C2(keyinput94), 
        .A(n6653), .ZN(n6664) );
  AOI22_X1 U7616 ( .A1(n6658), .A2(keyinput74), .B1(keyinput98), .B2(n6657), 
        .ZN(n6656) );
  OAI221_X1 U7617 ( .B1(n6658), .B2(keyinput74), .C1(n6657), .C2(keyinput98), 
        .A(n6656), .ZN(n6663) );
  INV_X1 U7618 ( .A(DATAI_26_), .ZN(n6661) );
  AOI22_X1 U7619 ( .A1(n6661), .A2(keyinput47), .B1(n6660), .B2(keyinput4), 
        .ZN(n6659) );
  OAI221_X1 U7620 ( .B1(n6661), .B2(keyinput47), .C1(n6660), .C2(keyinput4), 
        .A(n6659), .ZN(n6662) );
  NOR4_X1 U7621 ( .A1(n6665), .A2(n6664), .A3(n6663), .A4(n6662), .ZN(n6666)
         );
  NAND4_X1 U7622 ( .A1(n6669), .A2(n6668), .A3(n6667), .A4(n6666), .ZN(n6799)
         );
  INV_X1 U7623 ( .A(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n6671) );
  AOI22_X1 U7624 ( .A1(n3741), .A2(keyinput20), .B1(n6671), .B2(keyinput49), 
        .ZN(n6670) );
  OAI221_X1 U7625 ( .B1(n3741), .B2(keyinput20), .C1(n6671), .C2(keyinput49), 
        .A(n6670), .ZN(n6684) );
  AOI22_X1 U7626 ( .A1(n6674), .A2(keyinput102), .B1(keyinput96), .B2(n6673), 
        .ZN(n6672) );
  OAI221_X1 U7627 ( .B1(n6674), .B2(keyinput102), .C1(n6673), .C2(keyinput96), 
        .A(n6672), .ZN(n6683) );
  INV_X1 U7628 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n6676) );
  AOI22_X1 U7629 ( .A1(n6677), .A2(keyinput1), .B1(n6676), .B2(keyinput72), 
        .ZN(n6675) );
  OAI221_X1 U7630 ( .B1(n6677), .B2(keyinput1), .C1(n6676), .C2(keyinput72), 
        .A(n6675), .ZN(n6682) );
  INV_X1 U7631 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6679) );
  AOI22_X1 U7632 ( .A1(n6680), .A2(keyinput73), .B1(n6679), .B2(keyinput34), 
        .ZN(n6678) );
  OAI221_X1 U7633 ( .B1(n6680), .B2(keyinput73), .C1(n6679), .C2(keyinput34), 
        .A(n6678), .ZN(n6681) );
  NOR4_X1 U7634 ( .A1(n6684), .A2(n6683), .A3(n6682), .A4(n6681), .ZN(n6734)
         );
  AOI22_X1 U7635 ( .A1(n6687), .A2(keyinput64), .B1(n6686), .B2(keyinput70), 
        .ZN(n6685) );
  OAI221_X1 U7636 ( .B1(n6687), .B2(keyinput64), .C1(n6686), .C2(keyinput70), 
        .A(n6685), .ZN(n6700) );
  AOI22_X1 U7637 ( .A1(n6690), .A2(keyinput31), .B1(keyinput114), .B2(n6689), 
        .ZN(n6688) );
  OAI221_X1 U7638 ( .B1(n6690), .B2(keyinput31), .C1(n6689), .C2(keyinput114), 
        .A(n6688), .ZN(n6699) );
  INV_X1 U7639 ( .A(DATAI_22_), .ZN(n6693) );
  AOI22_X1 U7640 ( .A1(n6693), .A2(keyinput113), .B1(n6692), .B2(keyinput120), 
        .ZN(n6691) );
  OAI221_X1 U7641 ( .B1(n6693), .B2(keyinput113), .C1(n6692), .C2(keyinput120), 
        .A(n6691), .ZN(n6698) );
  AOI22_X1 U7642 ( .A1(n6696), .A2(keyinput100), .B1(keyinput107), .B2(n6695), 
        .ZN(n6694) );
  OAI221_X1 U7643 ( .B1(n6696), .B2(keyinput100), .C1(n6695), .C2(keyinput107), 
        .A(n6694), .ZN(n6697) );
  NOR4_X1 U7644 ( .A1(n6700), .A2(n6699), .A3(n6698), .A4(n6697), .ZN(n6733)
         );
  AOI22_X1 U7645 ( .A1(n6822), .A2(keyinput32), .B1(n6702), .B2(keyinput27), 
        .ZN(n6701) );
  OAI221_X1 U7646 ( .B1(n6822), .B2(keyinput32), .C1(n6702), .C2(keyinput27), 
        .A(n6701), .ZN(n6715) );
  AOI22_X1 U7647 ( .A1(n6705), .A2(keyinput42), .B1(n6704), .B2(keyinput91), 
        .ZN(n6703) );
  OAI221_X1 U7648 ( .B1(n6705), .B2(keyinput42), .C1(n6704), .C2(keyinput91), 
        .A(n6703), .ZN(n6714) );
  AOI22_X1 U7649 ( .A1(n6708), .A2(keyinput123), .B1(n6707), .B2(keyinput52), 
        .ZN(n6706) );
  OAI221_X1 U7650 ( .B1(n6708), .B2(keyinput123), .C1(n6707), .C2(keyinput52), 
        .A(n6706), .ZN(n6713) );
  AOI22_X1 U7651 ( .A1(n6711), .A2(keyinput80), .B1(keyinput29), .B2(n6710), 
        .ZN(n6709) );
  OAI221_X1 U7652 ( .B1(n6711), .B2(keyinput80), .C1(n6710), .C2(keyinput29), 
        .A(n6709), .ZN(n6712) );
  NOR4_X1 U7653 ( .A1(n6715), .A2(n6714), .A3(n6713), .A4(n6712), .ZN(n6732)
         );
  AOI22_X1 U7654 ( .A1(n6717), .A2(keyinput58), .B1(n6817), .B2(keyinput66), 
        .ZN(n6716) );
  OAI221_X1 U7655 ( .B1(n6717), .B2(keyinput58), .C1(n6817), .C2(keyinput66), 
        .A(n6716), .ZN(n6730) );
  INV_X1 U7656 ( .A(BS16_N), .ZN(n6719) );
  AOI22_X1 U7657 ( .A1(n6720), .A2(keyinput82), .B1(keyinput22), .B2(n6719), 
        .ZN(n6718) );
  OAI221_X1 U7658 ( .B1(n6720), .B2(keyinput82), .C1(n6719), .C2(keyinput22), 
        .A(n6718), .ZN(n6729) );
  AOI22_X1 U7659 ( .A1(n6723), .A2(keyinput15), .B1(keyinput51), .B2(n6722), 
        .ZN(n6721) );
  OAI221_X1 U7660 ( .B1(n6723), .B2(keyinput15), .C1(n6722), .C2(keyinput51), 
        .A(n6721), .ZN(n6728) );
  INV_X1 U7661 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n6725) );
  AOI22_X1 U7662 ( .A1(n6726), .A2(keyinput60), .B1(n6725), .B2(keyinput35), 
        .ZN(n6724) );
  OAI221_X1 U7663 ( .B1(n6726), .B2(keyinput60), .C1(n6725), .C2(keyinput35), 
        .A(n6724), .ZN(n6727) );
  NOR4_X1 U7664 ( .A1(n6730), .A2(n6729), .A3(n6728), .A4(n6727), .ZN(n6731)
         );
  NAND4_X1 U7665 ( .A1(n6734), .A2(n6733), .A3(n6732), .A4(n6731), .ZN(n6798)
         );
  AOI22_X1 U7666 ( .A1(n6737), .A2(keyinput46), .B1(n6736), .B2(keyinput43), 
        .ZN(n6735) );
  OAI221_X1 U7667 ( .B1(n6737), .B2(keyinput46), .C1(n6736), .C2(keyinput43), 
        .A(n6735), .ZN(n6749) );
  INV_X1 U7668 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n6739) );
  AOI22_X1 U7669 ( .A1(n6740), .A2(keyinput23), .B1(n6739), .B2(keyinput68), 
        .ZN(n6738) );
  OAI221_X1 U7670 ( .B1(n6740), .B2(keyinput23), .C1(n6739), .C2(keyinput68), 
        .A(n6738), .ZN(n6748) );
  INV_X1 U7671 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6742) );
  AOI22_X1 U7672 ( .A1(n6743), .A2(keyinput7), .B1(keyinput25), .B2(n6742), 
        .ZN(n6741) );
  OAI221_X1 U7673 ( .B1(n6743), .B2(keyinput7), .C1(n6742), .C2(keyinput25), 
        .A(n6741), .ZN(n6747) );
  INV_X1 U7674 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n6828) );
  AOI22_X1 U7675 ( .A1(n6828), .A2(keyinput67), .B1(keyinput44), .B2(n6745), 
        .ZN(n6744) );
  OAI221_X1 U7676 ( .B1(n6828), .B2(keyinput67), .C1(n6745), .C2(keyinput44), 
        .A(n6744), .ZN(n6746) );
  NOR4_X1 U7677 ( .A1(n6749), .A2(n6748), .A3(n6747), .A4(n6746), .ZN(n6796)
         );
  AOI22_X1 U7678 ( .A1(n3952), .A2(keyinput57), .B1(keyinput108), .B2(n6751), 
        .ZN(n6750) );
  OAI221_X1 U7679 ( .B1(n3952), .B2(keyinput57), .C1(n6751), .C2(keyinput108), 
        .A(n6750), .ZN(n6763) );
  INV_X1 U7680 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n6754) );
  AOI22_X1 U7681 ( .A1(n6754), .A2(keyinput28), .B1(keyinput87), .B2(n6753), 
        .ZN(n6752) );
  OAI221_X1 U7682 ( .B1(n6754), .B2(keyinput28), .C1(n6753), .C2(keyinput87), 
        .A(n6752), .ZN(n6762) );
  AOI22_X1 U7683 ( .A1(n6757), .A2(keyinput92), .B1(n6756), .B2(keyinput105), 
        .ZN(n6755) );
  OAI221_X1 U7684 ( .B1(n6757), .B2(keyinput92), .C1(n6756), .C2(keyinput105), 
        .A(n6755), .ZN(n6761) );
  AOI22_X1 U7685 ( .A1(n6759), .A2(keyinput6), .B1(n6827), .B2(keyinput18), 
        .ZN(n6758) );
  OAI221_X1 U7686 ( .B1(n6759), .B2(keyinput6), .C1(n6827), .C2(keyinput18), 
        .A(n6758), .ZN(n6760) );
  NOR4_X1 U7687 ( .A1(n6763), .A2(n6762), .A3(n6761), .A4(n6760), .ZN(n6795)
         );
  AOI22_X1 U7688 ( .A1(n6765), .A2(keyinput83), .B1(n3719), .B2(keyinput90), 
        .ZN(n6764) );
  OAI221_X1 U7689 ( .B1(n6765), .B2(keyinput83), .C1(n3719), .C2(keyinput90), 
        .A(n6764), .ZN(n6777) );
  AOI22_X1 U7690 ( .A1(n6768), .A2(keyinput112), .B1(n6767), .B2(keyinput54), 
        .ZN(n6766) );
  OAI221_X1 U7691 ( .B1(n6768), .B2(keyinput112), .C1(n6767), .C2(keyinput54), 
        .A(n6766), .ZN(n6776) );
  AOI22_X1 U7692 ( .A1(n5554), .A2(keyinput86), .B1(keyinput76), .B2(n6770), 
        .ZN(n6769) );
  OAI221_X1 U7693 ( .B1(n5554), .B2(keyinput86), .C1(n6770), .C2(keyinput76), 
        .A(n6769), .ZN(n6775) );
  INV_X1 U7694 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n6773) );
  AOI22_X1 U7695 ( .A1(n6773), .A2(keyinput117), .B1(keyinput5), .B2(n6772), 
        .ZN(n6771) );
  OAI221_X1 U7696 ( .B1(n6773), .B2(keyinput117), .C1(n6772), .C2(keyinput5), 
        .A(n6771), .ZN(n6774) );
  NOR4_X1 U7697 ( .A1(n6777), .A2(n6776), .A3(n6775), .A4(n6774), .ZN(n6794)
         );
  AOI22_X1 U7698 ( .A1(n6780), .A2(keyinput13), .B1(keyinput103), .B2(n6779), 
        .ZN(n6778) );
  OAI221_X1 U7699 ( .B1(n6780), .B2(keyinput13), .C1(n6779), .C2(keyinput103), 
        .A(n6778), .ZN(n6792) );
  INV_X1 U7700 ( .A(DATAI_16_), .ZN(n6782) );
  AOI22_X1 U7701 ( .A1(n6783), .A2(keyinput93), .B1(n6782), .B2(keyinput115), 
        .ZN(n6781) );
  OAI221_X1 U7702 ( .B1(n6783), .B2(keyinput93), .C1(n6782), .C2(keyinput115), 
        .A(n6781), .ZN(n6791) );
  AOI22_X1 U7703 ( .A1(n6786), .A2(keyinput110), .B1(n6785), .B2(keyinput109), 
        .ZN(n6784) );
  OAI221_X1 U7704 ( .B1(n6786), .B2(keyinput110), .C1(n6785), .C2(keyinput109), 
        .A(n6784), .ZN(n6790) );
  INV_X1 U7705 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6788) );
  AOI22_X1 U7706 ( .A1(n6826), .A2(keyinput81), .B1(keyinput116), .B2(n6788), 
        .ZN(n6787) );
  OAI221_X1 U7707 ( .B1(n6826), .B2(keyinput81), .C1(n6788), .C2(keyinput116), 
        .A(n6787), .ZN(n6789) );
  NOR4_X1 U7708 ( .A1(n6792), .A2(n6791), .A3(n6790), .A4(n6789), .ZN(n6793)
         );
  NAND4_X1 U7709 ( .A1(n6796), .A2(n6795), .A3(n6794), .A4(n6793), .ZN(n6797)
         );
  NOR4_X1 U7710 ( .A1(n6800), .A2(n6799), .A3(n6798), .A4(n6797), .ZN(n6801)
         );
  XNOR2_X1 U7711 ( .A(n6802), .B(n6801), .ZN(n6858) );
  NOR4_X1 U7712 ( .A1(EBX_REG_14__SCAN_IN), .A2(EAX_REG_14__SCAN_IN), .A3(
        DATAI_1_), .A4(DATAO_REG_14__SCAN_IN), .ZN(n6856) );
  NOR4_X1 U7713 ( .A1(EAX_REG_2__SCAN_IN), .A2(LWORD_REG_11__SCAN_IN), .A3(
        DATAO_REG_4__SCAN_IN), .A4(DATAO_REG_5__SCAN_IN), .ZN(n6855) );
  NAND4_X1 U7714 ( .A1(UWORD_REG_7__SCAN_IN), .A2(UWORD_REG_13__SCAN_IN), .A3(
        D_C_N_REG_SCAN_IN), .A4(ADDRESS_REG_29__SCAN_IN), .ZN(n6809) );
  NAND4_X1 U7715 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(UWORD_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(DATAWIDTH_REG_19__SCAN_IN), .ZN(
        n6808) );
  NOR4_X1 U7716 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .A3(EAX_REG_20__SCAN_IN), .A4(
        CODEFETCH_REG_SCAN_IN), .ZN(n6806) );
  NOR4_X1 U7717 ( .A1(EBX_REG_21__SCAN_IN), .A2(EBX_REG_4__SCAN_IN), .A3(
        PHYADDRPOINTER_REG_17__SCAN_IN), .A4(REIP_REG_7__SCAN_IN), .ZN(n6805)
         );
  NOR4_X1 U7718 ( .A1(EAX_REG_30__SCAN_IN), .A2(REIP_REG_23__SCAN_IN), .A3(
        REIP_REG_27__SCAN_IN), .A4(DATAI_11_), .ZN(n6804) );
  NOR4_X1 U7719 ( .A1(EAX_REG_21__SCAN_IN), .A2(EAX_REG_22__SCAN_IN), .A3(
        DATAI_26_), .A4(DATAI_22_), .ZN(n6803) );
  NAND4_X1 U7720 ( .A1(n6806), .A2(n6805), .A3(n6804), .A4(n6803), .ZN(n6807)
         );
  NOR3_X1 U7721 ( .A1(n6809), .A2(n6808), .A3(n6807), .ZN(n6854) );
  NAND4_X1 U7722 ( .A1(EBX_REG_10__SCAN_IN), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .A3(EBX_REG_25__SCAN_IN), .A4(REIP_REG_4__SCAN_IN), .ZN(n6852) );
  NAND4_X1 U7723 ( .A1(EBX_REG_17__SCAN_IN), .A2(DATAI_0_), .A3(DATAI_16_), 
        .A4(UWORD_REG_6__SCAN_IN), .ZN(n6851) );
  NAND4_X1 U7724 ( .A1(EBX_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A3(REIP_REG_12__SCAN_IN), .A4(
        REIP_REG_8__SCAN_IN), .ZN(n6810) );
  NOR3_X1 U7725 ( .A1(ADDRESS_REG_25__SCAN_IN), .A2(n5347), .A3(n6810), .ZN(
        n6816) );
  NOR4_X1 U7726 ( .A1(DATAO_REG_25__SCAN_IN), .A2(ADDRESS_REG_5__SCAN_IN), 
        .A3(ADDRESS_REG_1__SCAN_IN), .A4(REIP_REG_0__SCAN_IN), .ZN(n6814) );
  NOR4_X1 U7727 ( .A1(ADDRESS_REG_23__SCAN_IN), .A2(DATAWIDTH_REG_31__SCAN_IN), 
        .A3(UWORD_REG_12__SCAN_IN), .A4(DATAO_REG_11__SCAN_IN), .ZN(n6813) );
  NOR4_X1 U7728 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A3(PHYADDRPOINTER_REG_11__SCAN_IN), 
        .A4(EAX_REG_8__SCAN_IN), .ZN(n6812) );
  NOR4_X1 U7729 ( .A1(FLUSH_REG_SCAN_IN), .A2(BS16_N), .A3(
        BYTEENABLE_REG_3__SCAN_IN), .A4(HOLD), .ZN(n6811) );
  AND4_X1 U7730 ( .A1(n6814), .A2(n6813), .A3(n6812), .A4(n6811), .ZN(n6815)
         );
  NAND4_X1 U7731 ( .A1(EBX_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .A3(n6816), .A4(n6815), .ZN(n6850)
         );
  NAND4_X1 U7732 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(
        INSTQUEUE_REG_5__7__SCAN_IN), .A3(INSTQUEUE_REG_2__7__SCAN_IN), .A4(
        n6817), .ZN(n6818) );
  NOR4_X1 U7733 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUE_REG_1__7__SCAN_IN), .A3(n6819), .A4(n6818), .ZN(n6848) );
  NOR4_X1 U7734 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(
        INSTQUEUE_REG_11__4__SCAN_IN), .A3(INSTQUEUE_REG_12__4__SCAN_IN), .A4(
        n6820), .ZN(n6821) );
  NAND3_X1 U7735 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(
        INSTQUEUE_REG_4__0__SCAN_IN), .A3(n6821), .ZN(n6834) );
  NAND2_X1 U7736 ( .A1(n6823), .A2(n6822), .ZN(n6825) );
  NOR4_X1 U7737 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_21__SCAN_IN), .A3(n6825), .A4(n6824), .ZN(n6831) );
  NOR4_X1 U7738 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(
        INSTQUEUE_REG_15__1__SCAN_IN), .A3(n6827), .A4(n6826), .ZN(n6830) );
  NOR4_X1 U7739 ( .A1(INSTQUEUE_REG_2__5__SCAN_IN), .A2(
        INSTQUEUE_REG_14__5__SCAN_IN), .A3(INSTQUEUE_REG_5__5__SCAN_IN), .A4(
        n6828), .ZN(n6829) );
  NAND4_X1 U7740 ( .A1(n6832), .A2(n6831), .A3(n6830), .A4(n6829), .ZN(n6833)
         );
  NOR4_X1 U7741 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n6835), .A3(n6834), 
        .A4(n6833), .ZN(n6847) );
  NAND4_X1 U7742 ( .A1(ADDRESS_REG_10__SCAN_IN), .A2(BYTEENABLE_REG_1__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(REQUESTPENDING_REG_SCAN_IN), .ZN(n6839)
         );
  NAND4_X1 U7743 ( .A1(REIP_REG_26__SCAN_IN), .A2(ADDRESS_REG_7__SCAN_IN), 
        .A3(ADDRESS_REG_26__SCAN_IN), .A4(READREQUEST_REG_SCAN_IN), .ZN(n6838)
         );
  NAND4_X1 U7744 ( .A1(EAX_REG_4__SCAN_IN), .A2(EAX_REG_15__SCAN_IN), .A3(
        LWORD_REG_6__SCAN_IN), .A4(DATAO_REG_13__SCAN_IN), .ZN(n6837) );
  NAND4_X1 U7745 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_0__SCAN_IN), .A3(ADDRESS_REG_18__SCAN_IN), .A4(
        LWORD_REG_2__SCAN_IN), .ZN(n6836) );
  NOR4_X1 U7746 ( .A1(n6839), .A2(n6838), .A3(n6837), .A4(n6836), .ZN(n6846)
         );
  NAND4_X1 U7747 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(
        INSTQUEUE_REG_15__6__SCAN_IN), .A3(INSTQUEUE_REG_12__2__SCAN_IN), .A4(
        INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6844) );
  NAND4_X1 U7748 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(
        INSTQUEUE_REG_8__2__SCAN_IN), .A3(INSTQUEUE_REG_6__2__SCAN_IN), .A4(
        n6840), .ZN(n6843) );
  NAND4_X1 U7749 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        EAX_REG_26__SCAN_IN), .A3(DATAI_30_), .A4(DATAI_13_), .ZN(n6842) );
  NAND4_X1 U7750 ( .A1(REIP_REG_24__SCAN_IN), .A2(INSTQUEUE_REG_0__3__SCAN_IN), 
        .A3(EAX_REG_31__SCAN_IN), .A4(DATAI_4_), .ZN(n6841) );
  NOR4_X1 U7751 ( .A1(n6844), .A2(n6843), .A3(n6842), .A4(n6841), .ZN(n6845)
         );
  NAND4_X1 U7752 ( .A1(n6848), .A2(n6847), .A3(n6846), .A4(n6845), .ZN(n6849)
         );
  NOR4_X1 U7753 ( .A1(n6852), .A2(n6851), .A3(n6850), .A4(n6849), .ZN(n6853)
         );
  NAND4_X1 U7754 ( .A1(n6856), .A2(n6855), .A3(n6854), .A4(n6853), .ZN(n6857)
         );
  XNOR2_X1 U7755 ( .A(n6858), .B(n6857), .ZN(U3105) );
  NAND2_X2 U3581 ( .A1(n3261), .A2(n3260), .ZN(n3293) );
  AND4_X1 U3582 ( .A1(n3255), .A2(n3254), .A3(n3253), .A4(n3252), .ZN(n3261)
         );
  CLKBUF_X1 U3563 ( .A(n3103), .Z(n3975) );
  CLKBUF_X1 U3588 ( .A(n3443), .Z(n3105) );
  INV_X1 U3591 ( .A(n3293), .ZN(n3706) );
  CLKBUF_X1 U3592 ( .A(n5243), .Z(n5244) );
  CLKBUF_X1 U3645 ( .A(n5233), .Z(n5234) );
  CLKBUF_X1 U3679 ( .A(n4578), .Z(n3113) );
  CLKBUF_X1 U3979 ( .A(n4480), .Z(n3110) );
endmodule

