

module b17_C_SARLock_k_64_3 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, U355, U356, U357, U358, 
        U359, U360, U361, U362, U363, U364, U366, U367, U368, U369, U370, U371, 
        U372, U373, U374, U375, U347, U348, U349, U350, U351, U352, U353, U354, 
        U365, U376, U247, U246, U245, U244, U243, U242, U241, U240, U239, U238, 
        U237, U236, U235, U234, U233, U232, U231, U230, U229, U228, U227, U226, 
        U225, U224, U223, U222, U221, U220, U219, U218, U217, U216, U251, U252, 
        U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, 
        U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, 
        U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274, 
        P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, 
        P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, 
        P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, 
        P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, 
        P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, 
        P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, 
        P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, 
        P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, 
        P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, 
        P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, 
        P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, 
        P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, 
        P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, 
        P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, 
        P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, 
        P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, 
        P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, 
        P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, 
        P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, 
        P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, 
        P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, 
        P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, 
        P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, 
        P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, 
        P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, 
        P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, 
        P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, 
        P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, 
        P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, 
        P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, 
        P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, 
        P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, 
        P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, 
        P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, 
        P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, 
        P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, 
        P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, 
        P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, 
        P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, 
        P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, 
        P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, 
        P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, 
        P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, 
        P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, 
        P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, 
        P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, 
        P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, 
        P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, 
        P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, 
        P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, 
        P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, 
        P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, 
        P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, 
        P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, 
        P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, 
        P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, 
        P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, 
        P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, 
        P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, 
        P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, 
        P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, 
        P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, 
        P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, 
        P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, 
        P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, 
        P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, 
        P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, 
        P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, 
        P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, 
        P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, 
        P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, 
        P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, 
        P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, 
        P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, 
        P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, 
        P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, 
        P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, 
        P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, 
        P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, 
        P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, 
        P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, 
        P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, 
        P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, 
        P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, 
        P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, 
        P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, 
        P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, 
        P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, 
        P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, 
        P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, 
        P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, 
        P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, 
        P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, 
        P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, 
        P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, 
        P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, 
        P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, 
        P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, 
        P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, 
        P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, 
        P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, 
        P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, 
        P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, 
        P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, 
        P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, 
        P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, 
        P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, 
        P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, 
        P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, 
        P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, 
        P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, 
        P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, 
        P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, 
        P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, 
        P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, 
        P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, 
        P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, 
        P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, 
        P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, 
        P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, 
        P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, 
        P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, 
        P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, 
        P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, 
        P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, 
        P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, 
        P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, 
        P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, 
        P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, 
        P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, 
        P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, 
        P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, 
        P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, 
        P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, 
        P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, 
        P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, 
        P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, 
        P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, 
        P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, 
        P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, 
        P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, 
        P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, 
        P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, 
        P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, 
        P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, 
        P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, 
        P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, 
        P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, 
        P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, 
        P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, 
        P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, 
        P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, 
        P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, 
        P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, 
        P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, 
        P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, 
        P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, 
        P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, 
        P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, 
        P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, 
        P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, 
        P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, 
        P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, 
        P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, 
        P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, 
        P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, 
        P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, 
        P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, 
        P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, 
        P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, 
        P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, 
        P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, 
        P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, 
        P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, 
        P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, 
        P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, 
        P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, 
        P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, 
        P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, 
        P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, 
        P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19810,
         n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818,
         n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
         n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834,
         n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
         n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
         n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
         n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906,
         n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914,
         n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
         n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
         n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938,
         n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
         n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954,
         n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962,
         n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970,
         n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978,
         n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986,
         n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
         n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
         n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
         n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018,
         n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
         n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034,
         n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
         n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
         n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
         n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
         n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
         n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
         n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
         n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
         n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
         n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
         n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
         n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162,
         n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
         n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178,
         n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
         n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
         n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202,
         n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
         n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
         n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226,
         n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250,
         n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
         n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
         n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274,
         n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282,
         n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
         n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298,
         n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306,
         n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314,
         n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322,
         n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
         n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338,
         n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
         n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
         n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
         n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370,
         n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378,
         n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
         n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
         n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
         n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
         n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
         n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
         n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
         n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442,
         n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450,
         n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
         n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
         n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
         n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482,
         n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490,
         n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
         n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
         n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514,
         n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
         n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
         n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
         n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
         n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554,
         n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562,
         n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
         n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
         n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
         n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610,
         n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
         n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626,
         n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634,
         n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
         n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
         n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
         n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
         n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
         n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
         n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
         n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
         n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
         n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754,
         n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
         n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770,
         n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778,
         n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
         n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
         n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
         n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
         n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
         n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
         n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842,
         n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
         n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
         n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
         n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874,
         n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
         n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
         n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
         n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
         n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946,
         n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
         n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
         n20963, n20964, n20965, n20966;

  INV_X2 U11006 ( .A(n19810), .ZN(n19744) );
  NOR2_X1 U11007 ( .A1(n17600), .A2(n17929), .ZN(n17599) );
  AND2_X1 U11008 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16932), .ZN(n16917) );
  NAND2_X1 U11010 ( .A1(n17005), .A2(P3_EBX_REG_10__SCAN_IN), .ZN(n16982) );
  OAI211_X1 U11011 ( .C1(n20060), .C2(n12311), .A(n12141), .B(n12140), .ZN(
        n13536) );
  INV_X1 U11012 ( .A(n18702), .ZN(n18046) );
  BUF_X2 U11013 ( .A(n12900), .Z(n12993) );
  CLKBUF_X1 U11014 ( .A(n10725), .Z(n17001) );
  CLKBUF_X1 U11015 ( .A(n16723), .Z(n9575) );
  NOR2_X1 U11016 ( .A1(n17687), .A2(n17694), .ZN(n17686) );
  XNOR2_X1 U11017 ( .A(n11984), .B(n11983), .ZN(n20194) );
  CLKBUF_X2 U11018 ( .A(n15414), .Z(n9579) );
  AND2_X1 U11019 ( .A1(n11631), .A2(n10156), .ZN(n10172) );
  AND2_X1 U11020 ( .A1(n11631), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10120) );
  AND2_X1 U11021 ( .A1(n11616), .A2(n10156), .ZN(n10279) );
  INV_X2 U11022 ( .A(n16723), .ZN(n16988) );
  AND2_X1 U11023 ( .A1(n11622), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10273) );
  INV_X2 U11025 ( .A(n10008), .ZN(n17013) );
  BUF_X4 U11026 ( .A(n10873), .Z(n9571) );
  AND4_X1 U11027 ( .A1(n18661), .A2(n10687), .A3(n18671), .A4(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10873) );
  INV_X4 U11028 ( .A(n10740), .ZN(n17009) );
  CLKBUF_X1 U11029 ( .A(n15414), .Z(n9578) );
  INV_X2 U11030 ( .A(n10725), .ZN(n16955) );
  OR2_X1 U11031 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10701), .ZN(
        n10725) );
  CLKBUF_X1 U11032 ( .A(n12484), .Z(n12048) );
  CLKBUF_X1 U11033 ( .A(n12066), .Z(n12543) );
  CLKBUF_X1 U11034 ( .A(n12641), .Z(n12570) );
  OR2_X2 U11035 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16645) );
  INV_X1 U11036 ( .A(n13325), .ZN(n11957) );
  BUF_X1 U11037 ( .A(n11960), .Z(n20094) );
  AND2_X1 U11038 ( .A1(n10017), .A2(n11879), .ZN(n11960) );
  AND2_X1 U11039 ( .A1(n13424), .A2(n13570), .ZN(n11939) );
  AND2_X2 U11040 ( .A1(n11851), .A2(n11858), .ZN(n11892) );
  AND2_X2 U11041 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13425) );
  CLKBUF_X2 U11042 ( .A(n10072), .Z(n11740) );
  CLKBUF_X3 U11043 ( .A(n11656), .Z(n9573) );
  AND2_X1 U11044 ( .A1(n10059), .A2(n16022), .ZN(n11656) );
  CLKBUF_X1 U11045 ( .A(n19902), .Z(n9561) );
  NOR2_X1 U11046 ( .A1(n13062), .A2(n13061), .ZN(n19902) );
  NOR2_X1 U11047 ( .A1(n17357), .A2(n10914), .ZN(n9562) );
  NOR2_X1 U11048 ( .A1(n17357), .A2(n10914), .ZN(n10915) );
  BUF_X1 U11049 ( .A(n12146), .Z(n12571) );
  NOR2_X1 U11050 ( .A1(n13104), .A2(n16044), .ZN(n10537) );
  AND2_X2 U11051 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13355) );
  INV_X1 U11052 ( .A(n13575), .ZN(n12615) );
  AND2_X1 U11053 ( .A1(n12673), .A2(n13126), .ZN(n13418) );
  BUF_X1 U11054 ( .A(n11921), .Z(n13437) );
  NAND2_X1 U11055 ( .A1(n12120), .A2(n12119), .ZN(n12714) );
  AND2_X1 U11056 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10092) );
  OR2_X1 U11057 ( .A1(n11071), .A2(n11070), .ZN(n11072) );
  NAND2_X1 U11058 ( .A1(n13144), .A2(n13381), .ZN(n13433) );
  CLKBUF_X3 U11059 ( .A(n11927), .Z(n12634) );
  BUF_X1 U11060 ( .A(n11918), .Z(n12671) );
  AND2_X1 U11061 ( .A1(n11787), .A2(n10156), .ZN(n10271) );
  AND2_X1 U11062 ( .A1(n11782), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10145) );
  INV_X1 U11063 ( .A(n10009), .ZN(n17012) );
  INV_X1 U11064 ( .A(n15418), .ZN(n10884) );
  INV_X1 U11065 ( .A(n10959), .ZN(n10964) );
  OR2_X1 U11066 ( .A1(n13433), .A2(n20072), .ZN(n13138) );
  OR2_X1 U11067 ( .A1(n13832), .A2(n13967), .ZN(n13969) );
  INV_X1 U11069 ( .A(n10439), .ZN(n10288) );
  INV_X2 U11071 ( .A(n10797), .ZN(n16734) );
  NAND2_X1 U11072 ( .A1(n12901), .A2(n12993), .ZN(n13315) );
  BUF_X1 U11074 ( .A(n10571), .Z(n10677) );
  CLKBUF_X2 U11075 ( .A(n10531), .Z(n14096) );
  NOR2_X1 U11076 ( .A1(n14984), .A2(n9948), .ZN(n14143) );
  INV_X1 U11077 ( .A(n17597), .ZN(n17557) );
  INV_X1 U11078 ( .A(n11010), .ZN(n18059) );
  NOR2_X1 U11079 ( .A1(n13878), .A2(n13877), .ZN(n13920) );
  OR2_X1 U11080 ( .A1(n14213), .A2(n14212), .ZN(n14214) );
  INV_X1 U11081 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11846) );
  INV_X1 U11082 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15369) );
  INV_X1 U11083 ( .A(n16654), .ZN(n16613) );
  INV_X2 U11084 ( .A(n17011), .ZN(n16903) );
  NAND2_X1 U11086 ( .A1(n18511), .A2(n14059), .ZN(n18506) );
  INV_X1 U11087 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19611) );
  INV_X1 U11088 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18683) );
  CLKBUF_X3 U11089 ( .A(n10677), .Z(n9595) );
  NAND4_X1 U11090 ( .A1(n18661), .A2(n9675), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A4(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16723) );
  OR3_X1 U11091 ( .A1(n10053), .A2(n14925), .A3(n9700), .ZN(n9563) );
  AND3_X4 U11092 ( .A1(n15368), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9564) );
  CLKBUF_X3 U11093 ( .A(n10072), .Z(n11782) );
  AND2_X1 U11094 ( .A1(n10493), .A2(n10012), .ZN(n9565) );
  AND2_X1 U11095 ( .A1(n10526), .A2(n10523), .ZN(n9566) );
  NAND2_X2 U11096 ( .A1(n15028), .A2(n15029), .ZN(n15027) );
  OAI21_X2 U11097 ( .B1(n12894), .B2(n11977), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11986) );
  NOR2_X2 U11098 ( .A1(n17666), .A2(n17665), .ZN(n17664) );
  AOI21_X2 U11099 ( .B1(n15052), .B2(n15014), .A(n15013), .ZN(n15028) );
  AOI22_X1 U11100 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14124), .B1(n14157), 
        .B2(n16078), .ZN(n13685) );
  NOR2_X2 U11101 ( .A1(n10195), .A2(n9923), .ZN(n9922) );
  NAND2_X1 U11102 ( .A1(n13517), .A2(n12773), .ZN(n12777) );
  NAND2_X2 U11103 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18509) );
  OAI21_X2 U11104 ( .B1(n15154), .B2(n15150), .A(n15151), .ZN(n14990) );
  NAND2_X2 U11105 ( .A1(n11481), .A2(n11480), .ZN(n11484) );
  AND2_X1 U11107 ( .A1(n10092), .A2(n15369), .ZN(n9568) );
  BUF_X8 U11109 ( .A(n11892), .Z(n12591) );
  NAND2_X4 U11111 ( .A1(n10233), .A2(n10232), .ZN(n19085) );
  NAND2_X1 U11112 ( .A1(n11215), .A2(n19070), .ZN(n14098) );
  INV_X2 U11113 ( .A(n19070), .ZN(n10531) );
  NAND2_X2 U11114 ( .A1(n13355), .A2(n16022), .ZN(n10102) );
  NOR2_X2 U11116 ( .A1(n14025), .A2(n14026), .ZN(n14352) );
  XNOR2_X1 U11117 ( .A(n12097), .B(n12096), .ZN(n13595) );
  XNOR2_X2 U11118 ( .A(n10923), .B(n10793), .ZN(n17640) );
  BUF_X4 U11119 ( .A(n10744), .Z(n17025) );
  INV_X1 U11120 ( .A(n10725), .ZN(n9570) );
  XNOR2_X2 U11121 ( .A(n10563), .B(n10564), .ZN(n11036) );
  BUF_X2 U11122 ( .A(n11656), .Z(n9572) );
  INV_X2 U11123 ( .A(n17538), .ZN(n17611) );
  INV_X1 U11124 ( .A(n10886), .ZN(n9576) );
  NAND2_X2 U11125 ( .A1(n10688), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10886) );
  NOR2_X1 U11126 ( .A1(n10724), .A2(n10699), .ZN(n15414) );
  NOR2_X1 U11127 ( .A1(n15088), .A2(n15977), .ZN(n14944) );
  INV_X2 U11129 ( .A(n15076), .ZN(n11223) );
  OAI21_X1 U11130 ( .B1(n16083), .B2(n17844), .A(n9738), .ZN(n9737) );
  AOI21_X1 U11131 ( .B1(n9791), .B2(n9799), .A(n9628), .ZN(n9790) );
  AOI21_X1 U11132 ( .B1(n17557), .B2(n17341), .A(n16139), .ZN(n17326) );
  NOR2_X1 U11133 ( .A1(n17341), .A2(n16131), .ZN(n15448) );
  INV_X4 U11134 ( .A(n15651), .ZN(n15631) );
  AND2_X1 U11135 ( .A1(n17377), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10912) );
  INV_X1 U11136 ( .A(n17688), .ZN(n17680) );
  NOR2_X1 U11138 ( .A1(n17601), .A2(n17671), .ZN(n17693) );
  BUF_X2 U11140 ( .A(n17689), .Z(n9596) );
  INV_X1 U11141 ( .A(n17420), .ZN(n9580) );
  OR2_X1 U11142 ( .A1(n11045), .A2(n15355), .ZN(n11051) );
  INV_X2 U11143 ( .A(n18486), .ZN(n17999) );
  CLKBUF_X2 U11144 ( .A(n11027), .Z(n11037) );
  NOR2_X1 U11146 ( .A1(n17627), .A2(n17626), .ZN(n17625) );
  INV_X2 U11147 ( .A(n17176), .ZN(n18077) );
  INV_X1 U11148 ( .A(n9588), .ZN(n19060) );
  INV_X2 U11149 ( .A(n19065), .ZN(n10520) );
  AND2_X2 U11150 ( .A1(n10260), .A2(n10259), .ZN(n9588) );
  AND4_X1 U11151 ( .A1(n11938), .A2(n11937), .A3(n11936), .A4(n11935), .ZN(
        n11955) );
  CLKBUF_X1 U11152 ( .A(n10273), .Z(n11595) );
  CLKBUF_X2 U11153 ( .A(n10884), .Z(n16965) );
  INV_X1 U11154 ( .A(n9564), .ZN(n9581) );
  INV_X1 U11155 ( .A(n9571), .ZN(n16958) );
  CLKBUF_X2 U11156 ( .A(n12296), .Z(n12401) );
  BUF_X2 U11157 ( .A(n11939), .Z(n12646) );
  NOR3_X1 U11158 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n18509), .ZN(n10744) );
  INV_X2 U11160 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16022) );
  AOI211_X1 U11161 ( .C1(n19042), .C2(n14946), .A(n14945), .B(n14944), .ZN(
        n14947) );
  AOI211_X1 U11162 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n15091), .A(
        n15090), .B(n15089), .ZN(n15092) );
  XNOR2_X1 U11163 ( .A(n12849), .B(n12848), .ZN(n14076) );
  AOI21_X1 U11164 ( .B1(n9831), .B2(n9830), .A(n9829), .ZN(n15240) );
  MUX2_X1 U11165 ( .A(n12847), .B(n12846), .S(n15651), .Z(n12849) );
  OAI21_X1 U11166 ( .B1(n9795), .B2(n9792), .A(n9790), .ZN(n14103) );
  NOR2_X1 U11167 ( .A1(n14934), .A2(n11325), .ZN(n11331) );
  NAND2_X1 U11168 ( .A1(n9932), .A2(n11490), .ZN(n15320) );
  NAND2_X1 U11169 ( .A1(n14501), .A2(n15631), .ZN(n9905) );
  NAND2_X1 U11170 ( .A1(n9813), .A2(n11485), .ZN(n15992) );
  OAI21_X1 U11171 ( .B1(n15065), .B2(n15066), .A(n15011), .ZN(n15052) );
  INV_X1 U11172 ( .A(n14479), .ZN(n14410) );
  NAND2_X1 U11173 ( .A1(n14980), .A2(n9808), .ZN(n9806) );
  CLKBUF_X1 U11174 ( .A(n14524), .Z(n14547) );
  OAI21_X1 U11175 ( .B1(n9766), .B2(n11223), .A(n9765), .ZN(n9764) );
  NAND2_X1 U11176 ( .A1(n14816), .A2(n11707), .ZN(n11729) );
  XNOR2_X1 U11177 ( .A(n11176), .B(n11453), .ZN(n13852) );
  NAND2_X1 U11178 ( .A1(n13652), .A2(n11466), .ZN(n13718) );
  NAND2_X1 U11179 ( .A1(n11153), .A2(n13709), .ZN(n11176) );
  NAND2_X1 U11180 ( .A1(n14166), .A2(n14165), .ZN(n14164) );
  NOR2_X1 U11181 ( .A1(n17342), .A2(n10917), .ZN(n15447) );
  INV_X1 U11182 ( .A(n17342), .ZN(n16139) );
  OR2_X1 U11183 ( .A1(n14889), .A2(n11653), .ZN(n9995) );
  XNOR2_X1 U11184 ( .A(n9931), .B(n9930), .ZN(n14360) );
  NAND2_X1 U11185 ( .A1(n9562), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17341) );
  AND2_X1 U11186 ( .A1(n14568), .A2(n12830), .ZN(n12831) );
  AND2_X1 U11187 ( .A1(n14042), .A2(n9631), .ZN(n14044) );
  AND2_X1 U11188 ( .A1(n10913), .A2(n17557), .ZN(n10914) );
  OR2_X1 U11189 ( .A1(n14867), .A2(n14866), .ZN(n15847) );
  NAND2_X1 U11190 ( .A1(n9809), .A2(n11312), .ZN(n9807) );
  AND2_X1 U11191 ( .A1(n12804), .A2(n12803), .ZN(n15667) );
  AND2_X1 U11192 ( .A1(n11208), .A2(n11207), .ZN(n11472) );
  OR2_X1 U11193 ( .A1(n11335), .A2(n10196), .ZN(n14097) );
  OR2_X1 U11194 ( .A1(n11204), .A2(n11203), .ZN(n11208) );
  OR2_X1 U11195 ( .A1(n11328), .A2(n11327), .ZN(n11335) );
  OR2_X1 U11196 ( .A1(n15845), .A2(n14100), .ZN(n11332) );
  INV_X2 U11197 ( .A(n17554), .ZN(n17506) );
  NAND2_X1 U11198 ( .A1(n17433), .A2(n10911), .ZN(n17404) );
  NAND2_X1 U11199 ( .A1(n12163), .A2(n9858), .ZN(n12798) );
  NAND2_X1 U11200 ( .A1(n11528), .A2(n11527), .ZN(n13276) );
  OR2_X2 U11201 ( .A1(n9670), .A2(n16430), .ZN(n16873) );
  OAI21_X1 U11202 ( .B1(n13600), .B2(n12311), .A(n12093), .ZN(n12094) );
  AND2_X1 U11203 ( .A1(n11506), .A2(n11530), .ZN(n13277) );
  OR2_X1 U11204 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n9619), .ZN(n11321) );
  OR2_X1 U11205 ( .A1(n13302), .A2(n13301), .ZN(n11528) );
  CLKBUF_X1 U11206 ( .A(n11117), .Z(n11118) );
  NAND2_X1 U11207 ( .A1(n11273), .A2(n11298), .ZN(n11304) );
  OR2_X1 U11208 ( .A1(n11086), .A2(n11664), .ZN(n11087) );
  NOR2_X2 U11209 ( .A1(n20110), .A2(n20099), .ZN(n20661) );
  NAND2_X1 U11210 ( .A1(n11299), .A2(n14098), .ZN(n11273) );
  OR2_X1 U11211 ( .A1(n11514), .A2(n11513), .ZN(n11515) );
  NAND2_X1 U11212 ( .A1(n11514), .A2(n11513), .ZN(n11527) );
  INV_X1 U11213 ( .A(n17696), .ZN(n17601) );
  NOR2_X1 U11214 ( .A1(n11070), .A2(n11040), .ZN(n9823) );
  OR2_X1 U11215 ( .A1(n9599), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11299) );
  AOI21_X1 U11216 ( .B1(n17501), .B2(n17597), .A(n9754), .ZN(n9751) );
  NAND2_X1 U11217 ( .A1(n11511), .A2(n11510), .ZN(n11514) );
  NAND2_X2 U11218 ( .A1(n14428), .A2(n13383), .ZN(n14434) );
  NOR2_X1 U11219 ( .A1(n13803), .A2(n13805), .ZN(n13804) );
  NOR2_X1 U11220 ( .A1(n11040), .A2(n11519), .ZN(n11041) );
  CLKBUF_X1 U11221 ( .A(n13076), .Z(n20512) );
  OR2_X1 U11222 ( .A1(n14019), .A2(n14018), .ZN(n14025) );
  NOR2_X1 U11223 ( .A1(n17931), .A2(n10905), .ZN(n17541) );
  NAND2_X1 U11224 ( .A1(n10581), .A2(n10580), .ZN(n11026) );
  INV_X1 U11225 ( .A(n16630), .ZN(n16646) );
  NAND2_X1 U11226 ( .A1(n13283), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13282) );
  NOR2_X1 U11227 ( .A1(n15332), .A2(n9644), .ZN(n13820) );
  XNOR2_X1 U11228 ( .A(n11039), .B(n11038), .ZN(n11519) );
  AOI211_X2 U11229 ( .C1(n18555), .C2(n18400), .A(n18718), .B(n16285), .ZN(
        n16649) );
  NAND2_X1 U11230 ( .A1(n9863), .A2(n9862), .ZN(n11267) );
  INV_X1 U11231 ( .A(n11265), .ZN(n9863) );
  NOR2_X2 U11232 ( .A1(n13174), .A2(n19054), .ZN(n13164) );
  NAND2_X1 U11233 ( .A1(n11982), .A2(n11981), .ZN(n11984) );
  XNOR2_X1 U11234 ( .A(n10590), .B(n10588), .ZN(n11025) );
  NAND2_X1 U11235 ( .A1(n11236), .A2(n11243), .ZN(n11265) );
  AND2_X2 U11236 ( .A1(n17233), .A2(n17266), .ZN(n17263) );
  AOI21_X1 U11237 ( .B1(n10677), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10587), .ZN(n10588) );
  OAI21_X1 U11238 ( .B1(n16265), .B2(n10976), .A(n10975), .ZN(n18500) );
  NAND2_X1 U11239 ( .A1(n11244), .A2(n14098), .ZN(n11236) );
  NAND2_X2 U11240 ( .A1(n17271), .A2(n13092), .ZN(n16265) );
  AND2_X1 U11241 ( .A1(n10576), .A2(n10575), .ZN(n11033) );
  INV_X2 U11242 ( .A(n13232), .ZN(n9582) );
  NOR2_X1 U11243 ( .A1(n17049), .A2(n20934), .ZN(n17056) );
  NOR2_X1 U11244 ( .A1(n10936), .A2(n10935), .ZN(n10938) );
  XOR2_X1 U11245 ( .A(n17953), .B(n10794), .Z(n17626) );
  NOR2_X1 U11246 ( .A1(n10770), .A2(n9761), .ZN(n9760) );
  XOR2_X1 U11247 ( .A(n17183), .B(n10796), .Z(n10794) );
  NOR2_X1 U11248 ( .A1(n9942), .A2(n13610), .ZN(n9939) );
  OR2_X1 U11249 ( .A1(n10544), .A2(n13104), .ZN(n10512) );
  NAND2_X1 U11250 ( .A1(n15509), .A2(n15432), .ZN(n17049) );
  NOR2_X1 U11251 ( .A1(n15429), .A2(n18702), .ZN(n10960) );
  NOR2_X1 U11252 ( .A1(n17674), .A2(n10738), .ZN(n10755) );
  NAND2_X1 U11253 ( .A1(n10793), .A2(n10923), .ZN(n10796) );
  AND2_X1 U11254 ( .A1(n10506), .A2(n10505), .ZN(n11440) );
  AND2_X1 U11255 ( .A1(n13196), .A2(n13197), .ZN(n13195) );
  AND2_X1 U11256 ( .A1(n13004), .A2(n20094), .ZN(n12885) );
  CLKBUF_X1 U11257 ( .A(n11352), .Z(n19805) );
  AND2_X1 U11258 ( .A1(n11405), .A2(n9810), .ZN(n10545) );
  OR2_X1 U11259 ( .A1(n10624), .A2(n19699), .ZN(n10561) );
  MUX2_X1 U11260 ( .A(n11339), .B(n13735), .S(n14096), .Z(n11167) );
  INV_X2 U11261 ( .A(n10624), .ZN(n14107) );
  NAND2_X1 U11262 ( .A1(n13418), .A2(n13382), .ZN(n12897) );
  NAND2_X1 U11263 ( .A1(n9865), .A2(n9864), .ZN(n11381) );
  NOR2_X1 U11264 ( .A1(n16266), .A2(n18077), .ZN(n10959) );
  NOR2_X1 U11265 ( .A1(n18066), .A2(n11001), .ZN(n11003) );
  OR2_X1 U11266 ( .A1(n11963), .A2(n11962), .ZN(n15460) );
  AND2_X1 U11267 ( .A1(n11974), .A2(n11973), .ZN(n13144) );
  AND2_X1 U11268 ( .A1(n10537), .A2(n11406), .ZN(n10525) );
  NAND2_X1 U11269 ( .A1(n13063), .A2(n12993), .ZN(n12986) );
  NOR2_X1 U11270 ( .A1(n17479), .A2(n17478), .ZN(n16279) );
  AND2_X1 U11271 ( .A1(n11959), .A2(n13381), .ZN(n11995) );
  INV_X1 U11272 ( .A(n10957), .ZN(n18066) );
  INV_X1 U11273 ( .A(n11264), .ZN(n9862) );
  AND2_X1 U11274 ( .A1(n16044), .A2(n19048), .ZN(n19801) );
  INV_X1 U11275 ( .A(n17203), .ZN(n10929) );
  OAI211_X1 U11276 ( .C1(n20895), .C2(n17001), .A(n10832), .B(n10831), .ZN(
        n16266) );
  OAI211_X1 U11277 ( .C1(n10009), .C2(n18074), .A(n10872), .B(n10871), .ZN(
        n17060) );
  OAI211_X1 U11278 ( .C1(n10009), .C2(n18063), .A(n10852), .B(n10851), .ZN(
        n11010) );
  OAI211_X1 U11279 ( .C1(n10009), .C2(n18069), .A(n10862), .B(n10861), .ZN(
        n10957) );
  OR2_X1 U11280 ( .A1(n9742), .A2(n10733), .ZN(n17695) );
  OR2_X1 U11281 ( .A1(n10099), .A2(n10098), .ZN(n11114) );
  OAI211_X1 U11282 ( .C1(n17001), .C2(n20844), .A(n10753), .B(n10752), .ZN(
        n17193) );
  OR2_X1 U11283 ( .A1(n10155), .A2(n10154), .ZN(n10316) );
  OR2_X1 U11284 ( .A1(n10137), .A2(n10136), .ZN(n10311) );
  INV_X1 U11285 ( .A(n10496), .ZN(n11824) );
  AND3_X1 U11286 ( .A1(n20085), .A2(n20104), .A3(n12759), .ZN(n11973) );
  NAND2_X4 U11287 ( .A1(n20090), .A2(n12697), .ZN(n12901) );
  INV_X2 U11288 ( .A(n16151), .ZN(n16201) );
  OR2_X1 U11289 ( .A1(n16045), .A2(n16078), .ZN(n13104) );
  CLKBUF_X3 U11290 ( .A(n10498), .Z(n19070) );
  INV_X1 U11291 ( .A(n16045), .ZN(n19048) );
  AOI211_X2 U11292 ( .C1(n16893), .C2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n10881), .B(n10880), .ZN(n10882) );
  AND2_X1 U11293 ( .A1(n10520), .A2(n9588), .ZN(n11406) );
  NAND2_X1 U11294 ( .A1(n10720), .A2(n10719), .ZN(n10721) );
  CLKBUF_X1 U11295 ( .A(n11503), .Z(n13192) );
  NOR2_X1 U11296 ( .A1(n10031), .A2(n18820), .ZN(n10030) );
  AOI211_X1 U11297 ( .C1(n9571), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n10830), .B(n10829), .ZN(n10831) );
  NAND2_X1 U11298 ( .A1(n10016), .A2(n9611), .ZN(n11918) );
  NAND2_X1 U11299 ( .A1(n11898), .A2(n10014), .ZN(n11921) );
  NAND2_X1 U11300 ( .A1(n10220), .A2(n10219), .ZN(n11503) );
  NAND2_X1 U11301 ( .A1(n10071), .A2(n9879), .ZN(n10514) );
  NAND2_X2 U11302 ( .A1(n9882), .A2(n9881), .ZN(n16045) );
  INV_X2 U11303 ( .A(U212), .ZN(n16198) );
  NAND2_X1 U11304 ( .A1(n10077), .A2(n10156), .ZN(n9882) );
  NAND2_X1 U11305 ( .A1(n10070), .A2(n9880), .ZN(n9879) );
  NOR2_X2 U11306 ( .A1(n20068), .A2(n20067), .ZN(n20069) );
  AND4_X1 U11307 ( .A1(n11943), .A2(n11942), .A3(n11941), .A4(n11940), .ZN(
        n11954) );
  AND4_X1 U11308 ( .A1(n11947), .A2(n11946), .A3(n11945), .A4(n11944), .ZN(
        n11953) );
  AND4_X1 U11309 ( .A1(n11891), .A2(n11890), .A3(n11889), .A4(n11888), .ZN(
        n11898) );
  AND4_X1 U11310 ( .A1(n11883), .A2(n11882), .A3(n11881), .A4(n11880), .ZN(
        n10016) );
  AND4_X1 U11311 ( .A1(n11845), .A2(n11844), .A3(n11843), .A4(n11842), .ZN(
        n11868) );
  INV_X2 U11312 ( .A(U214), .ZN(n16199) );
  AND4_X1 U11313 ( .A1(n11850), .A2(n11849), .A3(n11848), .A4(n11847), .ZN(
        n11867) );
  NAND2_X2 U11314 ( .A1(n19744), .A2(n19698), .ZN(n19749) );
  AND4_X1 U11315 ( .A1(n10201), .A2(n10200), .A3(n10199), .A4(n10198), .ZN(
        n10202) );
  AND4_X1 U11316 ( .A1(n10206), .A2(n10205), .A3(n10204), .A4(n10203), .ZN(
        n10207) );
  AND4_X1 U11317 ( .A1(n11864), .A2(n11863), .A3(n11862), .A4(n11861), .ZN(
        n11865) );
  AND4_X1 U11318 ( .A1(n11857), .A2(n11856), .A3(n11855), .A4(n11854), .ZN(
        n11866) );
  BUF_X2 U11319 ( .A(n10884), .Z(n16893) );
  INV_X2 U11320 ( .A(n17233), .ZN(n17264) );
  AND2_X2 U11321 ( .A1(n11809), .A2(n10156), .ZN(n11547) );
  INV_X2 U11322 ( .A(n18586), .ZN(n9583) );
  NAND2_X2 U11323 ( .A1(n18712), .A2(n18580), .ZN(n18639) );
  INV_X2 U11324 ( .A(n16234), .ZN(U215) );
  AND4_X1 U11325 ( .A1(n10076), .A2(n10075), .A3(n10074), .A4(n10073), .ZN(
        n10077) );
  AND2_X1 U11326 ( .A1(n10064), .A2(n10063), .ZN(n10065) );
  AND2_X1 U11327 ( .A1(n10069), .A2(n10068), .ZN(n9880) );
  CLKBUF_X2 U11328 ( .A(n11922), .Z(n12469) );
  CLKBUF_X3 U11329 ( .A(n11928), .Z(n12396) );
  INV_X2 U11330 ( .A(n10009), .ZN(n16992) );
  INV_X2 U11331 ( .A(n19038), .ZN(n18765) );
  BUF_X2 U11332 ( .A(n11892), .Z(n12642) );
  CLKBUF_X3 U11333 ( .A(n11922), .Z(n12636) );
  CLKBUF_X2 U11334 ( .A(n11927), .Z(n12503) );
  INV_X2 U11335 ( .A(n19920), .ZN(n19930) );
  INV_X2 U11336 ( .A(n14713), .ZN(n19026) );
  INV_X4 U11337 ( .A(n10892), .ZN(n9585) );
  INV_X2 U11338 ( .A(n20035), .ZN(n20053) );
  INV_X2 U11339 ( .A(n10814), .ZN(n16991) );
  INV_X2 U11340 ( .A(n11709), .ZN(n11622) );
  AND2_X2 U11341 ( .A1(n11616), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10280) );
  BUF_X2 U11342 ( .A(n10246), .Z(n11809) );
  BUF_X2 U11343 ( .A(n10252), .Z(n11668) );
  AND2_X2 U11344 ( .A1(n11859), .A2(n11852), .ZN(n12614) );
  BUF_X2 U11345 ( .A(n10072), .Z(n11787) );
  AND2_X2 U11346 ( .A1(n11851), .A2(n13424), .ZN(n12641) );
  BUF_X2 U11347 ( .A(n11893), .Z(n12644) );
  BUF_X2 U11348 ( .A(n10252), .Z(n11631) );
  AND2_X1 U11349 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10689), .ZN(
        n10745) );
  CLKBUF_X2 U11350 ( .A(n10726), .Z(n10887) );
  INV_X2 U11351 ( .A(n16237), .ZN(n16239) );
  AND2_X2 U11352 ( .A1(n11810), .A2(n10156), .ZN(n10274) );
  INV_X2 U11353 ( .A(n18713), .ZN(n18712) );
  AND2_X1 U11354 ( .A1(n11840), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11851) );
  CLKBUF_X1 U11355 ( .A(n20632), .Z(n20618) );
  NAND3_X1 U11356 ( .A1(n10687), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10701) );
  AND2_X1 U11357 ( .A1(n10058), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10252) );
  AND2_X2 U11358 ( .A1(n12091), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11859) );
  AND2_X2 U11359 ( .A1(n10059), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10253) );
  NOR3_X4 U11360 ( .A1(n16645), .A2(n18661), .A3(n18671), .ZN(n10708) );
  AND2_X1 U11361 ( .A1(n10062), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10072) );
  NAND2_X1 U11362 ( .A1(n18671), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10724) );
  AND2_X1 U11363 ( .A1(n11846), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11852) );
  AND2_X2 U11364 ( .A1(n11860), .A2(n13425), .ZN(n12296) );
  INV_X4 U11365 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18661) );
  AND2_X1 U11366 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13570) );
  NOR2_X2 U11367 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10059) );
  AND2_X1 U11368 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13569) );
  NOR2_X1 U11369 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11853) );
  NOR2_X2 U11370 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11860) );
  NOR2_X2 U11371 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13424) );
  INV_X1 U11372 ( .A(n9868), .ZN(n9586) );
  NAND2_X1 U11373 ( .A1(n10493), .A2(n10012), .ZN(n10495) );
  NAND2_X1 U11374 ( .A1(n12868), .A2(n15624), .ZN(n12867) );
  NAND2_X1 U11375 ( .A1(n13322), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20038) );
  NAND2_X1 U11376 ( .A1(n20194), .A2(n12001), .ZN(n12077) );
  INV_X1 U11377 ( .A(n15369), .ZN(n9587) );
  NOR2_X2 U11378 ( .A1(n11404), .A2(n10513), .ZN(n11400) );
  NOR2_X1 U11379 ( .A1(n17621), .A2(n17943), .ZN(n17620) );
  NAND2_X1 U11380 ( .A1(n10901), .A2(n17929), .ZN(n17931) );
  NOR2_X2 U11381 ( .A1(n11267), .A2(n11262), .ZN(n11257) );
  NOR4_X1 U11382 ( .A1(n15013), .A2(n15247), .A3(n15009), .A4(n15004), .ZN(
        n11280) );
  NAND2_X2 U11383 ( .A1(n11170), .A2(n11152), .ZN(n11151) );
  INV_X1 U11384 ( .A(n13192), .ZN(n9589) );
  INV_X1 U11385 ( .A(n11503), .ZN(n10530) );
  INV_X1 U11386 ( .A(n10221), .ZN(n9590) );
  NAND2_X1 U11387 ( .A1(n10524), .A2(n9566), .ZN(n10528) );
  INV_X1 U11388 ( .A(n10221), .ZN(n10510) );
  NOR2_X2 U11389 ( .A1(n16082), .A2(n17699), .ZN(n17608) );
  NOR2_X2 U11390 ( .A1(n16119), .A2(n16118), .ZN(n16089) );
  NAND2_X2 U11391 ( .A1(n14824), .A2(n14823), .ZN(n11704) );
  NAND2_X1 U11392 ( .A1(n10567), .A2(n10566), .ZN(n9591) );
  NAND2_X1 U11393 ( .A1(n10567), .A2(n10566), .ZN(n11035) );
  NOR2_X4 U11394 ( .A1(n10901), .A2(n17929), .ZN(n10902) );
  NOR2_X2 U11395 ( .A1(n17620), .A2(n10810), .ZN(n10901) );
  BUF_X1 U11396 ( .A(n11507), .Z(n9592) );
  BUF_X2 U11397 ( .A(n11507), .Z(n9593) );
  XNOR2_X1 U11398 ( .A(n9591), .B(n11034), .ZN(n11507) );
  NAND2_X2 U11399 ( .A1(n11464), .A2(n11463), .ZN(n13652) );
  NOR2_X2 U11400 ( .A1(n17041), .A2(n17037), .ZN(n17040) );
  NAND2_X1 U11401 ( .A1(n10538), .A2(n10537), .ZN(n10624) );
  OAI21_X2 U11402 ( .B1(n14949), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14943), .ZN(n15088) );
  OR2_X2 U11403 ( .A1(n11061), .A2(n18875), .ZN(n11071) );
  NAND2_X1 U11404 ( .A1(n11035), .A2(n10578), .ZN(n10581) );
  AND2_X2 U11405 ( .A1(n9823), .A2(n11076), .ZN(n11119) );
  NOR2_X2 U11406 ( .A1(n15002), .A2(n15261), .ZN(n15939) );
  OAI21_X2 U11407 ( .B1(n11223), .B2(n9770), .A(n9768), .ZN(n15002) );
  INV_X1 U11408 ( .A(n11154), .ZN(n9870) );
  NOR2_X2 U11409 ( .A1(n16413), .A2(n16587), .ZN(n16462) );
  NOR2_X4 U11410 ( .A1(n10502), .A2(n10515), .ZN(n10538) );
  OR2_X4 U11411 ( .A1(n14983), .A2(n11312), .ZN(n14984) );
  OAI211_X2 U11412 ( .C1(n11479), .C2(n11478), .A(n11474), .B(n11477), .ZN(
        n13941) );
  OR2_X1 U11413 ( .A1(n11059), .A2(n11061), .ZN(n11122) );
  OR2_X1 U11414 ( .A1(n11061), .A2(n11060), .ZN(n11124) );
  OR2_X1 U11415 ( .A1(n11054), .A2(n11061), .ZN(n19100) );
  AND2_X1 U11416 ( .A1(n11061), .A2(n15355), .ZN(n11076) );
  NAND2_X1 U11417 ( .A1(n9806), .A2(n9620), .ZN(n14934) );
  NAND2_X1 U11418 ( .A1(n15631), .A2(n12865), .ZN(n9907) );
  OR2_X1 U11419 ( .A1(n12879), .A2(n13382), .ZN(n9692) );
  NAND2_X1 U11420 ( .A1(n11964), .A2(n15460), .ZN(n11965) );
  NOR2_X1 U11421 ( .A1(n13641), .A2(n13647), .ZN(n9788) );
  NAND2_X1 U11422 ( .A1(n9859), .A2(n14589), .ZN(n9900) );
  AND2_X1 U11423 ( .A1(n14553), .A2(n9860), .ZN(n9859) );
  NOR2_X1 U11424 ( .A1(n9901), .A2(n9861), .ZN(n9860) );
  INV_X1 U11425 ( .A(n13676), .ZN(n9971) );
  XNOR2_X1 U11426 ( .A(n12798), .B(n12209), .ZN(n12814) );
  INV_X1 U11427 ( .A(n12311), .ZN(n12336) );
  NAND2_X1 U11428 ( .A1(n12163), .A2(n9972), .ZN(n12205) );
  AND2_X1 U11429 ( .A1(n9894), .A2(n9605), .ZN(n9893) );
  NAND2_X1 U11430 ( .A1(n12133), .A2(n12134), .ZN(n12161) );
  NAND2_X1 U11431 ( .A1(n10530), .A2(n10498), .ZN(n10509) );
  NAND2_X1 U11432 ( .A1(n11218), .A2(n11209), .ZN(n10195) );
  INV_X1 U11433 ( .A(n14081), .ZN(n9957) );
  INV_X1 U11434 ( .A(n14092), .ZN(n9798) );
  NAND2_X1 U11435 ( .A1(n14978), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9808) );
  INV_X1 U11436 ( .A(n14992), .ZN(n11493) );
  NAND2_X1 U11437 ( .A1(n9769), .A2(n9654), .ZN(n9768) );
  INV_X1 U11438 ( .A(n9774), .ZN(n9769) );
  AOI21_X1 U11439 ( .B1(n9779), .B2(n9777), .A(n9775), .ZN(n9774) );
  INV_X1 U11440 ( .A(n15276), .ZN(n9775) );
  INV_X1 U11441 ( .A(n9654), .ZN(n9772) );
  INV_X1 U11442 ( .A(n9777), .ZN(n9776) );
  OR2_X1 U11443 ( .A1(n19085), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10005) );
  NAND2_X1 U11444 ( .A1(n11503), .A2(n10498), .ZN(n10496) );
  NAND2_X1 U11445 ( .A1(n16044), .A2(n10287), .ZN(n10439) );
  INV_X1 U11446 ( .A(n10718), .ZN(n10892) );
  NOR2_X1 U11447 ( .A1(n16645), .A2(n10698), .ZN(n10718) );
  INV_X1 U11448 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n16702) );
  NAND2_X1 U11449 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17612), .ZN(
        n10952) );
  INV_X1 U11450 ( .A(n18490), .ZN(n16080) );
  NAND2_X1 U11451 ( .A1(n13039), .A2(n13434), .ZN(n13326) );
  INV_X1 U11452 ( .A(n13063), .ZN(n13292) );
  NOR3_X1 U11453 ( .A1(n14602), .A2(n13021), .A3(n9929), .ZN(n9690) );
  AND2_X1 U11454 ( .A1(n20031), .A2(n14607), .ZN(n9929) );
  NAND2_X1 U11455 ( .A1(n15631), .A2(n12870), .ZN(n12871) );
  NAND2_X1 U11456 ( .A1(n12891), .A2(n13295), .ZN(n13012) );
  INV_X1 U11457 ( .A(n14094), .ZN(n14100) );
  OR2_X1 U11458 ( .A1(n11495), .A2(n16042), .ZN(n15223) );
  OR2_X1 U11459 ( .A1(n11495), .A2(n11419), .ZN(n15221) );
  OAI211_X1 U11460 ( .C1(n10797), .C2(n16724), .A(n10807), .B(n10806), .ZN(
        n16082) );
  CLKBUF_X1 U11461 ( .A(n20042), .Z(n20001) );
  NAND2_X1 U11462 ( .A1(n9741), .A2(n9740), .ZN(n16083) );
  NAND2_X1 U11463 ( .A1(n10921), .A2(n10922), .ZN(n9740) );
  CLKBUF_X1 U11464 ( .A(n11036), .Z(n11045) );
  NOR2_X1 U11465 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10062) );
  NAND2_X1 U11466 ( .A1(n9850), .A2(n9849), .ZN(n12081) );
  AOI21_X1 U11467 ( .B1(n9851), .B2(n12056), .A(n12060), .ZN(n9849) );
  AOI21_X1 U11468 ( .B1(n12057), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n9852), 
        .ZN(n9851) );
  CLKBUF_X1 U11469 ( .A(n12005), .Z(n12006) );
  INV_X1 U11470 ( .A(n11303), .ZN(n9918) );
  NOR2_X1 U11471 ( .A1(n10520), .A2(n9868), .ZN(n9867) );
  NOR2_X1 U11472 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10058) );
  NAND2_X1 U11473 ( .A1(n10768), .A2(n17193), .ZN(n10781) );
  INV_X1 U11474 ( .A(n18054), .ZN(n10972) );
  NAND2_X1 U11475 ( .A1(n18661), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10698) );
  INV_X1 U11476 ( .A(n10822), .ZN(n9674) );
  AND2_X1 U11477 ( .A1(n9985), .A2(n14292), .ZN(n9984) );
  AND2_X1 U11478 ( .A1(n14311), .A2(n12522), .ZN(n9985) );
  INV_X1 U11479 ( .A(n14326), .ZN(n12522) );
  NAND2_X1 U11480 ( .A1(n14349), .A2(n9978), .ZN(n9977) );
  INV_X1 U11481 ( .A(n9979), .ZN(n9978) );
  OR2_X1 U11482 ( .A1(n13832), .A2(n14008), .ZN(n12313) );
  NAND2_X1 U11483 ( .A1(n12163), .A2(n12162), .ZN(n12183) );
  INV_X1 U11484 ( .A(n13041), .ZN(n12658) );
  AOI21_X1 U11485 ( .B1(n12867), .B2(n14621), .A(n12866), .ZN(n14482) );
  NAND2_X1 U11486 ( .A1(n14655), .A2(n9652), .ZN(n9938) );
  INV_X1 U11487 ( .A(n14322), .ZN(n9935) );
  AND2_X1 U11488 ( .A1(n12835), .A2(n9660), .ZN(n9899) );
  NOR2_X1 U11489 ( .A1(n9946), .A2(n15595), .ZN(n9945) );
  INV_X1 U11490 ( .A(n14013), .ZN(n9946) );
  INV_X1 U11491 ( .A(n9609), .ZN(n9944) );
  NAND2_X1 U11492 ( .A1(n15662), .A2(n9889), .ZN(n9888) );
  INV_X1 U11493 ( .A(n12805), .ZN(n9890) );
  INV_X1 U11494 ( .A(n9888), .ZN(n9886) );
  AND2_X1 U11495 ( .A1(n9972), .A2(n12207), .ZN(n9858) );
  INV_X1 U11496 ( .A(n12206), .ZN(n12207) );
  NAND2_X1 U11497 ( .A1(n12766), .A2(n20038), .ZN(n12772) );
  OR2_X1 U11498 ( .A1(n12054), .A2(n12053), .ZN(n12760) );
  INV_X1 U11499 ( .A(n13051), .ZN(n12080) );
  NOR2_X1 U11500 ( .A1(n14721), .A2(n14722), .ZN(n11445) );
  NOR2_X1 U11501 ( .A1(n11764), .A2(n9841), .ZN(n9839) );
  NAND2_X1 U11502 ( .A1(n11706), .A2(n11701), .ZN(n11707) );
  INV_X1 U11503 ( .A(n11704), .ZN(n11706) );
  NAND2_X1 U11504 ( .A1(n11574), .A2(n9847), .ZN(n9846) );
  INV_X1 U11505 ( .A(n14836), .ZN(n9847) );
  NOR2_X1 U11506 ( .A1(n13789), .A2(n9726), .ZN(n9725) );
  INV_X1 U11507 ( .A(n15299), .ZN(n9726) );
  NAND2_X1 U11508 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n9700) );
  NOR2_X1 U11509 ( .A1(n14760), .A2(n9707), .ZN(n9706) );
  NOR2_X1 U11510 ( .A1(n15983), .A2(n9702), .ZN(n9701) );
  INV_X1 U11511 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n9702) );
  INV_X1 U11512 ( .A(n10544), .ZN(n10547) );
  INV_X1 U11513 ( .A(n14749), .ZN(n9967) );
  INV_X1 U11514 ( .A(n9768), .ZN(n9767) );
  NOR2_X1 U11515 ( .A1(n15209), .A2(n9735), .ZN(n9734) );
  INV_X1 U11516 ( .A(n13959), .ZN(n9735) );
  INV_X1 U11517 ( .A(n13926), .ZN(n9956) );
  INV_X1 U11518 ( .A(n9987), .ZN(n9780) );
  INV_X1 U11519 ( .A(n15993), .ZN(n9814) );
  INV_X1 U11520 ( .A(n15075), .ZN(n9815) );
  OR2_X1 U11521 ( .A1(n11482), .A2(n11483), .ZN(n11488) );
  NOR2_X1 U11522 ( .A1(n13706), .A2(n9954), .ZN(n9953) );
  INV_X1 U11523 ( .A(n13693), .ZN(n9785) );
  OR2_X1 U11524 ( .A1(n9788), .A2(n9783), .ZN(n9782) );
  NAND2_X1 U11525 ( .A1(n13693), .A2(n14094), .ZN(n9783) );
  NOR2_X1 U11526 ( .A1(n9727), .A2(n10308), .ZN(n9730) );
  NAND2_X1 U11527 ( .A1(n9811), .A2(n9870), .ZN(n11469) );
  NAND2_X1 U11528 ( .A1(n10570), .A2(n10569), .ZN(n11032) );
  BUF_X1 U11529 ( .A(n10426), .Z(n11638) );
  NAND2_X1 U11530 ( .A1(n11381), .A2(n9586), .ZN(n11413) );
  NAND2_X1 U11531 ( .A1(n9997), .A2(n10214), .ZN(n10220) );
  NAND2_X1 U11532 ( .A1(n10007), .A2(n9998), .ZN(n10219) );
  NOR3_X1 U11533 ( .A1(n11001), .A2(n11010), .A3(n17060), .ZN(n10963) );
  XNOR2_X1 U11534 ( .A(n10929), .B(n10754), .ZN(n10737) );
  AND2_X1 U11535 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n10794), .ZN(
        n10795) );
  OAI21_X1 U11536 ( .B1(n16141), .B2(n16082), .A(n17597), .ZN(n10808) );
  NOR2_X1 U11537 ( .A1(n10946), .A2(n17630), .ZN(n10949) );
  NOR2_X1 U11538 ( .A1(n17189), .A2(n10781), .ZN(n10793) );
  AND2_X1 U11539 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n10934), .ZN(
        n10936) );
  NOR2_X1 U11540 ( .A1(n10929), .A2(n10754), .ZN(n10768) );
  NOR4_X1 U11541 ( .A1(n10972), .A2(n11010), .A3(n10964), .A4(n10965), .ZN(
        n10973) );
  NAND2_X1 U11542 ( .A1(n10956), .A2(n18501), .ZN(n15429) );
  NOR2_X1 U11543 ( .A1(n10889), .A2(n9664), .ZN(n9663) );
  INV_X1 U11544 ( .A(n10893), .ZN(n10895) );
  OAI221_X1 U11545 ( .B1(n18513), .B2(n17269), .C1(n18513), .C2(n18702), .A(
        n14063), .ZN(n15511) );
  INV_X1 U11546 ( .A(n13271), .ZN(n20789) );
  NAND2_X1 U11547 ( .A1(n15531), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13053) );
  INV_X1 U11548 ( .A(n12137), .ZN(n12668) );
  INV_X1 U11549 ( .A(n12854), .ZN(n12611) );
  NAND2_X1 U11550 ( .A1(n12204), .A2(n12203), .ZN(n13676) );
  INV_X1 U11551 ( .A(n13672), .ZN(n12203) );
  XNOR2_X1 U11552 ( .A(n13282), .B(n12764), .ZN(n13322) );
  NAND2_X1 U11553 ( .A1(n9693), .A2(n12729), .ZN(n13434) );
  NAND2_X1 U11554 ( .A1(n12727), .A2(n12728), .ZN(n9693) );
  NAND2_X1 U11555 ( .A1(n14484), .A2(n13028), .ZN(n14206) );
  NOR2_X1 U11556 ( .A1(n9681), .A2(n9638), .ZN(n14068) );
  NAND2_X1 U11557 ( .A1(n9913), .A2(n9912), .ZN(n9906) );
  INV_X1 U11558 ( .A(n14501), .ZN(n9913) );
  NOR2_X1 U11559 ( .A1(n13018), .A2(n9680), .ZN(n9679) );
  INV_X1 U11560 ( .A(n13017), .ZN(n9680) );
  INV_X1 U11561 ( .A(n13539), .ZN(n9940) );
  NOR2_X1 U11562 ( .A1(n9878), .A2(n9877), .ZN(n9873) );
  OR2_X1 U11563 ( .A1(n13539), .A2(n9942), .ZN(n13618) );
  NOR2_X1 U11564 ( .A1(n13539), .A2(n13538), .ZN(n13616) );
  INV_X1 U11565 ( .A(n14689), .ZN(n14638) );
  OR2_X1 U11566 ( .A1(n13012), .A2(n13145), .ZN(n13023) );
  AND4_X1 U11567 ( .A1(n11951), .A2(n11950), .A3(n11949), .A4(n11948), .ZN(
        n11952) );
  NAND2_X1 U11568 ( .A1(n12056), .A2(n12102), .ZN(n9897) );
  AND2_X1 U11569 ( .A1(n12102), .A2(n20071), .ZN(n9891) );
  NAND2_X1 U11570 ( .A1(n9898), .A2(n9618), .ZN(n9896) );
  NAND2_X1 U11571 ( .A1(n12104), .A2(n20071), .ZN(n9898) );
  NAND2_X1 U11572 ( .A1(n12161), .A2(n12136), .ZN(n20060) );
  INV_X1 U11573 ( .A(n12697), .ZN(n20072) );
  INV_X2 U11574 ( .A(n11921), .ZN(n20085) );
  AOI21_X1 U11575 ( .B1(n20773), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20242), 
        .ZN(n20629) );
  INV_X1 U11576 ( .A(n13434), .ZN(n15484) );
  INV_X1 U11577 ( .A(n11214), .ZN(n9923) );
  OAI21_X1 U11578 ( .B1(n14797), .B2(n11778), .A(n14793), .ZN(n14788) );
  NOR4_X2 U11579 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A4(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10426) );
  XNOR2_X1 U11580 ( .A(n11704), .B(n11701), .ZN(n14818) );
  OR2_X2 U11581 ( .A1(n14891), .A2(n14892), .ZN(n14889) );
  AND2_X1 U11582 ( .A1(n14772), .A2(n14773), .ZN(n14775) );
  INV_X1 U11583 ( .A(n18883), .ZN(n9842) );
  NAND2_X1 U11584 ( .A1(n9724), .A2(n9725), .ZN(n15298) );
  INV_X1 U11585 ( .A(n15332), .ZN(n9724) );
  NOR2_X1 U11586 ( .A1(n14827), .A2(n14826), .ZN(n14825) );
  INV_X1 U11587 ( .A(n10045), .ZN(n10018) );
  AOI21_X1 U11588 ( .B1(n11026), .B2(n11025), .A(n10591), .ZN(n13721) );
  NAND2_X1 U11589 ( .A1(n9949), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9948) );
  AND2_X1 U11590 ( .A1(n14936), .A2(n11324), .ZN(n11325) );
  NOR2_X1 U11591 ( .A1(n14938), .A2(n9659), .ZN(n9801) );
  INV_X1 U11592 ( .A(n14933), .ZN(n9804) );
  INV_X1 U11593 ( .A(n14969), .ZN(n9805) );
  AOI22_X1 U11594 ( .A1(n14990), .A2(n14991), .B1(n11308), .B2(n11307), .ZN(
        n14980) );
  OR2_X1 U11595 ( .A1(n15993), .A2(n9934), .ZN(n9933) );
  OR2_X1 U11596 ( .A1(n15916), .A2(n15070), .ZN(n9831) );
  NAND2_X1 U11597 ( .A1(n15320), .A2(n15222), .ZN(n15916) );
  OR2_X1 U11598 ( .A1(n11242), .A2(n11241), .ZN(n9777) );
  NAND2_X1 U11599 ( .A1(n13768), .A2(n15331), .ZN(n15332) );
  AND2_X1 U11600 ( .A1(n9719), .A2(n9630), .ZN(n9718) );
  OR2_X1 U11601 ( .A1(n13743), .A2(n10325), .ZN(n9719) );
  NAND2_X1 U11602 ( .A1(n9717), .A2(n9715), .ZN(n15339) );
  AOI21_X1 U11603 ( .B1(n9718), .B2(n13743), .A(n9716), .ZN(n9715) );
  NAND2_X1 U11604 ( .A1(n13701), .A2(n9718), .ZN(n9717) );
  INV_X1 U11605 ( .A(n15340), .ZN(n9716) );
  NAND2_X1 U11606 ( .A1(n9827), .A2(n9825), .ZN(n13857) );
  NAND2_X1 U11607 ( .A1(n9826), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9825) );
  NAND2_X1 U11608 ( .A1(n13718), .A2(n9828), .ZN(n9827) );
  OAI22_X1 U11609 ( .A1(n13714), .A2(n13715), .B1(n14195), .B2(n13860), .ZN(
        n13853) );
  INV_X1 U11610 ( .A(n9789), .ZN(n9786) );
  OAI21_X1 U11611 ( .B1(n13654), .B2(n14094), .A(n13693), .ZN(n9789) );
  BUF_X4 U11612 ( .A(n10514), .Z(n16044) );
  NAND2_X1 U11613 ( .A1(n11398), .A2(n13133), .ZN(n11495) );
  NAND2_X1 U11614 ( .A1(n13163), .A2(n13162), .ZN(n19609) );
  NOR2_X1 U11615 ( .A1(n11008), .A2(n11007), .ZN(n18490) );
  NAND2_X1 U11616 ( .A1(n16798), .A2(P3_EBX_REG_25__SCAN_IN), .ZN(n16786) );
  NAND2_X1 U11617 ( .A1(n16891), .A2(n9669), .ZN(n9670) );
  NOR2_X1 U11618 ( .A1(n16875), .A2(n16453), .ZN(n9669) );
  NAND2_X1 U11619 ( .A1(n17040), .A2(P3_EBX_REG_5__SCAN_IN), .ZN(n17032) );
  INV_X1 U11620 ( .A(n10704), .ZN(n16935) );
  OAI211_X1 U11621 ( .C1(n10009), .C2(n20936), .A(n10780), .B(n10779), .ZN(
        n10923) );
  INV_X1 U11622 ( .A(n10735), .ZN(n9746) );
  AND2_X1 U11623 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n9745)
         );
  NOR2_X1 U11624 ( .A1(n17011), .A2(n18267), .ZN(n9744) );
  INV_X1 U11625 ( .A(n10734), .ZN(n9747) );
  NAND2_X1 U11626 ( .A1(n9755), .A2(n10904), .ZN(n9754) );
  NAND2_X1 U11627 ( .A1(n17557), .A2(n10903), .ZN(n10904) );
  OR2_X1 U11628 ( .A1(n17557), .A2(n9756), .ZN(n9755) );
  XOR2_X1 U11629 ( .A(n17965), .B(n10769), .Z(n17656) );
  NOR2_X1 U11630 ( .A1(n17657), .A2(n17656), .ZN(n17655) );
  NAND2_X1 U11631 ( .A1(n17695), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17694) );
  INV_X1 U11632 ( .A(n18523), .ZN(n18533) );
  NOR2_X1 U11633 ( .A1(n13325), .A2(n12697), .ZN(n13126) );
  NAND2_X1 U11634 ( .A1(n9926), .A2(n9925), .ZN(n9924) );
  INV_X1 U11635 ( .A(n14086), .ZN(n9925) );
  NAND2_X1 U11636 ( .A1(n9928), .A2(n9927), .ZN(n9926) );
  AOI21_X1 U11637 ( .B1(n9613), .B2(n13022), .A(n20891), .ZN(n9927) );
  INV_X1 U11638 ( .A(n12994), .ZN(n9930) );
  AND2_X1 U11639 ( .A1(n9854), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9853) );
  NOR2_X1 U11640 ( .A1(n14597), .A2(n9690), .ZN(n9689) );
  OR2_X1 U11641 ( .A1(n20046), .A2(n15729), .ZN(n20018) );
  NOR2_X1 U11642 ( .A1(n13012), .A2(n12899), .ZN(n20042) );
  OR2_X1 U11643 ( .A1(n13012), .A2(n12896), .ZN(n20050) );
  INV_X1 U11644 ( .A(n20390), .ZN(n20366) );
  INV_X1 U11645 ( .A(n11399), .ZN(n19800) );
  NAND2_X1 U11646 ( .A1(n9694), .A2(n9567), .ZN(n14744) );
  NAND2_X1 U11647 ( .A1(n14780), .A2(n15019), .ZN(n9694) );
  XNOR2_X1 U11648 ( .A(n14118), .B(n14117), .ZN(n15811) );
  AND2_X1 U11649 ( .A1(n13189), .A2(n14096), .ZN(n18926) );
  OR2_X1 U11650 ( .A1(n13368), .A2(n11822), .ZN(n11823) );
  XNOR2_X1 U11651 ( .A(n14106), .B(n14105), .ZN(n14919) );
  OAI21_X1 U11652 ( .B1(n14149), .B2(n14148), .A(n14147), .ZN(n14150) );
  INV_X1 U11653 ( .A(n15352), .ZN(n16011) );
  INV_X1 U11654 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19797) );
  INV_X1 U11655 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19788) );
  NOR2_X1 U11656 ( .A1(n19516), .A2(n19388), .ZN(n19436) );
  NAND4_X1 U11657 ( .A1(n16287), .A2(P3_EBX_REG_31__SCAN_IN), .A3(n18702), 
        .A4(n16267), .ZN(n16653) );
  NOR2_X1 U11658 ( .A1(n11016), .A2(n9739), .ZN(n9738) );
  NOR2_X1 U11659 ( .A1(n16100), .A2(n17835), .ZN(n9739) );
  NOR2_X1 U11660 ( .A1(n18023), .A2(n17844), .ZN(n17878) );
  OR2_X1 U11661 ( .A1(n12702), .A2(n12701), .ZN(n12705) );
  INV_X1 U11662 ( .A(n12885), .ZN(n11964) );
  INV_X1 U11663 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12675) );
  AND2_X2 U11664 ( .A1(n11851), .A2(n13425), .ZN(n11927) );
  NOR2_X1 U11665 ( .A1(n9974), .A2(n9973), .ZN(n9972) );
  INV_X1 U11666 ( .A(n12184), .ZN(n9974) );
  INV_X1 U11667 ( .A(n12162), .ZN(n9973) );
  NAND3_X1 U11668 ( .A1(n11972), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n12697), 
        .ZN(n12718) );
  NAND2_X1 U11669 ( .A1(n20094), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12120) );
  NAND2_X1 U11670 ( .A1(n20072), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12119) );
  NAND2_X1 U11671 ( .A1(n11962), .A2(n11976), .ZN(n11919) );
  INV_X1 U11672 ( .A(n12718), .ZN(n12723) );
  AND2_X1 U11673 ( .A1(n11985), .A2(n11979), .ZN(n11978) );
  INV_X1 U11674 ( .A(n10253), .ZN(n11709) );
  NOR2_X1 U11675 ( .A1(n16044), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10296) );
  AND2_X1 U11676 ( .A1(n11150), .A2(n11149), .ZN(n11179) );
  NAND2_X1 U11677 ( .A1(n9821), .A2(n9819), .ZN(n9818) );
  INV_X1 U11678 ( .A(n11071), .ZN(n9821) );
  NOR2_X1 U11679 ( .A1(n9824), .A2(n9820), .ZN(n9819) );
  NAND2_X1 U11680 ( .A1(n11076), .A2(n9624), .ZN(n9817) );
  AOI21_X1 U11681 ( .B1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n15401), .A(
        n11089), .ZN(n11091) );
  AND2_X1 U11682 ( .A1(n14711), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10557) );
  NAND2_X1 U11683 ( .A1(n11824), .A2(n19065), .ZN(n10518) );
  NAND2_X1 U11684 ( .A1(n10517), .A2(n10516), .ZN(n10519) );
  NAND2_X1 U11685 ( .A1(n11824), .A2(n9590), .ZN(n9864) );
  NAND2_X1 U11686 ( .A1(n11385), .A2(n10221), .ZN(n9865) );
  AOI22_X1 U11687 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(n9568), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10205) );
  INV_X1 U11688 ( .A(n13104), .ZN(n11377) );
  INV_X1 U11689 ( .A(n9667), .ZN(n9666) );
  OAI211_X1 U11690 ( .C1(n10009), .C2(n18057), .A(n9621), .B(n9668), .ZN(n9667) );
  NAND2_X1 U11691 ( .A1(n16988), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n9668) );
  AOI22_X1 U11692 ( .A1(n10887), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9571), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n9665) );
  AOI21_X1 U11693 ( .B1(n12006), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12007), .ZN(n12016) );
  NOR2_X1 U11694 ( .A1(n15632), .A2(n12834), .ZN(n12835) );
  NAND2_X1 U11695 ( .A1(n12362), .A2(n9980), .ZN(n9979) );
  INV_X1 U11696 ( .A(n14024), .ZN(n9980) );
  NAND2_X1 U11697 ( .A1(n12304), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12305) );
  INV_X1 U11698 ( .A(n12303), .ZN(n12304) );
  AND3_X1 U11699 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A3(n12176), .ZN(n12196) );
  INV_X1 U11700 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12091) );
  NOR2_X1 U11701 ( .A1(n12718), .A2(n12779), .ZN(n12720) );
  NAND2_X1 U11702 ( .A1(n15625), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12868) );
  NOR2_X1 U11703 ( .A1(n12979), .A2(n9937), .ZN(n9936) );
  INV_X1 U11704 ( .A(n14654), .ZN(n9937) );
  AND2_X1 U11705 ( .A1(n14580), .A2(n14577), .ZN(n14566) );
  OR2_X1 U11706 ( .A1(n13538), .A2(n9941), .ZN(n9942) );
  NAND2_X1 U11707 ( .A1(n13434), .A2(n9692), .ZN(n12880) );
  NAND2_X1 U11708 ( .A1(n12085), .A2(n12084), .ZN(n12086) );
  OR2_X1 U11709 ( .A1(n12081), .A2(n12083), .ZN(n12084) );
  OAI21_X1 U11710 ( .B1(n20790), .B2(n15802), .A(n20758), .ZN(n20070) );
  NOR2_X1 U11711 ( .A1(n9916), .A2(n9915), .ZN(n9914) );
  NAND2_X1 U11712 ( .A1(n9918), .A2(n9917), .ZN(n9916) );
  NOR2_X1 U11713 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(P2_EBX_REG_25__SCAN_IN), 
        .ZN(n9917) );
  NAND2_X1 U11714 ( .A1(n14098), .A2(n11321), .ZN(n11319) );
  NAND2_X1 U11715 ( .A1(n9904), .A2(n9903), .ZN(n9902) );
  INV_X1 U11716 ( .A(n11252), .ZN(n9903) );
  OR2_X1 U11717 ( .A1(n11276), .A2(n11275), .ZN(n11259) );
  NOR2_X1 U11718 ( .A1(n11151), .A2(n9920), .ZN(n11232) );
  NAND2_X1 U11719 ( .A1(n9922), .A2(n9653), .ZN(n9920) );
  INV_X1 U11720 ( .A(n11033), .ZN(n10577) );
  INV_X1 U11721 ( .A(n9810), .ZN(n10511) );
  CLKBUF_X1 U11722 ( .A(n11631), .Z(n11801) );
  INV_X1 U11723 ( .A(n14807), .ZN(n9841) );
  NOR2_X1 U11724 ( .A1(n9965), .A2(n9964), .ZN(n9963) );
  INV_X1 U11725 ( .A(n11436), .ZN(n9964) );
  NOR2_X1 U11726 ( .A1(n15933), .A2(n9705), .ZN(n9704) );
  INV_X1 U11727 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n9705) );
  NAND2_X1 U11728 ( .A1(n9709), .A2(n9602), .ZN(n9713) );
  NOR2_X1 U11729 ( .A1(n19046), .A2(n9711), .ZN(n9710) );
  INV_X1 U11730 ( .A(n10021), .ZN(n9709) );
  NAND2_X1 U11731 ( .A1(n10583), .A2(n10582), .ZN(n10590) );
  NOR2_X1 U11732 ( .A1(n9951), .A2(n9950), .ZN(n9949) );
  NAND2_X1 U11733 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n9951) );
  INV_X1 U11734 ( .A(n11490), .ZN(n9934) );
  AND2_X1 U11735 ( .A1(n9960), .A2(n9959), .ZN(n9958) );
  INV_X1 U11736 ( .A(n13524), .ZN(n9959) );
  AND2_X1 U11737 ( .A1(n13414), .A2(n13786), .ZN(n9960) );
  INV_X1 U11738 ( .A(n11472), .ZN(n11483) );
  NAND2_X1 U11739 ( .A1(n13716), .A2(n13860), .ZN(n9828) );
  INV_X1 U11740 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15368) );
  NAND2_X1 U11741 ( .A1(n10521), .A2(n11400), .ZN(n9832) );
  AND2_X1 U11742 ( .A1(n11401), .A2(n11406), .ZN(n10521) );
  INV_X1 U11743 ( .A(n11041), .ZN(n9824) );
  NAND2_X2 U11744 ( .A1(n10115), .A2(n10114), .ZN(n10498) );
  NAND2_X1 U11745 ( .A1(n10113), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10114) );
  NAND2_X1 U11746 ( .A1(n9675), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10699) );
  NOR3_X1 U11747 ( .A1(n17413), .A2(n17397), .A3(n16369), .ZN(n17366) );
  NOR2_X1 U11748 ( .A1(n17444), .A2(n17443), .ZN(n17396) );
  NAND2_X1 U11749 ( .A1(n17403), .A2(n17432), .ZN(n17433) );
  AND2_X1 U11750 ( .A1(n10906), .A2(n9757), .ZN(n9756) );
  NOR2_X1 U11751 ( .A1(n10942), .A2(n17636), .ZN(n10944) );
  INV_X1 U11752 ( .A(n18511), .ZN(n18515) );
  AOI211_X1 U11753 ( .C1(n16965), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n10850), .B(n10849), .ZN(n10851) );
  NOR2_X1 U11754 ( .A1(n9674), .A2(n9673), .ZN(n9672) );
  AOI211_X1 U11755 ( .C1(n16893), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n10820), .B(n10819), .ZN(n10821) );
  NOR2_X1 U11756 ( .A1(n10009), .A2(n20898), .ZN(n9673) );
  AOI211_X1 U11757 ( .C1(n16893), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n10860), .B(n10859), .ZN(n10861) );
  NOR2_X1 U11758 ( .A1(n14282), .A2(n14069), .ZN(n14247) );
  OR2_X1 U11759 ( .A1(n9977), .A2(n9976), .ZN(n9975) );
  INV_X1 U11760 ( .A(n14393), .ZN(n9976) );
  OR2_X1 U11761 ( .A1(n12606), .A2(n14487), .ZN(n12607) );
  OR2_X1 U11762 ( .A1(n12610), .A2(n12609), .ZN(n12854) );
  AND2_X1 U11763 ( .A1(n9984), .A2(n9983), .ZN(n9982) );
  INV_X1 U11764 ( .A(n14284), .ZN(n9983) );
  NAND2_X1 U11765 ( .A1(n12561), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12606) );
  NAND2_X1 U11766 ( .A1(n14325), .A2(n9984), .ZN(n14291) );
  AND2_X1 U11767 ( .A1(n14325), .A2(n9985), .ZN(n14309) );
  AND2_X1 U11768 ( .A1(n12515), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12516) );
  OR2_X1 U11769 ( .A1(n12521), .A2(n12520), .ZN(n14326) );
  NOR2_X1 U11770 ( .A1(n12448), .A2(n14528), .ZN(n12413) );
  OR2_X1 U11771 ( .A1(n14395), .A2(n14383), .ZN(n14447) );
  NOR2_X1 U11772 ( .A1(n12392), .A2(n14560), .ZN(n12393) );
  NAND2_X1 U11773 ( .A1(n12393), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12465) );
  NOR2_X1 U11774 ( .A1(n12358), .A2(n14033), .ZN(n12359) );
  NAND2_X1 U11775 ( .A1(n12359), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12392) );
  NOR2_X1 U11776 ( .A1(n20874), .A2(n12305), .ZN(n12339) );
  CLKBUF_X1 U11777 ( .A(n14000), .Z(n14023) );
  AND2_X1 U11778 ( .A1(n13976), .A2(n13975), .ZN(n13978) );
  AND2_X1 U11779 ( .A1(n12262), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12263) );
  NAND2_X1 U11780 ( .A1(n12263), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12303) );
  AND2_X1 U11781 ( .A1(n12244), .A2(n13834), .ZN(n9969) );
  NAND2_X1 U11782 ( .A1(n9971), .A2(n12244), .ZN(n9970) );
  OR2_X1 U11783 ( .A1(n9639), .A2(n13876), .ZN(n13906) );
  NAND2_X1 U11784 ( .A1(n12210), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12214) );
  AND2_X1 U11785 ( .A1(n12196), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12210) );
  AOI21_X1 U11786 ( .B1(n12797), .B2(n12336), .A(n12202), .ZN(n13672) );
  NAND2_X1 U11787 ( .A1(n12182), .A2(n12181), .ZN(n13608) );
  NOR2_X1 U11788 ( .A1(n12138), .A2(n19895), .ZN(n12176) );
  INV_X1 U11789 ( .A(n9690), .ZN(n9928) );
  NOR2_X1 U11790 ( .A1(n12872), .A2(n9855), .ZN(n9854) );
  NAND2_X1 U11791 ( .A1(n14247), .A2(n14225), .ZN(n14244) );
  NAND2_X1 U11792 ( .A1(n14307), .A2(n14298), .ZN(n14300) );
  OR2_X1 U11793 ( .A1(n14300), .A2(n14280), .ZN(n14282) );
  NAND2_X1 U11794 ( .A1(n14484), .A2(n15631), .ZN(n9911) );
  NOR2_X1 U11795 ( .A1(n9938), .A2(n12983), .ZN(n14307) );
  NAND2_X1 U11796 ( .A1(n14655), .A2(n9936), .ZN(n14380) );
  NAND2_X1 U11797 ( .A1(n12838), .A2(n15631), .ZN(n15624) );
  NAND2_X1 U11798 ( .A1(n14655), .A2(n14654), .ZN(n15530) );
  AND2_X1 U11799 ( .A1(n14390), .A2(n14389), .ZN(n14655) );
  NOR2_X1 U11800 ( .A1(n14399), .A2(n14335), .ZN(n14390) );
  NAND2_X1 U11801 ( .A1(n14352), .A2(n12955), .ZN(n14397) );
  INV_X1 U11802 ( .A(n12831), .ZN(n15632) );
  AND2_X1 U11803 ( .A1(n13013), .A2(n14685), .ZN(n9691) );
  INV_X1 U11804 ( .A(n13973), .ZN(n9943) );
  NAND2_X1 U11805 ( .A1(n9944), .A2(n9945), .ZN(n14015) );
  NOR2_X1 U11806 ( .A1(n9609), .A2(n15595), .ZN(n15594) );
  AND3_X1 U11807 ( .A1(n12937), .A2(n12962), .A3(n12936), .ZN(n13836) );
  AND2_X1 U11808 ( .A1(n15651), .A2(n12819), .ZN(n13911) );
  INV_X1 U11809 ( .A(n9885), .ZN(n9884) );
  OAI21_X1 U11810 ( .B1(n9888), .B2(n12807), .A(n15661), .ZN(n9885) );
  NAND2_X1 U11811 ( .A1(n12927), .A2(n10000), .ZN(n13878) );
  OR2_X1 U11812 ( .A1(n20029), .A2(n20030), .ZN(n15765) );
  INV_X1 U11813 ( .A(n12778), .ZN(n9878) );
  NAND2_X1 U11814 ( .A1(n13023), .A2(n15765), .ZN(n15785) );
  NAND2_X1 U11815 ( .A1(n12914), .A2(n12913), .ZN(n13539) );
  INV_X1 U11816 ( .A(n13081), .ZN(n12914) );
  INV_X1 U11817 ( .A(n20018), .ZN(n15762) );
  NAND2_X1 U11818 ( .A1(n12763), .A2(n12762), .ZN(n13283) );
  NAND2_X1 U11819 ( .A1(n9893), .A2(n9896), .ZN(n12763) );
  CLKBUF_X1 U11820 ( .A(n12104), .Z(n20195) );
  OR2_X1 U11821 ( .A1(n9569), .A2(n20061), .ZN(n20365) );
  INV_X1 U11822 ( .A(n20242), .ZN(n20112) );
  NAND2_X1 U11823 ( .A1(n13623), .A2(n20059), .ZN(n20480) );
  NAND2_X1 U11824 ( .A1(n9981), .A2(n12078), .ZN(n20540) );
  INV_X1 U11825 ( .A(n20479), .ZN(n20334) );
  INV_X1 U11826 ( .A(n20423), .ZN(n20577) );
  NOR2_X1 U11827 ( .A1(n20059), .A2(n13625), .ZN(n20624) );
  INV_X1 U11828 ( .A(n14915), .ZN(n9698) );
  NOR2_X1 U11829 ( .A1(n14915), .A2(n15826), .ZN(n9696) );
  NAND2_X1 U11830 ( .A1(n14719), .A2(n9567), .ZN(n15825) );
  NAND2_X1 U11831 ( .A1(n11319), .A2(n11320), .ZN(n11328) );
  NOR2_X1 U11832 ( .A1(n11261), .A2(n9902), .ZN(n11249) );
  NAND2_X1 U11833 ( .A1(n11257), .A2(n11255), .ZN(n11276) );
  OR2_X1 U11834 ( .A1(n11151), .A2(n9921), .ZN(n11231) );
  INV_X1 U11835 ( .A(n9922), .ZN(n9921) );
  NOR2_X1 U11836 ( .A1(n14079), .A2(n14078), .ZN(n11542) );
  AND2_X1 U11837 ( .A1(n13457), .A2(n13773), .ZN(n13775) );
  AND2_X1 U11838 ( .A1(n11445), .A2(n11446), .ZN(n10476) );
  OAI211_X1 U11839 ( .C1(n11730), .C2(n9841), .A(n9838), .B(n11764), .ZN(
        n14792) );
  NAND2_X1 U11840 ( .A1(n9840), .A2(n14808), .ZN(n9838) );
  NOR2_X1 U11841 ( .A1(n9722), .A2(n9655), .ZN(n9721) );
  NAND2_X1 U11842 ( .A1(n9834), .A2(n9651), .ZN(n9833) );
  INV_X1 U11843 ( .A(n9722), .ZN(n9720) );
  NAND2_X1 U11844 ( .A1(n14818), .A2(n14817), .ZN(n14816) );
  NAND2_X1 U11845 ( .A1(n14164), .A2(n9995), .ZN(n14824) );
  NAND2_X1 U11846 ( .A1(n9844), .A2(n15884), .ZN(n9843) );
  INV_X1 U11847 ( .A(n9846), .ZN(n9844) );
  NAND2_X1 U11848 ( .A1(n9845), .A2(n11574), .ZN(n15890) );
  INV_X1 U11849 ( .A(n15892), .ZN(n9845) );
  INV_X1 U11850 ( .A(n9725), .ZN(n9723) );
  AND2_X1 U11851 ( .A1(n10320), .A2(n10319), .ZN(n13724) );
  AND2_X1 U11852 ( .A1(n11530), .A2(n11529), .ZN(n11531) );
  INV_X1 U11853 ( .A(n15407), .ZN(n15405) );
  XNOR2_X1 U11854 ( .A(n9563), .B(n10019), .ZN(n14157) );
  NAND2_X1 U11855 ( .A1(n9963), .A2(n14105), .ZN(n9962) );
  NOR3_X1 U11856 ( .A1(n10053), .A2(n14925), .A3(n10052), .ZN(n10055) );
  NOR3_X1 U11857 ( .A1(n14811), .A2(n14801), .A3(n9961), .ZN(n14106) );
  INV_X1 U11858 ( .A(n9963), .ZN(n9961) );
  OR2_X1 U11859 ( .A1(n14810), .A2(n14813), .ZN(n14811) );
  NAND2_X1 U11860 ( .A1(n10047), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10046) );
  NOR2_X2 U11861 ( .A1(n10046), .A2(n14972), .ZN(n10048) );
  NAND2_X1 U11862 ( .A1(n10041), .A2(n9608), .ZN(n10045) );
  AND2_X1 U11863 ( .A1(n10033), .A2(n9703), .ZN(n10038) );
  AND2_X1 U11864 ( .A1(n9600), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9703) );
  NAND2_X1 U11865 ( .A1(n10038), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10042) );
  AND2_X1 U11866 ( .A1(n13800), .A2(n9640), .ZN(n13925) );
  NAND2_X1 U11867 ( .A1(n10033), .A2(n9600), .ZN(n10039) );
  NAND2_X1 U11868 ( .A1(n13800), .A2(n9636), .ZN(n14083) );
  NAND2_X1 U11869 ( .A1(n10033), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10036) );
  NOR2_X1 U11870 ( .A1(n10034), .A2(n15953), .ZN(n10033) );
  NAND2_X1 U11871 ( .A1(n10030), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10034) );
  NAND2_X1 U11872 ( .A1(n10020), .A2(n9603), .ZN(n10031) );
  INV_X1 U11873 ( .A(n10025), .ZN(n10020) );
  NAND2_X1 U11874 ( .A1(n10020), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10028) );
  OR2_X1 U11875 ( .A1(n9713), .A2(n9712), .ZN(n10025) );
  NAND2_X1 U11876 ( .A1(n9709), .A2(n9710), .ZN(n10023) );
  NAND2_X1 U11877 ( .A1(n13721), .A2(n13720), .ZN(n13722) );
  NAND2_X1 U11878 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n10022), .ZN(
        n10021) );
  NOR2_X1 U11879 ( .A1(n10021), .A2(n19046), .ZN(n10024) );
  AND2_X1 U11880 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10022) );
  NAND2_X1 U11881 ( .A1(n10547), .A2(n9598), .ZN(n10548) );
  INV_X1 U11882 ( .A(n14140), .ZN(n9793) );
  NAND2_X1 U11883 ( .A1(n9794), .A2(n9797), .ZN(n14137) );
  NAND2_X1 U11884 ( .A1(n9947), .A2(n9949), .ZN(n14943) );
  INV_X1 U11885 ( .A(n14984), .ZN(n9947) );
  NOR2_X1 U11886 ( .A1(n14811), .A2(n14801), .ZN(n14802) );
  AND2_X1 U11887 ( .A1(n14802), .A2(n14716), .ZN(n14718) );
  OR2_X1 U11888 ( .A1(n15832), .A2(n14100), .ZN(n14936) );
  XNOR2_X1 U11889 ( .A(n14935), .B(n14936), .ZN(n14951) );
  NAND2_X1 U11890 ( .A1(n14757), .A2(n9642), .ZN(n14827) );
  INV_X1 U11891 ( .A(n14176), .ZN(n9966) );
  NAND2_X1 U11892 ( .A1(n14757), .A2(n9633), .ZN(n14751) );
  AOI21_X1 U11893 ( .B1(n11297), .B2(n9767), .A(n11296), .ZN(n9765) );
  NOR2_X1 U11894 ( .A1(n15059), .A2(n14838), .ZN(n14839) );
  NOR2_X1 U11895 ( .A1(n9733), .A2(n14905), .ZN(n9732) );
  INV_X1 U11896 ( .A(n9734), .ZN(n9733) );
  NAND2_X1 U11897 ( .A1(n13929), .A2(n9734), .ZN(n15211) );
  AND2_X1 U11898 ( .A1(n9640), .A2(n13897), .ZN(n9955) );
  OR2_X1 U11899 ( .A1(n15057), .A2(n15056), .ZN(n15059) );
  OAI21_X1 U11900 ( .B1(n15249), .B2(n15246), .A(n15006), .ZN(n15237) );
  NAND2_X1 U11901 ( .A1(n13775), .A2(n9960), .ZN(n13785) );
  AND2_X1 U11902 ( .A1(n13775), .A2(n13414), .ZN(n13787) );
  INV_X1 U11903 ( .A(n11485), .ZN(n9816) );
  AOI21_X1 U11904 ( .B1(n11485), .B2(n9815), .A(n9814), .ZN(n9812) );
  NAND2_X1 U11905 ( .A1(n11223), .A2(n9987), .ZN(n15285) );
  NAND2_X1 U11906 ( .A1(n15074), .A2(n15075), .ZN(n9813) );
  AND2_X1 U11907 ( .A1(n10342), .A2(n10341), .ZN(n13769) );
  AND2_X1 U11908 ( .A1(n9953), .A2(n13447), .ZN(n9952) );
  NAND2_X1 U11909 ( .A1(n9784), .A2(n9781), .ZN(n13714) );
  AND2_X1 U11910 ( .A1(n9782), .A2(n9787), .ZN(n9781) );
  NAND2_X1 U11911 ( .A1(n13641), .A2(n13647), .ZN(n9787) );
  OR2_X1 U11912 ( .A1(n10315), .A2(n10314), .ZN(n13643) );
  XNOR2_X1 U11913 ( .A(n11033), .B(n11032), .ZN(n11034) );
  INV_X1 U11914 ( .A(n9832), .ZN(n11438) );
  NOR2_X1 U11915 ( .A1(n10286), .A2(n10285), .ZN(n13347) );
  AOI21_X1 U11916 ( .B1(n11519), .B2(n11520), .A(n11518), .ZN(n13132) );
  NAND2_X1 U11917 ( .A1(n10251), .A2(n10156), .ZN(n10260) );
  AND2_X1 U11918 ( .A1(n19770), .A2(n19782), .ZN(n19757) );
  OR2_X1 U11919 ( .A1(n19770), .A2(n19782), .ZN(n19515) );
  INV_X1 U11920 ( .A(n19516), .ZN(n19445) );
  INV_X1 U11921 ( .A(n19482), .ZN(n19543) );
  INV_X1 U11922 ( .A(n19762), .ZN(n19604) );
  NAND2_X1 U11923 ( .A1(n10226), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10233) );
  INV_X1 U11925 ( .A(n16756), .ZN(n17010) );
  AND2_X1 U11926 ( .A1(n10718), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n9749) );
  NOR2_X1 U11927 ( .A1(n10725), .A2(n16700), .ZN(n10702) );
  NOR2_X1 U11928 ( .A1(n10697), .A2(n10696), .ZN(n10703) );
  AND2_X1 U11929 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10696) );
  AOI21_X2 U11930 ( .B1(n15511), .B2(n15510), .A(n18552), .ZN(n15513) );
  NAND4_X1 U11931 ( .A1(n10974), .A2(n18066), .A3(n10963), .A4(n16266), .ZN(
        n17271) );
  NOR2_X1 U11932 ( .A1(n17714), .A2(n17374), .ZN(n15451) );
  NOR2_X1 U11933 ( .A1(n17714), .A2(n17365), .ZN(n16112) );
  AOI21_X1 U11934 ( .B1(n15495), .B2(n18662), .A(n15496), .ZN(n10919) );
  NAND2_X1 U11935 ( .A1(n17352), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17329) );
  NOR2_X1 U11936 ( .A1(n17742), .A2(n17735), .ZN(n17375) );
  INV_X1 U11937 ( .A(n17396), .ZN(n17413) );
  NAND2_X1 U11938 ( .A1(n17603), .A2(n16084), .ZN(n17531) );
  NOR2_X1 U11939 ( .A1(n17616), .A2(n17617), .ZN(n17603) );
  INV_X1 U11940 ( .A(n17628), .ZN(n17632) );
  AOI211_X1 U11941 ( .C1(n16965), .C2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n10840), .B(n10839), .ZN(n10841) );
  INV_X1 U11942 ( .A(n16112), .ZN(n17703) );
  NAND2_X1 U11943 ( .A1(n17836), .A2(n10907), .ZN(n17735) );
  NAND2_X1 U11944 ( .A1(n17403), .A2(n10910), .ZN(n17383) );
  INV_X1 U11945 ( .A(n9756), .ZN(n9753) );
  INV_X1 U11946 ( .A(n17891), .ZN(n17567) );
  INV_X1 U11947 ( .A(n18514), .ZN(n18524) );
  NOR2_X1 U11948 ( .A1(n10954), .A2(n17599), .ZN(n17891) );
  NOR2_X1 U11949 ( .A1(n10948), .A2(n10952), .ZN(n10954) );
  AOI21_X1 U11950 ( .B1(n10953), .B2(n10952), .A(n10951), .ZN(n17600) );
  NOR2_X1 U11951 ( .A1(n17953), .A2(n17631), .ZN(n17630) );
  OAI211_X1 U11952 ( .C1(n9763), .C2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n9759), .B(n9758), .ZN(n17627) );
  NOR2_X1 U11953 ( .A1(n10940), .A2(n17651), .ZN(n17638) );
  NOR2_X1 U11954 ( .A1(n17965), .A2(n17652), .ZN(n17651) );
  INV_X1 U11955 ( .A(n17994), .ZN(n17970) );
  XNOR2_X1 U11956 ( .A(n17203), .B(n18663), .ZN(n17687) );
  NOR2_X1 U11957 ( .A1(n10687), .A2(n18671), .ZN(n18499) );
  NOR2_X1 U11958 ( .A1(n18717), .A2(n15430), .ZN(n18497) );
  CLKBUF_X1 U11959 ( .A(n10008), .Z(n16987) );
  INV_X1 U11960 ( .A(n16266), .ZN(n18040) );
  NOR2_X1 U11961 ( .A1(n10897), .A2(n10896), .ZN(n18054) );
  NAND2_X1 U11962 ( .A1(n10890), .A2(n9663), .ZN(n10897) );
  NAND2_X1 U11963 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10894) );
  OAI22_X1 U11964 ( .A1(n16081), .A2(n18491), .B1(n16080), .B2(n17999), .ZN(
        n18545) );
  NAND2_X1 U11965 ( .A1(n13058), .A2(n13057), .ZN(n19852) );
  AND2_X1 U11966 ( .A1(n15531), .A2(n13049), .ZN(n19870) );
  INV_X1 U11967 ( .A(n14406), .ZN(n19914) );
  AND2_X2 U11968 ( .A1(n12731), .A2(n13295), .ZN(n14428) );
  AND2_X1 U11969 ( .A1(n14429), .A2(n13387), .ZN(n14038) );
  AND2_X1 U11970 ( .A1(n13328), .A2(n15479), .ZN(n19922) );
  NOR2_X1 U11971 ( .A1(n19922), .A2(n19930), .ZN(n19934) );
  BUF_X1 U11972 ( .A(n19934), .Z(n19945) );
  XOR2_X1 U11973 ( .A(n14448), .B(n14447), .Z(n15619) );
  AND2_X1 U11974 ( .A1(n12852), .A2(n13434), .ZN(n19990) );
  INV_X1 U11975 ( .A(n19990), .ZN(n19822) );
  NAND2_X1 U11976 ( .A1(n14068), .A2(n9641), .ZN(n14602) );
  XNOR2_X1 U11977 ( .A(n14209), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14610) );
  XNOR2_X1 U11978 ( .A(n9909), .B(n9908), .ZN(n14618) );
  INV_X1 U11979 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9908) );
  NAND2_X1 U11980 ( .A1(n9911), .A2(n9910), .ZN(n9909) );
  NAND2_X1 U11981 ( .A1(n14483), .A2(n15651), .ZN(n9910) );
  NAND2_X1 U11982 ( .A1(n9906), .A2(n15631), .ZN(n14495) );
  NOR2_X1 U11983 ( .A1(n9678), .A2(n13019), .ZN(n9677) );
  INV_X1 U11984 ( .A(n9679), .ZN(n9678) );
  NAND2_X1 U11985 ( .A1(n14649), .A2(n13017), .ZN(n14637) );
  NOR2_X1 U11986 ( .A1(n15693), .A2(n13026), .ZN(n15683) );
  NAND2_X1 U11987 ( .A1(n9601), .A2(n9691), .ZN(n15687) );
  AND2_X1 U11988 ( .A1(n14042), .A2(n12826), .ZN(n9857) );
  INV_X1 U11989 ( .A(n9691), .ZN(n15731) );
  NOR2_X1 U11990 ( .A1(n13012), .A2(n15462), .ZN(n15729) );
  NAND2_X1 U11991 ( .A1(n15669), .A2(n12805), .ZN(n9887) );
  NAND2_X1 U11992 ( .A1(n19986), .A2(n19985), .ZN(n19988) );
  NAND2_X1 U11993 ( .A1(n13634), .A2(n12778), .ZN(n19986) );
  NAND2_X1 U11994 ( .A1(n15762), .A2(n13023), .ZN(n20031) );
  INV_X1 U11995 ( .A(n15729), .ZN(n20055) );
  INV_X1 U11996 ( .A(n13023), .ZN(n20047) );
  NOR2_X1 U11997 ( .A1(n13012), .A2(n13011), .ZN(n20046) );
  AND2_X1 U11998 ( .A1(n9894), .A2(n9897), .ZN(n9892) );
  NOR2_X1 U12000 ( .A1(n20756), .A2(n15484), .ZN(n14696) );
  INV_X1 U12001 ( .A(n20142), .ZN(n20147) );
  NAND2_X1 U12002 ( .A1(n20207), .A2(n20577), .ZN(n20228) );
  INV_X1 U12003 ( .A(n20206), .ZN(n20230) );
  INV_X1 U12004 ( .A(n20348), .ZN(n20353) );
  OAI211_X1 U12005 ( .C1(n20384), .C2(n20756), .A(n20433), .B(n20369), .ZN(
        n20387) );
  INV_X1 U12006 ( .A(n20440), .ZN(n20623) );
  INV_X1 U12007 ( .A(n20443), .ZN(n20638) );
  INV_X1 U12008 ( .A(n20447), .ZN(n20644) );
  INV_X1 U12009 ( .A(n20450), .ZN(n20650) );
  INV_X1 U12010 ( .A(n20453), .ZN(n20656) );
  INV_X1 U12011 ( .A(n20456), .ZN(n20662) );
  INV_X1 U12012 ( .A(n20459), .ZN(n20668) );
  INV_X1 U12013 ( .A(n20673), .ZN(n20680) );
  INV_X1 U12014 ( .A(n9699), .ZN(n10057) );
  OAI21_X1 U12015 ( .B1(n15825), .B2(n9697), .A(n9695), .ZN(n9699) );
  AOI21_X1 U12016 ( .B1(n9567), .B2(n9696), .A(n18863), .ZN(n9695) );
  NAND2_X1 U12017 ( .A1(n9567), .A2(n9698), .ZN(n9697) );
  NAND2_X1 U12018 ( .A1(n15838), .A2(n15839), .ZN(n15837) );
  NAND2_X1 U12019 ( .A1(n15851), .A2(n15852), .ZN(n15850) );
  OR2_X1 U12020 ( .A1(n11305), .A2(n11309), .ZN(n14741) );
  NAND2_X1 U12021 ( .A1(n14743), .A2(n13685), .ZN(n14733) );
  NAND2_X1 U12022 ( .A1(n14733), .A2(n14734), .ZN(n14732) );
  NAND2_X1 U12023 ( .A1(n14744), .A2(n15915), .ZN(n14743) );
  NAND2_X1 U12024 ( .A1(n13685), .A2(n9996), .ZN(n14780) );
  AND2_X1 U12025 ( .A1(n18725), .A2(n10485), .ZN(n18853) );
  OR2_X1 U12026 ( .A1(n11151), .A2(n9919), .ZN(n11225) );
  NAND2_X1 U12027 ( .A1(n9922), .A2(n10611), .ZN(n9919) );
  INV_X1 U12028 ( .A(n18853), .ZN(n18866) );
  OR2_X1 U12029 ( .A1(n18725), .A2(n10682), .ZN(n18856) );
  NAND2_X1 U12030 ( .A1(n13410), .A2(n9637), .ZN(n18884) );
  INV_X1 U12031 ( .A(n19782), .ZN(n15396) );
  NOR2_X1 U12032 ( .A1(n14808), .A2(n14807), .ZN(n14806) );
  INV_X1 U12033 ( .A(n18926), .ZN(n14908) );
  NOR2_X1 U12034 ( .A1(n15332), .A2(n13789), .ZN(n15300) );
  AND2_X1 U12035 ( .A1(n18986), .A2(n18935), .ZN(n18966) );
  OR2_X1 U12036 ( .A1(n14106), .A2(n11437), .ZN(n15821) );
  NOR2_X1 U12037 ( .A1(n14718), .A2(n11436), .ZN(n11437) );
  OR2_X1 U12038 ( .A1(n14948), .A2(n14963), .ZN(n15109) );
  INV_X1 U12039 ( .A(n9831), .ZN(n15917) );
  INV_X1 U12040 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13187) );
  AND2_X1 U12041 ( .A1(n19047), .A2(n14133), .ZN(n19037) );
  AND2_X1 U12042 ( .A1(n16020), .A2(n15225), .ZN(n15293) );
  AOI211_X1 U12043 ( .C1(n15811), .C2(n16010), .A(n14121), .B(n9736), .ZN(
        n14125) );
  NOR2_X1 U12044 ( .A1(n15810), .A2(n15343), .ZN(n9736) );
  XNOR2_X1 U12045 ( .A(n14093), .B(n10013), .ZN(n14932) );
  AND2_X1 U12046 ( .A1(n9806), .A2(n9615), .ZN(n14958) );
  NAND2_X1 U12047 ( .A1(n15352), .A2(n15223), .ZN(n9830) );
  OR2_X1 U12048 ( .A1(n15251), .A2(n9656), .ZN(n9829) );
  NAND2_X1 U12049 ( .A1(n9773), .A2(n9777), .ZN(n15278) );
  NAND2_X1 U12050 ( .A1(n11223), .A2(n9778), .ZN(n9773) );
  NAND2_X1 U12051 ( .A1(n9714), .A2(n9718), .ZN(n15341) );
  OR2_X1 U12052 ( .A1(n13701), .A2(n13743), .ZN(n9714) );
  AND2_X1 U12053 ( .A1(n13701), .A2(n10325), .ZN(n13744) );
  INV_X1 U12054 ( .A(n11061), .ZN(n11498) );
  NAND2_X1 U12055 ( .A1(n9789), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13639) );
  NAND2_X1 U12056 ( .A1(n9786), .A2(n13647), .ZN(n13640) );
  INV_X1 U12057 ( .A(n19334), .ZN(n19792) );
  OR2_X1 U12058 ( .A1(n19770), .A2(n15396), .ZN(n19762) );
  XNOR2_X1 U12059 ( .A(n13132), .B(n13131), .ZN(n19782) );
  CLKBUF_X1 U12060 ( .A(n10555), .Z(n16047) );
  INV_X1 U12061 ( .A(n19107), .ZN(n19123) );
  NOR2_X1 U12062 ( .A1(n19388), .A2(n19310), .ZN(n19147) );
  INV_X1 U12063 ( .A(n19324), .ZN(n19333) );
  OAI21_X1 U12064 ( .B1(n19423), .B2(n19439), .A(n19609), .ZN(n19441) );
  NOR2_X1 U12065 ( .A1(n19482), .A2(n19515), .ZN(n19504) );
  INV_X1 U12066 ( .A(n19663), .ZN(n19637) );
  INV_X1 U12067 ( .A(n19640), .ZN(n19659) );
  NOR2_X1 U12068 ( .A1(n18487), .A2(n17270), .ZN(n18718) );
  INV_X1 U12069 ( .A(n16268), .ZN(n16587) );
  INV_X1 U12070 ( .A(n16607), .ZN(n16642) );
  INV_X1 U12071 ( .A(n16649), .ZN(n16657) );
  NAND2_X1 U12072 ( .A1(n16789), .A2(n9661), .ZN(n16778) );
  NOR2_X2 U12073 ( .A1(n16795), .A2(n16772), .ZN(n16798) );
  AND2_X1 U12074 ( .A1(n16948), .A2(P3_EBX_REG_13__SCAN_IN), .ZN(n16932) );
  AND2_X1 U12075 ( .A1(n16971), .A2(P3_EBX_REG_12__SCAN_IN), .ZN(n16948) );
  NOR2_X2 U12076 ( .A1(n16982), .A2(n16951), .ZN(n16971) );
  NAND2_X1 U12077 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .ZN(n9676) );
  NAND2_X1 U12078 ( .A1(n17048), .A2(P3_EBX_REG_3__SCAN_IN), .ZN(n17041) );
  NAND2_X1 U12079 ( .A1(n17056), .A2(P3_EBX_REG_1__SCAN_IN), .ZN(n17044) );
  INV_X1 U12080 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n20934) );
  INV_X1 U12081 ( .A(n17077), .ZN(n17074) );
  INV_X1 U12082 ( .A(n17091), .ZN(n17087) );
  NOR2_X1 U12083 ( .A1(n17176), .A2(n17096), .ZN(n17092) );
  NOR3_X1 U12084 ( .A1(n17137), .A2(n17102), .A3(n17059), .ZN(n17097) );
  INV_X1 U12085 ( .A(n17125), .ZN(n17121) );
  NAND2_X1 U12086 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17141), .ZN(n17137) );
  INV_X1 U12087 ( .A(n17103), .ZN(n17135) );
  INV_X1 U12088 ( .A(n17119), .ZN(n17136) );
  NAND4_X1 U12089 ( .A1(n17171), .A2(P3_EAX_REG_14__SCAN_IN), .A3(
        P3_EAX_REG_13__SCAN_IN), .A4(n17058), .ZN(n17147) );
  NAND2_X1 U12090 ( .A1(n18525), .A2(n15513), .ZN(n17190) );
  AOI211_X1 U12091 ( .C1(n16965), .C2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n10751), .B(n10750), .ZN(n10752) );
  NAND2_X1 U12092 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10719) );
  NAND2_X1 U12093 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17207), .ZN(n17206) );
  NAND2_X1 U12094 ( .A1(n9747), .A2(n9743), .ZN(n9742) );
  NOR3_X1 U12095 ( .A1(n9746), .A2(n9745), .A3(n9744), .ZN(n9743) );
  INV_X1 U12096 ( .A(n17202), .ZN(n17205) );
  CLKBUF_X1 U12097 ( .A(n17313), .Z(n17310) );
  INV_X1 U12099 ( .A(n17847), .ZN(n17758) );
  NAND2_X1 U12100 ( .A1(n17632), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17616) );
  NOR2_X1 U12101 ( .A1(n18046), .A2(n16248), .ZN(n17689) );
  NOR2_X1 U12102 ( .A1(n18702), .A2(n16248), .ZN(n17685) );
  INV_X1 U12103 ( .A(n9596), .ZN(n17699) );
  AND2_X1 U12104 ( .A1(n9751), .A2(n9750), .ZN(n17476) );
  INV_X1 U12105 ( .A(n9752), .ZN(n17487) );
  OAI21_X1 U12106 ( .B1(n17501), .B2(n9753), .A(n17597), .ZN(n9752) );
  NAND2_X1 U12107 ( .A1(n17567), .A2(n17804), .ZN(n17847) );
  NOR2_X1 U12108 ( .A1(n17501), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17521) );
  NOR2_X1 U12109 ( .A1(n18497), .A2(n18506), .ZN(n17907) );
  NAND2_X1 U12110 ( .A1(n9650), .A2(n17640), .ZN(n17639) );
  INV_X1 U12111 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18530) );
  NOR2_X1 U12112 ( .A1(n18039), .A2(n14066), .ZN(n18684) );
  CLKBUF_X1 U12113 ( .A(n16226), .Z(n16234) );
  AOI21_X1 U12114 ( .B1(n14360), .B2(n20001), .A(n9924), .ZN(n13030) );
  NOR3_X1 U12115 ( .A1(n9689), .A2(n14598), .A3(n9617), .ZN(n14600) );
  AOI21_X1 U12116 ( .B1(n15817), .B2(n18874), .A(n15816), .ZN(n15818) );
  AND2_X1 U12117 ( .A1(n11838), .A2(n11837), .ZN(n11839) );
  AOI21_X1 U12118 ( .B1(n14151), .B2(n16014), .A(n14150), .ZN(n14152) );
  AOI211_X1 U12119 ( .C1(n9662), .C2(n16541), .A(n17821), .B(n16540), .ZN(
        n16542) );
  AOI211_X1 U12120 ( .C1(n9662), .C2(n16609), .A(n17821), .B(n16608), .ZN(
        n16610) );
  NAND2_X1 U12121 ( .A1(n16891), .A2(P3_EBX_REG_16__SCAN_IN), .ZN(n16876) );
  NAND2_X1 U12122 ( .A1(n9737), .A2(n18006), .ZN(n11024) );
  AOI21_X1 U12123 ( .B1(n16146), .B2(n16145), .A(n16144), .ZN(n16147) );
  AND3_X1 U12124 ( .A1(n10692), .A2(n10691), .A3(n10690), .ZN(n9597) );
  INV_X4 U12125 ( .A(n10886), .ZN(n10704) );
  NAND2_X2 U12126 ( .A1(n16141), .A2(n16082), .ZN(n17597) );
  INV_X1 U12128 ( .A(n12102), .ZN(n9852) );
  AND2_X1 U12129 ( .A1(n10546), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9598) );
  NAND2_X1 U12130 ( .A1(n9892), .A2(n9896), .ZN(n12758) );
  OR3_X1 U12131 ( .A1(n11261), .A2(n9902), .A3(P2_EBX_REG_20__SCAN_IN), .ZN(
        n9599) );
  AND2_X1 U12132 ( .A1(n9704), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9600) );
  NAND2_X1 U12133 ( .A1(n20031), .A2(n13015), .ZN(n9601) );
  INV_X1 U12134 ( .A(n10649), .ZN(n10584) );
  INV_X1 U12135 ( .A(n19085), .ZN(n9868) );
  AND2_X1 U12136 ( .A1(n9710), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9602) );
  AND2_X1 U12137 ( .A1(n9701), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9603) );
  INV_X1 U12138 ( .A(n9800), .ZN(n9799) );
  NOR2_X1 U12139 ( .A1(n9804), .A2(n9801), .ZN(n9800) );
  AND2_X1 U12140 ( .A1(n9933), .A2(n11492), .ZN(n9604) );
  AND2_X1 U12141 ( .A1(n9897), .A2(n9895), .ZN(n9605) );
  NOR2_X1 U12142 ( .A1(n10702), .A2(n9748), .ZN(n9606) );
  AND2_X1 U12143 ( .A1(n10041), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9607) );
  AND2_X1 U12144 ( .A1(n9706), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9608) );
  OR2_X1 U12145 ( .A1(n13392), .A2(n9728), .ZN(n13644) );
  OR2_X1 U12146 ( .A1(n13918), .A2(n13836), .ZN(n9609) );
  NAND2_X1 U12147 ( .A1(n14589), .A2(n13988), .ZN(n14041) );
  OR2_X2 U12148 ( .A1(n10701), .A2(n18661), .ZN(n10797) );
  OR3_X1 U12149 ( .A1(n14811), .A2(n14801), .A3(n9962), .ZN(n9610) );
  NAND2_X1 U12150 ( .A1(n9796), .A2(n9800), .ZN(n14093) );
  NOR2_X1 U12151 ( .A1(n14000), .A2(n14024), .ZN(n14022) );
  NOR2_X1 U12152 ( .A1(n14000), .A2(n9979), .ZN(n14050) );
  AND2_X1 U12153 ( .A1(n14325), .A2(n12522), .ZN(n14308) );
  AND4_X1 U12154 ( .A1(n11887), .A2(n11886), .A3(n11885), .A4(n11884), .ZN(
        n9611) );
  INV_X2 U12155 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10156) );
  AND2_X1 U12156 ( .A1(n9900), .A2(n9899), .ZN(n9612) );
  AND2_X1 U12157 ( .A1(n14649), .A2(n9679), .ZN(n9613) );
  INV_X1 U12158 ( .A(n13381), .ZN(n20109) );
  NOR2_X1 U12159 ( .A1(n14788), .A2(n14787), .ZN(n14786) );
  INV_X1 U12160 ( .A(n10741), .ZN(n17006) );
  NOR2_X1 U12161 ( .A1(n14000), .A2(n9977), .ZN(n14347) );
  AND2_X1 U12162 ( .A1(n14680), .A2(n14579), .ZN(n9614) );
  INV_X1 U12163 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9675) );
  NAND2_X1 U12164 ( .A1(n9806), .A2(n9807), .ZN(n14967) );
  AND2_X1 U12165 ( .A1(n9805), .A2(n9807), .ZN(n9615) );
  AND4_X1 U12166 ( .A1(n11907), .A2(n11906), .A3(n11905), .A4(n11904), .ZN(
        n9616) );
  NAND2_X1 U12167 ( .A1(n10510), .A2(n19085), .ZN(n10513) );
  AND2_X1 U12168 ( .A1(n14599), .A2(n20001), .ZN(n9617) );
  NAND2_X1 U12169 ( .A1(n10821), .A2(n9672), .ZN(n11001) );
  INV_X1 U12170 ( .A(n11001), .ZN(n9671) );
  NAND2_X1 U12171 ( .A1(n9900), .A2(n12835), .ZN(n14546) );
  AND2_X1 U12172 ( .A1(n12057), .A2(n9852), .ZN(n9618) );
  NAND2_X1 U12173 ( .A1(n11273), .A2(n9914), .ZN(n9619) );
  AND2_X1 U12174 ( .A1(n9615), .A2(n14960), .ZN(n9620) );
  OR2_X1 U12175 ( .A1(n16962), .A2(n20910), .ZN(n9621) );
  AND2_X1 U12176 ( .A1(n9958), .A2(n15273), .ZN(n9622) );
  AND3_X1 U12177 ( .A1(n10079), .A2(n10078), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9623) );
  AND2_X1 U12178 ( .A1(n14168), .A2(n9720), .ZN(n14856) );
  INV_X1 U12179 ( .A(n9803), .ZN(n9802) );
  NOR2_X1 U12180 ( .A1(n11330), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9803) );
  AND2_X1 U12181 ( .A1(n11043), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n9624) );
  AND3_X1 U12182 ( .A1(n9822), .A2(n9818), .A3(n9817), .ZN(n9625) );
  OR2_X1 U12183 ( .A1(n12725), .A2(n12724), .ZN(n9626) );
  NAND2_X1 U12184 ( .A1(n14484), .A2(n9854), .ZN(n9627) );
  NAND2_X1 U12185 ( .A1(n14168), .A2(n14169), .ZN(n14167) );
  XNOR2_X1 U12186 ( .A(n11482), .B(n11472), .ZN(n11471) );
  AND2_X1 U12187 ( .A1(n14325), .A2(n9982), .ZN(n12853) );
  NOR2_X1 U12188 ( .A1(n14984), .A2(n9951), .ZN(n14948) );
  NAND2_X1 U12189 ( .A1(n14138), .A2(n14136), .ZN(n9628) );
  INV_X1 U12190 ( .A(n9792), .ZN(n9791) );
  NAND2_X1 U12191 ( .A1(n9797), .A2(n9793), .ZN(n9792) );
  INV_X1 U12192 ( .A(n9779), .ZN(n9778) );
  OR2_X1 U12193 ( .A1(n11241), .A2(n9780), .ZN(n9779) );
  OR2_X1 U12194 ( .A1(n14167), .A2(n14881), .ZN(n9629) );
  INV_X4 U12195 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18671) );
  OR2_X1 U12196 ( .A1(n14100), .A2(n10439), .ZN(n9630) );
  NAND2_X1 U12197 ( .A1(n11180), .A2(n11179), .ZN(n11482) );
  AND2_X1 U12198 ( .A1(n9614), .A2(n12826), .ZN(n9631) );
  NAND2_X1 U12199 ( .A1(n20031), .A2(n13026), .ZN(n9632) );
  INV_X1 U12200 ( .A(n12786), .ZN(n9877) );
  AND2_X2 U12201 ( .A1(n13570), .A2(n13425), .ZN(n12022) );
  NAND2_X1 U12202 ( .A1(n13410), .A2(n11541), .ZN(n14077) );
  INV_X1 U12203 ( .A(n13988), .ZN(n9901) );
  XNOR2_X1 U12204 ( .A(n9610), .B(n14112), .ZN(n15810) );
  NOR2_X1 U12205 ( .A1(n15892), .A2(n9846), .ZN(n14835) );
  NOR2_X1 U12206 ( .A1(n10042), .A2(n15043), .ZN(n10041) );
  NAND2_X1 U12207 ( .A1(n13800), .A2(n13802), .ZN(n13801) );
  NAND2_X1 U12208 ( .A1(n14757), .A2(n14758), .ZN(n14748) );
  NAND2_X1 U12209 ( .A1(n13929), .A2(n13959), .ZN(n13958) );
  NAND2_X1 U12210 ( .A1(n14649), .A2(n9677), .ZN(n9681) );
  AND2_X1 U12211 ( .A1(n14758), .A2(n9967), .ZN(n9633) );
  AND2_X1 U12212 ( .A1(n10033), .A2(n9704), .ZN(n9634) );
  AND2_X1 U12213 ( .A1(n10020), .A2(n9701), .ZN(n9635) );
  AND2_X1 U12214 ( .A1(n13802), .A2(n9957), .ZN(n9636) );
  AND2_X1 U12215 ( .A1(n11541), .A2(n11542), .ZN(n9637) );
  NOR2_X1 U12216 ( .A1(n13927), .A2(n13928), .ZN(n13929) );
  AND2_X1 U12217 ( .A1(n20031), .A2(n13020), .ZN(n9638) );
  NOR2_X1 U12218 ( .A1(n13613), .A2(n13614), .ZN(n13607) );
  AND2_X1 U12219 ( .A1(n13775), .A2(n9958), .ZN(n13525) );
  INV_X1 U12220 ( .A(n12779), .ZN(n9895) );
  NAND2_X1 U12221 ( .A1(n9887), .A2(n12807), .ZN(n15660) );
  AND2_X1 U12222 ( .A1(n14839), .A2(n14769), .ZN(n14757) );
  NOR2_X1 U12223 ( .A1(n9970), .A2(n13675), .ZN(n13833) );
  NAND2_X1 U12224 ( .A1(n17475), .A2(n17597), .ZN(n17403) );
  AND2_X1 U12225 ( .A1(n13929), .A2(n9732), .ZN(n14772) );
  OR2_X1 U12226 ( .A1(n13675), .A2(n13676), .ZN(n9639) );
  AND2_X1 U12227 ( .A1(n9636), .A2(n9956), .ZN(n9640) );
  OR2_X1 U12228 ( .A1(n13022), .A2(n13028), .ZN(n9641) );
  AND2_X1 U12229 ( .A1(n9633), .A2(n9966), .ZN(n9642) );
  NOR2_X1 U12230 ( .A1(n12120), .A2(n12079), .ZN(n9643) );
  INV_X1 U12231 ( .A(n11976), .ZN(n13382) );
  NAND2_X1 U12232 ( .A1(n12671), .A2(n13381), .ZN(n11976) );
  OR2_X1 U12233 ( .A1(n9723), .A2(n15272), .ZN(n9644) );
  NAND2_X1 U12234 ( .A1(n14168), .A2(n9721), .ZN(n14721) );
  OR2_X1 U12235 ( .A1(n12723), .A2(n12721), .ZN(n9645) );
  AND2_X1 U12236 ( .A1(n9945), .A2(n9943), .ZN(n9646) );
  NOR2_X1 U12237 ( .A1(n9788), .A2(n9785), .ZN(n9647) );
  INV_X1 U12238 ( .A(n12134), .ZN(n13625) );
  NAND2_X1 U12239 ( .A1(n12132), .A2(n12131), .ZN(n12134) );
  AND2_X1 U12240 ( .A1(n9637), .A2(n9842), .ZN(n9648) );
  INV_X1 U12241 ( .A(n9771), .ZN(n9770) );
  NOR2_X1 U12242 ( .A1(n9776), .A2(n9772), .ZN(n9771) );
  NAND2_X1 U12243 ( .A1(n10525), .A2(n10511), .ZN(n10649) );
  NAND2_X1 U12244 ( .A1(n13820), .A2(n13821), .ZN(n13803) );
  NOR2_X1 U12245 ( .A1(n13448), .A2(n13456), .ZN(n13457) );
  NAND2_X1 U12246 ( .A1(n13775), .A2(n9622), .ZN(n13816) );
  NOR2_X1 U12247 ( .A1(n13392), .A2(n9729), .ZN(n13700) );
  OR2_X1 U12248 ( .A1(n10053), .A2(n10052), .ZN(n9649) );
  INV_X1 U12249 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20071) );
  AND2_X1 U12250 ( .A1(n13410), .A2(n9648), .ZN(n13895) );
  NOR2_X1 U12251 ( .A1(n15339), .A2(n13769), .ZN(n13768) );
  NOR2_X1 U12252 ( .A1(n17655), .A2(n10770), .ZN(n9650) );
  INV_X1 U12253 ( .A(n11298), .ZN(n9915) );
  XNOR2_X1 U12254 ( .A(n12772), .B(n20029), .ZN(n13515) );
  AND2_X1 U12255 ( .A1(n11764), .A2(n9841), .ZN(n9651) );
  AND2_X1 U12256 ( .A1(n9936), .A2(n9935), .ZN(n9652) );
  NAND2_X1 U12257 ( .A1(n9940), .A2(n9939), .ZN(n15779) );
  INV_X1 U12258 ( .A(n15779), .ZN(n12927) );
  NAND2_X1 U12259 ( .A1(n10041), .A2(n9706), .ZN(n9708) );
  AND2_X1 U12260 ( .A1(n10611), .A2(n10614), .ZN(n9653) );
  NAND2_X1 U12261 ( .A1(n11248), .A2(n11247), .ZN(n9654) );
  NAND2_X1 U12262 ( .A1(n14857), .A2(n14865), .ZN(n9655) );
  INV_X1 U12263 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n9762) );
  AND2_X1 U12264 ( .A1(n15224), .A2(n15252), .ZN(n9656) );
  AND2_X1 U12265 ( .A1(n13721), .A2(n9953), .ZN(n9657) );
  NOR2_X1 U12266 ( .A1(n13392), .A2(n10308), .ZN(n9658) );
  INV_X1 U12267 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n9707) );
  INV_X1 U12268 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n9820) );
  INV_X1 U12269 ( .A(n12865), .ZN(n9912) );
  AND2_X1 U12270 ( .A1(n11324), .A2(n11326), .ZN(n9659) );
  NOR2_X1 U12271 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n9660) );
  INV_X1 U12272 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n9757) );
  INV_X1 U12273 ( .A(n14119), .ZN(n9950) );
  INV_X1 U12274 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9711) );
  INV_X1 U12275 ( .A(n13028), .ZN(n9855) );
  AND2_X1 U12276 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n9661) );
  INV_X1 U12277 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n9712) );
  OR2_X1 U12278 ( .A1(n19761), .A2(n19334), .ZN(n19482) );
  OR2_X1 U12279 ( .A1(n19761), .A2(n19792), .ZN(n19516) );
  AOI22_X2 U12280 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19079), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19078), .ZN(n19621) );
  AOI22_X2 U12281 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19079), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19078), .ZN(n19627) );
  AOI22_X2 U12282 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19079), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19078), .ZN(n19653) );
  NOR3_X2 U12283 ( .A1(n18400), .A2(n18530), .A3(n18167), .ZN(n18141) );
  AOI22_X2 U12284 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20114), .B1(DATAI_26_), 
        .B2(n20069), .ZN(n20648) );
  NOR3_X2 U12285 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18400), .A3(
        n18258), .ZN(n18230) );
  INV_X1 U12286 ( .A(n11250), .ZN(n9904) );
  CLKBUF_X1 U12287 ( .A(n18557), .Z(n9662) );
  NOR4_X1 U12288 ( .A1(n18664), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .A4(P3_STATEBS16_REG_SCAN_IN), .ZN(n18557)
         );
  AOI22_X2 U12289 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20114), .B1(DATAI_24_), 
        .B2(n20069), .ZN(n20636) );
  AOI22_X2 U12290 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19078), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19079), .ZN(n19633) );
  NAND3_X1 U12291 ( .A1(n10888), .A2(n9666), .A3(n9665), .ZN(n9664) );
  INV_X1 U12292 ( .A(n9670), .ZN(n16890) );
  NOR2_X4 U12293 ( .A1(n16873), .A2(n16847), .ZN(n16861) );
  NOR2_X4 U12294 ( .A1(n16786), .A2(n16773), .ZN(n16789) );
  OAI22_X2 U12295 ( .A1(n15430), .A2(n16080), .B1(n15428), .B2(n15429), .ZN(
        n15509) );
  AND2_X2 U12296 ( .A1(n18054), .A2(n9671), .ZN(n18501) );
  AND2_X2 U12297 ( .A1(n17026), .A2(P3_EBX_REG_8__SCAN_IN), .ZN(n16985) );
  NOR2_X2 U12298 ( .A1(n17032), .A2(n9676), .ZN(n17026) );
  NAND2_X1 U12299 ( .A1(n9682), .A2(n9626), .ZN(n12726) );
  NAND2_X1 U12300 ( .A1(n9683), .A2(n9645), .ZN(n9682) );
  NAND2_X1 U12301 ( .A1(n9685), .A2(n9684), .ZN(n9683) );
  NAND2_X1 U12302 ( .A1(n12720), .A2(n12719), .ZN(n9684) );
  NAND2_X1 U12303 ( .A1(n9687), .A2(n9686), .ZN(n9685) );
  NAND2_X1 U12304 ( .A1(n12718), .A2(n12719), .ZN(n9686) );
  NAND2_X1 U12305 ( .A1(n9688), .A2(n12717), .ZN(n9687) );
  NAND3_X1 U12306 ( .A1(n12712), .A2(n12710), .A3(n12711), .ZN(n9688) );
  NAND3_X1 U12307 ( .A1(n9601), .A2(n9691), .A3(n9632), .ZN(n15679) );
  NAND2_X1 U12308 ( .A1(n15825), .A2(n15826), .ZN(n15824) );
  NAND2_X1 U12309 ( .A1(n15824), .A2(n9567), .ZN(n10056) );
  INV_X1 U12310 ( .A(n9708), .ZN(n10044) );
  INV_X1 U12311 ( .A(n9713), .ZN(n10026) );
  NAND3_X1 U12312 ( .A1(n10460), .A2(n10463), .A3(n14169), .ZN(n9722) );
  INV_X1 U12313 ( .A(n13643), .ZN(n9727) );
  INV_X1 U12314 ( .A(n9730), .ZN(n9728) );
  NAND2_X1 U12315 ( .A1(n9731), .A2(n9730), .ZN(n9729) );
  INV_X1 U12316 ( .A(n13724), .ZN(n9731) );
  NOR2_X1 U12317 ( .A1(n13391), .A2(n13390), .ZN(n13392) );
  NAND3_X1 U12318 ( .A1(n10918), .A2(n10920), .A3(n11022), .ZN(n9741) );
  NAND4_X1 U12319 ( .A1(n10700), .A2(n9606), .A3(n10703), .A4(n9597), .ZN(
        n17203) );
  OR2_X1 U12320 ( .A1(n10693), .A2(n9749), .ZN(n9748) );
  NAND2_X1 U12321 ( .A1(n9580), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9750) );
  NAND3_X1 U12322 ( .A1(n9751), .A2(n17819), .A3(n9750), .ZN(n17475) );
  NAND2_X1 U12323 ( .A1(n9760), .A2(n17656), .ZN(n9758) );
  NAND2_X1 U12324 ( .A1(n9760), .A2(n17657), .ZN(n9759) );
  NOR2_X1 U12325 ( .A1(n17640), .A2(n9762), .ZN(n9761) );
  INV_X1 U12326 ( .A(n17640), .ZN(n9763) );
  NAND2_X1 U12327 ( .A1(n11297), .A2(n9771), .ZN(n9766) );
  INV_X1 U12328 ( .A(n9764), .ZN(n15154) );
  NAND2_X1 U12329 ( .A1(n13654), .A2(n9647), .ZN(n9784) );
  INV_X1 U12330 ( .A(n11331), .ZN(n9795) );
  NAND2_X1 U12331 ( .A1(n11331), .A2(n9802), .ZN(n9796) );
  OR2_X1 U12332 ( .A1(n11331), .A2(n9799), .ZN(n9794) );
  AOI21_X2 U12333 ( .B1(n9800), .B2(n9803), .A(n9798), .ZN(n9797) );
  INV_X1 U12334 ( .A(n14978), .ZN(n9809) );
  NAND2_X1 U12335 ( .A1(n10500), .A2(n10499), .ZN(n9810) );
  NOR2_X1 U12336 ( .A1(n9810), .A2(n11408), .ZN(n11822) );
  AND2_X1 U12337 ( .A1(n15373), .A2(n9810), .ZN(n11419) );
  NAND3_X1 U12338 ( .A1(n9811), .A2(n9870), .A3(n10316), .ZN(n11467) );
  INV_X1 U12339 ( .A(n11155), .ZN(n9811) );
  OAI21_X1 U12340 ( .B1(n9816), .B2(n15074), .A(n9812), .ZN(n9932) );
  XNOR2_X2 U12341 ( .A(n11484), .B(n15342), .ZN(n15074) );
  NOR2_X2 U12342 ( .A1(n11071), .A2(n9824), .ZN(n19205) );
  NAND3_X1 U12343 ( .A1(n9823), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A3(
        n11076), .ZN(n9822) );
  AND2_X2 U12344 ( .A1(n11076), .A2(n11043), .ZN(n11134) );
  INV_X1 U12345 ( .A(n13716), .ZN(n9826) );
  NAND2_X1 U12346 ( .A1(n13854), .A2(n13857), .ZN(n11475) );
  NAND4_X1 U12347 ( .A1(n9832), .A2(n10555), .A3(n10533), .A4(n10534), .ZN(
        n10535) );
  NAND2_X1 U12348 ( .A1(n13353), .A2(n9832), .ZN(n15378) );
  AOI22_X1 U12349 ( .A1(n9573), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(n9564), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10078) );
  AND2_X2 U12350 ( .A1(n11364), .A2(n11399), .ZN(n11404) );
  OR2_X2 U12351 ( .A1(n16045), .A2(n10514), .ZN(n11399) );
  NAND3_X1 U12352 ( .A1(n9837), .A2(n9835), .A3(n9833), .ZN(n14799) );
  INV_X1 U12353 ( .A(n14808), .ZN(n9834) );
  OAI21_X1 U12354 ( .B1(n11730), .B2(n9839), .A(n9836), .ZN(n9835) );
  NAND2_X1 U12355 ( .A1(n11730), .A2(n11763), .ZN(n9836) );
  NAND3_X1 U12356 ( .A1(n9840), .A2(n11763), .A3(n14808), .ZN(n9837) );
  INV_X1 U12357 ( .A(n11730), .ZN(n9840) );
  NOR2_X2 U12358 ( .A1(n15892), .A2(n9843), .ZN(n15886) );
  NAND2_X1 U12359 ( .A1(n9848), .A2(n11502), .ZN(n11505) );
  NAND2_X1 U12360 ( .A1(n11061), .A2(n11520), .ZN(n9848) );
  NAND2_X1 U12361 ( .A1(n12104), .A2(n9851), .ZN(n9850) );
  OR2_X2 U12362 ( .A1(n12867), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14501) );
  NAND2_X1 U12363 ( .A1(n14484), .A2(n9853), .ZN(n9856) );
  OAI21_X2 U12364 ( .B1(n14473), .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n9856), .ZN(n12873) );
  XNOR2_X1 U12365 ( .A(n14581), .B(n9857), .ZN(n15732) );
  NAND2_X4 U12366 ( .A1(n12798), .A2(n12751), .ZN(n15651) );
  NOR2_X1 U12367 ( .A1(n15631), .A2(n13014), .ZN(n9861) );
  AND2_X2 U12368 ( .A1(n10245), .A2(n10244), .ZN(n10493) );
  NAND2_X1 U12369 ( .A1(n12757), .A2(n12756), .ZN(n12764) );
  NAND2_X1 U12370 ( .A1(n11381), .A2(n9867), .ZN(n9866) );
  NAND2_X1 U12371 ( .A1(n9866), .A2(n9869), .ZN(n10544) );
  NAND3_X1 U12372 ( .A1(n10500), .A2(n10499), .A3(n10520), .ZN(n9869) );
  OAI21_X1 U12373 ( .B1(n13634), .B2(n9876), .A(n9871), .ZN(n15673) );
  AOI21_X1 U12374 ( .B1(n9878), .B2(n19985), .A(n9877), .ZN(n9871) );
  NAND2_X1 U12375 ( .A1(n9874), .A2(n9872), .ZN(n15675) );
  NAND2_X1 U12376 ( .A1(n13634), .A2(n9873), .ZN(n9872) );
  AND2_X1 U12377 ( .A1(n15672), .A2(n9875), .ZN(n9874) );
  NAND2_X1 U12378 ( .A1(n9876), .A2(n12786), .ZN(n9875) );
  INV_X1 U12379 ( .A(n19985), .ZN(n9876) );
  NAND3_X1 U12380 ( .A1(n9623), .A2(n10080), .A3(n10081), .ZN(n9881) );
  NAND2_X1 U12381 ( .A1(n15669), .A2(n9886), .ZN(n9883) );
  NAND2_X1 U12382 ( .A1(n9883), .A2(n9884), .ZN(n13910) );
  NAND2_X1 U12383 ( .A1(n9890), .A2(n12807), .ZN(n9889) );
  NAND2_X1 U12384 ( .A1(n12104), .A2(n9891), .ZN(n9894) );
  OR2_X2 U12385 ( .A1(n11261), .A2(n11252), .ZN(n11254) );
  NAND3_X2 U12386 ( .A1(n9905), .A2(n12869), .A3(n9907), .ZN(n14484) );
  NOR2_X1 U12387 ( .A1(n11304), .A2(n11303), .ZN(n11309) );
  NOR3_X2 U12388 ( .A1(n11304), .A2(n11303), .A3(P2_EBX_REG_24__SCAN_IN), .ZN(
        n11316) );
  NOR2_X2 U12389 ( .A1(n11151), .A2(n10195), .ZN(n11215) );
  MUX2_X1 U12390 ( .A(n14250), .B(n12993), .S(n14244), .Z(n9931) );
  OAI21_X2 U12391 ( .B1(n15992), .B2(n9934), .A(n9604), .ZN(n14992) );
  INV_X1 U12392 ( .A(n9938), .ZN(n14323) );
  INV_X1 U12393 ( .A(n13615), .ZN(n9941) );
  NAND2_X1 U12394 ( .A1(n9944), .A2(n9646), .ZN(n14019) );
  NOR2_X2 U12395 ( .A1(n14984), .A2(n15115), .ZN(n14971) );
  NAND2_X1 U12396 ( .A1(n13721), .A2(n9952), .ZN(n13448) );
  INV_X1 U12397 ( .A(n13720), .ZN(n9954) );
  NAND2_X1 U12398 ( .A1(n13800), .A2(n9955), .ZN(n15057) );
  INV_X1 U12399 ( .A(n14716), .ZN(n9965) );
  INV_X1 U12400 ( .A(n13675), .ZN(n9968) );
  NAND3_X1 U12401 ( .A1(n9971), .A2(n9969), .A3(n9968), .ZN(n13832) );
  NOR2_X2 U12402 ( .A1(n14000), .A2(n9975), .ZN(n14441) );
  NAND2_X1 U12403 ( .A1(n20540), .A2(n12077), .ZN(n13051) );
  INV_X1 U12404 ( .A(n20194), .ZN(n9981) );
  NAND2_X1 U12405 ( .A1(n15886), .A2(n14832), .ZN(n14891) );
  AOI22_X1 U12406 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n11120), .B1(
        n19419), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11109) );
  NOR3_X4 U12407 ( .A1(n11333), .A2(n14100), .A3(n15115), .ZN(n14968) );
  AOI211_X2 U12408 ( .C1(n19042), .C2(n15849), .A(n14965), .B(n14964), .ZN(
        n14966) );
  NAND2_X1 U12409 ( .A1(n13277), .A2(n13276), .ZN(n13275) );
  AOI211_X2 U12410 ( .C1(n15112), .C2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15111), .B(n15110), .ZN(n15113) );
  NAND2_X1 U12411 ( .A1(n13278), .A2(n11055), .ZN(n11187) );
  NAND2_X1 U12412 ( .A1(n13278), .A2(n11050), .ZN(n11189) );
  NAND2_X1 U12413 ( .A1(n13278), .A2(n11044), .ZN(n11123) );
  NAND2_X1 U12414 ( .A1(n10011), .A2(n14152), .ZN(n14153) );
  OAI211_X1 U12415 ( .C1(n14218), .C2(n19995), .A(n14217), .B(n14216), .ZN(
        n14219) );
  INV_X1 U12416 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11840) );
  NOR2_X1 U12417 ( .A1(n11187), .A2(n11092), .ZN(n11095) );
  NAND2_X1 U12418 ( .A1(n11452), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13855) );
  CLKBUF_X1 U12419 ( .A(n13051), .Z(n20571) );
  INV_X1 U12420 ( .A(n14792), .ZN(n11778) );
  INV_X1 U12421 ( .A(n11986), .ZN(n11983) );
  NAND2_X1 U12422 ( .A1(n12033), .A2(n12031), .ZN(n12078) );
  NAND2_X1 U12423 ( .A1(n11988), .A2(n11987), .ZN(n12033) );
  OR2_X1 U12424 ( .A1(n14206), .A2(n15631), .ZN(n14207) );
  NAND2_X1 U12425 ( .A1(n14125), .A2(n10010), .ZN(n14126) );
  NAND2_X1 U12426 ( .A1(n12135), .A2(n12088), .ZN(n13600) );
  INV_X1 U12427 ( .A(n11467), .ZN(n11180) );
  XNOR2_X1 U12428 ( .A(n11467), .B(n11179), .ZN(n11452) );
  NAND2_X1 U12429 ( .A1(n13515), .A2(n13516), .ZN(n13517) );
  NOR2_X2 U12430 ( .A1(n14484), .A2(n12871), .ZN(n14205) );
  NOR2_X2 U12431 ( .A1(n14372), .A2(n14373), .ZN(n14325) );
  NAND2_X1 U12432 ( .A1(n14441), .A2(n12468), .ZN(n14372) );
  NAND2_X1 U12433 ( .A1(n14825), .A2(n14819), .ZN(n14810) );
  NAND2_X1 U12434 ( .A1(n12996), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11985) );
  NOR2_X1 U12435 ( .A1(n11123), .A2(n11663), .ZN(n11098) );
  CLKBUF_X1 U12436 ( .A(n12674), .Z(n15793) );
  XNOR2_X1 U12437 ( .A(n14104), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14161) );
  AOI21_X1 U12438 ( .B1(n14161), .B2(n16011), .A(n14126), .ZN(n14127) );
  NAND2_X1 U12439 ( .A1(n11963), .A2(n12759), .ZN(n11989) );
  OAI21_X1 U12440 ( .B1(n13277), .B2(n13276), .A(n13275), .ZN(n19761) );
  NAND2_X1 U12441 ( .A1(n13275), .A2(n11531), .ZN(n13410) );
  NOR2_X2 U12442 ( .A1(n13816), .A2(n13817), .ZN(n13800) );
  NOR3_X2 U12443 ( .A1(n17382), .A2(n17404), .A3(n17756), .ZN(n17377) );
  OR2_X2 U12444 ( .A1(n12087), .A2(n12086), .ZN(n12135) );
  AOI21_X2 U12445 ( .B1(n12080), .B2(n20071), .A(n9643), .ZN(n12752) );
  AOI21_X1 U12446 ( .B1(n14921), .B2(n16011), .A(n14153), .ZN(n14154) );
  AOI21_X2 U12447 ( .B1(n13969), .B2(n12313), .A(n12312), .ZN(n13970) );
  AND2_X1 U12448 ( .A1(n13577), .A2(n20099), .ZN(n12673) );
  NAND2_X1 U12449 ( .A1(n20104), .A2(n11971), .ZN(n11963) );
  AND2_X2 U12450 ( .A1(n11971), .A2(n11960), .ZN(n13000) );
  INV_X1 U12451 ( .A(n11971), .ZN(n20099) );
  CLKBUF_X1 U12452 ( .A(n12882), .Z(n13142) );
  INV_X1 U12453 ( .A(n17199), .ZN(n17172) );
  AND2_X1 U12454 ( .A1(n17597), .A2(n17727), .ZN(n9986) );
  AND2_X1 U12455 ( .A1(n11222), .A2(n11221), .ZN(n9987) );
  AND2_X1 U12456 ( .A1(n11254), .A2(n11250), .ZN(n9988) );
  OR2_X1 U12457 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20074), .ZN(n9989) );
  OR2_X1 U12458 ( .A1(n17972), .A2(n11022), .ZN(n9990) );
  OR2_X1 U12459 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17581), .ZN(
        n9991) );
  OR2_X1 U12460 ( .A1(n13315), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9992) );
  OR2_X1 U12461 ( .A1(n13315), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9993) );
  INV_X1 U12462 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10739) );
  AND2_X1 U12463 ( .A1(n10649), .A2(n15369), .ZN(n9994) );
  OR2_X1 U12464 ( .A1(n14781), .A2(n15035), .ZN(n9996) );
  AND3_X1 U12465 ( .A1(n10211), .A2(n10156), .A3(n10210), .ZN(n9997) );
  INV_X1 U12466 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10723) );
  AND2_X1 U12467 ( .A1(n10218), .A2(n10217), .ZN(n9998) );
  INV_X1 U12468 ( .A(n11705), .ZN(n11701) );
  NOR2_X1 U12469 ( .A1(n17699), .A2(n17179), .ZN(n17538) );
  OAI211_X2 U12470 ( .C1(n10797), .C2(n16702), .A(n10842), .B(n10841), .ZN(
        n18702) );
  OR2_X1 U12471 ( .A1(n13315), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9999) );
  AND2_X1 U12472 ( .A1(n13678), .A2(n15778), .ZN(n10000) );
  OAI21_X1 U12473 ( .B1(n15631), .B2(n12841), .A(n14520), .ZN(n12842) );
  AND2_X1 U12474 ( .A1(n11728), .A2(n11761), .ZN(n10001) );
  INV_X1 U12475 ( .A(n15234), .ZN(n16015) );
  INV_X1 U12476 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12864) );
  OR3_X1 U12477 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17422), .ZN(n10002) );
  INV_X1 U12478 ( .A(n10296), .ZN(n10453) );
  AND3_X1 U12479 ( .A1(n10061), .A2(n10060), .A3(n10156), .ZN(n10003) );
  OR2_X1 U12480 ( .A1(n10299), .A2(n13195), .ZN(n10004) );
  INV_X1 U12481 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20507) );
  AND2_X1 U12482 ( .A1(n10509), .A2(n9588), .ZN(n10006) );
  AND3_X1 U12483 ( .A1(n10216), .A2(n10215), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10007) );
  OR2_X1 U12484 ( .A1(n10698), .A2(n18509), .ZN(n10008) );
  OR2_X2 U12485 ( .A1(n16645), .A2(n10695), .ZN(n10009) );
  INV_X1 U12486 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20773) );
  INV_X1 U12487 ( .A(n14022), .ZN(n14051) );
  OR3_X1 U12488 ( .A1(n14149), .A2(n15293), .A3(n14124), .ZN(n10010) );
  OR2_X1 U12489 ( .A1(n15348), .A2(n14144), .ZN(n10011) );
  AND4_X1 U12490 ( .A1(n10221), .A2(n19085), .A3(n10498), .A4(n19060), .ZN(
        n10012) );
  AND2_X1 U12491 ( .A1(n14092), .A2(n14136), .ZN(n10013) );
  AND4_X1 U12492 ( .A1(n11897), .A2(n11896), .A3(n11895), .A4(n11894), .ZN(
        n10014) );
  AND4_X1 U12493 ( .A1(n11903), .A2(n11902), .A3(n11901), .A4(n11900), .ZN(
        n10015) );
  AND4_X1 U12494 ( .A1(n11872), .A2(n11871), .A3(n11870), .A4(n11869), .ZN(
        n10017) );
  INV_X1 U12495 ( .A(n15460), .ZN(n13427) );
  OAI22_X1 U12496 ( .A1(n11189), .A2(n11102), .B1(n19100), .B2(n11101), .ZN(
        n11103) );
  AOI21_X1 U12497 ( .B1(n12714), .B2(n13325), .A(n12695), .ZN(n12706) );
  AND4_X1 U12498 ( .A1(n11133), .A2(n11132), .A3(n11131), .A4(n11130), .ZN(
        n11145) );
  NAND2_X1 U12499 ( .A1(n11138), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11104) );
  OAI21_X1 U12500 ( .B1(n13138), .B2(n12874), .A(n12897), .ZN(n11977) );
  INV_X1 U12501 ( .A(n10515), .ZN(n10516) );
  OR3_X1 U12502 ( .A1(n12684), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n20058), .ZN(n12721) );
  AND3_X1 U12503 ( .A1(n12076), .A2(n12075), .A3(n12074), .ZN(n12082) );
  AOI22_X1 U12504 ( .A1(n12067), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11927), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11887) );
  AND2_X1 U12505 ( .A1(n14711), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10522) );
  INV_X1 U12506 ( .A(n15985), .ZN(n11221) );
  AND2_X1 U12507 ( .A1(n11091), .A2(n11090), .ZN(n11111) );
  NAND2_X1 U12508 ( .A1(n10289), .A2(n10288), .ZN(n10292) );
  NOR2_X1 U12509 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18509), .ZN(
        n10688) );
  INV_X1 U12510 ( .A(n11963), .ZN(n12883) );
  OR2_X1 U12511 ( .A1(n12043), .A2(n12042), .ZN(n12811) );
  INV_X1 U12512 ( .A(n11960), .ZN(n11972) );
  AND2_X1 U12513 ( .A1(n11729), .A2(n10001), .ZN(n11730) );
  AND2_X1 U12514 ( .A1(n10213), .A2(n10212), .ZN(n10214) );
  INV_X1 U12515 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11326) );
  AND2_X1 U12516 ( .A1(n12683), .A2(n12682), .ZN(n12694) );
  INV_X1 U12517 ( .A(n14052), .ZN(n12362) );
  AND2_X1 U12518 ( .A1(n12560), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12561) );
  INV_X1 U12519 ( .A(n13075), .ZN(n12110) );
  NAND2_X1 U12520 ( .A1(n12839), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12840) );
  INV_X1 U12521 ( .A(n13433), .ZN(n12692) );
  NAND2_X1 U12522 ( .A1(n13000), .A2(n20072), .ZN(n11969) );
  NAND2_X1 U12523 ( .A1(n20357), .A2(n20071), .ZN(n12132) );
  OR2_X1 U12524 ( .A1(n10171), .A2(n10170), .ZN(n10321) );
  AND2_X1 U12525 ( .A1(n11540), .A2(n18895), .ZN(n11541) );
  INV_X1 U12526 ( .A(n10309), .ZN(n14116) );
  NAND2_X1 U12527 ( .A1(n14775), .A2(n14761), .ZN(n14745) );
  INV_X1 U12528 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11312) );
  OR2_X1 U12529 ( .A1(n10126), .A2(n10125), .ZN(n11112) );
  NOR3_X1 U12530 ( .A1(n18661), .A2(n18671), .A3(n18509), .ZN(n10726) );
  INV_X2 U12531 ( .A(n10745), .ZN(n16962) );
  INV_X1 U12532 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10916) );
  AND2_X1 U12533 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n10769), .ZN(
        n10770) );
  INV_X1 U12534 ( .A(n12973), .ZN(n12992) );
  AND2_X1 U12535 ( .A1(n14442), .A2(n14440), .ZN(n12468) );
  OR2_X1 U12536 ( .A1(n12607), .A2(n14271), .ZN(n12663) );
  INV_X1 U12537 ( .A(n12661), .ZN(n12626) );
  INV_X1 U12538 ( .A(n12214), .ZN(n12240) );
  NAND2_X1 U12539 ( .A1(n12823), .A2(n12822), .ZN(n13989) );
  INV_X1 U12540 ( .A(n13080), .ZN(n12913) );
  NAND2_X1 U12541 ( .A1(n12118), .A2(n12117), .ZN(n20234) );
  INV_X1 U12542 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13942) );
  INV_X2 U12543 ( .A(n10584), .ZN(n14110) );
  INV_X1 U12544 ( .A(n11763), .ZN(n11764) );
  INV_X1 U12545 ( .A(n15893), .ZN(n11574) );
  OR2_X1 U12546 ( .A1(n10194), .A2(n10193), .ZN(n11205) );
  AND4_X1 U12547 ( .A1(n15307), .A2(n15284), .A3(n15321), .A4(n15289), .ZN(
        n11242) );
  INV_X1 U12548 ( .A(n15226), .ZN(n15330) );
  NAND2_X1 U12549 ( .A1(n11454), .A2(n11453), .ZN(n13854) );
  AND3_X1 U12550 ( .A1(n11418), .A2(n11417), .A3(n11416), .ZN(n15373) );
  OR2_X1 U12551 ( .A1(n9593), .A2(n11519), .ZN(n11042) );
  NAND2_X1 U12552 ( .A1(n16266), .A2(n18700), .ZN(n15431) );
  NOR2_X1 U12553 ( .A1(n17329), .A2(n16085), .ZN(n17331) );
  NOR2_X1 U12554 ( .A1(n17531), .A2(n17493), .ZN(n17489) );
  NOR2_X1 U12555 ( .A1(n18564), .A2(n17601), .ZN(n17445) );
  NOR2_X1 U12556 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17557), .ZN(
        n17470) );
  OR2_X1 U12557 ( .A1(n17557), .A2(n9991), .ZN(n10905) );
  AOI21_X1 U12558 ( .B1(n10972), .B2(n10971), .A(n10982), .ZN(n10975) );
  NAND2_X1 U12559 ( .A1(n10895), .A2(n10894), .ZN(n10896) );
  INV_X1 U12560 ( .A(n12465), .ZN(n12412) );
  NAND2_X1 U12561 ( .A1(n12240), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12246) );
  OR2_X1 U12562 ( .A1(n13062), .A2(n13054), .ZN(n19897) );
  INV_X1 U12563 ( .A(n20784), .ZN(n13044) );
  NAND2_X1 U12564 ( .A1(n13073), .A2(n12112), .ZN(n13535) );
  NAND2_X1 U12565 ( .A1(n12516), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12559) );
  NOR2_X1 U12566 ( .A1(n12246), .A2(n12245), .ZN(n12262) );
  INV_X1 U12567 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n19895) );
  OR2_X1 U12568 ( .A1(n19990), .A2(n12856), .ZN(n14592) );
  NAND2_X1 U12569 ( .A1(n15675), .A2(n12796), .ZN(n15669) );
  INV_X1 U12570 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20429) );
  OR2_X1 U12571 ( .A1(n20059), .A2(n12134), .ZN(n20272) );
  INV_X1 U12572 ( .A(n12758), .ZN(n20061) );
  OR2_X1 U12573 ( .A1(n9569), .A2(n12758), .ZN(n20402) );
  NAND3_X1 U12574 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20071), .A3(n20070), 
        .ZN(n20110) );
  NAND2_X1 U12575 ( .A1(n10514), .A2(n16045), .ZN(n11364) );
  NAND2_X1 U12576 ( .A1(n9565), .A2(n16045), .ZN(n10555) );
  XNOR2_X1 U12577 ( .A(n15363), .B(n11523), .ZN(n13131) );
  AND2_X1 U12578 ( .A1(n11375), .A2(n10267), .ZN(n11383) );
  NAND2_X1 U12579 ( .A1(n10504), .A2(n10503), .ZN(n11352) );
  OR2_X1 U12580 ( .A1(n11495), .A2(n11444), .ZN(n15348) );
  AND2_X1 U12581 ( .A1(n15223), .A2(n15221), .ZN(n15225) );
  INV_X1 U12582 ( .A(n19335), .ZN(n19388) );
  AND2_X1 U12583 ( .A1(n19609), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19086) );
  CLKBUF_X3 U12584 ( .A(n16268), .Z(n16617) );
  NOR2_X1 U12585 ( .A1(n18046), .A2(n15431), .ZN(n15432) );
  AOI211_X1 U12586 ( .C1(n16965), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n10870), .B(n10869), .ZN(n10871) );
  INV_X1 U12587 ( .A(n16093), .ZN(n16094) );
  INV_X1 U12588 ( .A(n17366), .ZN(n17370) );
  NAND2_X1 U12589 ( .A1(n17829), .A2(n10902), .ZN(n17523) );
  AOI21_X1 U12590 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17445), .A(
        n18434), .ZN(n17527) );
  XNOR2_X1 U12591 ( .A(n10737), .B(n10723), .ZN(n17675) );
  INV_X1 U12592 ( .A(n15451), .ZN(n17702) );
  NAND2_X1 U12593 ( .A1(n10909), .A2(n10002), .ZN(n10910) );
  NOR2_X1 U12594 ( .A1(n18506), .A2(n18524), .ZN(n17994) );
  NOR2_X1 U12595 ( .A1(n17183), .A2(n10796), .ZN(n16141) );
  NOR2_X1 U12596 ( .A1(n17638), .A2(n17637), .ZN(n17636) );
  INV_X1 U12597 ( .A(n12900), .ZN(n14243) );
  OR2_X1 U12598 ( .A1(n13139), .A2(n19815), .ZN(n13125) );
  NAND2_X1 U12599 ( .A1(n12449), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12448) );
  AND2_X1 U12600 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n12412), .ZN(
        n12449) );
  AND2_X1 U12601 ( .A1(n15531), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19866) );
  AND2_X1 U12602 ( .A1(n15531), .A2(n13052), .ZN(n19907) );
  NAND2_X1 U12603 ( .A1(n13044), .A2(n13043), .ZN(n15531) );
  INV_X1 U12604 ( .A(n14247), .ZN(n14227) );
  INV_X1 U12605 ( .A(n14401), .ZN(n19913) );
  INV_X1 U12606 ( .A(n13331), .ZN(n19966) );
  NAND2_X1 U12607 ( .A1(n12413), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12514) );
  AOI21_X1 U12608 ( .B1(n14003), .B2(n14002), .A(n14001), .ZN(n15641) );
  INV_X1 U12609 ( .A(n14592), .ZN(n19984) );
  AND2_X1 U12610 ( .A1(n14592), .A2(n12859), .ZN(n15647) );
  NAND2_X1 U12611 ( .A1(n14208), .A2(n14207), .ZN(n14209) );
  AND2_X1 U12612 ( .A1(n15683), .A2(n13027), .ZN(n14651) );
  NOR2_X1 U12613 ( .A1(n15784), .A2(n13024), .ZN(n15702) );
  INV_X1 U12614 ( .A(n20050), .ZN(n20036) );
  NAND2_X1 U12615 ( .A1(n20071), .A2(n20070), .ZN(n20242) );
  INV_X1 U12616 ( .A(n14696), .ZN(n20758) );
  INV_X1 U12617 ( .A(n20187), .ZN(n20152) );
  AND2_X1 U12618 ( .A1(n20060), .A2(n20059), .ZN(n20207) );
  INV_X1 U12619 ( .A(n20228), .ZN(n20223) );
  AND2_X1 U12620 ( .A1(n20207), .A2(n20334), .ZN(n20261) );
  INV_X1 U12621 ( .A(n20295), .ZN(n20287) );
  INV_X1 U12622 ( .A(n20317), .ZN(n20319) );
  INV_X1 U12623 ( .A(n20422), .ZN(n20386) );
  INV_X1 U12624 ( .A(n20272), .ZN(n20335) );
  INV_X1 U12625 ( .A(n20437), .ZN(n20462) );
  INV_X1 U12626 ( .A(n20496), .ZN(n20500) );
  OAI22_X1 U12627 ( .A1(n20517), .A2(n20516), .B1(n20574), .B2(n20515), .ZN(
        n20533) );
  INV_X1 U12628 ( .A(n20365), .ZN(n20505) );
  INV_X1 U12629 ( .A(n20402), .ZN(n20546) );
  INV_X1 U12630 ( .A(n20684), .ZN(n20670) );
  INV_X1 U12631 ( .A(n20465), .ZN(n20678) );
  INV_X1 U12632 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n13584) );
  NOR2_X1 U12633 ( .A1(n14919), .A2(n18856), .ZN(n10683) );
  NAND2_X1 U12634 ( .A1(n14720), .A2(n14942), .ZN(n14719) );
  NAND2_X1 U12635 ( .A1(n15875), .A2(n15876), .ZN(n15874) );
  INV_X1 U12636 ( .A(n9567), .ZN(n18849) );
  INV_X1 U12637 ( .A(n18821), .ZN(n18879) );
  NAND2_X1 U12638 ( .A1(n11515), .A2(n11527), .ZN(n13302) );
  NOR2_X1 U12639 ( .A1(n15363), .A2(n13194), .ZN(n19334) );
  INV_X2 U12640 ( .A(n10514), .ZN(n19054) );
  AND2_X1 U12641 ( .A1(n13819), .A2(n13818), .ZN(n20957) );
  OR2_X1 U12642 ( .A1(n15319), .A2(n15265), .ZN(n15283) );
  NAND2_X1 U12643 ( .A1(n15320), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15319) );
  OAI21_X1 U12644 ( .B1(n15400), .B2(n15403), .A(n15399), .ZN(n19091) );
  INV_X1 U12645 ( .A(n19126), .ZN(n19116) );
  OR2_X1 U12646 ( .A1(n19134), .A2(n19549), .ZN(n19153) );
  OAI21_X1 U12647 ( .B1(n19208), .B2(n19207), .A(n19206), .ZN(n19231) );
  AND2_X1 U12648 ( .A1(n19236), .A2(n19759), .ZN(n19240) );
  AND2_X1 U12649 ( .A1(n19761), .A2(n19792), .ZN(n19274) );
  OR3_X1 U12650 ( .A1(n19281), .A2(n19549), .A3(n19280), .ZN(n19299) );
  INV_X1 U12651 ( .A(n19327), .ZN(n19330) );
  OAI21_X1 U12652 ( .B1(n19344), .B2(n19341), .A(n19609), .ZN(n19374) );
  INV_X1 U12653 ( .A(n19393), .ZN(n19413) );
  AND2_X1 U12654 ( .A1(n19770), .A2(n15396), .ZN(n19335) );
  INV_X1 U12655 ( .A(n19477), .ZN(n19466) );
  OAI21_X1 U12656 ( .B1(n19487), .B2(n19486), .A(n19485), .ZN(n19505) );
  AND2_X1 U12657 ( .A1(n19512), .A2(n19510), .ZN(n19538) );
  OAI21_X1 U12658 ( .B1(n19555), .B2(n19554), .A(n19553), .ZN(n19594) );
  INV_X1 U12659 ( .A(n19609), .ZN(n19549) );
  INV_X1 U12660 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n16078) );
  NAND2_X1 U12661 ( .A1(n18040), .A2(n18702), .ZN(n10958) );
  NOR2_X1 U12662 ( .A1(n18513), .A2(n16265), .ZN(n18487) );
  OR2_X1 U12663 ( .A1(n16320), .A2(P3_EBX_REG_28__SCAN_IN), .ZN(n16321) );
  NOR2_X1 U12664 ( .A1(n16296), .A2(n16358), .ZN(n16335) );
  NOR2_X1 U12665 ( .A1(n16294), .A2(n16470), .ZN(n16424) );
  NOR2_X1 U12666 ( .A1(n16646), .A2(n16293), .ZN(n16471) );
  INV_X1 U12667 ( .A(n16653), .ZN(n16600) );
  NAND2_X1 U12668 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17074), .ZN(n17073) );
  NAND2_X1 U12669 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17087), .ZN(n17086) );
  INV_X1 U12670 ( .A(n17120), .ZN(n17116) );
  NOR2_X1 U12671 ( .A1(n17206), .A2(n17145), .ZN(n17171) );
  INV_X1 U12672 ( .A(n17190), .ZN(n17204) );
  OAI211_X1 U12673 ( .C1(n16096), .C2(n17700), .A(n16095), .B(n16094), .ZN(
        n16097) );
  NOR2_X1 U12674 ( .A1(n17370), .A2(n17371), .ZN(n17352) );
  NOR2_X1 U12675 ( .A1(n17850), .A2(n17523), .ZN(n17836) );
  NOR2_X2 U12676 ( .A1(n18664), .A2(n17650), .ZN(n17554) );
  INV_X1 U12677 ( .A(n17693), .ZN(n17650) );
  OR2_X1 U12678 ( .A1(n16143), .A2(n16142), .ZN(n16144) );
  OR2_X1 U12679 ( .A1(n16138), .A2(n16137), .ZN(n16146) );
  OR2_X1 U12680 ( .A1(n17356), .A2(n17847), .ZN(n17365) );
  NOR2_X1 U12681 ( .A1(n18023), .A2(n17701), .ZN(n17769) );
  NOR2_X1 U12682 ( .A1(n17882), .A2(n18023), .ZN(n17914) );
  INV_X1 U12683 ( .A(n18007), .ZN(n17982) );
  INV_X1 U12684 ( .A(n18006), .ZN(n18023) );
  NAND2_X1 U12685 ( .A1(n13125), .A2(n13326), .ZN(n20784) );
  INV_X1 U12686 ( .A(n19866), .ZN(n19894) );
  INV_X1 U12687 ( .A(n9561), .ZN(n15586) );
  INV_X1 U12688 ( .A(n19870), .ZN(n15609) );
  INV_X1 U12689 ( .A(n19907), .ZN(n19890) );
  NOR2_X1 U12690 ( .A1(n12747), .A2(n12746), .ZN(n12748) );
  OR2_X1 U12691 ( .A1(n13978), .A2(n13977), .ZN(n15593) );
  INV_X1 U12692 ( .A(n19922), .ZN(n19947) );
  INV_X1 U12693 ( .A(n19974), .ZN(n13466) );
  OAI21_X1 U12694 ( .B1(n13978), .B2(n13971), .A(n14002), .ZN(n14586) );
  INV_X1 U12695 ( .A(n15647), .ZN(n19995) );
  INV_X1 U12696 ( .A(n13319), .ZN(n20067) );
  NAND2_X1 U12697 ( .A1(n15744), .A2(n15785), .ZN(n15784) );
  NAND2_X1 U12698 ( .A1(n20207), .A2(n20505), .ZN(n20142) );
  NAND2_X1 U12699 ( .A1(n20207), .A2(n20546), .ZN(n20187) );
  NAND2_X1 U12700 ( .A1(n20335), .A2(n20505), .ZN(n20295) );
  NAND2_X1 U12701 ( .A1(n20335), .A2(n20546), .ZN(n20317) );
  NAND2_X1 U12702 ( .A1(n20335), .A2(n20577), .ZN(n20348) );
  NAND2_X1 U12703 ( .A1(n20335), .A2(n20334), .ZN(n20390) );
  OR2_X1 U12704 ( .A1(n20480), .A2(n20365), .ZN(n20422) );
  OR2_X1 U12705 ( .A1(n20480), .A2(n20423), .ZN(n20496) );
  OR2_X1 U12706 ( .A1(n20480), .A2(n20479), .ZN(n20537) );
  OR2_X1 U12707 ( .A1(n13097), .A2(n16076), .ZN(n18725) );
  NOR2_X1 U12708 ( .A1(n10684), .A2(n10683), .ZN(n10685) );
  OR2_X1 U12709 ( .A1(n18725), .A2(n10270), .ZN(n18871) );
  OR2_X1 U12710 ( .A1(n18725), .A2(n10481), .ZN(n18858) );
  XNOR2_X1 U12711 ( .A(n13302), .B(n13301), .ZN(n19770) );
  AND2_X1 U12712 ( .A1(n11823), .A2(n13133), .ZN(n18956) );
  INV_X1 U12713 ( .A(n18958), .ZN(n18990) );
  NAND2_X1 U12714 ( .A1(n13103), .A2(n19682), .ZN(n19028) );
  AOI21_X1 U12715 ( .B1(n14161), .B2(n13164), .A(n14160), .ZN(n14162) );
  INV_X1 U12716 ( .A(n19037), .ZN(n15997) );
  INV_X1 U12717 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19046) );
  OR2_X1 U12718 ( .A1(n11495), .A2(n11439), .ZN(n15343) );
  INV_X1 U12719 ( .A(n19147), .ZN(n19156) );
  NAND2_X1 U12720 ( .A1(n19274), .A2(n19757), .ZN(n19194) );
  OR2_X1 U12721 ( .A1(n19310), .A2(n19452), .ZN(n19235) );
  NAND2_X1 U12722 ( .A1(n19274), .A2(n19195), .ZN(n19273) );
  OR2_X1 U12723 ( .A1(n19310), .A2(n19515), .ZN(n19302) );
  AND2_X1 U12724 ( .A1(n19306), .A2(n19305), .ZN(n19327) );
  OR2_X1 U12725 ( .A1(n19310), .A2(n19762), .ZN(n19377) );
  AND2_X1 U12726 ( .A1(n19382), .A2(n19381), .ZN(n19393) );
  NAND2_X1 U12727 ( .A1(n19543), .A2(n19335), .ZN(n19416) );
  INV_X1 U12728 ( .A(n19436), .ZN(n19444) );
  NAND2_X1 U12729 ( .A1(n19543), .A2(n19757), .ZN(n19477) );
  NAND2_X1 U12730 ( .A1(n19445), .A2(n19757), .ZN(n19508) );
  INV_X1 U12731 ( .A(n19504), .ZN(n19542) );
  NAND2_X1 U12732 ( .A1(n19445), .A2(n19604), .ZN(n19640) );
  NAND2_X1 U12733 ( .A1(n19543), .A2(n19604), .ZN(n19663) );
  NAND2_X1 U12734 ( .A1(n18700), .A2(n18545), .ZN(n16248) );
  NAND2_X1 U12735 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n16471), .ZN(n16470) );
  NAND2_X1 U12736 ( .A1(n16657), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n16607) );
  NOR2_X1 U12737 ( .A1(n16667), .A2(n16666), .ZN(n16770) );
  INV_X1 U12738 ( .A(n10792), .ZN(n17183) );
  AND2_X1 U12739 ( .A1(n15513), .A2(P3_EAX_REG_0__SCAN_IN), .ZN(n17207) );
  INV_X1 U12740 ( .A(n17231), .ZN(n17236) );
  NAND2_X1 U12741 ( .A1(n17268), .A2(n14062), .ZN(n17266) );
  INV_X1 U12742 ( .A(n17320), .ZN(n17315) );
  INV_X1 U12743 ( .A(n17608), .ZN(n17568) );
  OAI21_X1 U12744 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18699), .A(n16248), 
        .ZN(n17696) );
  INV_X1 U12745 ( .A(n17685), .ZN(n17700) );
  INV_X1 U12746 ( .A(n17878), .ZN(n17939) );
  INV_X1 U12747 ( .A(n18020), .ZN(n18015) );
  INV_X1 U12748 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n20898) );
  OAI21_X1 U12749 ( .B1(n14076), .B2(n19822), .A(n12863), .ZN(P1_U2971) );
  INV_X1 U12750 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15983) );
  INV_X1 U12751 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18820) );
  INV_X1 U12752 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15953) );
  INV_X1 U12753 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15933) );
  INV_X1 U12754 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15067) );
  INV_X1 U12755 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15043) );
  INV_X1 U12756 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14760) );
  AND2_X2 U12757 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n10018), .ZN(
        n10047) );
  INV_X1 U12758 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14972) );
  NAND2_X1 U12759 ( .A1(n10048), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10051) );
  INV_X1 U12760 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15831) );
  OR2_X2 U12761 ( .A1(n10051), .A2(n15831), .ZN(n10053) );
  INV_X1 U12762 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10052) );
  INV_X1 U12763 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14925) );
  XNOR2_X1 U12764 ( .A(n10055), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14915) );
  INV_X1 U12765 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14124) );
  INV_X1 U12766 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10019) );
  AOI21_X1 U12767 ( .B1(n14972), .B2(n10046), .A(n10048), .ZN(n14974) );
  INV_X1 U12768 ( .A(n14974), .ZN(n15863) );
  OAI21_X1 U12769 ( .B1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n9607), .A(
        n9708), .ZN(n15019) );
  OAI21_X1 U12770 ( .B1(n10038), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n10042), .ZN(n15062) );
  INV_X1 U12771 ( .A(n15062), .ZN(n18764) );
  OAI21_X1 U12772 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n9634), .A(
        n10039), .ZN(n15925) );
  INV_X1 U12773 ( .A(n15925), .ZN(n10037) );
  OAI21_X1 U12774 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n10033), .A(
        n10036), .ZN(n15946) );
  INV_X1 U12775 ( .A(n15946), .ZN(n10035) );
  OAI21_X1 U12776 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n10030), .A(
        n10034), .ZN(n18813) );
  INV_X1 U12777 ( .A(n18813), .ZN(n10032) );
  OAI21_X1 U12778 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n9635), .A(
        n10031), .ZN(n15973) );
  INV_X1 U12779 ( .A(n15973), .ZN(n10029) );
  OAI21_X1 U12780 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n10020), .A(
        n10028), .ZN(n15996) );
  INV_X1 U12781 ( .A(n15996), .ZN(n10027) );
  AOI21_X1 U12782 ( .B1(n13942), .B2(n10023), .A(n10026), .ZN(n13944) );
  AOI21_X1 U12783 ( .B1(n19046), .B2(n10021), .A(n10024), .ZN(n19036) );
  INV_X1 U12784 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13734) );
  AOI21_X1 U12785 ( .B1(n13187), .B2(n13734), .A(n10022), .ZN(n13731) );
  AOI22_X1 U12786 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16078), .ZN(n15354) );
  AOI22_X1 U12787 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n13187), .B2(n16078), .ZN(
        n13848) );
  NAND2_X1 U12788 ( .A1(n15354), .A2(n13848), .ZN(n13847) );
  NOR2_X1 U12789 ( .A1(n13731), .A2(n13847), .ZN(n13686) );
  OAI21_X1 U12790 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n10022), .A(
        n10021), .ZN(n13687) );
  NAND2_X1 U12791 ( .A1(n13686), .A2(n13687), .ZN(n14188) );
  NOR2_X1 U12792 ( .A1(n19036), .A2(n14188), .ZN(n13703) );
  OAI21_X1 U12793 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n10024), .A(
        n10023), .ZN(n13868) );
  NAND2_X1 U12794 ( .A1(n13703), .A2(n13868), .ZN(n13745) );
  NOR2_X1 U12795 ( .A1(n13944), .A2(n13745), .ZN(n18848) );
  OAI21_X1 U12796 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n10026), .A(
        n10025), .ZN(n18851) );
  NAND2_X1 U12797 ( .A1(n18848), .A2(n18851), .ZN(n13766) );
  NOR2_X1 U12798 ( .A1(n10027), .A2(n13766), .ZN(n18836) );
  AOI21_X1 U12799 ( .B1(n15983), .B2(n10028), .A(n9635), .ZN(n15974) );
  INV_X1 U12800 ( .A(n15974), .ZN(n18837) );
  NAND2_X1 U12801 ( .A1(n18836), .A2(n18837), .ZN(n13782) );
  NOR2_X1 U12802 ( .A1(n10029), .A2(n13782), .ZN(n18831) );
  AOI21_X1 U12803 ( .B1(n18820), .B2(n10031), .A(n10030), .ZN(n15961) );
  INV_X1 U12804 ( .A(n15961), .ZN(n18834) );
  NAND2_X1 U12805 ( .A1(n18831), .A2(n18834), .ZN(n18829) );
  NOR2_X1 U12806 ( .A1(n10032), .A2(n18829), .ZN(n13815) );
  AOI21_X1 U12807 ( .B1(n15953), .B2(n10034), .A(n10033), .ZN(n15947) );
  INV_X1 U12808 ( .A(n15947), .ZN(n13829) );
  NAND2_X1 U12809 ( .A1(n13815), .A2(n13829), .ZN(n13814) );
  NOR2_X1 U12810 ( .A1(n10035), .A2(n13814), .ZN(n18797) );
  AOI21_X1 U12811 ( .B1(n15933), .B2(n10036), .A(n9634), .ZN(n15926) );
  INV_X1 U12812 ( .A(n15926), .ZN(n18798) );
  NAND2_X1 U12813 ( .A1(n18797), .A2(n18798), .ZN(n13922) );
  NOR2_X1 U12814 ( .A1(n10037), .A2(n13922), .ZN(n18778) );
  AOI21_X1 U12815 ( .B1(n15067), .B2(n10039), .A(n10038), .ZN(n10040) );
  INV_X1 U12816 ( .A(n10040), .ZN(n18796) );
  NAND2_X1 U12817 ( .A1(n18778), .A2(n18796), .ZN(n18777) );
  NOR2_X1 U12818 ( .A1(n18764), .A2(n18777), .ZN(n18750) );
  AOI21_X1 U12819 ( .B1(n15043), .B2(n10042), .A(n10041), .ZN(n15045) );
  INV_X1 U12820 ( .A(n15045), .ZN(n18752) );
  NAND2_X1 U12821 ( .A1(n18750), .A2(n18752), .ZN(n14781) );
  INV_X1 U12822 ( .A(n10041), .ZN(n10043) );
  AOI21_X1 U12823 ( .B1(n10043), .B2(n9707), .A(n9607), .ZN(n15035) );
  OAI21_X1 U12824 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n10044), .A(
        n10045), .ZN(n15915) );
  INV_X1 U12825 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14994) );
  AOI21_X1 U12826 ( .B1(n14994), .B2(n10045), .A(n10047), .ZN(n14996) );
  INV_X1 U12827 ( .A(n14996), .ZN(n14734) );
  NAND2_X1 U12828 ( .A1(n13685), .A2(n14732), .ZN(n15875) );
  OAI21_X1 U12829 ( .B1(n10047), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n10046), .ZN(n15876) );
  NAND2_X1 U12830 ( .A1(n9567), .A2(n15874), .ZN(n15862) );
  NAND2_X1 U12831 ( .A1(n15863), .A2(n15862), .ZN(n15861) );
  NAND2_X1 U12832 ( .A1(n15861), .A2(n9567), .ZN(n15851) );
  OR2_X1 U12833 ( .A1(n10048), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10049) );
  NAND2_X1 U12834 ( .A1(n10051), .A2(n10049), .ZN(n15852) );
  NAND2_X1 U12835 ( .A1(n13685), .A2(n15850), .ZN(n15838) );
  INV_X1 U12836 ( .A(n10053), .ZN(n10050) );
  AOI21_X1 U12837 ( .B1(n15831), .B2(n10051), .A(n10050), .ZN(n14955) );
  INV_X1 U12838 ( .A(n14955), .ZN(n15839) );
  NAND2_X1 U12839 ( .A1(n13685), .A2(n15837), .ZN(n14720) );
  NAND2_X1 U12840 ( .A1(n10053), .A2(n10052), .ZN(n10054) );
  NAND2_X1 U12841 ( .A1(n9649), .A2(n10054), .ZN(n14942) );
  AOI21_X1 U12842 ( .B1(n14925), .B2(n9649), .A(n10055), .ZN(n14927) );
  INV_X1 U12843 ( .A(n14927), .ZN(n15826) );
  NAND2_X1 U12844 ( .A1(n14915), .A2(n10056), .ZN(n15819) );
  INV_X1 U12845 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19665) );
  INV_X1 U12846 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19544) );
  NAND4_X1 U12847 ( .A1(n16078), .A2(n19665), .A3(n19544), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n18863) );
  INV_X1 U12848 ( .A(n18863), .ZN(n19673) );
  NAND2_X1 U12849 ( .A1(n15819), .A2(n10057), .ZN(n10686) );
  AOI22_X1 U12850 ( .A1(n10253), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10061) );
  AOI22_X1 U12851 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(n9564), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10060) );
  NAND2_X2 U12852 ( .A1(n13355), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10108) );
  INV_X2 U12853 ( .A(n10102), .ZN(n10246) );
  AOI22_X1 U12854 ( .A1(n11616), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10246), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10064) );
  AND2_X4 U12855 ( .A1(n10092), .A2(n15369), .ZN(n11810) );
  AOI22_X1 U12856 ( .A1(n11810), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11740), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10063) );
  NAND2_X1 U12857 ( .A1(n10003), .A2(n10065), .ZN(n10071) );
  AOI22_X1 U12858 ( .A1(n10253), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10067) );
  AOI22_X1 U12859 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(n9564), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10066) );
  AND3_X1 U12860 ( .A1(n10067), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10066), .ZN(n10070) );
  AOI22_X1 U12861 ( .A1(n9568), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10069) );
  AOI22_X1 U12862 ( .A1(n11659), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10246), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10068) );
  INV_X2 U12863 ( .A(n10108), .ZN(n11616) );
  AOI22_X1 U12864 ( .A1(n11616), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10246), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10076) );
  AOI22_X1 U12865 ( .A1(n10253), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10075) );
  AOI22_X1 U12866 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(n9564), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10074) );
  AOI22_X1 U12867 ( .A1(n11810), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11787), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10073) );
  AOI22_X1 U12868 ( .A1(n10253), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11631), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10079) );
  AOI22_X1 U12869 ( .A1(n11810), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11740), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10081) );
  AOI22_X1 U12870 ( .A1(n11616), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10246), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10080) );
  MUX2_X1 U12871 ( .A(n19788), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n11359) );
  NAND2_X1 U12872 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19797), .ZN(
        n11160) );
  INV_X1 U12873 ( .A(n11160), .ZN(n10082) );
  NAND2_X1 U12874 ( .A1(n11359), .A2(n10082), .ZN(n10084) );
  NAND2_X1 U12875 ( .A1(n19788), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10083) );
  NAND2_X1 U12876 ( .A1(n10084), .A2(n10083), .ZN(n10139) );
  XNOR2_X1 U12877 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10138) );
  INV_X1 U12878 ( .A(n10138), .ZN(n10085) );
  XNOR2_X1 U12879 ( .A(n10139), .B(n10085), .ZN(n11356) );
  AND2_X1 U12880 ( .A1(n11399), .A2(n11356), .ZN(n11366) );
  INV_X1 U12881 ( .A(n11366), .ZN(n10101) );
  AOI22_X1 U12882 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n11547), .B1(
        n10279), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10089) );
  AND2_X2 U12883 ( .A1(n11809), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10165) );
  AOI22_X1 U12884 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10280), .B1(
        n10165), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10088) );
  AND2_X2 U12885 ( .A1(n9564), .A2(n10156), .ZN(n11640) );
  AND2_X2 U12886 ( .A1(n9564), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10369) );
  AOI22_X1 U12887 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n11640), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10087) );
  AOI22_X1 U12888 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10274), .B1(
        n10145), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10086) );
  NAND4_X1 U12889 ( .A1(n10089), .A2(n10088), .A3(n10087), .A4(n10086), .ZN(
        n10099) );
  NAND2_X1 U12890 ( .A1(n10273), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10091) );
  INV_X1 U12891 ( .A(n9573), .ZN(n11712) );
  AND2_X2 U12892 ( .A1(n9573), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10272) );
  NAND2_X1 U12893 ( .A1(n10272), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10090) );
  AND2_X1 U12894 ( .A1(n10091), .A2(n10090), .ZN(n10097) );
  AOI22_X1 U12895 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10271), .B1(
        n10172), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10096) );
  AND2_X4 U12896 ( .A1(n11622), .A2(n10156), .ZN(n11637) );
  AOI22_X1 U12897 ( .A1(n11637), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10095) );
  INV_X1 U12898 ( .A(n10092), .ZN(n10093) );
  NOR2_X1 U12899 ( .A1(n10093), .A2(n10156), .ZN(n13356) );
  AND2_X2 U12900 ( .A1(n13356), .A2(n15369), .ZN(n11639) );
  AOI22_X1 U12901 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n11638), .ZN(n10094) );
  NAND4_X1 U12902 ( .A1(n10097), .A2(n10096), .A3(n10095), .A4(n10094), .ZN(
        n10098) );
  NAND2_X1 U12903 ( .A1(n19800), .A2(n11114), .ZN(n10100) );
  NAND2_X1 U12904 ( .A1(n10101), .A2(n10100), .ZN(n11339) );
  INV_X1 U12905 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13735) );
  AOI22_X1 U12906 ( .A1(n11616), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10246), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10106) );
  AOI22_X1 U12907 ( .A1(n10253), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10105) );
  AOI22_X1 U12908 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(n9564), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10104) );
  AOI22_X1 U12909 ( .A1(n11810), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11787), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10103) );
  NAND4_X1 U12910 ( .A1(n10106), .A2(n10105), .A3(n10104), .A4(n10103), .ZN(
        n10107) );
  NAND2_X1 U12911 ( .A1(n10107), .A2(n10156), .ZN(n10115) );
  AOI22_X1 U12912 ( .A1(n10253), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10112) );
  AOI22_X1 U12913 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(n9564), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10111) );
  INV_X2 U12914 ( .A(n10108), .ZN(n11659) );
  AOI22_X1 U12915 ( .A1(n11659), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10246), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10110) );
  AOI22_X1 U12916 ( .A1(n11810), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10109) );
  NAND4_X1 U12917 ( .A1(n10112), .A2(n10111), .A3(n10110), .A4(n10109), .ZN(
        n10113) );
  AOI22_X1 U12918 ( .A1(n10272), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11637), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10119) );
  AOI22_X1 U12919 ( .A1(n10274), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10118) );
  AOI22_X1 U12920 ( .A1(n11547), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10279), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10117) );
  AOI22_X1 U12921 ( .A1(n10165), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10280), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10116) );
  NAND4_X1 U12922 ( .A1(n10119), .A2(n10118), .A3(n10117), .A4(n10116), .ZN(
        n10126) );
  AOI22_X1 U12923 ( .A1(n10273), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10124) );
  AOI22_X1 U12924 ( .A1(n11640), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10271), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10123) );
  AOI22_X1 U12925 ( .A1(n10145), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10172), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10122) );
  AOI22_X1 U12926 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10121) );
  NAND4_X1 U12927 ( .A1(n10124), .A2(n10123), .A3(n10122), .A4(n10121), .ZN(
        n10125) );
  NOR2_X1 U12928 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), 
        .ZN(n10127) );
  MUX2_X1 U12929 ( .A(n11112), .B(n10127), .S(n14096), .Z(n11166) );
  NAND2_X1 U12930 ( .A1(n11167), .A2(n11166), .ZN(n11165) );
  AOI22_X1 U12931 ( .A1(n10272), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10273), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10131) );
  AOI22_X1 U12932 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10130) );
  AOI22_X1 U12933 ( .A1(n10145), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10129) );
  AOI22_X1 U12934 ( .A1(n11637), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10172), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10128) );
  NAND4_X1 U12935 ( .A1(n10131), .A2(n10130), .A3(n10129), .A4(n10128), .ZN(
        n10137) );
  AOI22_X1 U12936 ( .A1(n10165), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11547), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10135) );
  AOI22_X1 U12937 ( .A1(n10279), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10280), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10134) );
  AOI22_X1 U12938 ( .A1(n11640), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10133) );
  AOI22_X1 U12939 ( .A1(n10274), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10271), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10132) );
  NAND4_X1 U12940 ( .A1(n10135), .A2(n10134), .A3(n10133), .A4(n10132), .ZN(
        n10136) );
  NAND2_X1 U12941 ( .A1(n10139), .A2(n10138), .ZN(n10141) );
  INV_X1 U12942 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19779) );
  NAND2_X1 U12943 ( .A1(n19779), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10140) );
  NAND2_X1 U12944 ( .A1(n10141), .A2(n10140), .ZN(n10159) );
  XNOR2_X1 U12945 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10158) );
  INV_X1 U12946 ( .A(n10158), .ZN(n10142) );
  XNOR2_X1 U12947 ( .A(n10159), .B(n10142), .ZN(n11369) );
  MUX2_X1 U12948 ( .A(n10311), .B(n11369), .S(n11399), .Z(n11344) );
  INV_X1 U12949 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10143) );
  MUX2_X1 U12950 ( .A(n11344), .B(n10143), .S(n10531), .Z(n10144) );
  INV_X1 U12951 ( .A(n10144), .ZN(n11158) );
  NOR2_X2 U12952 ( .A1(n11165), .A2(n11158), .ZN(n11157) );
  AOI22_X1 U12953 ( .A1(n11637), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10273), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10149) );
  AOI22_X1 U12954 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10148) );
  AOI22_X1 U12955 ( .A1(n10369), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10172), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10147) );
  AOI22_X1 U12956 ( .A1(n10145), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10271), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10146) );
  NAND4_X1 U12957 ( .A1(n10149), .A2(n10148), .A3(n10147), .A4(n10146), .ZN(
        n10155) );
  AOI22_X1 U12958 ( .A1(n11547), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10280), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10153) );
  AOI22_X1 U12959 ( .A1(n10165), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10279), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10152) );
  AOI22_X1 U12960 ( .A1(n10274), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11640), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10151) );
  AOI22_X1 U12961 ( .A1(n10272), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10150) );
  NAND4_X1 U12962 ( .A1(n10153), .A2(n10152), .A3(n10151), .A4(n10150), .ZN(
        n10154) );
  NOR2_X1 U12963 ( .A1(n10156), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10157) );
  AOI21_X1 U12964 ( .B1(n10159), .B2(n10158), .A(n10157), .ZN(n10263) );
  INV_X1 U12965 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15508) );
  NOR2_X1 U12966 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15508), .ZN(
        n10160) );
  NAND2_X1 U12967 ( .A1(n10263), .A2(n10160), .ZN(n11368) );
  MUX2_X1 U12968 ( .A(n10316), .B(n11368), .S(n11399), .Z(n11343) );
  INV_X1 U12969 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n18922) );
  MUX2_X1 U12970 ( .A(n11343), .B(n18922), .S(n14096), .Z(n11171) );
  AND2_X2 U12971 ( .A1(n11157), .A2(n11171), .ZN(n11170) );
  AOI22_X1 U12972 ( .A1(n10272), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11595), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10164) );
  AOI22_X1 U12973 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U12974 ( .A1(n11637), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10162) );
  AOI22_X1 U12975 ( .A1(n11640), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10161) );
  NAND4_X1 U12976 ( .A1(n10164), .A2(n10163), .A3(n10162), .A4(n10161), .ZN(
        n10171) );
  AOI22_X1 U12977 ( .A1(n10165), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10279), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10169) );
  AOI22_X1 U12978 ( .A1(n11547), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10280), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10168) );
  AOI22_X1 U12979 ( .A1(n10145), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10172), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10167) );
  AOI22_X1 U12980 ( .A1(n10274), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10271), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10166) );
  NAND4_X1 U12981 ( .A1(n10169), .A2(n10168), .A3(n10167), .A4(n10166), .ZN(
        n10170) );
  INV_X1 U12982 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n14181) );
  MUX2_X1 U12983 ( .A(n10321), .B(n14181), .S(n14096), .Z(n11152) );
  AOI22_X1 U12984 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n11547), .B1(
        n10279), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10176) );
  AOI22_X1 U12985 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10280), .B1(
        n10165), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10175) );
  AOI22_X1 U12986 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n11640), .B1(
        n10145), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U12987 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10274), .B1(
        n10172), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10173) );
  NAND4_X1 U12988 ( .A1(n10176), .A2(n10175), .A3(n10174), .A4(n10173), .ZN(
        n10184) );
  NAND2_X1 U12989 ( .A1(n10273), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10178) );
  NAND2_X1 U12990 ( .A1(n10272), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10177) );
  AND2_X1 U12991 ( .A1(n10178), .A2(n10177), .ZN(n10182) );
  AOI22_X1 U12992 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n10369), .B1(
        n10271), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10181) );
  AOI22_X1 U12993 ( .A1(n11637), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10180) );
  AOI22_X1 U12994 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n11638), .ZN(n10179) );
  NAND4_X1 U12995 ( .A1(n10182), .A2(n10181), .A3(n10180), .A4(n10179), .ZN(
        n10183) );
  OR2_X2 U12996 ( .A1(n10184), .A2(n10183), .ZN(n14094) );
  INV_X1 U12997 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n10602) );
  MUX2_X1 U12998 ( .A(n14094), .B(n10602), .S(n14096), .Z(n11218) );
  AOI22_X1 U12999 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n11547), .B1(
        n10165), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10188) );
  AOI22_X1 U13000 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10280), .B1(
        n10279), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10187) );
  AOI22_X1 U13001 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n10369), .B1(
        n10271), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10186) );
  AOI22_X1 U13002 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10274), .B1(
        n10172), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10185) );
  NAND4_X1 U13003 ( .A1(n10188), .A2(n10187), .A3(n10186), .A4(n10185), .ZN(
        n10194) );
  AOI22_X1 U13004 ( .A1(n10272), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11640), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10192) );
  AOI22_X1 U13005 ( .A1(n10273), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10145), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10191) );
  AOI22_X1 U13006 ( .A1(n11637), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10190) );
  AOI22_X1 U13007 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n10426), .ZN(n10189) );
  NAND4_X1 U13008 ( .A1(n10192), .A2(n10191), .A3(n10190), .A4(n10189), .ZN(
        n10193) );
  INV_X1 U13009 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n10599) );
  MUX2_X1 U13010 ( .A(n11205), .B(n10599), .S(n14096), .Z(n11209) );
  NAND2_X1 U13011 ( .A1(n14096), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11214) );
  INV_X1 U13012 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13528) );
  NAND2_X1 U13013 ( .A1(n11232), .A2(n13528), .ZN(n11244) );
  NAND2_X1 U13014 ( .A1(n14096), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11243) );
  INV_X1 U13015 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10622) );
  NOR2_X1 U13016 ( .A1(n19070), .A2(n10622), .ZN(n11264) );
  INV_X1 U13017 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n13807) );
  NOR2_X1 U13018 ( .A1(n19070), .A2(n13807), .ZN(n11262) );
  NAND2_X1 U13019 ( .A1(n14096), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11255) );
  INV_X1 U13020 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n18886) );
  NOR2_X1 U13021 ( .A1(n19070), .A2(n18886), .ZN(n11275) );
  INV_X1 U13022 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n18781) );
  NOR2_X1 U13023 ( .A1(n19070), .A2(n18781), .ZN(n11258) );
  OR2_X2 U13024 ( .A1(n11259), .A2(n11258), .ZN(n11261) );
  INV_X1 U13025 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n18767) );
  NOR2_X1 U13026 ( .A1(n19070), .A2(n18767), .ZN(n11252) );
  INV_X1 U13027 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n18754) );
  NOR2_X1 U13028 ( .A1(n19070), .A2(n18754), .ZN(n11250) );
  INV_X1 U13029 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n14771) );
  NAND2_X1 U13030 ( .A1(n14096), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11298) );
  INV_X1 U13031 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10656) );
  NOR2_X1 U13032 ( .A1(n19070), .A2(n10656), .ZN(n11303) );
  INV_X1 U13033 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10660) );
  INV_X1 U13034 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n14821) );
  NAND2_X1 U13035 ( .A1(n14096), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11320) );
  INV_X1 U13036 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n14725) );
  NOR2_X1 U13037 ( .A1(n19070), .A2(n14725), .ZN(n11327) );
  NAND2_X1 U13038 ( .A1(n14096), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11336) );
  INV_X1 U13039 ( .A(n11336), .ZN(n10196) );
  NAND2_X1 U13040 ( .A1(n14096), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10197) );
  XNOR2_X1 U13041 ( .A(n14097), .B(n10197), .ZN(n14095) );
  AOI22_X1 U13042 ( .A1(n9564), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11787), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10201) );
  AOI22_X1 U13043 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(n9568), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10200) );
  AOI22_X1 U13044 ( .A1(n11616), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10246), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10199) );
  AOI22_X1 U13045 ( .A1(n10253), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11631), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10198) );
  NAND2_X1 U13046 ( .A1(n10202), .A2(n10156), .ZN(n10209) );
  AOI22_X1 U13047 ( .A1(n11616), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10246), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10206) );
  AOI22_X1 U13048 ( .A1(n10253), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9564), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10204) );
  AOI22_X1 U13049 ( .A1(n11740), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11631), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10203) );
  NAND2_X1 U13050 ( .A1(n10207), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10208) );
  NAND2_X2 U13051 ( .A1(n10209), .A2(n10208), .ZN(n10221) );
  AOI22_X1 U13052 ( .A1(n10253), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11631), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10211) );
  AOI22_X1 U13053 ( .A1(n11616), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10246), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10210) );
  AOI22_X1 U13054 ( .A1(n11810), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11740), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10213) );
  AOI22_X1 U13055 ( .A1(n9573), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(n9564), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10212) );
  AOI22_X1 U13056 ( .A1(n10253), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11631), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10216) );
  AOI22_X1 U13057 ( .A1(n11616), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10246), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10215) );
  AOI22_X1 U13058 ( .A1(n11810), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10218) );
  AOI22_X1 U13059 ( .A1(n9573), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9564), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10217) );
  NAND2_X1 U13060 ( .A1(n10221), .A2(n10530), .ZN(n10497) );
  AOI22_X1 U13061 ( .A1(n9573), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(n9564), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10225) );
  AOI22_X1 U13062 ( .A1(n11659), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10246), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10224) );
  AOI22_X1 U13063 ( .A1(n10253), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10223) );
  AOI22_X1 U13064 ( .A1(n11810), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10222) );
  NAND4_X1 U13065 ( .A1(n10225), .A2(n10224), .A3(n10223), .A4(n10222), .ZN(
        n10226) );
  AOI22_X1 U13066 ( .A1(n10253), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11631), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10230) );
  AOI22_X1 U13067 ( .A1(n11659), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10246), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10229) );
  AOI22_X1 U13068 ( .A1(n9573), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(n9564), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10228) );
  AOI22_X1 U13069 ( .A1(n11810), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11787), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10227) );
  NAND4_X1 U13070 ( .A1(n10230), .A2(n10229), .A3(n10228), .A4(n10227), .ZN(
        n10231) );
  NAND2_X1 U13071 ( .A1(n10231), .A2(n10156), .ZN(n10232) );
  NAND2_X1 U13072 ( .A1(n10497), .A2(n10513), .ZN(n10245) );
  AOI22_X1 U13073 ( .A1(n11659), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10246), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10237) );
  AOI22_X1 U13074 ( .A1(n10253), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10236) );
  AOI22_X1 U13075 ( .A1(n9573), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(n9564), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10235) );
  AOI22_X1 U13076 ( .A1(n11810), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11787), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10234) );
  NAND4_X1 U13077 ( .A1(n10237), .A2(n10236), .A3(n10235), .A4(n10234), .ZN(
        n10243) );
  AOI22_X1 U13078 ( .A1(n11659), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10246), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10241) );
  AOI22_X1 U13079 ( .A1(n10253), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11631), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10240) );
  AOI22_X1 U13080 ( .A1(n9573), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(n9564), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10239) );
  AOI22_X1 U13081 ( .A1(n9568), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11787), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10238) );
  NAND4_X1 U13082 ( .A1(n10241), .A2(n10240), .A3(n10239), .A4(n10238), .ZN(
        n10242) );
  MUX2_X2 U13083 ( .A(n10243), .B(n10242), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n19065) );
  NAND2_X1 U13084 ( .A1(n10496), .A2(n19065), .ZN(n10244) );
  AOI22_X1 U13085 ( .A1(n9573), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(n9564), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10250) );
  AOI22_X1 U13086 ( .A1(n11659), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10246), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10249) );
  AOI22_X1 U13087 ( .A1(n10253), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11631), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10248) );
  AOI22_X1 U13088 ( .A1(n11810), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11740), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10247) );
  NAND4_X1 U13089 ( .A1(n10250), .A2(n10249), .A3(n10248), .A4(n10247), .ZN(
        n10251) );
  AOI22_X1 U13090 ( .A1(n9573), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(n9564), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10257) );
  AOI22_X1 U13091 ( .A1(n9568), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11787), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10256) );
  AOI22_X1 U13092 ( .A1(n11616), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10246), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10255) );
  AOI22_X1 U13093 ( .A1(n10253), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10254) );
  NAND4_X1 U13094 ( .A1(n10257), .A2(n10256), .A3(n10255), .A4(n10254), .ZN(
        n10258) );
  NAND2_X1 U13095 ( .A1(n10258), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10259) );
  NAND4_X2 U13096 ( .A1(n10221), .A2(n9588), .A3(n19085), .A4(n19065), .ZN(
        n10502) );
  INV_X1 U13097 ( .A(n10498), .ZN(n10261) );
  NAND2_X2 U13098 ( .A1(n10261), .A2(n11503), .ZN(n10515) );
  NAND2_X1 U13099 ( .A1(n10538), .A2(n19048), .ZN(n10552) );
  NAND2_X1 U13100 ( .A1(n16047), .A2(n10552), .ZN(n16036) );
  NAND2_X1 U13101 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15508), .ZN(
        n10262) );
  NAND2_X1 U13102 ( .A1(n10263), .A2(n10262), .ZN(n10265) );
  INV_X1 U13103 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15445) );
  NAND2_X1 U13104 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n15445), .ZN(
        n10264) );
  NAND2_X1 U13105 ( .A1(n10265), .A2(n10264), .ZN(n11375) );
  XNOR2_X1 U13106 ( .A(n11359), .B(n11160), .ZN(n11357) );
  NAND3_X1 U13107 ( .A1(n11369), .A2(n11356), .A3(n11368), .ZN(n11348) );
  INV_X1 U13108 ( .A(n11348), .ZN(n10266) );
  NAND2_X1 U13109 ( .A1(n11357), .A2(n10266), .ZN(n10267) );
  NAND2_X1 U13110 ( .A1(n16036), .A2(n11383), .ZN(n13097) );
  INV_X1 U13111 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n19668) );
  NAND2_X1 U13112 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19668), .ZN(n10482) );
  INV_X1 U13113 ( .A(n10482), .ZN(n10268) );
  NAND2_X1 U13114 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10268), .ZN(n16076) );
  NAND2_X1 U13115 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19669) );
  INV_X1 U13116 ( .A(n19669), .ZN(n19690) );
  NOR2_X1 U13117 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19690), .ZN(n10681) );
  INV_X1 U13118 ( .A(n10681), .ZN(n10269) );
  NAND3_X1 U13119 ( .A1(n19800), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n10269), 
        .ZN(n10270) );
  INV_X1 U13120 ( .A(n18871), .ZN(n18786) );
  AOI22_X1 U13121 ( .A1(n10271), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10172), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10278) );
  AOI22_X1 U13122 ( .A1(n10272), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11639), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10277) );
  AOI22_X1 U13123 ( .A1(n10273), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10276) );
  AOI22_X1 U13124 ( .A1(n10274), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10145), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10275) );
  NAND4_X1 U13125 ( .A1(n10278), .A2(n10277), .A3(n10276), .A4(n10275), .ZN(
        n10286) );
  AOI22_X1 U13126 ( .A1(n10279), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10284) );
  AOI22_X1 U13127 ( .A1(n11547), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10280), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10283) );
  AOI22_X1 U13128 ( .A1(n11637), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10165), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10282) );
  AOI22_X1 U13129 ( .A1(n11640), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10281) );
  NAND4_X1 U13130 ( .A1(n10284), .A2(n10283), .A3(n10282), .A4(n10281), .ZN(
        n10285) );
  INV_X1 U13131 ( .A(n13347), .ZN(n10289) );
  AND2_X1 U13132 ( .A1(n10498), .A2(n19611), .ZN(n10287) );
  MUX2_X1 U13133 ( .A(n19085), .B(n19797), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10290) );
  NAND2_X1 U13134 ( .A1(n10296), .A2(n11824), .ZN(n10302) );
  AND2_X1 U13135 ( .A1(n10290), .A2(n10302), .ZN(n10291) );
  NAND2_X1 U13136 ( .A1(n10292), .A2(n10291), .ZN(n13196) );
  NAND4_X1 U13137 ( .A1(n10531), .A2(n16044), .A3(n19085), .A4(n19611), .ZN(
        n10303) );
  INV_X1 U13138 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18865) );
  INV_X1 U13139 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13351) );
  NAND2_X1 U13140 ( .A1(n9868), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n10293) );
  OAI211_X1 U13141 ( .C1(n16044), .C2(n13351), .A(n10293), .B(n19611), .ZN(
        n10294) );
  INV_X1 U13142 ( .A(n10294), .ZN(n10295) );
  OAI21_X1 U13143 ( .B1(n10303), .B2(n18865), .A(n10295), .ZN(n13197) );
  INV_X1 U13144 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15366) );
  INV_X1 U13145 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19024) );
  INV_X1 U13146 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19699) );
  OAI222_X1 U13147 ( .A1(n10453), .A2(n15366), .B1(n10005), .B2(n19024), .C1(
        n10303), .C2(n19699), .ZN(n10299) );
  XNOR2_X1 U13148 ( .A(n13195), .B(n10299), .ZN(n13306) );
  INV_X1 U13149 ( .A(n11112), .ZN(n11458) );
  NAND2_X1 U13150 ( .A1(n10496), .A2(n19085), .ZN(n10297) );
  MUX2_X1 U13151 ( .A(n10297), .B(n19788), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10298) );
  OAI21_X1 U13152 ( .B1(n11458), .B2(n10439), .A(n10298), .ZN(n13307) );
  OAI21_X1 U13153 ( .B1(n13306), .B2(n13307), .A(n10004), .ZN(n10300) );
  INV_X1 U13154 ( .A(n10300), .ZN(n10307) );
  NAND2_X1 U13155 ( .A1(n10288), .A2(n11114), .ZN(n10301) );
  OAI211_X1 U13156 ( .C1(n19611), .C2(n19779), .A(n10302), .B(n10301), .ZN(
        n10306) );
  XNOR2_X1 U13157 ( .A(n10307), .B(n10306), .ZN(n13391) );
  INV_X1 U13158 ( .A(n10303), .ZN(n10309) );
  INV_X1 U13159 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19701) );
  INV_X2 U13160 ( .A(n10453), .ZN(n10466) );
  NAND2_X1 U13161 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10305) );
  INV_X2 U13162 ( .A(n10005), .ZN(n14113) );
  NAND2_X1 U13163 ( .A1(n14113), .A2(P2_EAX_REG_2__SCAN_IN), .ZN(n10304) );
  OAI211_X1 U13164 ( .C1(n14116), .C2(n19701), .A(n10305), .B(n10304), .ZN(
        n13390) );
  NOR2_X1 U13165 ( .A1(n10307), .A2(n10306), .ZN(n10308) );
  INV_X1 U13166 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n13657) );
  NAND2_X1 U13167 ( .A1(n14113), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n10310) );
  OAI21_X1 U13168 ( .B1(n14116), .B2(n13657), .A(n10310), .ZN(n10315) );
  INV_X1 U13169 ( .A(n10311), .ZN(n11083) );
  NAND2_X1 U13170 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10313) );
  NAND2_X1 U13171 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10312) );
  OAI211_X1 U13172 ( .C1(n11083), .C2(n10439), .A(n10313), .B(n10312), .ZN(
        n10314) );
  INV_X1 U13173 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n10317) );
  INV_X1 U13174 ( .A(n10316), .ZN(n11468) );
  OAI22_X1 U13175 ( .A1(n14116), .A2(n10317), .B1(n10439), .B2(n11468), .ZN(
        n10318) );
  INV_X1 U13176 ( .A(n10318), .ZN(n10320) );
  AOI22_X1 U13177 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n14113), .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n10319) );
  INV_X1 U13178 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n13861) );
  INV_X1 U13179 ( .A(n10321), .ZN(n11148) );
  OAI22_X1 U13180 ( .A1(n14116), .A2(n13861), .B1(n10439), .B2(n11148), .ZN(
        n10322) );
  INV_X1 U13181 ( .A(n10322), .ZN(n10324) );
  AOI22_X1 U13182 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n14113), .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n10323) );
  NAND2_X1 U13183 ( .A1(n10324), .A2(n10323), .ZN(n13702) );
  NAND2_X1 U13184 ( .A1(n13700), .A2(n13702), .ZN(n13701) );
  NAND2_X1 U13185 ( .A1(n10288), .A2(n11205), .ZN(n10325) );
  INV_X1 U13186 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19707) );
  NAND2_X1 U13187 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10327) );
  NAND2_X1 U13188 ( .A1(n14113), .A2(P2_EAX_REG_6__SCAN_IN), .ZN(n10326) );
  OAI211_X1 U13189 ( .C1(n14116), .C2(n19707), .A(n10327), .B(n10326), .ZN(
        n10328) );
  INV_X1 U13190 ( .A(n10328), .ZN(n13743) );
  INV_X1 U13191 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15342) );
  INV_X1 U13192 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19012) );
  INV_X1 U13193 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19709) );
  OAI222_X1 U13194 ( .A1(n15342), .A2(n10453), .B1(n10005), .B2(n19012), .C1(
        n14116), .C2(n19709), .ZN(n15340) );
  INV_X1 U13195 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n10339) );
  AOI22_X1 U13196 ( .A1(n11547), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10280), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10332) );
  AOI22_X1 U13197 ( .A1(n10165), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10279), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10331) );
  AOI22_X1 U13198 ( .A1(n10369), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10145), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10330) );
  AOI22_X1 U13199 ( .A1(n10274), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10172), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10329) );
  NAND4_X1 U13200 ( .A1(n10332), .A2(n10331), .A3(n10330), .A4(n10329), .ZN(
        n10338) );
  AOI22_X1 U13201 ( .A1(n11595), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U13202 ( .A1(n10272), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11640), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10335) );
  AOI22_X1 U13203 ( .A1(n11637), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10271), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10334) );
  AOI22_X1 U13204 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10333) );
  NAND4_X1 U13205 ( .A1(n10336), .A2(n10335), .A3(n10334), .A4(n10333), .ZN(
        n10337) );
  OR2_X1 U13206 ( .A1(n10338), .A2(n10337), .ZN(n11534) );
  INV_X1 U13207 ( .A(n11534), .ZN(n18914) );
  OAI22_X1 U13208 ( .A1(n14116), .A2(n10339), .B1(n10439), .B2(n18914), .ZN(
        n10340) );
  INV_X1 U13209 ( .A(n10340), .ZN(n10342) );
  AOI22_X1 U13210 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n14113), .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n10341) );
  AOI22_X1 U13211 ( .A1(n10272), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11595), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10346) );
  AOI22_X1 U13212 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10345) );
  AOI22_X1 U13213 ( .A1(n11637), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10344) );
  AOI22_X1 U13214 ( .A1(n11640), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10343) );
  NAND4_X1 U13215 ( .A1(n10346), .A2(n10345), .A3(n10344), .A4(n10343), .ZN(
        n10352) );
  AOI22_X1 U13216 ( .A1(n10165), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10279), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10350) );
  AOI22_X1 U13217 ( .A1(n11547), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10280), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10349) );
  AOI22_X1 U13218 ( .A1(n10145), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10172), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10348) );
  AOI22_X1 U13219 ( .A1(n10274), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10271), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10347) );
  NAND4_X1 U13220 ( .A1(n10350), .A2(n10349), .A3(n10348), .A4(n10347), .ZN(
        n10351) );
  NOR2_X1 U13221 ( .A1(n10352), .A2(n10351), .ZN(n11532) );
  AOI22_X1 U13222 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n14113), .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n10354) );
  NAND2_X1 U13223 ( .A1(n10309), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n10353) );
  OAI211_X1 U13224 ( .C1(n11532), .C2(n10439), .A(n10354), .B(n10353), .ZN(
        n15331) );
  INV_X1 U13225 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n10365) );
  AOI22_X1 U13226 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n11637), .B1(
        n11595), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10358) );
  AOI22_X1 U13227 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n10426), .ZN(n10357) );
  AOI22_X1 U13228 ( .A1(n10272), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10356) );
  AOI22_X1 U13229 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10271), .B1(
        n10145), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10355) );
  NAND4_X1 U13230 ( .A1(n10358), .A2(n10357), .A3(n10356), .A4(n10355), .ZN(
        n10364) );
  AOI22_X1 U13231 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n11547), .B1(
        n10279), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10362) );
  AOI22_X1 U13232 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10280), .B1(
        n10165), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10361) );
  AOI22_X1 U13233 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11640), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10360) );
  AOI22_X1 U13234 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n10274), .B1(
        n10172), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10359) );
  NAND4_X1 U13235 ( .A1(n10362), .A2(n10361), .A3(n10360), .A4(n10359), .ZN(
        n10363) );
  NOR2_X1 U13236 ( .A1(n10364), .A2(n10363), .ZN(n18905) );
  OAI22_X1 U13237 ( .A1(n14116), .A2(n10365), .B1(n10439), .B2(n18905), .ZN(
        n10366) );
  INV_X1 U13238 ( .A(n10366), .ZN(n10368) );
  AOI22_X1 U13239 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n14113), .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n10367) );
  AND2_X1 U13240 ( .A1(n10368), .A2(n10367), .ZN(n13789) );
  AOI22_X1 U13241 ( .A1(n10272), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11595), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10377) );
  AOI22_X1 U13242 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10376) );
  AOI22_X1 U13243 ( .A1(n11637), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10375) );
  INV_X1 U13244 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10372) );
  INV_X1 U13245 ( .A(n10369), .ZN(n10371) );
  INV_X1 U13246 ( .A(n11640), .ZN(n10370) );
  INV_X1 U13247 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11062) );
  OAI22_X1 U13248 ( .A1(n10372), .A2(n10371), .B1(n10370), .B2(n11062), .ZN(
        n10373) );
  INV_X1 U13249 ( .A(n10373), .ZN(n10374) );
  NAND4_X1 U13250 ( .A1(n10377), .A2(n10376), .A3(n10375), .A4(n10374), .ZN(
        n10383) );
  AOI22_X1 U13251 ( .A1(n10165), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10279), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10381) );
  AOI22_X1 U13252 ( .A1(n11547), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10280), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10380) );
  AOI22_X1 U13253 ( .A1(n10145), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10172), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10379) );
  AOI22_X1 U13254 ( .A1(n10274), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10271), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10378) );
  NAND4_X1 U13255 ( .A1(n10381), .A2(n10380), .A3(n10379), .A4(n10378), .ZN(
        n10382) );
  OR2_X1 U13256 ( .A1(n10383), .A2(n10382), .ZN(n18897) );
  AOI22_X1 U13257 ( .A1(n10309), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n10288), 
        .B2(n18897), .ZN(n10385) );
  AOI22_X1 U13258 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n14113), .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n10384) );
  NAND2_X1 U13259 ( .A1(n10385), .A2(n10384), .ZN(n15299) );
  INV_X1 U13260 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n10397) );
  AOI22_X1 U13261 ( .A1(n11637), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11595), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10389) );
  AOI22_X1 U13262 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10388) );
  AOI22_X1 U13263 ( .A1(n10272), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10387) );
  AOI22_X1 U13264 ( .A1(n11640), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10386) );
  NAND4_X1 U13265 ( .A1(n10389), .A2(n10388), .A3(n10387), .A4(n10386), .ZN(
        n10395) );
  AOI22_X1 U13266 ( .A1(n10165), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11547), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10393) );
  AOI22_X1 U13267 ( .A1(n10279), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10280), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10392) );
  AOI22_X1 U13268 ( .A1(n10145), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10172), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10391) );
  AOI22_X1 U13269 ( .A1(n10274), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10271), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10390) );
  NAND4_X1 U13270 ( .A1(n10393), .A2(n10392), .A3(n10391), .A4(n10390), .ZN(
        n10394) );
  OR2_X1 U13271 ( .A1(n10395), .A2(n10394), .ZN(n18896) );
  INV_X1 U13272 ( .A(n18896), .ZN(n10396) );
  OAI22_X1 U13273 ( .A1(n14116), .A2(n10397), .B1(n10439), .B2(n10396), .ZN(
        n10398) );
  INV_X1 U13274 ( .A(n10398), .ZN(n10400) );
  AOI22_X1 U13275 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n14113), .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n10399) );
  AND2_X1 U13276 ( .A1(n10400), .A2(n10399), .ZN(n15272) );
  AOI22_X1 U13277 ( .A1(n10272), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11595), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10404) );
  AOI22_X1 U13278 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10403) );
  AOI22_X1 U13279 ( .A1(n11637), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10402) );
  AOI22_X1 U13280 ( .A1(n10369), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10145), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10401) );
  NAND4_X1 U13281 ( .A1(n10404), .A2(n10403), .A3(n10402), .A4(n10401), .ZN(
        n10410) );
  AOI22_X1 U13282 ( .A1(n11547), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10279), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10408) );
  AOI22_X1 U13283 ( .A1(n10165), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10280), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10407) );
  AOI22_X1 U13284 ( .A1(n11640), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10271), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10406) );
  AOI22_X1 U13285 ( .A1(n10274), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10172), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10405) );
  NAND4_X1 U13286 ( .A1(n10408), .A2(n10407), .A3(n10406), .A4(n10405), .ZN(
        n10409) );
  OR2_X1 U13287 ( .A1(n10410), .A2(n10409), .ZN(n11540) );
  INV_X1 U13288 ( .A(n11540), .ZN(n20961) );
  AOI22_X1 U13289 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n14113), .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n10412) );
  NAND2_X1 U13290 ( .A1(n10309), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n10411) );
  OAI211_X1 U13291 ( .C1(n20961), .C2(n10439), .A(n10412), .B(n10411), .ZN(
        n13821) );
  INV_X1 U13292 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n10423) );
  AOI22_X1 U13293 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n11637), .B1(
        n11595), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10416) );
  AOI22_X1 U13294 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n10426), .ZN(n10415) );
  AOI22_X1 U13295 ( .A1(n10272), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10414) );
  AOI22_X1 U13296 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11640), .B1(
        n10271), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10413) );
  NAND4_X1 U13297 ( .A1(n10416), .A2(n10415), .A3(n10414), .A4(n10413), .ZN(
        n10422) );
  AOI22_X1 U13298 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n11547), .B1(
        n10165), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10420) );
  AOI22_X1 U13299 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10280), .B1(
        n10279), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10419) );
  AOI22_X1 U13300 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n10369), .B1(
        n10145), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10418) );
  AOI22_X1 U13301 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n10274), .B1(
        n10172), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10417) );
  NAND4_X1 U13302 ( .A1(n10420), .A2(n10419), .A3(n10418), .A4(n10417), .ZN(
        n10421) );
  OR2_X1 U13303 ( .A1(n10422), .A2(n10421), .ZN(n18890) );
  INV_X1 U13304 ( .A(n18890), .ZN(n14079) );
  OAI22_X1 U13305 ( .A1(n14116), .A2(n10423), .B1(n10439), .B2(n14079), .ZN(
        n10425) );
  INV_X1 U13306 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15935) );
  NOR2_X1 U13307 ( .A1(n10453), .A2(n15935), .ZN(n10424) );
  AOI211_X1 U13308 ( .C1(n14113), .C2(P2_EAX_REG_14__SCAN_IN), .A(n10425), .B(
        n10424), .ZN(n13805) );
  AOI22_X1 U13309 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n10272), .B1(
        n11595), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10430) );
  AOI22_X1 U13310 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n10426), .ZN(n10429) );
  AOI22_X1 U13311 ( .A1(n11637), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10428) );
  AOI22_X1 U13312 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11640), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10427) );
  NAND4_X1 U13313 ( .A1(n10430), .A2(n10429), .A3(n10428), .A4(n10427), .ZN(
        n10436) );
  AOI22_X1 U13314 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n10165), .B1(
        n10279), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10434) );
  AOI22_X1 U13315 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10280), .B1(
        n11547), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10433) );
  AOI22_X1 U13316 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10172), .B1(
        n10145), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10432) );
  AOI22_X1 U13317 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n10274), .B1(
        n10271), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10431) );
  NAND4_X1 U13318 ( .A1(n10434), .A2(n10433), .A3(n10432), .A4(n10431), .ZN(
        n10435) );
  NOR2_X1 U13319 ( .A1(n10436), .A2(n10435), .ZN(n14078) );
  AOI22_X1 U13320 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        n14113), .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n10438) );
  NAND2_X1 U13321 ( .A1(n10309), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n10437) );
  OAI211_X1 U13322 ( .C1(n14078), .C2(n10439), .A(n10438), .B(n10437), .ZN(
        n15255) );
  NAND2_X1 U13323 ( .A1(n13804), .A2(n15255), .ZN(n13927) );
  AOI22_X1 U13324 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n14113), .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n10441) );
  NAND2_X1 U13325 ( .A1(n10309), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n10440) );
  AND2_X1 U13326 ( .A1(n10441), .A2(n10440), .ZN(n13928) );
  INV_X1 U13327 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19721) );
  NAND2_X1 U13328 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10443) );
  NAND2_X1 U13329 ( .A1(n14113), .A2(P2_EAX_REG_17__SCAN_IN), .ZN(n10442) );
  OAI211_X1 U13330 ( .C1(n14116), .C2(n19721), .A(n10443), .B(n10442), .ZN(
        n13959) );
  INV_X1 U13331 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19723) );
  NAND2_X1 U13332 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10445) );
  NAND2_X1 U13333 ( .A1(n14113), .A2(P2_EAX_REG_18__SCAN_IN), .ZN(n10444) );
  OAI211_X1 U13334 ( .C1(n14116), .C2(n19723), .A(n10445), .B(n10444), .ZN(
        n10446) );
  INV_X1 U13335 ( .A(n10446), .ZN(n15209) );
  INV_X1 U13336 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19725) );
  NAND2_X1 U13337 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10448) );
  NAND2_X1 U13338 ( .A1(n14113), .A2(P2_EAX_REG_19__SCAN_IN), .ZN(n10447) );
  OAI211_X1 U13339 ( .C1(n14116), .C2(n19725), .A(n10448), .B(n10447), .ZN(
        n10449) );
  INV_X1 U13340 ( .A(n10449), .ZN(n14905) );
  INV_X1 U13341 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n10452) );
  NAND2_X1 U13342 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10451) );
  NAND2_X1 U13343 ( .A1(n14113), .A2(P2_EAX_REG_20__SCAN_IN), .ZN(n10450) );
  OAI211_X1 U13344 ( .C1(n14116), .C2(n10452), .A(n10451), .B(n10450), .ZN(
        n14773) );
  INV_X1 U13345 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19728) );
  INV_X1 U13346 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n14899) );
  INV_X1 U13347 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15168) );
  OAI222_X1 U13348 ( .A1(n14116), .A2(n19728), .B1(n10005), .B2(n14899), .C1(
        n15168), .C2(n10453), .ZN(n14761) );
  AOI22_X1 U13349 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B1(
        n14113), .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n10455) );
  NAND2_X1 U13350 ( .A1(n10309), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n10454) );
  AND2_X1 U13351 ( .A1(n10455), .A2(n10454), .ZN(n14746) );
  NOR2_X2 U13352 ( .A1(n14745), .A2(n14746), .ZN(n14168) );
  INV_X1 U13353 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19731) );
  NAND2_X1 U13354 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10457) );
  NAND2_X1 U13355 ( .A1(n14113), .A2(P2_EAX_REG_23__SCAN_IN), .ZN(n10456) );
  OAI211_X1 U13356 ( .C1(n14116), .C2(n19731), .A(n10457), .B(n10456), .ZN(
        n14169) );
  INV_X1 U13357 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19733) );
  NAND2_X1 U13358 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10459) );
  NAND2_X1 U13359 ( .A1(n14113), .A2(P2_EAX_REG_24__SCAN_IN), .ZN(n10458) );
  OAI211_X1 U13360 ( .C1(n14116), .C2(n19733), .A(n10459), .B(n10458), .ZN(
        n10460) );
  INV_X1 U13361 ( .A(n10460), .ZN(n14881) );
  INV_X1 U13362 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19735) );
  NAND2_X1 U13363 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10462) );
  NAND2_X1 U13364 ( .A1(n14113), .A2(P2_EAX_REG_25__SCAN_IN), .ZN(n10461) );
  OAI211_X1 U13365 ( .C1(n14116), .C2(n19735), .A(n10462), .B(n10461), .ZN(
        n10463) );
  INV_X1 U13366 ( .A(n10463), .ZN(n14872) );
  INV_X1 U13367 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19739) );
  NAND2_X1 U13368 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10465) );
  NAND2_X1 U13369 ( .A1(n14113), .A2(P2_EAX_REG_27__SCAN_IN), .ZN(n10464) );
  OAI211_X1 U13370 ( .C1(n14116), .C2(n19739), .A(n10465), .B(n10464), .ZN(
        n14857) );
  INV_X1 U13371 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n14961) );
  NAND2_X1 U13372 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10468) );
  NAND2_X1 U13373 ( .A1(n14113), .A2(P2_EAX_REG_26__SCAN_IN), .ZN(n10467) );
  OAI211_X1 U13374 ( .C1(n14116), .C2(n14961), .A(n10468), .B(n10467), .ZN(
        n14865) );
  INV_X1 U13375 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19740) );
  NAND2_X1 U13376 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10470) );
  NAND2_X1 U13377 ( .A1(n14113), .A2(P2_EAX_REG_28__SCAN_IN), .ZN(n10469) );
  OAI211_X1 U13378 ( .C1(n14116), .C2(n19740), .A(n10470), .B(n10469), .ZN(
        n10471) );
  INV_X1 U13379 ( .A(n10471), .ZN(n14722) );
  INV_X1 U13380 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19743) );
  NAND2_X1 U13381 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10473) );
  NAND2_X1 U13382 ( .A1(n14113), .A2(P2_EAX_REG_29__SCAN_IN), .ZN(n10472) );
  OAI211_X1 U13383 ( .C1(n14116), .C2(n19743), .A(n10473), .B(n10472), .ZN(
        n11446) );
  INV_X1 U13384 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n14146) );
  NAND2_X1 U13385 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10475) );
  NAND2_X1 U13386 ( .A1(n14113), .A2(P2_EAX_REG_30__SCAN_IN), .ZN(n10474) );
  OAI211_X1 U13387 ( .C1(n14116), .C2(n14146), .A(n10475), .B(n10474), .ZN(
        n10477) );
  NAND2_X1 U13388 ( .A1(n10476), .A2(n10477), .ZN(n14118) );
  INV_X1 U13389 ( .A(n10476), .ZN(n10479) );
  INV_X1 U13390 ( .A(n10477), .ZN(n10478) );
  NAND2_X1 U13391 ( .A1(n10479), .A2(n10478), .ZN(n10480) );
  NAND2_X1 U13392 ( .A1(n14118), .A2(n10480), .ZN(n14144) );
  INV_X1 U13393 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n18723) );
  INV_X1 U13394 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19698) );
  NOR2_X1 U13395 ( .A1(n18723), .A2(n19698), .ZN(n19689) );
  NOR2_X1 U13396 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19691) );
  NOR3_X1 U13397 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19689), .A3(n19691), 
        .ZN(n19682) );
  NAND2_X1 U13398 ( .A1(n19669), .A2(n19682), .ZN(n13371) );
  INV_X1 U13399 ( .A(n13371), .ZN(n11380) );
  NAND3_X1 U13400 ( .A1(n19801), .A2(n19544), .A3(n11380), .ZN(n10481) );
  NOR2_X2 U13401 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19759) );
  AND2_X1 U13402 ( .A1(n19759), .A2(n19668), .ZN(n14200) );
  AND2_X2 U13403 ( .A1(n14200), .A2(n16078), .ZN(n19038) );
  NOR3_X1 U13404 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10482), .A3(n19611), 
        .ZN(n16061) );
  INV_X1 U13405 ( .A(n16061), .ZN(n10483) );
  NAND2_X1 U13406 ( .A1(n18863), .A2(n10483), .ZN(n10484) );
  NOR2_X1 U13407 ( .A1(n19038), .A2(n10484), .ZN(n10485) );
  INV_X1 U13408 ( .A(n10538), .ZN(n10506) );
  INV_X1 U13409 ( .A(n16076), .ZN(n13133) );
  NAND3_X1 U13410 ( .A1(n10538), .A2(n13133), .A3(n11383), .ZN(n13101) );
  OR2_X1 U13411 ( .A1(n13101), .A2(n16045), .ZN(n13094) );
  INV_X1 U13412 ( .A(n13094), .ZN(n13154) );
  INV_X1 U13413 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n15881) );
  OAI21_X1 U13414 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n19690), .A(n15881), 
        .ZN(n10486) );
  NOR2_X1 U13415 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n13371), .ZN(n16065) );
  AOI21_X1 U13416 ( .B1(n19054), .B2(n10486), .A(n16065), .ZN(n10487) );
  NAND2_X1 U13417 ( .A1(n13154), .A2(n10487), .ZN(n18864) );
  INV_X1 U13418 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n10680) );
  NAND2_X1 U13419 ( .A1(n18866), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18821) );
  INV_X1 U13420 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10488) );
  OAI22_X1 U13421 ( .A1(n18864), .A2(n10680), .B1(n18821), .B2(n10488), .ZN(
        n10489) );
  AOI21_X1 U13422 ( .B1(n18853), .B2(P2_REIP_REG_30__SCAN_IN), .A(n10489), 
        .ZN(n10490) );
  OAI21_X1 U13423 ( .B1(n14144), .B2(n18858), .A(n10490), .ZN(n10491) );
  AOI21_X1 U13424 ( .B1(n14095), .B2(n18786), .A(n10491), .ZN(n10492) );
  INV_X1 U13425 ( .A(n10492), .ZN(n10684) );
  NAND2_X1 U13426 ( .A1(n10493), .A2(n10006), .ZN(n10494) );
  NAND2_X1 U13427 ( .A1(n10495), .A2(n10494), .ZN(n11403) );
  AND2_X1 U13428 ( .A1(n10496), .A2(n16044), .ZN(n11405) );
  INV_X1 U13429 ( .A(n10497), .ZN(n10500) );
  NOR2_X1 U13430 ( .A1(n19085), .A2(n10498), .ZN(n10499) );
  NAND2_X1 U13431 ( .A1(n11403), .A2(n10545), .ZN(n10501) );
  NOR2_X1 U13432 ( .A1(n19048), .A2(n16078), .ZN(n14705) );
  NAND2_X1 U13433 ( .A1(n10501), .A2(n14705), .ZN(n10508) );
  INV_X1 U13434 ( .A(n10502), .ZN(n10504) );
  INV_X1 U13435 ( .A(n10509), .ZN(n10503) );
  NAND3_X1 U13436 ( .A1(n11352), .A2(n9588), .A3(n19054), .ZN(n10505) );
  NAND2_X1 U13437 ( .A1(n11440), .A2(n11377), .ZN(n10507) );
  AND2_X2 U13438 ( .A1(n10508), .A2(n10507), .ZN(n10536) );
  NAND2_X1 U13439 ( .A1(n10509), .A2(n10515), .ZN(n11385) );
  NAND2_X2 U13440 ( .A1(n10536), .A2(n10512), .ZN(n10568) );
  INV_X1 U13441 ( .A(n10568), .ZN(n10524) );
  AND2_X1 U13442 ( .A1(n10514), .A2(n10520), .ZN(n10517) );
  NAND2_X1 U13443 ( .A1(n10519), .A2(n10518), .ZN(n11401) );
  NOR2_X1 U13444 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n14711) );
  AOI21_X1 U13445 ( .B1(n11438), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10522), 
        .ZN(n10526) );
  INV_X1 U13446 ( .A(n10525), .ZN(n10523) );
  NAND2_X1 U13447 ( .A1(n10526), .A2(n9994), .ZN(n10527) );
  NAND2_X1 U13448 ( .A1(n10528), .A2(n10527), .ZN(n11028) );
  INV_X1 U13449 ( .A(n11028), .ZN(n10551) );
  INV_X1 U13450 ( .A(n11364), .ZN(n10529) );
  NAND2_X1 U13451 ( .A1(n11406), .A2(n10529), .ZN(n11408) );
  NAND3_X1 U13452 ( .A1(n10531), .A2(n19085), .A3(n10530), .ZN(n10532) );
  NOR2_X1 U13453 ( .A1(n11408), .A2(n10532), .ZN(n10553) );
  INV_X1 U13454 ( .A(n10553), .ZN(n10534) );
  NAND2_X1 U13455 ( .A1(n10538), .A2(n19801), .ZN(n10533) );
  AND2_X2 U13456 ( .A1(n10535), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10571) );
  NAND2_X1 U13457 ( .A1(n10571), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10550) );
  INV_X1 U13458 ( .A(n10536), .ZN(n10543) );
  OR2_X1 U13459 ( .A1(n10624), .A2(n18865), .ZN(n10541) );
  NAND2_X1 U13460 ( .A1(n10584), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10540) );
  INV_X1 U13461 ( .A(n14711), .ZN(n16066) );
  NAND2_X1 U13462 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10539) );
  NAND4_X1 U13463 ( .A1(n10541), .A2(n10540), .A3(n16066), .A4(n10539), .ZN(
        n10542) );
  NOR2_X1 U13464 ( .A1(n10543), .A2(n10542), .ZN(n10549) );
  INV_X1 U13465 ( .A(n10545), .ZN(n10546) );
  NAND3_X1 U13466 ( .A1(n10550), .A2(n10549), .A3(n10548), .ZN(n11029) );
  NAND2_X1 U13467 ( .A1(n10551), .A2(n11029), .ZN(n11027) );
  NAND2_X1 U13468 ( .A1(n10568), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10559) );
  INV_X1 U13469 ( .A(n10552), .ZN(n10554) );
  NOR2_X1 U13470 ( .A1(n10554), .A2(n10553), .ZN(n10556) );
  NAND2_X1 U13471 ( .A1(n10556), .A2(n10555), .ZN(n15379) );
  AOI21_X1 U13472 ( .B1(n15379), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10557), 
        .ZN(n10558) );
  NAND2_X1 U13473 ( .A1(n10559), .A2(n10558), .ZN(n10563) );
  NAND2_X1 U13474 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10560) );
  OAI211_X1 U13475 ( .C1(n10649), .C2(n13135), .A(n10561), .B(n10560), .ZN(
        n10562) );
  AOI21_X2 U13476 ( .B1(n10571), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n10562), .ZN(n10564) );
  NAND2_X1 U13477 ( .A1(n11027), .A2(n11036), .ZN(n10567) );
  INV_X1 U13478 ( .A(n10563), .ZN(n10565) );
  NAND2_X1 U13479 ( .A1(n10565), .A2(n10564), .ZN(n10566) );
  NAND2_X1 U13480 ( .A1(n10568), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10570) );
  AOI21_X1 U13481 ( .B1(n16078), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10569) );
  NAND2_X1 U13482 ( .A1(n10571), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10576) );
  NAND2_X1 U13483 ( .A1(n10584), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10573) );
  NAND2_X1 U13484 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10572) );
  OAI211_X1 U13485 ( .C1(n10624), .C2(n19701), .A(n10573), .B(n10572), .ZN(
        n10574) );
  INV_X1 U13486 ( .A(n10574), .ZN(n10575) );
  NAND2_X1 U13487 ( .A1(n11032), .A2(n10577), .ZN(n10578) );
  INV_X1 U13488 ( .A(n11032), .ZN(n10579) );
  NAND2_X1 U13489 ( .A1(n10579), .A2(n11033), .ZN(n10580) );
  NAND2_X1 U13490 ( .A1(n10568), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10583) );
  NAND2_X1 U13491 ( .A1(n14711), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10582) );
  NAND2_X1 U13492 ( .A1(n10584), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10586) );
  NAND2_X1 U13493 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10585) );
  OAI211_X1 U13494 ( .C1(n10624), .C2(n13657), .A(n10586), .B(n10585), .ZN(
        n10587) );
  INV_X1 U13495 ( .A(n10588), .ZN(n10589) );
  NOR2_X1 U13496 ( .A1(n10590), .A2(n10589), .ZN(n10591) );
  NAND2_X1 U13497 ( .A1(n10677), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10593) );
  AOI22_X1 U13498 ( .A1(n14107), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10592) );
  OAI211_X1 U13499 ( .C1(n14110), .C2(n18922), .A(n10593), .B(n10592), .ZN(
        n13720) );
  NAND2_X1 U13500 ( .A1(n14107), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n10595) );
  NAND2_X1 U13501 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10594) );
  OAI211_X1 U13502 ( .C1(n14181), .C2(n14110), .A(n10595), .B(n10594), .ZN(
        n10596) );
  AOI21_X1 U13503 ( .B1(n9595), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n10596), .ZN(n13706) );
  NAND2_X1 U13504 ( .A1(n9595), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10598) );
  AOI22_X1 U13505 ( .A1(n14107), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10597) );
  OAI211_X1 U13506 ( .C1(n14110), .C2(n10599), .A(n10598), .B(n10597), .ZN(
        n13447) );
  NAND2_X1 U13507 ( .A1(n14107), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n10601) );
  NAND2_X1 U13508 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10600) );
  OAI211_X1 U13509 ( .C1(n10602), .C2(n14110), .A(n10601), .B(n10600), .ZN(
        n10603) );
  AOI21_X1 U13510 ( .B1(n9595), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n10603), .ZN(n13456) );
  NAND2_X1 U13511 ( .A1(n9595), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10608) );
  INV_X1 U13512 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n13771) );
  NAND2_X1 U13513 ( .A1(n14107), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10605) );
  NAND2_X1 U13514 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10604) );
  OAI211_X1 U13515 ( .C1(n13771), .C2(n14110), .A(n10605), .B(n10604), .ZN(
        n10606) );
  INV_X1 U13516 ( .A(n10606), .ZN(n10607) );
  NAND2_X1 U13517 ( .A1(n10608), .A2(n10607), .ZN(n13773) );
  INV_X1 U13518 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10611) );
  NAND2_X1 U13519 ( .A1(n9595), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10610) );
  AOI22_X1 U13520 ( .A1(n14107), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10609) );
  OAI211_X1 U13521 ( .C1(n10611), .C2(n14110), .A(n10610), .B(n10609), .ZN(
        n13414) );
  INV_X1 U13522 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n10614) );
  NAND2_X1 U13523 ( .A1(n9595), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10613) );
  AOI22_X1 U13524 ( .A1(n14107), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n10612) );
  OAI211_X1 U13525 ( .C1(n10614), .C2(n14110), .A(n10613), .B(n10612), .ZN(
        n13786) );
  NAND2_X1 U13526 ( .A1(n14107), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n10616) );
  NAND2_X1 U13527 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10615) );
  OAI211_X1 U13528 ( .C1(n13528), .C2(n14110), .A(n10616), .B(n10615), .ZN(
        n10617) );
  AOI21_X1 U13529 ( .B1(n9595), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n10617), .ZN(n13524) );
  INV_X1 U13530 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n18808) );
  NAND2_X1 U13531 ( .A1(n9595), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10619) );
  AOI22_X1 U13532 ( .A1(n14107), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n10618) );
  OAI211_X1 U13533 ( .C1(n18808), .C2(n14110), .A(n10619), .B(n10618), .ZN(
        n15273) );
  NAND2_X1 U13534 ( .A1(n14107), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n10621) );
  NAND2_X1 U13535 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10620) );
  OAI211_X1 U13536 ( .C1(n10622), .C2(n14110), .A(n10621), .B(n10620), .ZN(
        n10623) );
  AOI21_X1 U13537 ( .B1(n9595), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n10623), .ZN(n13817) );
  NAND2_X1 U13538 ( .A1(n9595), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10629) );
  NAND2_X1 U13539 ( .A1(n14107), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n10626) );
  NAND2_X1 U13540 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10625) );
  OAI211_X1 U13541 ( .C1(n13807), .C2(n14110), .A(n10626), .B(n10625), .ZN(
        n10627) );
  INV_X1 U13542 ( .A(n10627), .ZN(n10628) );
  NAND2_X1 U13543 ( .A1(n10629), .A2(n10628), .ZN(n13802) );
  INV_X1 U13544 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n10632) );
  NAND2_X1 U13545 ( .A1(n14107), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n10631) );
  NAND2_X1 U13546 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10630) );
  OAI211_X1 U13547 ( .C1(n10632), .C2(n14110), .A(n10631), .B(n10630), .ZN(
        n10633) );
  AOI21_X1 U13548 ( .B1(n9595), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n10633), .ZN(n14081) );
  NAND2_X1 U13549 ( .A1(n14107), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n10635) );
  NAND2_X1 U13550 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10634) );
  OAI211_X1 U13551 ( .C1(n18886), .C2(n14110), .A(n10635), .B(n10634), .ZN(
        n10636) );
  AOI21_X1 U13552 ( .B1(n9595), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n10636), .ZN(n13926) );
  NAND2_X1 U13553 ( .A1(n9595), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10638) );
  AOI22_X1 U13554 ( .A1(n14107), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n10637) );
  OAI211_X1 U13555 ( .C1(n14110), .C2(n18781), .A(n10638), .B(n10637), .ZN(
        n13897) );
  NAND2_X1 U13556 ( .A1(n14107), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n10640) );
  NAND2_X1 U13557 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10639) );
  OAI211_X1 U13558 ( .C1(n18767), .C2(n14110), .A(n10640), .B(n10639), .ZN(
        n10641) );
  AOI21_X1 U13559 ( .B1(n9595), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n10641), .ZN(n15056) );
  NAND2_X1 U13560 ( .A1(n14107), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n10643) );
  NAND2_X1 U13561 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10642) );
  OAI211_X1 U13562 ( .C1(n18754), .C2(n14110), .A(n10643), .B(n10642), .ZN(
        n10644) );
  AOI21_X1 U13563 ( .B1(n9595), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n10644), .ZN(n14838) );
  NAND2_X1 U13564 ( .A1(n9595), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10646) );
  AOI22_X1 U13565 ( .A1(n14107), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n10645) );
  OAI211_X1 U13566 ( .C1(n14110), .C2(n14771), .A(n10646), .B(n10645), .ZN(
        n14769) );
  INV_X1 U13567 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n11270) );
  NAND2_X1 U13568 ( .A1(n9595), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10648) );
  AOI22_X1 U13569 ( .A1(n14107), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n10647) );
  OAI211_X1 U13570 ( .C1(n14110), .C2(n11270), .A(n10648), .B(n10647), .ZN(
        n14758) );
  INV_X1 U13571 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n10652) );
  NAND2_X1 U13572 ( .A1(n14107), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n10651) );
  NAND2_X1 U13573 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10650) );
  OAI211_X1 U13574 ( .C1(n10652), .C2(n14110), .A(n10651), .B(n10650), .ZN(
        n10653) );
  AOI21_X1 U13575 ( .B1(n9595), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n10653), .ZN(n14749) );
  NAND2_X1 U13576 ( .A1(n14107), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n10655) );
  NAND2_X1 U13577 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10654) );
  OAI211_X1 U13578 ( .C1(n10656), .C2(n14110), .A(n10655), .B(n10654), .ZN(
        n10657) );
  AOI21_X1 U13579 ( .B1(n9595), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n10657), .ZN(n14176) );
  NAND2_X1 U13580 ( .A1(n14107), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n10659) );
  NAND2_X1 U13581 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10658) );
  OAI211_X1 U13582 ( .C1(n10660), .C2(n14110), .A(n10659), .B(n10658), .ZN(
        n10661) );
  AOI21_X1 U13583 ( .B1(n9595), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n10661), .ZN(n14826) );
  NAND2_X1 U13584 ( .A1(n10677), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10663) );
  AOI22_X1 U13585 ( .A1(n14107), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n10662) );
  OAI211_X1 U13586 ( .C1(n14110), .C2(n14821), .A(n10663), .B(n10662), .ZN(
        n14819) );
  INV_X1 U13587 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n10666) );
  NAND2_X1 U13588 ( .A1(n14107), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n10665) );
  NAND2_X1 U13589 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10664) );
  OAI211_X1 U13590 ( .C1(n10666), .C2(n14110), .A(n10665), .B(n10664), .ZN(
        n10667) );
  AOI21_X1 U13591 ( .B1(n10677), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n10667), .ZN(n14813) );
  INV_X1 U13592 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n10670) );
  NAND2_X1 U13593 ( .A1(n14107), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n10669) );
  NAND2_X1 U13594 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10668) );
  OAI211_X1 U13595 ( .C1(n14110), .C2(n10670), .A(n10669), .B(n10668), .ZN(
        n10671) );
  AOI21_X1 U13596 ( .B1(n9595), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n10671), .ZN(n14801) );
  NAND2_X1 U13597 ( .A1(n9595), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10673) );
  AOI22_X1 U13598 ( .A1(n14107), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n10672) );
  OAI211_X1 U13599 ( .C1(n14110), .C2(n14725), .A(n10673), .B(n10672), .ZN(
        n14716) );
  INV_X1 U13600 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n10676) );
  NAND2_X1 U13601 ( .A1(n10677), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10675) );
  AOI22_X1 U13602 ( .A1(n14107), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n10674) );
  OAI211_X1 U13603 ( .C1(n14110), .C2(n10676), .A(n10675), .B(n10674), .ZN(
        n11436) );
  NAND2_X1 U13604 ( .A1(n9595), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10679) );
  AOI22_X1 U13605 ( .A1(n14107), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n10678) );
  OAI211_X1 U13606 ( .C1(n14110), .C2(n10680), .A(n10679), .B(n10678), .ZN(
        n14105) );
  NAND2_X1 U13607 ( .A1(n19800), .A2(n10681), .ZN(n10682) );
  NAND2_X1 U13608 ( .A1(n10686), .A2(n10685), .ZN(P2_U2825) );
  INV_X1 U13609 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18662) );
  INV_X1 U13610 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17714) );
  INV_X1 U13611 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17742) );
  INV_X1 U13612 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17850) );
  NAND2_X1 U13613 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17560) );
  INV_X1 U13614 ( .A(n17560), .ZN(n17895) );
  NAND2_X1 U13615 ( .A1(n17895), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17881) );
  INV_X1 U13616 ( .A(n17881), .ZN(n17542) );
  NAND2_X1 U13617 ( .A1(n17542), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17853) );
  INV_X1 U13618 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17857) );
  NOR2_X1 U13619 ( .A1(n17853), .A2(n17857), .ZN(n17851) );
  INV_X1 U13620 ( .A(n17851), .ZN(n17515) );
  INV_X1 U13621 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17860) );
  NOR2_X1 U13622 ( .A1(n17515), .A2(n17860), .ZN(n17829) );
  INV_X1 U13623 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16879) );
  NAND3_X2 U13624 ( .A1(n18683), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n18499), .ZN(n15418) );
  INV_X1 U13625 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16701) );
  OAI22_X1 U13626 ( .A1(n10797), .A2(n16879), .B1(n15418), .B2(n16701), .ZN(
        n10693) );
  AOI22_X1 U13627 ( .A1(n17025), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10692) );
  NOR3_X1 U13628 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n9675), .ZN(n10689) );
  AOI22_X1 U13629 ( .A1(n10745), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9571), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10691) );
  NOR2_X2 U13630 ( .A1(n16645), .A2(n10724), .ZN(n16990) );
  AOI22_X1 U13631 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10726), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10690) );
  INV_X2 U13632 ( .A(n10708), .ZN(n10814) );
  INV_X1 U13633 ( .A(n10740), .ZN(n10758) );
  AOI22_X1 U13634 ( .A1(n10758), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n15414), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10694) );
  OAI21_X1 U13635 ( .B1(n10814), .B2(n16702), .A(n10694), .ZN(n10697) );
  NAND2_X1 U13636 ( .A1(n18661), .A2(n18671), .ZN(n10695) );
  AOI22_X1 U13637 ( .A1(n17013), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10709), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10700) );
  INV_X1 U13638 ( .A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n16700) );
  INV_X1 U13639 ( .A(n10726), .ZN(n10741) );
  AOI22_X1 U13640 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n16734), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10715) );
  INV_X1 U13641 ( .A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n20868) );
  NAND2_X1 U13642 ( .A1(n9570), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10706) );
  NAND2_X1 U13643 ( .A1(n9576), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10705) );
  AND2_X1 U13644 ( .A1(n10706), .A2(n10705), .ZN(n10707) );
  OAI21_X1 U13645 ( .B1(n16958), .B2(n20868), .A(n10707), .ZN(n10713) );
  INV_X1 U13646 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18309) );
  AOI22_X1 U13647 ( .A1(n10758), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10708), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10711) );
  INV_X1 U13648 ( .A(n16723), .ZN(n10709) );
  AOI22_X1 U13649 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10709), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10710) );
  OAI211_X1 U13650 ( .C1(n16962), .C2(n18309), .A(n10711), .B(n10710), .ZN(
        n10712) );
  AOI211_X1 U13651 ( .C1(n16965), .C2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n10713), .B(n10712), .ZN(n10714) );
  OAI211_X1 U13652 ( .C1(n10741), .C2(n20898), .A(n10715), .B(n10714), .ZN(
        n10722) );
  INV_X1 U13653 ( .A(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16862) );
  AOI22_X1 U13654 ( .A1(n17025), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9577), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10716) );
  OAI21_X1 U13655 ( .B1(n16987), .B2(n16862), .A(n10716), .ZN(n10717) );
  INV_X1 U13656 ( .A(n10717), .ZN(n10720) );
  NOR2_X2 U13657 ( .A1(n10722), .A2(n10721), .ZN(n10754) );
  INV_X1 U13658 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18663) );
  OR2_X2 U13659 ( .A1(n16645), .A2(n10724), .ZN(n17011) );
  INV_X1 U13660 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18267) );
  AOI22_X1 U13661 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10735) );
  INV_X1 U13662 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18303) );
  AOI22_X1 U13663 ( .A1(n17009), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9578), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10728) );
  AOI22_X1 U13664 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n10726), .B1(
        P3_INSTQUEUE_REG_13__0__SCAN_IN), .B2(n10708), .ZN(n10727) );
  OAI211_X1 U13665 ( .C1(n18303), .C2(n16962), .A(n10728), .B(n10727), .ZN(
        n10734) );
  AOI22_X1 U13666 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n17013), .B1(
        P3_INSTQUEUE_REG_12__0__SCAN_IN), .B2(n10704), .ZN(n10732) );
  AOI22_X1 U13667 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__0__SCAN_IN), .B2(n10709), .ZN(n10731) );
  AOI22_X1 U13668 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n17025), .B1(
        n16734), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10730) );
  NAND2_X1 U13669 ( .A1(n16965), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10729) );
  NAND4_X1 U13670 ( .A1(n10732), .A2(n10731), .A3(n10730), .A4(n10729), .ZN(
        n10733) );
  NOR2_X1 U13671 ( .A1(n18663), .A2(n17203), .ZN(n10736) );
  NOR2_X1 U13672 ( .A1(n17686), .A2(n10736), .ZN(n17676) );
  NOR2_X1 U13673 ( .A1(n17675), .A2(n17676), .ZN(n17674) );
  NOR2_X1 U13674 ( .A1(n10723), .A2(n10737), .ZN(n10738) );
  XNOR2_X1 U13675 ( .A(n10755), .B(n10739), .ZN(n17666) );
  INV_X1 U13676 ( .A(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n20844) );
  AOI22_X1 U13677 ( .A1(n17009), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10753) );
  INV_X1 U13678 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16850) );
  AOI22_X1 U13679 ( .A1(n17013), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10743) );
  AOI22_X1 U13680 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10887), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10742) );
  OAI211_X1 U13681 ( .C1(n16958), .C2(n16850), .A(n10743), .B(n10742), .ZN(
        n10751) );
  AOI22_X1 U13682 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9579), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10749) );
  AOI22_X1 U13683 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10748) );
  AOI22_X1 U13684 ( .A1(n16734), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17025), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10747) );
  NAND2_X1 U13685 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10746) );
  NAND4_X1 U13686 ( .A1(n10749), .A2(n10748), .A3(n10747), .A4(n10746), .ZN(
        n10750) );
  XNOR2_X1 U13687 ( .A(n17193), .B(n10768), .ZN(n17665) );
  NOR2_X1 U13688 ( .A1(n10755), .A2(n10739), .ZN(n10756) );
  NOR2_X2 U13689 ( .A1(n17664), .A2(n10756), .ZN(n17657) );
  INV_X1 U13690 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17965) );
  INV_X1 U13691 ( .A(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16936) );
  INV_X1 U13692 ( .A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16934) );
  OAI22_X1 U13693 ( .A1(n9575), .A2(n16936), .B1(n10814), .B2(n16934), .ZN(
        n10767) );
  INV_X1 U13694 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16834) );
  AOI22_X1 U13695 ( .A1(n16734), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10765) );
  INV_X1 U13696 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18063) );
  AOI22_X1 U13697 ( .A1(n9578), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10757) );
  OAI21_X1 U13698 ( .B1(n10741), .B2(n18063), .A(n10757), .ZN(n10763) );
  AOI22_X1 U13699 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10761) );
  AOI22_X1 U13700 ( .A1(n10758), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9585), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10760) );
  AOI22_X1 U13701 ( .A1(n16893), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9571), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10759) );
  NAND3_X1 U13702 ( .A1(n10761), .A2(n10760), .A3(n10759), .ZN(n10762) );
  AOI211_X1 U13703 ( .C1(n17025), .C2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n10763), .B(n10762), .ZN(n10764) );
  OAI211_X1 U13704 ( .C1(n10009), .C2(n16834), .A(n10765), .B(n10764), .ZN(
        n10766) );
  AOI211_X4 U13705 ( .C1(n16955), .C2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A(
        n10767), .B(n10766), .ZN(n17189) );
  INV_X1 U13706 ( .A(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n20936) );
  AOI22_X1 U13707 ( .A1(n9579), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10780) );
  INV_X1 U13708 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n18319) );
  AOI22_X1 U13709 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U13710 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17025), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10771) );
  OAI211_X1 U13711 ( .C1(n16962), .C2(n18319), .A(n10772), .B(n10771), .ZN(
        n10778) );
  AOI22_X1 U13712 ( .A1(n10887), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10776) );
  AOI22_X1 U13713 ( .A1(n17009), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10775) );
  AOI22_X1 U13714 ( .A1(n16734), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10774) );
  NAND2_X1 U13715 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10773) );
  NAND4_X1 U13716 ( .A1(n10776), .A2(n10775), .A3(n10774), .A4(n10773), .ZN(
        n10777) );
  AOI211_X1 U13717 ( .C1(n16965), .C2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n10778), .B(n10777), .ZN(n10779) );
  INV_X1 U13718 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17953) );
  INV_X1 U13719 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18286) );
  AOI22_X1 U13720 ( .A1(n16734), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10791) );
  INV_X1 U13721 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18323) );
  AOI22_X1 U13722 ( .A1(n17009), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9577), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10783) );
  AOI22_X1 U13723 ( .A1(n17025), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10782) );
  OAI211_X1 U13724 ( .C1(n16962), .C2(n18323), .A(n10783), .B(n10782), .ZN(
        n10789) );
  AOI22_X1 U13725 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10887), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10787) );
  AOI22_X1 U13726 ( .A1(n16988), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10786) );
  AOI22_X1 U13727 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10785) );
  NAND2_X1 U13728 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n10784) );
  NAND4_X1 U13729 ( .A1(n10787), .A2(n10786), .A3(n10785), .A4(n10784), .ZN(
        n10788) );
  AOI211_X1 U13730 ( .C1(n16965), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n10789), .B(n10788), .ZN(n10790) );
  OAI211_X1 U13731 ( .C1(n17011), .C2(n18286), .A(n10791), .B(n10790), .ZN(
        n10792) );
  NOR2_X2 U13732 ( .A1(n17625), .A2(n10795), .ZN(n10809) );
  INV_X1 U13733 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16724) );
  AOI22_X1 U13734 ( .A1(n17013), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10807) );
  INV_X1 U13735 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16764) );
  AOI22_X1 U13736 ( .A1(n9578), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10887), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10799) );
  AOI22_X1 U13737 ( .A1(n17009), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9585), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10798) );
  OAI211_X1 U13738 ( .C1(n16958), .C2(n16764), .A(n10799), .B(n10798), .ZN(
        n10805) );
  AOI22_X1 U13739 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10803) );
  AOI22_X1 U13740 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17025), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10802) );
  AOI22_X1 U13741 ( .A1(n16955), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10801) );
  NAND2_X1 U13742 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10800) );
  NAND4_X1 U13743 ( .A1(n10803), .A2(n10802), .A3(n10801), .A4(n10800), .ZN(
        n10804) );
  AOI211_X1 U13744 ( .C1(n16965), .C2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n10805), .B(n10804), .ZN(n10806) );
  XNOR2_X1 U13745 ( .A(n10809), .B(n10808), .ZN(n17621) );
  INV_X1 U13746 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17943) );
  NOR2_X1 U13747 ( .A1(n10809), .A2(n10808), .ZN(n10810) );
  INV_X1 U13748 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17929) );
  NAND2_X1 U13749 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17811) );
  INV_X1 U13750 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17812) );
  NOR2_X1 U13751 ( .A1(n17811), .A2(n17812), .ZN(n17441) );
  INV_X1 U13752 ( .A(n17441), .ZN(n17773) );
  INV_X1 U13753 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17800) );
  INV_X1 U13754 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17787) );
  NOR2_X1 U13755 ( .A1(n17800), .A2(n17787), .ZN(n17778) );
  NAND2_X1 U13756 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17778), .ZN(
        n17766) );
  NOR2_X1 U13757 ( .A1(n17773), .A2(n17766), .ZN(n17764) );
  INV_X1 U13758 ( .A(n17764), .ZN(n17424) );
  INV_X1 U13759 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17427) );
  NOR2_X1 U13760 ( .A1(n17424), .A2(n17427), .ZN(n17751) );
  NAND2_X1 U13761 ( .A1(n17751), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17389) );
  INV_X1 U13762 ( .A(n17389), .ZN(n10907) );
  NAND2_X1 U13763 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17375), .ZN(
        n17374) );
  NAND2_X1 U13764 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16124) );
  INV_X1 U13765 ( .A(n16124), .ZN(n16113) );
  NAND2_X1 U13766 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16113), .ZN(
        n15498) );
  INV_X1 U13767 ( .A(n15498), .ZN(n11021) );
  NAND3_X1 U13768 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15451), .A3(
        n11021), .ZN(n10811) );
  XNOR2_X1 U13769 ( .A(n18662), .B(n10811), .ZN(n16100) );
  AOI22_X1 U13770 ( .A1(n16955), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10822) );
  INV_X1 U13771 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18274) );
  AOI22_X1 U13772 ( .A1(n17025), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10813) );
  AOI22_X1 U13773 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9579), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10812) );
  OAI211_X1 U13774 ( .C1(n16962), .C2(n18274), .A(n10813), .B(n10812), .ZN(
        n10820) );
  AOI22_X1 U13775 ( .A1(n17010), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10818) );
  AOI22_X1 U13776 ( .A1(n17009), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9585), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10817) );
  AOI22_X1 U13777 ( .A1(n16734), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10887), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10816) );
  NAND2_X1 U13778 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n10815) );
  NAND4_X1 U13779 ( .A1(n10818), .A2(n10817), .A3(n10816), .A4(n10815), .ZN(
        n10819) );
  INV_X1 U13780 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n20895) );
  AOI22_X1 U13781 ( .A1(n16893), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10887), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10832) );
  AOI22_X1 U13782 ( .A1(n17013), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10824) );
  AOI22_X1 U13783 ( .A1(n16991), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10823) );
  OAI211_X1 U13784 ( .C1(n16962), .C2(n18267), .A(n10824), .B(n10823), .ZN(
        n10830) );
  AOI22_X1 U13785 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17012), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10828) );
  AOI22_X1 U13786 ( .A1(n17009), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9585), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10827) );
  AOI22_X1 U13787 ( .A1(n17025), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9579), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10826) );
  NAND2_X1 U13788 ( .A1(n16734), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10825) );
  NAND4_X1 U13789 ( .A1(n10828), .A2(n10827), .A3(n10826), .A4(n10825), .ZN(
        n10829) );
  AOI22_X1 U13790 ( .A1(n17013), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10842) );
  INV_X1 U13791 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18271) );
  AOI22_X1 U13792 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17012), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10834) );
  AOI22_X1 U13793 ( .A1(n17009), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10887), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10833) );
  OAI211_X1 U13794 ( .C1(n16962), .C2(n18271), .A(n10834), .B(n10833), .ZN(
        n10840) );
  AOI22_X1 U13795 ( .A1(n17025), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9579), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10838) );
  AOI22_X1 U13796 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10837) );
  AOI22_X1 U13797 ( .A1(n16955), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10836) );
  NAND2_X1 U13798 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10835) );
  NAND4_X1 U13799 ( .A1(n10838), .A2(n10837), .A3(n10836), .A4(n10835), .ZN(
        n10839) );
  NAND2_X1 U13800 ( .A1(n9671), .A2(n10958), .ZN(n10966) );
  AOI22_X1 U13801 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16734), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10852) );
  INV_X1 U13802 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n18280) );
  AOI22_X1 U13803 ( .A1(n10887), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17010), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10844) );
  AOI22_X1 U13804 ( .A1(n17025), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10843) );
  OAI211_X1 U13805 ( .C1(n16962), .C2(n18280), .A(n10844), .B(n10843), .ZN(
        n10850) );
  AOI22_X1 U13806 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10848) );
  AOI22_X1 U13807 ( .A1(n17009), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9578), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10847) );
  AOI22_X1 U13808 ( .A1(n16955), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10846) );
  NAND2_X1 U13809 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10845) );
  NAND4_X1 U13810 ( .A1(n10848), .A2(n10847), .A3(n10846), .A4(n10845), .ZN(
        n10849) );
  INV_X1 U13811 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18069) );
  AOI22_X1 U13812 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10862) );
  INV_X1 U13813 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18283) );
  AOI22_X1 U13814 ( .A1(n17009), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9579), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10854) );
  AOI22_X1 U13815 ( .A1(n10887), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10853) );
  OAI211_X1 U13816 ( .C1(n16962), .C2(n18283), .A(n10854), .B(n10853), .ZN(
        n10860) );
  AOI22_X1 U13817 ( .A1(n17013), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10858) );
  AOI22_X1 U13818 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17010), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U13819 ( .A1(n16734), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17025), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10856) );
  NAND2_X1 U13820 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10855) );
  NAND4_X1 U13821 ( .A1(n10858), .A2(n10857), .A3(n10856), .A4(n10855), .ZN(
        n10859) );
  INV_X1 U13822 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18074) );
  AOI22_X1 U13823 ( .A1(n16734), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10872) );
  AOI22_X1 U13824 ( .A1(n17009), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10864) );
  AOI22_X1 U13825 ( .A1(n9577), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10863) );
  OAI211_X1 U13826 ( .C1(n16962), .C2(n18286), .A(n10864), .B(n10863), .ZN(
        n10870) );
  AOI22_X1 U13827 ( .A1(n10887), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10868) );
  AOI22_X1 U13828 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17025), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10867) );
  AOI22_X1 U13829 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10866) );
  NAND2_X1 U13830 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10865) );
  NAND4_X1 U13831 ( .A1(n10868), .A2(n10867), .A3(n10866), .A4(n10865), .ZN(
        n10869) );
  INV_X1 U13832 ( .A(n17060), .ZN(n18071) );
  NAND2_X1 U13833 ( .A1(n10957), .A2(n18071), .ZN(n15512) );
  INV_X1 U13834 ( .A(n15512), .ZN(n18525) );
  NOR2_X1 U13835 ( .A1(n18071), .A2(n10957), .ZN(n10956) );
  INV_X1 U13836 ( .A(n10956), .ZN(n10898) );
  INV_X1 U13837 ( .A(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n20923) );
  AOI22_X1 U13838 ( .A1(n16955), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9571), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10883) );
  INV_X1 U13839 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18293) );
  AOI22_X1 U13840 ( .A1(n16988), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10875) );
  AOI22_X1 U13841 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10726), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10874) );
  OAI211_X1 U13842 ( .C1(n16962), .C2(n18293), .A(n10875), .B(n10874), .ZN(
        n10881) );
  AOI22_X1 U13843 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9585), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10879) );
  AOI22_X1 U13844 ( .A1(n17009), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10744), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10878) );
  AOI22_X1 U13845 ( .A1(n9577), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10877) );
  NAND2_X1 U13846 ( .A1(n16734), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10876) );
  NAND4_X1 U13847 ( .A1(n10879), .A2(n10878), .A3(n10877), .A4(n10876), .ZN(
        n10880) );
  OAI211_X4 U13848 ( .C1(n10886), .C2(n20923), .A(n10883), .B(n10882), .ZN(
        n17176) );
  INV_X1 U13849 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18057) );
  AOI22_X1 U13850 ( .A1(n16734), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10890) );
  INV_X1 U13851 ( .A(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16961) );
  AOI22_X1 U13852 ( .A1(n10884), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10885) );
  OAI21_X1 U13853 ( .B1(n10886), .B2(n16961), .A(n10885), .ZN(n10889) );
  INV_X1 U13854 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n20910) );
  AOI22_X1 U13855 ( .A1(n17025), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9579), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10888) );
  INV_X1 U13856 ( .A(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16954) );
  AOI22_X1 U13857 ( .A1(n17009), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10891) );
  OAI21_X1 U13858 ( .B1(n10892), .B2(n16954), .A(n10891), .ZN(n10893) );
  NOR2_X2 U13859 ( .A1(n18077), .A2(n18054), .ZN(n10974) );
  OAI211_X1 U13860 ( .C1(n18059), .C2(n18525), .A(n10898), .B(n10974), .ZN(
        n10899) );
  NOR2_X1 U13861 ( .A1(n10966), .A2(n10899), .ZN(n10980) );
  NAND2_X1 U13862 ( .A1(n9671), .A2(n18702), .ZN(n10900) );
  NOR2_X1 U13863 ( .A1(n18071), .A2(n10900), .ZN(n11014) );
  NAND2_X1 U13864 ( .A1(n10980), .A2(n11014), .ZN(n18491) );
  NOR2_X1 U13865 ( .A1(n16082), .A2(n18491), .ZN(n17890) );
  INV_X1 U13866 ( .A(n17890), .ZN(n17835) );
  INV_X1 U13867 ( .A(n18491), .ZN(n17991) );
  NAND2_X1 U13868 ( .A1(n17991), .A2(n16082), .ZN(n17844) );
  AOI22_X1 U13869 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17597), .B1(
        n17557), .B2(n18662), .ZN(n10920) );
  INV_X1 U13870 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15496) );
  NAND2_X1 U13871 ( .A1(n17829), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16106) );
  OAI21_X2 U13872 ( .B1(n10902), .B2(n17597), .A(n17931), .ZN(n17572) );
  NOR2_X2 U13873 ( .A1(n16106), .A2(n17572), .ZN(n17420) );
  INV_X1 U13874 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10903) );
  INV_X1 U13875 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17913) );
  INV_X1 U13876 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17571) );
  NAND2_X1 U13877 ( .A1(n17913), .A2(n17571), .ZN(n17581) );
  NAND2_X1 U13878 ( .A1(n17541), .A2(n17857), .ZN(n17501) );
  NOR2_X1 U13879 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10906) );
  INV_X1 U13880 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17819) );
  NAND2_X1 U13881 ( .A1(n17420), .A2(n10907), .ZN(n10909) );
  NAND2_X1 U13882 ( .A1(n17470), .A2(n17800), .ZN(n10908) );
  NOR2_X1 U13883 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n10908), .ZN(
        n17434) );
  INV_X1 U13884 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17775) );
  NAND2_X1 U13885 ( .A1(n17434), .A2(n17775), .ZN(n17422) );
  NOR2_X2 U13886 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17383), .ZN(
        n17382) );
  INV_X1 U13887 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17756) );
  INV_X1 U13888 ( .A(n17811), .ZN(n17806) );
  NAND2_X1 U13889 ( .A1(n17806), .A2(n17420), .ZN(n17432) );
  NOR2_X1 U13890 ( .A1(n17766), .A2(n17427), .ZN(n17720) );
  AND2_X1 U13891 ( .A1(n17720), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10911) );
  INV_X1 U13892 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17727) );
  OR2_X1 U13893 ( .A1(n17557), .A2(n17382), .ZN(n17376) );
  OAI21_X2 U13894 ( .B1(n10912), .B2(n9986), .A(n17376), .ZN(n17358) );
  NOR2_X2 U13895 ( .A1(n17358), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17357) );
  INV_X1 U13896 ( .A(n10912), .ZN(n10913) );
  NAND2_X1 U13897 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17557), .ZN(
        n16131) );
  NAND2_X1 U13898 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15448), .ZN(
        n15495) );
  OR2_X2 U13899 ( .A1(n10915), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17342) );
  NAND2_X1 U13900 ( .A1(n17597), .A2(n10916), .ZN(n10917) );
  INV_X1 U13901 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n20920) );
  NAND2_X1 U13902 ( .A1(n15447), .A2(n20920), .ZN(n15494) );
  NAND2_X1 U13903 ( .A1(n17597), .A2(n15494), .ZN(n10922) );
  OAI211_X1 U13904 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n15496), .A(
        n15495), .B(n10922), .ZN(n10918) );
  NAND2_X1 U13905 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n15496), .ZN(
        n11022) );
  NOR2_X1 U13906 ( .A1(n10920), .A2(n10919), .ZN(n10921) );
  INV_X1 U13907 ( .A(n17751), .ZN(n17410) );
  NAND2_X1 U13908 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17721) );
  NOR2_X1 U13909 ( .A1(n17410), .A2(n17721), .ZN(n17723) );
  NAND2_X1 U13910 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17723), .ZN(
        n17356) );
  NAND2_X1 U13911 ( .A1(n17695), .A2(n17203), .ZN(n10926) );
  NAND2_X1 U13912 ( .A1(n10754), .A2(n10926), .ZN(n10925) );
  NAND2_X1 U13913 ( .A1(n10925), .A2(n17193), .ZN(n10937) );
  NOR2_X1 U13914 ( .A1(n17189), .A2(n10937), .ZN(n10924) );
  NAND2_X1 U13915 ( .A1(n10924), .A2(n10923), .ZN(n10943) );
  NOR2_X1 U13916 ( .A1(n17183), .A2(n10943), .ZN(n10947) );
  NAND2_X1 U13917 ( .A1(n10947), .A2(n16082), .ZN(n10948) );
  INV_X1 U13918 ( .A(n10923), .ZN(n17186) );
  XNOR2_X1 U13919 ( .A(n10924), .B(n17186), .ZN(n10941) );
  AND2_X1 U13920 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n10941), .ZN(
        n10942) );
  XOR2_X1 U13921 ( .A(n10925), .B(n17193), .Z(n10934) );
  XOR2_X1 U13922 ( .A(n10926), .B(n10754), .Z(n10927) );
  NOR2_X1 U13923 ( .A1(n10927), .A2(n10723), .ZN(n10933) );
  XOR2_X1 U13924 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n10927), .Z(
        n17678) );
  INV_X1 U13925 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18680) );
  NOR2_X1 U13926 ( .A1(n10929), .A2(n18680), .ZN(n10931) );
  INV_X1 U13927 ( .A(n17695), .ZN(n10930) );
  NAND3_X1 U13928 ( .A1(n10930), .A2(n10929), .A3(n18680), .ZN(n10928) );
  OAI221_X1 U13929 ( .B1(n10931), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n10930), .C2(n10929), .A(n10928), .ZN(n17677) );
  NOR2_X1 U13930 ( .A1(n17678), .A2(n17677), .ZN(n10932) );
  NOR2_X1 U13931 ( .A1(n10933), .A2(n10932), .ZN(n17663) );
  XOR2_X1 U13932 ( .A(n10739), .B(n10934), .Z(n17662) );
  NOR2_X1 U13933 ( .A1(n17663), .A2(n17662), .ZN(n10935) );
  XNOR2_X1 U13934 ( .A(n10937), .B(n17189), .ZN(n10939) );
  NOR2_X1 U13935 ( .A1(n10938), .A2(n10939), .ZN(n10940) );
  XNOR2_X1 U13936 ( .A(n10939), .B(n10938), .ZN(n17652) );
  XNOR2_X1 U13937 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n10941), .ZN(
        n17637) );
  XNOR2_X1 U13938 ( .A(n10943), .B(n17183), .ZN(n10945) );
  NOR2_X1 U13939 ( .A1(n10944), .A2(n10945), .ZN(n10946) );
  XNOR2_X1 U13940 ( .A(n10945), .B(n10944), .ZN(n17631) );
  XNOR2_X1 U13941 ( .A(n10947), .B(n16082), .ZN(n10950) );
  NAND2_X1 U13942 ( .A1(n10949), .A2(n10950), .ZN(n17612) );
  INV_X1 U13943 ( .A(n10948), .ZN(n10953) );
  OR2_X1 U13944 ( .A1(n10950), .A2(n10949), .ZN(n17613) );
  OAI21_X1 U13945 ( .B1(n10953), .B2(n10952), .A(n17613), .ZN(n10951) );
  INV_X1 U13946 ( .A(n16106), .ZN(n17804) );
  NAND3_X1 U13947 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16112), .A3(
        n11021), .ZN(n10955) );
  XNOR2_X1 U13948 ( .A(n18662), .B(n10955), .ZN(n16096) );
  NAND2_X1 U13949 ( .A1(n18046), .A2(n16266), .ZN(n10961) );
  NAND2_X1 U13950 ( .A1(n10958), .A2(n10961), .ZN(n18717) );
  NOR2_X1 U13951 ( .A1(n18059), .A2(n17060), .ZN(n18502) );
  NAND3_X1 U13952 ( .A1(n10974), .A2(n11003), .A3(n18502), .ZN(n15430) );
  NAND2_X1 U13953 ( .A1(n10957), .A2(n17060), .ZN(n10965) );
  NAND2_X1 U13954 ( .A1(n10973), .A2(n11001), .ZN(n10984) );
  NAND2_X1 U13955 ( .A1(n17271), .A2(n10984), .ZN(n16247) );
  INV_X1 U13956 ( .A(n16247), .ZN(n16242) );
  OR2_X2 U13957 ( .A1(n10958), .A2(n16242), .ZN(n13092) );
  AOI21_X4 U13958 ( .B1(n10960), .B2(n10959), .A(n16265), .ZN(n18511) );
  AOI21_X1 U13959 ( .B1(n17176), .B2(n15512), .A(n10961), .ZN(n10981) );
  INV_X1 U13960 ( .A(n10981), .ZN(n10962) );
  OAI21_X1 U13961 ( .B1(n11003), .B2(n10963), .A(n10962), .ZN(n10971) );
  NOR2_X1 U13962 ( .A1(n11001), .A2(n10965), .ZN(n11009) );
  NOR2_X1 U13963 ( .A1(n10963), .A2(n11009), .ZN(n10970) );
  AOI22_X1 U13964 ( .A1(n18054), .A2(n10964), .B1(n18059), .B2(n18525), .ZN(
        n10969) );
  NAND2_X1 U13965 ( .A1(n17176), .A2(n10965), .ZN(n10967) );
  AOI22_X1 U13966 ( .A1(n10967), .A2(n11010), .B1(n10966), .B2(n10965), .ZN(
        n10968) );
  OAI211_X1 U13967 ( .C1(n10970), .C2(n16266), .A(n10969), .B(n10968), .ZN(
        n10982) );
  NAND2_X1 U13968 ( .A1(n10973), .A2(n10975), .ZN(n14059) );
  OR2_X1 U13969 ( .A1(n18046), .A2(n10974), .ZN(n10976) );
  AOI21_X4 U13970 ( .B1(n18501), .B2(n18511), .A(n18500), .ZN(n18514) );
  NOR2_X4 U13971 ( .A1(n18702), .A2(n17926), .ZN(n18486) );
  NAND3_X1 U13972 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n11021), .A3(
        n18662), .ZN(n10979) );
  NOR2_X1 U13973 ( .A1(n17356), .A2(n17714), .ZN(n17708) );
  INV_X1 U13974 ( .A(n18497), .ZN(n18519) );
  AOI21_X1 U13975 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n17968) );
  NAND3_X1 U13976 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10978) );
  NOR2_X1 U13977 ( .A1(n17968), .A2(n10978), .ZN(n17924) );
  NAND2_X1 U13978 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17925) );
  NOR2_X1 U13979 ( .A1(n17925), .A2(n17929), .ZN(n10977) );
  NAND2_X1 U13980 ( .A1(n17924), .A2(n10977), .ZN(n17852) );
  NOR2_X1 U13981 ( .A1(n17852), .A2(n16106), .ZN(n17807) );
  INV_X1 U13982 ( .A(n17807), .ZN(n17719) );
  INV_X1 U13983 ( .A(n10977), .ZN(n17802) );
  INV_X1 U13984 ( .A(n10978), .ZN(n17801) );
  NAND3_X1 U13985 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n17801), .ZN(n17922) );
  NOR2_X1 U13986 ( .A1(n17802), .A2(n17922), .ZN(n17868) );
  INV_X1 U13987 ( .A(n17868), .ZN(n17904) );
  NOR2_X1 U13988 ( .A1(n16106), .A2(n17904), .ZN(n11018) );
  INV_X1 U13989 ( .A(n11018), .ZN(n17760) );
  INV_X1 U13990 ( .A(n18506), .ZN(n18526) );
  NAND2_X1 U13991 ( .A1(n18526), .A2(n18680), .ZN(n18011) );
  NAND2_X1 U13992 ( .A1(n18011), .A2(n17970), .ZN(n17988) );
  OAI22_X1 U13993 ( .A1(n18519), .A2(n17719), .B1(n17760), .B2(n17988), .ZN(
        n17722) );
  NAND2_X1 U13994 ( .A1(n17708), .A2(n17722), .ZN(n15454) );
  OAI22_X1 U13995 ( .A1(n16096), .A2(n17999), .B1(n10979), .B2(n15454), .ZN(
        n11016) );
  INV_X1 U13996 ( .A(n10980), .ZN(n10983) );
  AOI211_X1 U13997 ( .C1(n10984), .C2(n10983), .A(n10982), .B(n10981), .ZN(
        n14065) );
  NOR2_X1 U13998 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18683), .ZN(
        n10991) );
  AOI21_X1 U13999 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n18683), .A(
        n10991), .ZN(n11005) );
  OAI22_X1 U14000 ( .A1(n10687), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n18530), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10990) );
  INV_X1 U14001 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18539) );
  INV_X1 U14002 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18535) );
  AOI22_X1 U14003 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18535), .B1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18671), .ZN(n10992) );
  INV_X1 U14004 ( .A(n10990), .ZN(n11004) );
  NAND2_X1 U14005 ( .A1(n11004), .A2(n10991), .ZN(n10985) );
  OAI21_X1 U14006 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n10687), .A(
        n10985), .ZN(n10993) );
  NAND2_X1 U14007 ( .A1(n10992), .A2(n10993), .ZN(n10986) );
  OAI21_X1 U14008 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18671), .A(
        n10986), .ZN(n10987) );
  NAND2_X1 U14009 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10987), .ZN(
        n10995) );
  OAI22_X1 U14010 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18539), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n10987), .ZN(n10996) );
  AOI21_X1 U14011 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n10995), .A(
        n10996), .ZN(n10988) );
  AOI21_X1 U14012 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18539), .A(
        n10988), .ZN(n10997) );
  NAND2_X1 U14013 ( .A1(n10991), .A2(n10990), .ZN(n10989) );
  OAI211_X1 U14014 ( .C1(n10991), .C2(n10990), .A(n10997), .B(n10989), .ZN(
        n11000) );
  XNOR2_X1 U14015 ( .A(n10993), .B(n10992), .ZN(n10999) );
  NOR2_X1 U14016 ( .A1(n18539), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10994) );
  AOI22_X1 U14017 ( .A1(n10996), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(
        n10995), .B2(n10994), .ZN(n11006) );
  INV_X1 U14018 ( .A(n11006), .ZN(n10998) );
  OAI21_X1 U14019 ( .B1(n10999), .B2(n10998), .A(n10997), .ZN(n11007) );
  OAI21_X1 U14020 ( .B1(n11005), .B2(n11000), .A(n11007), .ZN(n18492) );
  NAND2_X1 U14021 ( .A1(n11007), .A2(n11000), .ZN(n18488) );
  INV_X1 U14022 ( .A(n18488), .ZN(n14060) );
  INV_X1 U14023 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18578) );
  NAND2_X1 U14024 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18578), .ZN(n18713) );
  AND2_X1 U14025 ( .A1(n18712), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18586) );
  NOR2_X1 U14026 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18566) );
  NOR3_X1 U14027 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18586), .A3(n18566), 
        .ZN(n18701) );
  XNOR2_X1 U14028 ( .A(n18046), .B(n11001), .ZN(n11002) );
  NAND2_X1 U14029 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18697) );
  OAI21_X1 U14030 ( .B1(n18701), .B2(n11002), .A(n18697), .ZN(n16246) );
  NOR3_X1 U14031 ( .A1(n11003), .A2(n14060), .A3(n16246), .ZN(n11013) );
  AND3_X1 U14032 ( .A1(n11006), .A2(n11005), .A3(n11004), .ZN(n11008) );
  OAI21_X1 U14033 ( .B1(n11010), .B2(n11009), .A(n18490), .ZN(n11011) );
  INV_X1 U14034 ( .A(n11011), .ZN(n11012) );
  AOI211_X1 U14035 ( .C1(n11014), .C2(n18492), .A(n11013), .B(n11012), .ZN(
        n11015) );
  INV_X1 U14036 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18715) );
  INV_X1 U14037 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18664) );
  NAND2_X1 U14038 ( .A1(n18664), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n16284) );
  NOR2_X1 U14039 ( .A1(n18715), .A2(n16284), .ZN(n18700) );
  INV_X1 U14040 ( .A(n18700), .ZN(n18552) );
  AOI21_X2 U14041 ( .B1(n14065), .B2(n11015), .A(n18552), .ZN(n18006) );
  INV_X1 U14042 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18705) );
  NOR2_X1 U14043 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18716) );
  NAND3_X1 U14044 ( .A1(n18705), .A2(n18715), .A3(n18716), .ZN(n18017) );
  INV_X1 U14045 ( .A(n17909), .ZN(n17815) );
  CLKBUF_X1 U14046 ( .A(n18017), .Z(n17909) );
  NAND2_X1 U14047 ( .A1(n17909), .A2(n18023), .ZN(n18007) );
  AOI21_X1 U14048 ( .B1(n17807), .B2(n17708), .A(n18519), .ZN(n17706) );
  NOR2_X1 U14049 ( .A1(n18680), .A2(n17904), .ZN(n17917) );
  NAND2_X1 U14050 ( .A1(n17804), .A2(n17917), .ZN(n17827) );
  INV_X1 U14051 ( .A(n17827), .ZN(n11017) );
  AND2_X1 U14052 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17708), .ZN(
        n16130) );
  AOI21_X1 U14053 ( .B1(n11017), .B2(n16130), .A(n18514), .ZN(n11020) );
  AOI21_X1 U14054 ( .B1(n17708), .B2(n11018), .A(n18526), .ZN(n11019) );
  NOR4_X1 U14055 ( .A1(n17982), .A2(n17706), .A3(n11020), .A4(n11019), .ZN(
        n15450) );
  INV_X1 U14056 ( .A(n17926), .ZN(n17744) );
  NOR2_X1 U14057 ( .A1(n18023), .A2(n17744), .ZN(n18012) );
  INV_X1 U14058 ( .A(n18012), .ZN(n17972) );
  OAI22_X1 U14059 ( .A1(n17815), .A2(n15450), .B1(n11021), .B2(n17972), .ZN(
        n15501) );
  AOI22_X1 U14060 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n17815), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n15501), .ZN(n11023) );
  NAND3_X1 U14061 ( .A1(n11024), .A2(n11023), .A3(n9990), .ZN(P3_U2831) );
  XNOR2_X2 U14062 ( .A(n11026), .B(n11025), .ZN(n11061) );
  INV_X1 U14063 ( .A(n11029), .ZN(n11030) );
  NAND2_X1 U14064 ( .A1(n11028), .A2(n11030), .ZN(n11031) );
  NAND2_X2 U14065 ( .A1(n11037), .A2(n11031), .ZN(n15355) );
  INV_X1 U14066 ( .A(n11036), .ZN(n11039) );
  INV_X1 U14067 ( .A(n11037), .ZN(n11038) );
  NOR2_X2 U14068 ( .A1(n11071), .A2(n11042), .ZN(n15401) );
  INV_X1 U14069 ( .A(n9593), .ZN(n11040) );
  AND2_X2 U14070 ( .A1(n11076), .A2(n11041), .ZN(n11138) );
  AOI22_X1 U14071 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n15401), .B1(
        n11138), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11069) );
  INV_X1 U14072 ( .A(n11042), .ZN(n11043) );
  AOI22_X1 U14073 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19205), .B1(
        n11134), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11068) );
  INV_X2 U14074 ( .A(n11498), .ZN(n13278) );
  INV_X1 U14075 ( .A(n15355), .ZN(n18875) );
  NAND2_X1 U14076 ( .A1(n18875), .A2(n11045), .ZN(n11048) );
  OR2_X1 U14077 ( .A1(n9593), .A2(n11048), .ZN(n11059) );
  INV_X1 U14078 ( .A(n11059), .ZN(n11044) );
  INV_X1 U14079 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11718) );
  INV_X1 U14080 ( .A(n11051), .ZN(n11046) );
  NAND2_X1 U14081 ( .A1(n9593), .A2(n11046), .ZN(n11056) );
  INV_X1 U14082 ( .A(n11056), .ZN(n11047) );
  NAND2_X1 U14083 ( .A1(n11061), .A2(n11047), .ZN(n11086) );
  INV_X1 U14084 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11719) );
  OAI22_X1 U14085 ( .A1(n11123), .A2(n11718), .B1(n11086), .B2(n11719), .ZN(
        n11053) );
  INV_X1 U14086 ( .A(n11048), .ZN(n11049) );
  NAND2_X1 U14087 ( .A1(n9593), .A2(n11049), .ZN(n11060) );
  INV_X1 U14088 ( .A(n11060), .ZN(n11050) );
  INV_X1 U14089 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11710) );
  OR2_X2 U14090 ( .A1(n9593), .A2(n11051), .ZN(n11054) );
  OAI22_X1 U14091 ( .A1(n11189), .A2(n10372), .B1(n11710), .B2(n19100), .ZN(
        n11052) );
  NOR2_X1 U14092 ( .A1(n11053), .A2(n11052), .ZN(n11067) );
  INV_X1 U14093 ( .A(n11054), .ZN(n11055) );
  INV_X1 U14094 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11058) );
  OR2_X1 U14095 ( .A1(n11061), .A2(n11056), .ZN(n11121) );
  INV_X1 U14096 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11057) );
  OAI22_X1 U14097 ( .A1(n11187), .A2(n11058), .B1(n11121), .B2(n11057), .ZN(
        n11065) );
  INV_X1 U14098 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11063) );
  OAI22_X1 U14099 ( .A1(n11063), .A2(n11122), .B1(n11124), .B2(n11062), .ZN(
        n11064) );
  NOR2_X1 U14100 ( .A1(n11065), .A2(n11064), .ZN(n11066) );
  AND4_X2 U14101 ( .A1(n11069), .A2(n11068), .A3(n11067), .A4(n11066), .ZN(
        n11082) );
  INV_X1 U14102 ( .A(n11519), .ZN(n11070) );
  NOR2_X2 U14103 ( .A1(n11072), .A2(n15388), .ZN(n11120) );
  NAND2_X1 U14104 ( .A1(n11120), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11074) );
  NOR2_X2 U14105 ( .A1(n11072), .A2(n11040), .ZN(n11117) );
  NAND2_X1 U14106 ( .A1(n11117), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11073) );
  NAND2_X1 U14107 ( .A1(n11074), .A2(n11073), .ZN(n11080) );
  AOI21_X1 U14108 ( .B1(n11119), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n16044), .ZN(n11078) );
  NOR2_X1 U14109 ( .A1(n11070), .A2(n15388), .ZN(n11075) );
  AND2_X2 U14110 ( .A1(n11076), .A2(n11075), .ZN(n19419) );
  NAND2_X1 U14111 ( .A1(n19419), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11077) );
  NAND2_X1 U14112 ( .A1(n11078), .A2(n11077), .ZN(n11079) );
  NOR2_X1 U14113 ( .A1(n11080), .A2(n11079), .ZN(n11081) );
  NAND2_X1 U14114 ( .A1(n11082), .A2(n11081), .ZN(n11085) );
  NAND2_X1 U14115 ( .A1(n11083), .A2(n16044), .ZN(n11084) );
  NAND2_X1 U14116 ( .A1(n11085), .A2(n11084), .ZN(n11154) );
  INV_X1 U14117 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11088) );
  INV_X1 U14118 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11664) );
  OAI211_X1 U14119 ( .C1(n11124), .C2(n11088), .A(n11087), .B(n19054), .ZN(
        n11089) );
  NAND2_X1 U14120 ( .A1(n11117), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11090) );
  INV_X1 U14121 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11092) );
  INV_X1 U14122 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11093) );
  NOR2_X1 U14123 ( .A1(n11122), .A2(n11093), .ZN(n11094) );
  NOR2_X1 U14124 ( .A1(n11095), .A2(n11094), .ZN(n11100) );
  INV_X1 U14125 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11663) );
  INV_X1 U14126 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11096) );
  NOR2_X1 U14127 ( .A1(n11121), .A2(n11096), .ZN(n11097) );
  NOR2_X1 U14128 ( .A1(n11098), .A2(n11097), .ZN(n11099) );
  NAND2_X1 U14129 ( .A1(n11100), .A2(n11099), .ZN(n11107) );
  INV_X1 U14130 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11102) );
  INV_X1 U14131 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11101) );
  INV_X1 U14132 ( .A(n11103), .ZN(n11105) );
  NAND2_X1 U14133 ( .A1(n11105), .A2(n11104), .ZN(n11106) );
  NOR2_X1 U14134 ( .A1(n11107), .A2(n11106), .ZN(n11110) );
  INV_X1 U14135 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11108) );
  NAND4_X1 U14136 ( .A1(n11111), .A2(n11110), .A3(n9625), .A4(n11109), .ZN(
        n11116) );
  OR2_X1 U14137 ( .A1(n13347), .A2(n19054), .ZN(n11457) );
  INV_X1 U14138 ( .A(n11457), .ZN(n11113) );
  NAND2_X1 U14139 ( .A1(n11113), .A2(n11112), .ZN(n11455) );
  INV_X1 U14140 ( .A(n11114), .ZN(n11456) );
  NAND2_X1 U14141 ( .A1(n11455), .A2(n11456), .ZN(n11115) );
  NAND2_X1 U14142 ( .A1(n11116), .A2(n11115), .ZN(n11155) );
  AOI22_X1 U14143 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n11118), .B1(
        n11119), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11147) );
  AOI22_X1 U14144 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19129), .B1(
        n19419), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11146) );
  INV_X1 U14145 ( .A(n11121), .ZN(n19241) );
  INV_X1 U14146 ( .A(n11187), .ZN(n19384) );
  AOI22_X1 U14147 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19241), .B1(
        n19384), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11133) );
  INV_X1 U14148 ( .A(n11122), .ZN(n19164) );
  INV_X1 U14149 ( .A(n11123), .ZN(n19448) );
  AOI22_X1 U14150 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19164), .B1(
        n19448), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11132) );
  INV_X1 U14151 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11126) );
  INV_X1 U14152 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11125) );
  OAI22_X1 U14153 ( .A1(n11126), .A2(n19100), .B1(n11124), .B2(n11125), .ZN(
        n11127) );
  INV_X1 U14154 ( .A(n11127), .ZN(n11131) );
  INV_X1 U14155 ( .A(n11086), .ZN(n11129) );
  INV_X1 U14156 ( .A(n11189), .ZN(n11128) );
  AOI22_X1 U14157 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n11129), .B1(
        n11128), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11130) );
  INV_X1 U14158 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11137) );
  INV_X1 U14159 ( .A(n19205), .ZN(n19197) );
  INV_X1 U14160 ( .A(n11134), .ZN(n11136) );
  INV_X1 U14161 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11135) );
  OAI22_X1 U14162 ( .A1(n11137), .A2(n19197), .B1(n11136), .B2(n11135), .ZN(
        n11143) );
  INV_X1 U14163 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13450) );
  INV_X1 U14164 ( .A(n15401), .ZN(n11141) );
  INV_X1 U14165 ( .A(n11138), .ZN(n11140) );
  INV_X1 U14166 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11139) );
  OAI22_X1 U14167 ( .A1(n13450), .A2(n11141), .B1(n11140), .B2(n11139), .ZN(
        n11142) );
  NOR2_X1 U14168 ( .A1(n11143), .A2(n11142), .ZN(n11144) );
  NAND4_X1 U14169 ( .A1(n11147), .A2(n11146), .A3(n11145), .A4(n11144), .ZN(
        n11150) );
  NAND2_X1 U14170 ( .A1(n11148), .A2(n16044), .ZN(n11149) );
  NAND2_X1 U14171 ( .A1(n11452), .A2(n14100), .ZN(n11153) );
  OAI21_X1 U14172 ( .B1(n11170), .B2(n11152), .A(n11151), .ZN(n13709) );
  INV_X1 U14173 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11453) );
  NAND2_X1 U14174 ( .A1(n11155), .A2(n11154), .ZN(n11156) );
  NAND2_X2 U14175 ( .A1(n11469), .A2(n11156), .ZN(n13654) );
  INV_X1 U14176 ( .A(n11157), .ZN(n11173) );
  NAND2_X1 U14177 ( .A1(n11158), .A2(n11165), .ZN(n11159) );
  NAND2_X1 U14178 ( .A1(n11173), .A2(n11159), .ZN(n13693) );
  OAI21_X1 U14179 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19797), .A(
        n11160), .ZN(n11360) );
  MUX2_X1 U14180 ( .A(n11360), .B(n13347), .S(n19800), .Z(n11342) );
  INV_X1 U14181 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n11161) );
  MUX2_X1 U14182 ( .A(n11342), .B(n11161), .S(n14096), .Z(n18872) );
  OR2_X1 U14183 ( .A1(n18872), .A2(n13351), .ZN(n13345) );
  INV_X1 U14184 ( .A(n11166), .ZN(n11163) );
  INV_X1 U14185 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13135) );
  NAND3_X1 U14186 ( .A1(n14096), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n11162) );
  NAND2_X1 U14187 ( .A1(n11163), .A2(n11162), .ZN(n13843) );
  NOR2_X1 U14188 ( .A1(n13345), .A2(n13843), .ZN(n11164) );
  NAND2_X1 U14189 ( .A1(n13345), .A2(n13843), .ZN(n13183) );
  OAI21_X1 U14190 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n11164), .A(
        n13183), .ZN(n13169) );
  OAI21_X1 U14191 ( .B1(n11167), .B2(n11166), .A(n11165), .ZN(n11168) );
  INV_X1 U14192 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13399) );
  XNOR2_X1 U14193 ( .A(n11168), .B(n13399), .ZN(n13168) );
  OR2_X1 U14194 ( .A1(n13169), .A2(n13168), .ZN(n13171) );
  INV_X1 U14195 ( .A(n11168), .ZN(n13737) );
  NAND2_X1 U14196 ( .A1(n13737), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11169) );
  AND2_X1 U14197 ( .A1(n13171), .A2(n11169), .ZN(n13641) );
  INV_X1 U14198 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13647) );
  INV_X1 U14199 ( .A(n11170), .ZN(n11175) );
  INV_X1 U14200 ( .A(n11171), .ZN(n11172) );
  NAND2_X1 U14201 ( .A1(n11173), .A2(n11172), .ZN(n11174) );
  NAND2_X1 U14202 ( .A1(n11175), .A2(n11174), .ZN(n14195) );
  INV_X1 U14203 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13860) );
  XNOR2_X1 U14204 ( .A(n14195), .B(n13860), .ZN(n13715) );
  NAND2_X1 U14205 ( .A1(n13852), .A2(n13853), .ZN(n11178) );
  NAND2_X1 U14206 ( .A1(n11176), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11177) );
  NAND2_X1 U14207 ( .A1(n11178), .A2(n11177), .ZN(n13940) );
  NAND2_X1 U14208 ( .A1(n19419), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11184) );
  NAND2_X1 U14209 ( .A1(n19129), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11183) );
  NAND2_X1 U14210 ( .A1(n11118), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11182) );
  NAND2_X1 U14211 ( .A1(n11119), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11181) );
  NAND4_X1 U14212 ( .A1(n11184), .A2(n11183), .A3(n11182), .A4(n11181), .ZN(
        n11204) );
  AOI22_X1 U14213 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n15401), .B1(
        n11138), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11202) );
  AOI22_X1 U14214 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19205), .B1(
        n11134), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11201) );
  INV_X1 U14215 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11186) );
  INV_X1 U14216 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11185) );
  OAI22_X1 U14217 ( .A1(n11186), .A2(n11124), .B1(n11121), .B2(n11185), .ZN(
        n11192) );
  INV_X1 U14218 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11190) );
  INV_X1 U14219 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11188) );
  OAI22_X1 U14220 ( .A1(n11190), .A2(n11187), .B1(n11189), .B2(n11188), .ZN(
        n11191) );
  NOR2_X1 U14221 ( .A1(n11192), .A2(n11191), .ZN(n11200) );
  INV_X1 U14222 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11194) );
  INV_X1 U14223 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11193) );
  OAI22_X1 U14224 ( .A1(n11194), .A2(n11123), .B1(n19100), .B2(n11193), .ZN(
        n11198) );
  INV_X1 U14225 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11196) );
  INV_X1 U14226 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11195) );
  OAI22_X1 U14227 ( .A1(n11196), .A2(n11122), .B1(n11086), .B2(n11195), .ZN(
        n11197) );
  NOR2_X1 U14228 ( .A1(n11198), .A2(n11197), .ZN(n11199) );
  NAND4_X1 U14229 ( .A1(n11202), .A2(n11201), .A3(n11200), .A4(n11199), .ZN(
        n11203) );
  INV_X1 U14230 ( .A(n11205), .ZN(n11206) );
  NAND2_X1 U14231 ( .A1(n11206), .A2(n16044), .ZN(n11207) );
  NAND2_X1 U14232 ( .A1(n11471), .A2(n14100), .ZN(n11210) );
  INV_X1 U14233 ( .A(n11209), .ZN(n11217) );
  XNOR2_X1 U14234 ( .A(n11151), .B(n11217), .ZN(n13748) );
  NAND2_X1 U14235 ( .A1(n11210), .A2(n13748), .ZN(n11211) );
  INV_X1 U14236 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13949) );
  XNOR2_X1 U14237 ( .A(n11211), .B(n13949), .ZN(n13939) );
  NAND2_X1 U14238 ( .A1(n13940), .A2(n13939), .ZN(n11213) );
  NAND2_X1 U14239 ( .A1(n11211), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11212) );
  NAND2_X1 U14240 ( .A1(n11213), .A2(n11212), .ZN(n15076) );
  OR2_X1 U14241 ( .A1(n11215), .A2(n11214), .ZN(n11216) );
  NAND2_X1 U14242 ( .A1(n11231), .A2(n11216), .ZN(n13778) );
  OR2_X1 U14243 ( .A1(n13778), .A2(n14100), .ZN(n11228) );
  INV_X1 U14244 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11486) );
  NOR2_X1 U14245 ( .A1(n11228), .A2(n11486), .ZN(n15989) );
  INV_X1 U14246 ( .A(n15989), .ZN(n11222) );
  NOR2_X1 U14247 ( .A1(n11151), .A2(n11217), .ZN(n11220) );
  INV_X1 U14248 ( .A(n11218), .ZN(n11219) );
  XNOR2_X1 U14249 ( .A(n11220), .B(n11219), .ZN(n11229) );
  AND2_X1 U14250 ( .A1(n11229), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15985) );
  NAND3_X1 U14251 ( .A1(n11225), .A2(n14096), .A3(P2_EBX_REG_10__SCAN_IN), 
        .ZN(n11224) );
  OAI211_X1 U14252 ( .C1(n11225), .C2(P2_EBX_REG_10__SCAN_IN), .A(n14098), .B(
        n11224), .ZN(n13796) );
  OR2_X1 U14253 ( .A1(n13796), .A2(n14100), .ZN(n11227) );
  INV_X1 U14254 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11226) );
  NAND2_X1 U14255 ( .A1(n11227), .A2(n11226), .ZN(n15307) );
  NAND2_X1 U14256 ( .A1(n11228), .A2(n11486), .ZN(n15987) );
  INV_X1 U14257 ( .A(n11229), .ZN(n18855) );
  NAND2_X1 U14258 ( .A1(n18855), .A2(n15342), .ZN(n15986) );
  AND2_X1 U14259 ( .A1(n15987), .A2(n15986), .ZN(n15284) );
  NAND2_X1 U14260 ( .A1(n14096), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11230) );
  XNOR2_X1 U14261 ( .A(n11231), .B(n11230), .ZN(n18839) );
  NAND2_X1 U14262 ( .A1(n18839), .A2(n14094), .ZN(n11239) );
  INV_X1 U14263 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15329) );
  NAND2_X1 U14264 ( .A1(n11239), .A2(n15329), .ZN(n15321) );
  INV_X1 U14265 ( .A(n11232), .ZN(n11233) );
  NAND2_X1 U14266 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n11233), .ZN(n11234) );
  NOR2_X1 U14267 ( .A1(n19070), .A2(n11234), .ZN(n11235) );
  OR2_X1 U14268 ( .A1(n11236), .A2(n11235), .ZN(n18826) );
  OR2_X1 U14269 ( .A1(n18826), .A2(n14100), .ZN(n11237) );
  INV_X1 U14270 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15295) );
  NAND2_X1 U14271 ( .A1(n11237), .A2(n15295), .ZN(n15289) );
  NAND2_X1 U14272 ( .A1(n14094), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11238) );
  OR2_X1 U14273 ( .A1(n13796), .A2(n11238), .ZN(n15306) );
  OR2_X1 U14274 ( .A1(n11239), .A2(n15329), .ZN(n15322) );
  AND2_X1 U14275 ( .A1(n15306), .A2(n15322), .ZN(n15286) );
  NAND2_X1 U14276 ( .A1(n14094), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11240) );
  OR2_X1 U14277 ( .A1(n18826), .A2(n11240), .ZN(n15288) );
  NAND2_X1 U14278 ( .A1(n15286), .A2(n15288), .ZN(n11241) );
  INV_X1 U14279 ( .A(n11243), .ZN(n11245) );
  NAND2_X1 U14280 ( .A1(n11245), .A2(n11244), .ZN(n11246) );
  NAND2_X1 U14281 ( .A1(n11265), .A2(n11246), .ZN(n18809) );
  OR2_X1 U14282 ( .A1(n18809), .A2(n14100), .ZN(n11248) );
  INV_X1 U14283 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11247) );
  OR2_X1 U14284 ( .A1(n11248), .A2(n11247), .ZN(n15276) );
  NOR2_X2 U14285 ( .A1(n11249), .A2(n9988), .ZN(n18756) );
  NAND2_X1 U14286 ( .A1(n18756), .A2(n14094), .ZN(n11251) );
  INV_X1 U14287 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15200) );
  NAND2_X1 U14288 ( .A1(n11251), .A2(n15200), .ZN(n15039) );
  NAND2_X1 U14289 ( .A1(n11261), .A2(n11252), .ZN(n11253) );
  NAND2_X1 U14290 ( .A1(n11254), .A2(n11253), .ZN(n11284) );
  INV_X1 U14291 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15207) );
  OAI21_X1 U14292 ( .B1(n11284), .B2(n14100), .A(n15207), .ZN(n15050) );
  NAND2_X1 U14293 ( .A1(n15039), .A2(n15050), .ZN(n15013) );
  INV_X1 U14294 ( .A(n11255), .ZN(n11256) );
  XNOR2_X1 U14295 ( .A(n11257), .B(n11256), .ZN(n11289) );
  AOI21_X1 U14296 ( .B1(n11289), .B2(n14094), .A(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15247) );
  NAND2_X1 U14297 ( .A1(n11259), .A2(n11258), .ZN(n11260) );
  AND2_X1 U14298 ( .A1(n11261), .A2(n11260), .ZN(n18787) );
  AOI21_X1 U14299 ( .B1(n18787), .B2(n14094), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15009) );
  INV_X1 U14300 ( .A(n11262), .ZN(n11263) );
  XNOR2_X1 U14301 ( .A(n11267), .B(n11263), .ZN(n13797) );
  NAND2_X1 U14302 ( .A1(n13797), .A2(n14094), .ZN(n11287) );
  NAND2_X1 U14303 ( .A1(n11287), .A2(n15935), .ZN(n15940) );
  NAND2_X1 U14304 ( .A1(n11265), .A2(n11264), .ZN(n11266) );
  NAND2_X1 U14305 ( .A1(n11267), .A2(n11266), .ZN(n13828) );
  OR2_X1 U14306 ( .A1(n13828), .A2(n14100), .ZN(n11269) );
  INV_X1 U14307 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11268) );
  NAND2_X1 U14308 ( .A1(n11269), .A2(n11268), .ZN(n15937) );
  NAND2_X1 U14309 ( .A1(n15940), .A2(n15937), .ZN(n15004) );
  NOR2_X1 U14310 ( .A1(n19070), .A2(n11270), .ZN(n11271) );
  AND2_X1 U14311 ( .A1(n9599), .A2(n11271), .ZN(n11272) );
  NOR2_X1 U14312 ( .A1(n11273), .A2(n11272), .ZN(n14766) );
  NAND2_X1 U14313 ( .A1(n14766), .A2(n14094), .ZN(n11274) );
  NAND2_X1 U14314 ( .A1(n11274), .A2(n15168), .ZN(n15001) );
  INV_X1 U14315 ( .A(n11275), .ZN(n11277) );
  MUX2_X1 U14316 ( .A(P2_EBX_REG_16__SCAN_IN), .B(n11277), .S(n11276), .Z(
        n11278) );
  NAND2_X1 U14317 ( .A1(n11278), .A2(n14098), .ZN(n13938) );
  OR2_X1 U14318 ( .A1(n13938), .A2(n14100), .ZN(n11286) );
  XNOR2_X1 U14319 ( .A(n11286), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15007) );
  NOR2_X1 U14320 ( .A1(n19070), .A2(n14771), .ZN(n11279) );
  XNOR2_X1 U14321 ( .A(n11249), .B(n11279), .ZN(n14784) );
  NAND2_X1 U14322 ( .A1(n14784), .A2(n14094), .ZN(n11294) );
  INV_X1 U14323 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15188) );
  NAND2_X1 U14324 ( .A1(n11294), .A2(n15188), .ZN(n15029) );
  AND4_X1 U14325 ( .A1(n11280), .A2(n15001), .A3(n15007), .A4(n15029), .ZN(
        n11297) );
  AND2_X1 U14326 ( .A1(n14094), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11281) );
  NAND2_X1 U14327 ( .A1(n14766), .A2(n11281), .ZN(n15000) );
  INV_X1 U14328 ( .A(n18756), .ZN(n11283) );
  NAND2_X1 U14329 ( .A1(n14094), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11282) );
  OR2_X1 U14330 ( .A1(n11283), .A2(n11282), .ZN(n15038) );
  INV_X1 U14331 ( .A(n11284), .ZN(n18769) );
  AND2_X1 U14332 ( .A1(n14094), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11285) );
  NAND2_X1 U14333 ( .A1(n18769), .A2(n11285), .ZN(n15049) );
  NAND2_X1 U14334 ( .A1(n15038), .A2(n15049), .ZN(n15012) );
  INV_X1 U14335 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15239) );
  OR2_X1 U14336 ( .A1(n11286), .A2(n15239), .ZN(n15008) );
  OR2_X1 U14337 ( .A1(n11287), .A2(n15935), .ZN(n15941) );
  NAND2_X1 U14338 ( .A1(n14094), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11288) );
  OR2_X1 U14339 ( .A1(n13828), .A2(n11288), .ZN(n15003) );
  AND2_X1 U14340 ( .A1(n15941), .A2(n15003), .ZN(n11292) );
  INV_X1 U14341 ( .A(n11289), .ZN(n18802) );
  INV_X1 U14342 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15252) );
  OR3_X1 U14343 ( .A1(n18802), .A2(n14100), .A3(n15252), .ZN(n15005) );
  INV_X1 U14344 ( .A(n18787), .ZN(n11291) );
  NAND2_X1 U14345 ( .A1(n14094), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11290) );
  OR2_X1 U14346 ( .A1(n11291), .A2(n11290), .ZN(n15010) );
  NAND4_X1 U14347 ( .A1(n15008), .A2(n11292), .A3(n15005), .A4(n15010), .ZN(
        n11293) );
  NOR2_X1 U14348 ( .A1(n15012), .A2(n11293), .ZN(n11295) );
  OR2_X1 U14349 ( .A1(n11294), .A2(n15188), .ZN(n15031) );
  NAND3_X1 U14350 ( .A1(n15000), .A2(n11295), .A3(n15031), .ZN(n11296) );
  NAND2_X1 U14351 ( .A1(n11299), .A2(n9915), .ZN(n11300) );
  AND2_X1 U14352 ( .A1(n11304), .A2(n11300), .ZN(n14742) );
  NAND2_X1 U14353 ( .A1(n14742), .A2(n14094), .ZN(n11301) );
  INV_X1 U14354 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15162) );
  AND2_X1 U14355 ( .A1(n11301), .A2(n15162), .ZN(n15150) );
  INV_X1 U14356 ( .A(n11301), .ZN(n11302) );
  NAND2_X1 U14357 ( .A1(n11302), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15151) );
  AND2_X1 U14358 ( .A1(n11304), .A2(n11303), .ZN(n11305) );
  NOR2_X1 U14359 ( .A1(n14741), .A2(n14100), .ZN(n11306) );
  INV_X1 U14360 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15139) );
  XNOR2_X1 U14361 ( .A(n11306), .B(n15139), .ZN(n14991) );
  NOR2_X1 U14362 ( .A1(n14100), .A2(n15139), .ZN(n11308) );
  INV_X1 U14363 ( .A(n14741), .ZN(n11307) );
  NAND2_X1 U14364 ( .A1(n14096), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11310) );
  MUX2_X1 U14365 ( .A(n11310), .B(P2_EBX_REG_24__SCAN_IN), .S(n11309), .Z(
        n11311) );
  NAND2_X1 U14366 ( .A1(n11311), .A2(n14098), .ZN(n15869) );
  NOR2_X1 U14367 ( .A1(n15869), .A2(n14100), .ZN(n14978) );
  NOR2_X1 U14368 ( .A1(n11316), .A2(n14821), .ZN(n11313) );
  NAND2_X1 U14369 ( .A1(n14096), .A2(n11313), .ZN(n11314) );
  NAND2_X1 U14370 ( .A1(n14098), .A2(n11314), .ZN(n11315) );
  AOI21_X1 U14371 ( .B1(n11316), .B2(n14821), .A(n11315), .ZN(n15857) );
  AOI21_X1 U14372 ( .B1(n15857), .B2(n14094), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14969) );
  NAND2_X1 U14373 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n9619), .ZN(n11317) );
  NOR2_X1 U14374 ( .A1(n19070), .A2(n11317), .ZN(n11318) );
  OR2_X1 U14375 ( .A1(n11319), .A2(n11318), .ZN(n15845) );
  XNOR2_X1 U14376 ( .A(n11332), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14960) );
  INV_X1 U14377 ( .A(n11320), .ZN(n11322) );
  NAND2_X1 U14378 ( .A1(n11322), .A2(n11321), .ZN(n11323) );
  NAND2_X1 U14379 ( .A1(n11328), .A2(n11323), .ZN(n15832) );
  INV_X1 U14380 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11324) );
  NAND2_X1 U14381 ( .A1(n11328), .A2(n11327), .ZN(n11329) );
  AND2_X1 U14382 ( .A1(n11335), .A2(n11329), .ZN(n14729) );
  NAND2_X1 U14383 ( .A1(n14729), .A2(n14094), .ZN(n14938) );
  INV_X1 U14384 ( .A(n14938), .ZN(n11330) );
  INV_X1 U14385 ( .A(n11332), .ZN(n11334) );
  INV_X1 U14386 ( .A(n15857), .ZN(n11333) );
  INV_X1 U14387 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15115) );
  AOI21_X1 U14388 ( .B1(n11334), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n14968), .ZN(n14933) );
  INV_X1 U14389 ( .A(n11335), .ZN(n11337) );
  XNOR2_X1 U14390 ( .A(n11337), .B(n11336), .ZN(n11338) );
  INV_X1 U14391 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11494) );
  OAI21_X1 U14392 ( .B1(n11338), .B2(n14100), .A(n11494), .ZN(n14092) );
  INV_X1 U14393 ( .A(n11338), .ZN(n15820) );
  NAND3_X1 U14394 ( .A1(n15820), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14094), .ZN(n14136) );
  INV_X1 U14395 ( .A(n11359), .ZN(n11341) );
  INV_X1 U14396 ( .A(n11339), .ZN(n11340) );
  OAI21_X1 U14397 ( .B1(n11342), .B2(n11341), .A(n11340), .ZN(n11346) );
  NAND2_X1 U14398 ( .A1(n11344), .A2(n11343), .ZN(n11355) );
  INV_X1 U14399 ( .A(n11355), .ZN(n11345) );
  NAND2_X1 U14400 ( .A1(n11346), .A2(n11345), .ZN(n11347) );
  NAND2_X1 U14401 ( .A1(n11347), .A2(n11375), .ZN(n19802) );
  INV_X1 U14402 ( .A(n19801), .ZN(n13100) );
  OAI21_X1 U14403 ( .B1(n11360), .B2(n11348), .A(n11383), .ZN(n11349) );
  INV_X1 U14404 ( .A(n11349), .ZN(n11351) );
  OR2_X1 U14405 ( .A1(n13356), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n16043) );
  INV_X1 U14406 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n11350) );
  OAI21_X1 U14407 ( .B1(n10369), .B2(n16043), .A(n11350), .ZN(n19789) );
  MUX2_X1 U14408 ( .A(n11351), .B(n19789), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n16063) );
  INV_X1 U14409 ( .A(n16063), .ZN(n19799) );
  OAI22_X1 U14410 ( .A1(n19802), .A2(n13100), .B1(n16044), .B2(n19799), .ZN(
        n11354) );
  INV_X1 U14411 ( .A(n19805), .ZN(n11353) );
  NAND2_X1 U14412 ( .A1(n11354), .A2(n11353), .ZN(n13099) );
  NAND2_X1 U14413 ( .A1(n11355), .A2(n11399), .ZN(n11372) );
  AOI21_X1 U14414 ( .B1(n13104), .B2(n19054), .A(n11356), .ZN(n11367) );
  INV_X1 U14415 ( .A(n11356), .ZN(n11363) );
  INV_X1 U14416 ( .A(n11360), .ZN(n11358) );
  OAI211_X1 U14417 ( .C1(n19054), .C2(n11358), .A(n16045), .B(n11357), .ZN(
        n11362) );
  OAI21_X1 U14418 ( .B1(n11360), .B2(n11341), .A(n19800), .ZN(n11361) );
  OAI211_X1 U14419 ( .C1(n11364), .C2(n11363), .A(n11362), .B(n11361), .ZN(
        n11365) );
  OAI21_X1 U14420 ( .B1(n11367), .B2(n11366), .A(n11365), .ZN(n11370) );
  NAND3_X1 U14421 ( .A1(n11370), .A2(n11369), .A3(n11368), .ZN(n11371) );
  NAND2_X1 U14422 ( .A1(n11372), .A2(n11371), .ZN(n11374) );
  AND2_X1 U14423 ( .A1(n11375), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11373) );
  NAND2_X1 U14424 ( .A1(n11374), .A2(n11373), .ZN(n11379) );
  INV_X1 U14425 ( .A(n11375), .ZN(n11378) );
  NOR2_X1 U14426 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n11376) );
  AOI21_X1 U14427 ( .B1(n11378), .B2(n11377), .A(n11376), .ZN(n13159) );
  NAND2_X1 U14428 ( .A1(n11379), .A2(n13159), .ZN(n16041) );
  NAND2_X1 U14429 ( .A1(n16041), .A2(n19054), .ZN(n13372) );
  NAND2_X1 U14430 ( .A1(n19060), .A2(n11380), .ZN(n11395) );
  OAI211_X1 U14431 ( .C1(n19048), .C2(n16041), .A(n13372), .B(n9590), .ZN(
        n11394) );
  NAND2_X1 U14432 ( .A1(n11381), .A2(n9588), .ZN(n13373) );
  NAND2_X1 U14433 ( .A1(n16047), .A2(n13373), .ZN(n11392) );
  MUX2_X1 U14434 ( .A(n10538), .B(n19060), .S(n16044), .Z(n11382) );
  NAND3_X1 U14435 ( .A1(n11382), .A2(n11383), .A3(n19669), .ZN(n11391) );
  INV_X1 U14436 ( .A(n11383), .ZN(n16035) );
  NOR2_X1 U14437 ( .A1(n16035), .A2(n13371), .ZN(n11384) );
  NAND2_X1 U14438 ( .A1(n10538), .A2(n11384), .ZN(n11390) );
  NAND2_X1 U14439 ( .A1(n11385), .A2(n19085), .ZN(n11386) );
  NAND2_X1 U14440 ( .A1(n11386), .A2(n19801), .ZN(n11414) );
  OAI22_X1 U14441 ( .A1(n19054), .A2(n10513), .B1(n9868), .B2(n16045), .ZN(
        n11387) );
  NAND2_X1 U14442 ( .A1(n11387), .A2(n19065), .ZN(n11388) );
  NAND2_X1 U14443 ( .A1(n11388), .A2(n9588), .ZN(n11389) );
  AND3_X1 U14444 ( .A1(n11390), .A2(n11414), .A3(n11389), .ZN(n13366) );
  AND3_X1 U14445 ( .A1(n11392), .A2(n11391), .A3(n13366), .ZN(n11393) );
  OAI211_X1 U14446 ( .C1(n13372), .C2(n11395), .A(n11394), .B(n11393), .ZN(
        n11396) );
  INV_X1 U14447 ( .A(n11396), .ZN(n11397) );
  NAND2_X1 U14448 ( .A1(n13099), .A2(n11397), .ZN(n11398) );
  OR3_X1 U14449 ( .A1(n11495), .A2(n19805), .A3(n11399), .ZN(n15234) );
  NAND2_X1 U14450 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15265) );
  INV_X1 U14451 ( .A(n15265), .ZN(n15294) );
  NAND2_X1 U14452 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15294), .ZN(
        n15227) );
  NOR2_X1 U14453 ( .A1(n11268), .A2(n11247), .ZN(n16004) );
  NAND2_X1 U14454 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16004), .ZN(
        n16002) );
  NOR2_X1 U14455 ( .A1(n15227), .A2(n16002), .ZN(n15222) );
  NAND4_X1 U14456 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n15222), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15212) );
  NOR2_X1 U14457 ( .A1(n15207), .A2(n15212), .ZN(n15185) );
  AND3_X1 U14458 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(n15185), .ZN(n15017) );
  NOR2_X1 U14459 ( .A1(n11453), .A2(n13860), .ZN(n13859) );
  INV_X1 U14460 ( .A(n13859), .ZN(n11422) );
  NAND2_X1 U14461 ( .A1(n11401), .A2(n11400), .ZN(n15356) );
  NAND3_X1 U14462 ( .A1(n16044), .A2(n9588), .A3(n19070), .ZN(n11402) );
  NOR2_X1 U14463 ( .A1(n15356), .A2(n11402), .ZN(n11819) );
  INV_X1 U14464 ( .A(n11819), .ZN(n16042) );
  NAND2_X1 U14465 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13398) );
  NOR2_X1 U14466 ( .A1(n13399), .A2(n13398), .ZN(n11427) );
  INV_X1 U14467 ( .A(n11427), .ZN(n11421) );
  NAND2_X1 U14468 ( .A1(n13399), .A2(n13398), .ZN(n11426) );
  INV_X1 U14469 ( .A(n11426), .ZN(n11420) );
  MUX2_X1 U14470 ( .A(n11403), .B(n9588), .S(n19048), .Z(n11418) );
  INV_X1 U14471 ( .A(n11404), .ZN(n11411) );
  OAI21_X1 U14472 ( .B1(n10511), .B2(n11405), .A(n11411), .ZN(n11407) );
  NAND2_X1 U14473 ( .A1(n11407), .A2(n11406), .ZN(n11410) );
  INV_X1 U14474 ( .A(n11822), .ZN(n11409) );
  OAI211_X1 U14475 ( .C1(n10221), .C2(n11411), .A(n11410), .B(n11409), .ZN(
        n11412) );
  INV_X1 U14476 ( .A(n11412), .ZN(n11417) );
  NAND2_X1 U14477 ( .A1(n11413), .A2(n19054), .ZN(n15357) );
  NAND2_X1 U14478 ( .A1(n15357), .A2(n11414), .ZN(n11415) );
  NAND2_X1 U14479 ( .A1(n11415), .A2(n19065), .ZN(n11416) );
  AOI211_X1 U14480 ( .C1(n15223), .C2(n11421), .A(n11420), .B(n15225), .ZN(
        n13648) );
  NAND2_X1 U14481 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13648), .ZN(
        n13858) );
  NOR2_X1 U14482 ( .A1(n11422), .A2(n13858), .ZN(n13950) );
  NAND2_X1 U14483 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13950), .ZN(
        n11425) );
  INV_X1 U14484 ( .A(n11425), .ZN(n16009) );
  NAND3_X1 U14485 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n16009), .ZN(n15226) );
  NAND2_X1 U14486 ( .A1(n15017), .A2(n15330), .ZN(n15171) );
  NOR2_X1 U14487 ( .A1(n15168), .A2(n15171), .ZN(n15140) );
  AND2_X1 U14488 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11432) );
  INV_X1 U14489 ( .A(n11432), .ZN(n15128) );
  NOR2_X1 U14490 ( .A1(n15128), .A2(n11312), .ZN(n11423) );
  NAND2_X1 U14491 ( .A1(n15140), .A2(n11423), .ZN(n15121) );
  AND2_X1 U14492 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11434) );
  INV_X1 U14493 ( .A(n11434), .ZN(n11424) );
  NOR2_X1 U14494 ( .A1(n15121), .A2(n11424), .ZN(n15081) );
  INV_X1 U14495 ( .A(n15081), .ZN(n15099) );
  AND2_X1 U14496 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14119) );
  AOI21_X1 U14497 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n11425), .ZN(n11430) );
  OR2_X1 U14498 ( .A1(n15223), .A2(n11426), .ZN(n13404) );
  OR2_X1 U14499 ( .A1(n15221), .A2(n11427), .ZN(n11428) );
  NAND2_X1 U14500 ( .A1(n11495), .A2(n18765), .ZN(n13396) );
  AND3_X1 U14501 ( .A1(n13404), .A2(n11428), .A3(n13396), .ZN(n13646) );
  OR2_X1 U14502 ( .A1(n15225), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11429) );
  AND2_X1 U14503 ( .A1(n13646), .A2(n11429), .ZN(n13862) );
  OAI221_X1 U14504 ( .B1(n15225), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(
        n15225), .C2(n13859), .A(n13862), .ZN(n15345) );
  NOR2_X1 U14505 ( .A1(n11430), .A2(n15345), .ZN(n16020) );
  NAND2_X1 U14506 ( .A1(n15017), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11491) );
  INV_X1 U14507 ( .A(n11491), .ZN(n15018) );
  AND2_X1 U14508 ( .A1(n16020), .A2(n15018), .ZN(n11431) );
  OR2_X1 U14509 ( .A1(n15293), .A2(n11431), .ZN(n15169) );
  OAI211_X1 U14510 ( .C1(n15293), .C2(n11432), .A(n15169), .B(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15133) );
  INV_X1 U14511 ( .A(n15293), .ZN(n11433) );
  NAND2_X1 U14512 ( .A1(n15133), .A2(n11433), .ZN(n15116) );
  OAI21_X1 U14513 ( .B1(n15293), .B2(n11434), .A(n15116), .ZN(n15101) );
  INV_X1 U14514 ( .A(n15101), .ZN(n11435) );
  OAI21_X1 U14515 ( .B1(n15099), .B2(n14119), .A(n11435), .ZN(n15091) );
  AOI21_X1 U14516 ( .B1(n16044), .B2(n15379), .A(n11438), .ZN(n11439) );
  NAND2_X1 U14517 ( .A1(n19038), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n14924) );
  INV_X1 U14518 ( .A(n11440), .ZN(n11442) );
  INV_X1 U14519 ( .A(n15356), .ZN(n11441) );
  NAND2_X1 U14520 ( .A1(n11442), .A2(n11441), .ZN(n16037) );
  NAND2_X1 U14521 ( .A1(n16036), .A2(n19054), .ZN(n11443) );
  AND2_X1 U14522 ( .A1(n16037), .A2(n11443), .ZN(n11444) );
  INV_X1 U14523 ( .A(n15348), .ZN(n16010) );
  INV_X1 U14524 ( .A(n11445), .ZN(n14724) );
  INV_X1 U14525 ( .A(n11446), .ZN(n11447) );
  AND2_X1 U14526 ( .A1(n14724), .A2(n11447), .ZN(n11448) );
  NOR2_X1 U14527 ( .A1(n10476), .A2(n11448), .ZN(n15822) );
  NAND2_X1 U14528 ( .A1(n16010), .A2(n15822), .ZN(n11449) );
  OAI211_X1 U14529 ( .C1(n15821), .C2(n15343), .A(n14924), .B(n11449), .ZN(
        n11451) );
  NOR3_X1 U14530 ( .A1(n15099), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n9950), .ZN(n11450) );
  AOI211_X1 U14531 ( .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15091), .A(
        n11451), .B(n11450), .ZN(n11497) );
  INV_X1 U14532 ( .A(n11452), .ZN(n11454) );
  INV_X1 U14533 ( .A(n13654), .ZN(n11464) );
  XOR2_X1 U14534 ( .A(n11456), .B(n11455), .Z(n13167) );
  NAND2_X1 U14535 ( .A1(n11457), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13346) );
  XNOR2_X1 U14536 ( .A(n13347), .B(n11458), .ZN(n11459) );
  NOR2_X1 U14537 ( .A1(n13346), .A2(n11459), .ZN(n11460) );
  XNOR2_X1 U14538 ( .A(n13346), .B(n11459), .ZN(n13181) );
  NOR2_X1 U14539 ( .A1(n15366), .A2(n13181), .ZN(n13180) );
  NOR2_X1 U14540 ( .A1(n11460), .A2(n13180), .ZN(n11461) );
  XOR2_X1 U14541 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11461), .Z(
        n13166) );
  NOR2_X1 U14542 ( .A1(n13167), .A2(n13166), .ZN(n13165) );
  NOR2_X1 U14543 ( .A1(n11461), .A2(n13399), .ZN(n11462) );
  OR2_X1 U14544 ( .A1(n13165), .A2(n11462), .ZN(n11465) );
  XNOR2_X1 U14545 ( .A(n11465), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13653) );
  INV_X1 U14546 ( .A(n13653), .ZN(n11463) );
  NAND2_X1 U14547 ( .A1(n11465), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11466) );
  NAND2_X1 U14548 ( .A1(n11469), .A2(n11468), .ZN(n11470) );
  NAND2_X1 U14549 ( .A1(n11467), .A2(n11470), .ZN(n13716) );
  NAND2_X1 U14550 ( .A1(n11475), .A2(n13855), .ZN(n11479) );
  INV_X1 U14551 ( .A(n11471), .ZN(n11478) );
  INV_X1 U14552 ( .A(n13855), .ZN(n11473) );
  NAND2_X1 U14553 ( .A1(n11473), .A2(n11483), .ZN(n11474) );
  INV_X1 U14554 ( .A(n11475), .ZN(n11476) );
  NAND2_X1 U14555 ( .A1(n11476), .A2(n11478), .ZN(n11477) );
  NAND2_X1 U14556 ( .A1(n13941), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11481) );
  NAND2_X1 U14557 ( .A1(n11479), .A2(n11471), .ZN(n11480) );
  XNOR2_X1 U14558 ( .A(n11488), .B(n14094), .ZN(n15075) );
  NAND2_X1 U14559 ( .A1(n11484), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11485) );
  NOR2_X1 U14560 ( .A1(n11488), .A2(n14100), .ZN(n11487) );
  XNOR2_X1 U14561 ( .A(n11487), .B(n11486), .ZN(n15993) );
  INV_X1 U14562 ( .A(n11488), .ZN(n11489) );
  NAND3_X1 U14563 ( .A1(n11489), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n14094), .ZN(n11490) );
  NOR2_X1 U14564 ( .A1(n11491), .A2(n15162), .ZN(n11492) );
  NAND2_X1 U14565 ( .A1(n11493), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14983) );
  AOI21_X1 U14566 ( .B1(n11494), .B2(n14943), .A(n14143), .ZN(n14930) );
  OR3_X1 U14567 ( .A1(n11495), .A2(n19805), .A3(n13100), .ZN(n15352) );
  NAND2_X1 U14568 ( .A1(n14930), .A2(n16011), .ZN(n11496) );
  OAI211_X1 U14569 ( .C1(n14932), .C2(n15234), .A(n11497), .B(n11496), .ZN(
        P2_U3017) );
  AND2_X1 U14570 ( .A1(n16078), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n11520) );
  NAND2_X1 U14571 ( .A1(n9589), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11499) );
  NAND2_X1 U14572 ( .A1(n11499), .A2(n19611), .ZN(n11521) );
  NOR2_X1 U14573 ( .A1(n19779), .A2(n19788), .ZN(n15398) );
  NAND2_X1 U14574 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15398), .ZN(
        n11508) );
  NAND2_X1 U14575 ( .A1(n11508), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11501) );
  INV_X1 U14576 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19769) );
  NAND2_X1 U14577 ( .A1(n19769), .A2(n15398), .ZN(n19309) );
  INV_X1 U14578 ( .A(n19309), .ZN(n11500) );
  NAND2_X1 U14579 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11500), .ZN(
        n19340) );
  NAND2_X1 U14580 ( .A1(n11501), .A2(n19340), .ZN(n19478) );
  AOI22_X1 U14581 ( .A1(n11521), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n19759), .B2(n19478), .ZN(n11502) );
  NAND3_X1 U14582 ( .A1(n13192), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n19054), 
        .ZN(n11536) );
  INV_X1 U14583 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19069) );
  NOR2_X1 U14584 ( .A1(n11536), .A2(n19069), .ZN(n11504) );
  OR2_X1 U14585 ( .A1(n11505), .A2(n11504), .ZN(n11506) );
  NAND2_X1 U14586 ( .A1(n11505), .A2(n11504), .ZN(n11530) );
  NAND2_X1 U14587 ( .A1(n9592), .A2(n11520), .ZN(n11511) );
  NAND2_X1 U14588 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19157) );
  NAND2_X1 U14589 ( .A1(n19157), .A2(n19779), .ZN(n11509) );
  AND2_X1 U14590 ( .A1(n11509), .A2(n11508), .ZN(n19200) );
  AOI22_X1 U14591 ( .A1(n11521), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19759), .B2(n19200), .ZN(n11510) );
  INV_X1 U14592 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11512) );
  NOR2_X1 U14593 ( .A1(n11536), .A2(n11512), .ZN(n11513) );
  NAND2_X1 U14594 ( .A1(n11521), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11517) );
  NAND2_X1 U14595 ( .A1(n19788), .A2(n19797), .ZN(n19336) );
  NAND2_X1 U14596 ( .A1(n19157), .A2(n19336), .ZN(n19199) );
  INV_X1 U14597 ( .A(n19199), .ZN(n11516) );
  NAND2_X1 U14598 ( .A1(n11516), .A2(n19759), .ZN(n19418) );
  NAND2_X1 U14599 ( .A1(n11517), .A2(n19418), .ZN(n11518) );
  INV_X1 U14600 ( .A(n11520), .ZN(n13177) );
  AOI22_X1 U14601 ( .A1(n11521), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19759), .B2(n19797), .ZN(n11522) );
  OAI21_X2 U14602 ( .B1(n15355), .B2(n13177), .A(n11522), .ZN(n15363) );
  INV_X1 U14603 ( .A(n11536), .ZN(n11761) );
  NAND2_X1 U14604 ( .A1(n11761), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11523) );
  NAND2_X1 U14605 ( .A1(n13132), .A2(n13131), .ZN(n11526) );
  INV_X1 U14606 ( .A(n15363), .ZN(n11524) );
  NAND2_X1 U14607 ( .A1(n11524), .A2(n11523), .ZN(n11525) );
  NAND2_X1 U14608 ( .A1(n11526), .A2(n11525), .ZN(n13301) );
  NAND2_X1 U14609 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n9589), .ZN(
        n11529) );
  AND2_X1 U14610 ( .A1(n18897), .A2(n18896), .ZN(n11539) );
  INV_X1 U14611 ( .A(n18905), .ZN(n11538) );
  INV_X1 U14612 ( .A(n11532), .ZN(n13413) );
  INV_X1 U14613 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11533) );
  NAND2_X1 U14614 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13451) );
  NOR2_X1 U14615 ( .A1(n11533), .A2(n13451), .ZN(n18910) );
  AND2_X1 U14616 ( .A1(n11534), .A2(n18910), .ZN(n11537) );
  INV_X1 U14617 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11535) );
  NOR2_X1 U14618 ( .A1(n11536), .A2(n11535), .ZN(n18909) );
  AND2_X1 U14619 ( .A1(n11537), .A2(n18909), .ZN(n13411) );
  AND2_X1 U14620 ( .A1(n13413), .A2(n13411), .ZN(n13412) );
  AND2_X1 U14621 ( .A1(n11538), .A2(n13412), .ZN(n13523) );
  AND2_X1 U14622 ( .A1(n11539), .A2(n13523), .ZN(n18895) );
  AOI22_X1 U14623 ( .A1(n10272), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11595), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11546) );
  AOI22_X1 U14624 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11545) );
  AOI22_X1 U14625 ( .A1(n11637), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11544) );
  AOI22_X1 U14626 ( .A1(n11640), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11543) );
  NAND4_X1 U14627 ( .A1(n11546), .A2(n11545), .A3(n11544), .A4(n11543), .ZN(
        n11553) );
  AOI22_X1 U14628 ( .A1(n10165), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10279), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U14629 ( .A1(n11547), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10280), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11550) );
  AOI22_X1 U14630 ( .A1(n10145), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10172), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11549) );
  AOI22_X1 U14631 ( .A1(n10274), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10271), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11548) );
  NAND4_X1 U14632 ( .A1(n11551), .A2(n11550), .A3(n11549), .A4(n11548), .ZN(
        n11552) );
  NOR2_X1 U14633 ( .A1(n11553), .A2(n11552), .ZN(n18883) );
  AOI22_X1 U14634 ( .A1(n10272), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11595), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U14635 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11556) );
  AOI22_X1 U14636 ( .A1(n11637), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11555) );
  AOI22_X1 U14637 ( .A1(n11640), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11554) );
  NAND4_X1 U14638 ( .A1(n11557), .A2(n11556), .A3(n11555), .A4(n11554), .ZN(
        n11563) );
  AOI22_X1 U14639 ( .A1(n10165), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10279), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11561) );
  AOI22_X1 U14640 ( .A1(n11547), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10280), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11560) );
  AOI22_X1 U14641 ( .A1(n10145), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10172), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11559) );
  AOI22_X1 U14642 ( .A1(n10274), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10271), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11558) );
  NAND4_X1 U14643 ( .A1(n11561), .A2(n11560), .A3(n11559), .A4(n11558), .ZN(
        n11562) );
  OR2_X1 U14644 ( .A1(n11563), .A2(n11562), .ZN(n13896) );
  NAND2_X1 U14645 ( .A1(n13895), .A2(n13896), .ZN(n15892) );
  AOI22_X1 U14646 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n11595), .B1(
        n10272), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11567) );
  AOI22_X1 U14647 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__2__SCAN_IN), .B2(n11638), .ZN(n11566) );
  AOI22_X1 U14648 ( .A1(n11637), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11565) );
  AOI22_X1 U14649 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10369), .B1(
        n11640), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11564) );
  NAND4_X1 U14650 ( .A1(n11567), .A2(n11566), .A3(n11565), .A4(n11564), .ZN(
        n11573) );
  AOI22_X1 U14651 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n10279), .B1(
        n10165), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11571) );
  AOI22_X1 U14652 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10280), .B1(
        n11547), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U14653 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10172), .B1(
        n10145), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U14654 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n10274), .B1(
        n10271), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11568) );
  NAND4_X1 U14655 ( .A1(n11571), .A2(n11570), .A3(n11569), .A4(n11568), .ZN(
        n11572) );
  NOR2_X1 U14656 ( .A1(n11573), .A2(n11572), .ZN(n15893) );
  AOI22_X1 U14657 ( .A1(n10272), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11595), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U14658 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11577) );
  AOI22_X1 U14659 ( .A1(n11637), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11576) );
  AOI22_X1 U14660 ( .A1(n11640), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11575) );
  NAND4_X1 U14661 ( .A1(n11578), .A2(n11577), .A3(n11576), .A4(n11575), .ZN(
        n11584) );
  AOI22_X1 U14662 ( .A1(n10165), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10279), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U14663 ( .A1(n11547), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10280), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11581) );
  AOI22_X1 U14664 ( .A1(n10145), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10172), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11580) );
  AOI22_X1 U14665 ( .A1(n10274), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10271), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11579) );
  NAND4_X1 U14666 ( .A1(n11582), .A2(n11581), .A3(n11580), .A4(n11579), .ZN(
        n11583) );
  NOR2_X1 U14667 ( .A1(n11584), .A2(n11583), .ZN(n14836) );
  AOI22_X1 U14668 ( .A1(n10272), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11595), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11588) );
  AOI22_X1 U14669 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11587) );
  AOI22_X1 U14670 ( .A1(n11637), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11586) );
  AOI22_X1 U14671 ( .A1(n11640), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11585) );
  NAND4_X1 U14672 ( .A1(n11588), .A2(n11587), .A3(n11586), .A4(n11585), .ZN(
        n11594) );
  AOI22_X1 U14673 ( .A1(n10165), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10279), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11592) );
  AOI22_X1 U14674 ( .A1(n11547), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10280), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11591) );
  AOI22_X1 U14675 ( .A1(n10145), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10172), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11590) );
  AOI22_X1 U14676 ( .A1(n10274), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10271), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11589) );
  NAND4_X1 U14677 ( .A1(n11592), .A2(n11591), .A3(n11590), .A4(n11589), .ZN(
        n11593) );
  OR2_X1 U14678 ( .A1(n11594), .A2(n11593), .ZN(n15884) );
  AOI22_X1 U14679 ( .A1(n10272), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11595), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11599) );
  AOI22_X1 U14680 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11638), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11598) );
  AOI22_X1 U14681 ( .A1(n11637), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11597) );
  AOI22_X1 U14682 ( .A1(n11640), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10369), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11596) );
  NAND4_X1 U14683 ( .A1(n11599), .A2(n11598), .A3(n11597), .A4(n11596), .ZN(
        n11605) );
  AOI22_X1 U14684 ( .A1(n10165), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10279), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11603) );
  AOI22_X1 U14685 ( .A1(n11547), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10280), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11602) );
  AOI22_X1 U14686 ( .A1(n10145), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10172), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11601) );
  AOI22_X1 U14687 ( .A1(n10274), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10271), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11600) );
  NAND4_X1 U14688 ( .A1(n11603), .A2(n11602), .A3(n11601), .A4(n11600), .ZN(
        n11604) );
  OR2_X1 U14689 ( .A1(n11605), .A2(n11604), .ZN(n14832) );
  AOI22_X1 U14690 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n11595), .B1(
        n10272), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11609) );
  AOI22_X1 U14691 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__6__SCAN_IN), .B2(n11638), .ZN(n11608) );
  AOI22_X1 U14692 ( .A1(n11637), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11607) );
  AOI22_X1 U14693 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10369), .B1(
        n11640), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11606) );
  NAND4_X1 U14694 ( .A1(n11609), .A2(n11608), .A3(n11607), .A4(n11606), .ZN(
        n11615) );
  AOI22_X1 U14695 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n10279), .B1(
        n10165), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11613) );
  AOI22_X1 U14696 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10280), .B1(
        n11547), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11612) );
  AOI22_X1 U14697 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10172), .B1(
        n10145), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11611) );
  AOI22_X1 U14698 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n10274), .B1(
        n10271), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11610) );
  NAND4_X1 U14699 ( .A1(n11613), .A2(n11612), .A3(n11611), .A4(n11610), .ZN(
        n11614) );
  NOR2_X1 U14700 ( .A1(n11615), .A2(n11614), .ZN(n14892) );
  INV_X1 U14701 ( .A(n11616), .ZN(n11747) );
  INV_X1 U14702 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11618) );
  INV_X1 U14703 ( .A(n11809), .ZN(n11745) );
  INV_X1 U14704 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11617) );
  OAI22_X1 U14705 ( .A1(n11747), .A2(n11618), .B1(n11745), .B2(n11617), .ZN(
        n11621) );
  INV_X1 U14706 ( .A(n11810), .ZN(n11751) );
  INV_X1 U14707 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11619) );
  INV_X1 U14708 ( .A(n11668), .ZN(n11736) );
  INV_X1 U14709 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n19558) );
  OAI22_X1 U14710 ( .A1(n11751), .A2(n11619), .B1(n11736), .B2(n19558), .ZN(
        n11620) );
  NOR2_X1 U14711 ( .A1(n11621), .A2(n11620), .ZN(n11625) );
  XNOR2_X1 U14712 ( .A(n10156), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11803) );
  INV_X1 U14713 ( .A(n11712), .ZN(n11805) );
  AOI22_X1 U14714 ( .A1(n11805), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11622), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11624) );
  INV_X1 U14715 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n19391) );
  AOI22_X1 U14716 ( .A1(n9564), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11740), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11623) );
  NAND4_X1 U14717 ( .A1(n11625), .A2(n11803), .A3(n11624), .A4(n11623), .ZN(
        n11636) );
  INV_X1 U14718 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11627) );
  INV_X1 U14719 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11626) );
  OAI22_X1 U14720 ( .A1(n11747), .A2(n11627), .B1(n11745), .B2(n11626), .ZN(
        n11630) );
  INV_X1 U14721 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11628) );
  INV_X1 U14722 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n19106) );
  OAI22_X1 U14723 ( .A1(n11751), .A2(n11628), .B1(n9581), .B2(n19106), .ZN(
        n11629) );
  NOR2_X1 U14724 ( .A1(n11630), .A2(n11629), .ZN(n11634) );
  AOI22_X1 U14725 ( .A1(n11622), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11633) );
  INV_X1 U14726 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n20829) );
  AOI22_X1 U14727 ( .A1(n11805), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11740), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11632) );
  INV_X1 U14728 ( .A(n11803), .ZN(n11806) );
  NAND4_X1 U14729 ( .A1(n11634), .A2(n11633), .A3(n11632), .A4(n11806), .ZN(
        n11635) );
  AND2_X1 U14730 ( .A1(n11636), .A2(n11635), .ZN(n11651) );
  NAND2_X1 U14731 ( .A1(n19054), .A2(n11651), .ZN(n11654) );
  AOI22_X1 U14732 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n11637), .B1(
        n10272), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U14733 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n11638), .ZN(n11643) );
  AOI22_X1 U14734 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n11640), .B1(
        n10145), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11642) );
  AOI22_X1 U14735 ( .A1(n11595), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10271), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11641) );
  NAND4_X1 U14736 ( .A1(n11644), .A2(n11643), .A3(n11642), .A4(n11641), .ZN(
        n11650) );
  AOI22_X1 U14737 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n11547), .B1(
        n10165), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11648) );
  AOI22_X1 U14738 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10280), .B1(
        n10279), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11647) );
  AOI22_X1 U14739 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10369), .B1(
        n10120), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U14740 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n10274), .B1(
        n10172), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11645) );
  NAND4_X1 U14741 ( .A1(n11648), .A2(n11647), .A3(n11646), .A4(n11645), .ZN(
        n11649) );
  NOR2_X1 U14742 ( .A1(n11650), .A2(n11649), .ZN(n11677) );
  XOR2_X1 U14743 ( .A(n11654), .B(n11677), .Z(n11652) );
  XNOR2_X2 U14744 ( .A(n14889), .B(n11652), .ZN(n14166) );
  INV_X1 U14745 ( .A(n11651), .ZN(n11675) );
  NOR2_X1 U14746 ( .A1(n19054), .A2(n11675), .ZN(n14165) );
  INV_X1 U14747 ( .A(n11652), .ZN(n11653) );
  NOR2_X1 U14748 ( .A1(n11677), .A2(n11654), .ZN(n11674) );
  INV_X1 U14749 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19059) );
  INV_X1 U14750 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11655) );
  OAI22_X1 U14751 ( .A1(n11709), .A2(n19059), .B1(n11736), .B2(n11655), .ZN(
        n11658) );
  OAI22_X1 U14752 ( .A1(n11712), .A2(n9820), .B1(n9581), .B2(n11101), .ZN(
        n11657) );
  NOR2_X1 U14753 ( .A1(n11658), .A2(n11657), .ZN(n11662) );
  AOI22_X1 U14754 ( .A1(n11810), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11661) );
  AOI22_X1 U14755 ( .A1(n11659), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11809), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11660) );
  NAND4_X1 U14756 ( .A1(n11662), .A2(n11661), .A3(n11660), .A4(n11806), .ZN(
        n11673) );
  OAI22_X1 U14757 ( .A1(n11747), .A2(n11663), .B1(n11745), .B2(n11102), .ZN(
        n11667) );
  INV_X1 U14758 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11665) );
  INV_X1 U14759 ( .A(n11787), .ZN(n11749) );
  OAI22_X1 U14760 ( .A1(n11751), .A2(n11665), .B1(n11749), .B2(n11664), .ZN(
        n11666) );
  NOR2_X1 U14761 ( .A1(n11667), .A2(n11666), .ZN(n11671) );
  AOI22_X1 U14762 ( .A1(n11622), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11668), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11670) );
  AOI22_X1 U14763 ( .A1(n11805), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9564), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11669) );
  NAND4_X1 U14764 ( .A1(n11671), .A2(n11803), .A3(n11670), .A4(n11669), .ZN(
        n11672) );
  NAND2_X1 U14765 ( .A1(n11673), .A2(n11672), .ZN(n11676) );
  XNOR2_X1 U14766 ( .A(n11674), .B(n11676), .ZN(n14823) );
  NOR2_X1 U14767 ( .A1(n11676), .A2(n11675), .ZN(n11679) );
  INV_X1 U14768 ( .A(n11677), .ZN(n11678) );
  AND2_X1 U14769 ( .A1(n11679), .A2(n11678), .ZN(n11700) );
  INV_X1 U14770 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11681) );
  INV_X1 U14771 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11680) );
  OAI22_X1 U14772 ( .A1(n11747), .A2(n11681), .B1(n11745), .B2(n11680), .ZN(
        n11685) );
  INV_X1 U14773 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11683) );
  INV_X1 U14774 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11682) );
  OAI22_X1 U14775 ( .A1(n11751), .A2(n11683), .B1(n11749), .B2(n11682), .ZN(
        n11684) );
  NOR2_X1 U14776 ( .A1(n11685), .A2(n11684), .ZN(n11688) );
  AOI22_X1 U14777 ( .A1(n11622), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U14778 ( .A1(n11805), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9564), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11686) );
  NAND4_X1 U14779 ( .A1(n11688), .A2(n11687), .A3(n11686), .A4(n11806), .ZN(
        n11699) );
  INV_X1 U14780 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11690) );
  INV_X1 U14781 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11689) );
  OAI22_X1 U14782 ( .A1(n11747), .A2(n11690), .B1(n11745), .B2(n11689), .ZN(
        n11694) );
  INV_X1 U14783 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11692) );
  INV_X1 U14784 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11691) );
  OAI22_X1 U14785 ( .A1(n11751), .A2(n11692), .B1(n11749), .B2(n11691), .ZN(
        n11693) );
  NOR2_X1 U14786 ( .A1(n11694), .A2(n11693), .ZN(n11697) );
  AOI22_X1 U14787 ( .A1(n11622), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U14788 ( .A1(n11805), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9564), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11695) );
  NAND4_X1 U14789 ( .A1(n11697), .A2(n11803), .A3(n11696), .A4(n11695), .ZN(
        n11698) );
  AND2_X1 U14790 ( .A1(n11699), .A2(n11698), .ZN(n11702) );
  NAND2_X1 U14791 ( .A1(n11700), .A2(n11702), .ZN(n11731) );
  OAI211_X1 U14792 ( .C1(n11700), .C2(n11702), .A(n11761), .B(n11731), .ZN(
        n11705) );
  INV_X1 U14793 ( .A(n11702), .ZN(n11703) );
  NOR2_X1 U14794 ( .A1(n19054), .A2(n11703), .ZN(n14817) );
  INV_X1 U14795 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11708) );
  OAI22_X1 U14796 ( .A1(n11709), .A2(n19069), .B1(n11736), .B2(n11708), .ZN(
        n11714) );
  INV_X1 U14797 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11711) );
  OAI22_X1 U14798 ( .A1(n11712), .A2(n11711), .B1(n9581), .B2(n11710), .ZN(
        n11713) );
  NOR2_X1 U14799 ( .A1(n11714), .A2(n11713), .ZN(n11717) );
  AOI22_X1 U14800 ( .A1(n11810), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11716) );
  AOI22_X1 U14801 ( .A1(n11659), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11809), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11715) );
  NAND4_X1 U14802 ( .A1(n11717), .A2(n11716), .A3(n11715), .A4(n11806), .ZN(
        n11727) );
  OAI22_X1 U14803 ( .A1(n11747), .A2(n11718), .B1(n11745), .B2(n10372), .ZN(
        n11722) );
  INV_X1 U14804 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11720) );
  OAI22_X1 U14805 ( .A1(n11751), .A2(n11720), .B1(n11749), .B2(n11719), .ZN(
        n11721) );
  NOR2_X1 U14806 ( .A1(n11722), .A2(n11721), .ZN(n11725) );
  AOI22_X1 U14807 ( .A1(n11622), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11724) );
  AOI22_X1 U14808 ( .A1(n11805), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9564), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11723) );
  NAND4_X1 U14809 ( .A1(n11725), .A2(n11803), .A3(n11724), .A4(n11723), .ZN(
        n11726) );
  AND2_X1 U14810 ( .A1(n11727), .A2(n11726), .ZN(n11732) );
  XNOR2_X1 U14811 ( .A(n11731), .B(n11732), .ZN(n11728) );
  XNOR2_X2 U14812 ( .A(n11729), .B(n10001), .ZN(n14808) );
  NAND2_X1 U14813 ( .A1(n16044), .A2(n11732), .ZN(n14807) );
  INV_X1 U14814 ( .A(n11731), .ZN(n11733) );
  NAND2_X1 U14815 ( .A1(n11733), .A2(n11732), .ZN(n11760) );
  INV_X1 U14816 ( .A(n11760), .ZN(n11762) );
  INV_X1 U14817 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n19321) );
  INV_X1 U14818 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11734) );
  OAI22_X1 U14819 ( .A1(n19321), .A2(n11745), .B1(n11747), .B2(n11734), .ZN(
        n11739) );
  INV_X1 U14820 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11737) );
  INV_X1 U14821 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11735) );
  OAI22_X1 U14822 ( .A1(n11751), .A2(n11737), .B1(n11736), .B2(n11735), .ZN(
        n11738) );
  NOR2_X1 U14823 ( .A1(n11739), .A2(n11738), .ZN(n11743) );
  AOI22_X1 U14824 ( .A1(n11622), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9564), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11742) );
  AOI22_X1 U14825 ( .A1(n11805), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11740), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11741) );
  NAND4_X1 U14826 ( .A1(n11743), .A2(n11742), .A3(n11741), .A4(n11806), .ZN(
        n11758) );
  INV_X1 U14827 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11746) );
  INV_X1 U14828 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11744) );
  OAI22_X1 U14829 ( .A1(n11747), .A2(n11746), .B1(n11745), .B2(n11744), .ZN(
        n11753) );
  INV_X1 U14830 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11750) );
  INV_X1 U14831 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11748) );
  OAI22_X1 U14832 ( .A1(n11751), .A2(n11750), .B1(n11749), .B2(n11748), .ZN(
        n11752) );
  NOR2_X1 U14833 ( .A1(n11753), .A2(n11752), .ZN(n11756) );
  AOI22_X1 U14834 ( .A1(n11622), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11755) );
  AOI22_X1 U14835 ( .A1(n11805), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9564), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11754) );
  NAND4_X1 U14836 ( .A1(n11756), .A2(n11803), .A3(n11755), .A4(n11754), .ZN(
        n11757) );
  NAND2_X1 U14837 ( .A1(n11758), .A2(n11757), .ZN(n11759) );
  INV_X1 U14838 ( .A(n11759), .ZN(n11765) );
  OR2_X1 U14839 ( .A1(n11760), .A2(n11759), .ZN(n14791) );
  OAI211_X1 U14840 ( .C1(n11762), .C2(n11765), .A(n14791), .B(n11761), .ZN(
        n11763) );
  NAND2_X1 U14841 ( .A1(n16044), .A2(n11765), .ZN(n14798) );
  NOR2_X2 U14842 ( .A1(n14799), .A2(n14798), .ZN(n14797) );
  AOI22_X1 U14843 ( .A1(n11659), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11809), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11767) );
  AOI22_X1 U14844 ( .A1(n11810), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11787), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11766) );
  NAND2_X1 U14845 ( .A1(n11767), .A2(n11766), .ZN(n11777) );
  AOI22_X1 U14846 ( .A1(n11805), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9564), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11769) );
  AOI22_X1 U14847 ( .A1(n11622), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11768) );
  NAND3_X1 U14848 ( .A1(n11769), .A2(n11768), .A3(n11806), .ZN(n11776) );
  AOI22_X1 U14849 ( .A1(n11805), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9564), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11771) );
  AOI22_X1 U14850 ( .A1(n11622), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11770) );
  NAND3_X1 U14851 ( .A1(n11771), .A2(n11770), .A3(n11803), .ZN(n11775) );
  AOI22_X1 U14852 ( .A1(n11659), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11809), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11773) );
  AOI22_X1 U14853 ( .A1(n11810), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11740), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11772) );
  NAND2_X1 U14854 ( .A1(n11773), .A2(n11772), .ZN(n11774) );
  OAI22_X1 U14855 ( .A1(n11777), .A2(n11776), .B1(n11775), .B2(n11774), .ZN(
        n11779) );
  INV_X1 U14856 ( .A(n11779), .ZN(n14793) );
  NOR3_X1 U14857 ( .A1(n14791), .A2(n16044), .A3(n11779), .ZN(n11796) );
  AOI22_X1 U14858 ( .A1(n11805), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11810), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11781) );
  AOI22_X1 U14859 ( .A1(n11616), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11809), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11780) );
  NAND2_X1 U14860 ( .A1(n11781), .A2(n11780), .ZN(n11793) );
  AOI22_X1 U14861 ( .A1(n11622), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11784) );
  AOI22_X1 U14862 ( .A1(n9564), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11783) );
  NAND3_X1 U14863 ( .A1(n11784), .A2(n11783), .A3(n11806), .ZN(n11792) );
  AOI22_X1 U14864 ( .A1(n11805), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11810), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11786) );
  AOI22_X1 U14865 ( .A1(n11659), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11809), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11785) );
  NAND2_X1 U14866 ( .A1(n11786), .A2(n11785), .ZN(n11791) );
  AOI22_X1 U14867 ( .A1(n11622), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11789) );
  AOI22_X1 U14868 ( .A1(n9564), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11787), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11788) );
  NAND3_X1 U14869 ( .A1(n11789), .A2(n11788), .A3(n11803), .ZN(n11790) );
  OAI22_X1 U14870 ( .A1(n11793), .A2(n11792), .B1(n11791), .B2(n11790), .ZN(
        n11794) );
  INV_X1 U14871 ( .A(n11794), .ZN(n11795) );
  NAND2_X1 U14872 ( .A1(n11796), .A2(n11795), .ZN(n11797) );
  OAI21_X1 U14873 ( .B1(n11796), .B2(n11795), .A(n11797), .ZN(n14787) );
  INV_X1 U14874 ( .A(n11797), .ZN(n11798) );
  NOR2_X1 U14875 ( .A1(n14786), .A2(n11798), .ZN(n11818) );
  AOI22_X1 U14876 ( .A1(n11659), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11809), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11800) );
  AOI22_X1 U14877 ( .A1(n11810), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11740), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11799) );
  NAND2_X1 U14878 ( .A1(n11800), .A2(n11799), .ZN(n11816) );
  AOI22_X1 U14879 ( .A1(n11805), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11622), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11804) );
  AOI22_X1 U14880 ( .A1(n9564), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11802) );
  NAND3_X1 U14881 ( .A1(n11804), .A2(n11803), .A3(n11802), .ZN(n11815) );
  AOI22_X1 U14882 ( .A1(n11805), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11782), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11808) );
  AOI22_X1 U14883 ( .A1(n11622), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11801), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11807) );
  NAND3_X1 U14884 ( .A1(n11808), .A2(n11807), .A3(n11806), .ZN(n11814) );
  AOI22_X1 U14885 ( .A1(n11659), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11809), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11812) );
  AOI22_X1 U14886 ( .A1(n11810), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9564), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11811) );
  NAND2_X1 U14887 ( .A1(n11812), .A2(n11811), .ZN(n11813) );
  OAI22_X1 U14888 ( .A1(n11816), .A2(n11815), .B1(n11814), .B2(n11813), .ZN(
        n11817) );
  XNOR2_X1 U14889 ( .A(n11818), .B(n11817), .ZN(n14204) );
  OR3_X1 U14890 ( .A1(n13097), .A2(n11404), .A3(n19690), .ZN(n11821) );
  NAND2_X1 U14891 ( .A1(n16041), .A2(n11819), .ZN(n11820) );
  NAND2_X1 U14892 ( .A1(n11821), .A2(n11820), .ZN(n13368) );
  NAND2_X1 U14893 ( .A1(n18956), .A2(n11824), .ZN(n18986) );
  AND2_X1 U14894 ( .A1(n18956), .A2(n9586), .ZN(n13189) );
  NOR4_X1 U14895 ( .A1(P2_ADDRESS_REG_17__SCAN_IN), .A2(
        P2_ADDRESS_REG_16__SCAN_IN), .A3(P2_ADDRESS_REG_15__SCAN_IN), .A4(
        P2_ADDRESS_REG_14__SCAN_IN), .ZN(n11828) );
  NOR4_X1 U14896 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_19__SCAN_IN), .A4(
        P2_ADDRESS_REG_18__SCAN_IN), .ZN(n11827) );
  NOR4_X1 U14897 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n11826) );
  NOR4_X1 U14898 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n11825) );
  NAND4_X1 U14899 ( .A1(n11828), .A2(n11827), .A3(n11826), .A4(n11825), .ZN(
        n11833) );
  NOR4_X1 U14900 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n11831) );
  NOR4_X1 U14901 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n11830) );
  NOR4_X1 U14902 ( .A1(P2_ADDRESS_REG_13__SCAN_IN), .A2(
        P2_ADDRESS_REG_11__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n11829) );
  INV_X1 U14903 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19703) );
  NAND4_X1 U14904 ( .A1(n11831), .A2(n11830), .A3(n11829), .A4(n19703), .ZN(
        n11832) );
  OAI21_X1 U14905 ( .B1(n11833), .B2(n11832), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n15407) );
  INV_X1 U14906 ( .A(n15405), .ZN(n13263) );
  MUX2_X1 U14907 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n13263), .Z(n19030) );
  NAND2_X1 U14908 ( .A1(n18956), .A2(n9868), .ZN(n18935) );
  INV_X1 U14909 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n11834) );
  OAI22_X1 U14910 ( .A1(n14144), .A2(n18935), .B1(n18956), .B2(n11834), .ZN(
        n11835) );
  AOI21_X1 U14911 ( .B1(n18926), .B2(n19030), .A(n11835), .ZN(n11838) );
  INV_X1 U14912 ( .A(n13189), .ZN(n11836) );
  NOR3_X4 U14913 ( .A1(n11836), .A2(n13192), .A3(n13263), .ZN(n18928) );
  NOR3_X2 U14914 ( .A1(n11836), .A2(n13192), .A3(n15405), .ZN(n18927) );
  AOI22_X1 U14915 ( .A1(n18928), .A2(BUF1_REG_30__SCAN_IN), .B1(n18927), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n11837) );
  OAI21_X1 U14916 ( .B1(n14204), .B2(n18986), .A(n11839), .ZN(P2_U2889) );
  AND2_X2 U14917 ( .A1(n11859), .A2(n13424), .ZN(n12484) );
  NAND2_X1 U14918 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11845) );
  INV_X1 U14919 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11841) );
  AND2_X2 U14920 ( .A1(n11841), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11858) );
  NAND2_X1 U14921 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11844) );
  NAND2_X1 U14922 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11843) );
  AND2_X4 U14923 ( .A1(n11858), .A2(n13570), .ZN(n12633) );
  NAND2_X1 U14924 ( .A1(n12633), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11842) );
  AND2_X2 U14925 ( .A1(n11859), .A2(n13425), .ZN(n12067) );
  NAND2_X1 U14926 ( .A1(n12067), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11850) );
  NAND2_X1 U14927 ( .A1(n12614), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11849) );
  AND2_X2 U14928 ( .A1(n11858), .A2(n11860), .ZN(n12146) );
  NAND2_X1 U14929 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11848) );
  NAND2_X1 U14930 ( .A1(n12022), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11847) );
  NAND2_X1 U14931 ( .A1(n12641), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11857) );
  AND2_X2 U14932 ( .A1(n11852), .A2(n11860), .ZN(n11928) );
  NAND2_X1 U14933 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11856) );
  AND2_X2 U14934 ( .A1(n13569), .A2(n11853), .ZN(n11893) );
  BUF_X4 U14935 ( .A(n11893), .Z(n12544) );
  NAND2_X1 U14936 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11855) );
  AND3_X4 U14937 ( .A1(n13569), .A2(n11846), .A3(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12635) );
  NAND2_X1 U14938 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11854) );
  AND2_X2 U14939 ( .A1(n11859), .A2(n11858), .ZN(n11922) );
  NAND2_X1 U14940 ( .A1(n11922), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11864) );
  AND2_X2 U14941 ( .A1(n11860), .A2(n13424), .ZN(n12066) );
  NAND2_X1 U14942 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11863) );
  NAND2_X1 U14943 ( .A1(n12296), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11862) );
  NAND2_X1 U14944 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11861) );
  NAND4_X4 U14945 ( .A1(n11868), .A2(n11867), .A3(n11866), .A4(n11865), .ZN(
        n11971) );
  AOI22_X1 U14946 ( .A1(n12067), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11927), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11872) );
  AOI22_X1 U14947 ( .A1(n12614), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11939), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11871) );
  AOI22_X1 U14948 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11870) );
  AOI22_X1 U14949 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12022), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11869) );
  AOI22_X1 U14950 ( .A1(n11922), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12066), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11874) );
  AOI22_X1 U14951 ( .A1(n12641), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11928), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11873) );
  NAND2_X1 U14952 ( .A1(n11874), .A2(n11873), .ZN(n11878) );
  AOI22_X1 U14953 ( .A1(n12642), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11876) );
  AOI22_X1 U14954 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11893), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11875) );
  NAND2_X1 U14955 ( .A1(n11876), .A2(n11875), .ZN(n11877) );
  NOR2_X1 U14956 ( .A1(n11878), .A2(n11877), .ZN(n11879) );
  AOI22_X1 U14957 ( .A1(n12641), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11928), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11883) );
  AOI22_X1 U14958 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11882) );
  AOI22_X1 U14959 ( .A1(n11922), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12066), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11881) );
  AOI22_X1 U14960 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12644), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11880) );
  AOI22_X1 U14961 ( .A1(n12614), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11939), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11886) );
  AOI22_X1 U14962 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11885) );
  AOI22_X1 U14963 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12022), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11884) );
  NAND2_X1 U14964 ( .A1(n11918), .A2(n11971), .ZN(n11899) );
  AOI22_X1 U14965 ( .A1(n12641), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12396), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U14966 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11890) );
  AOI22_X1 U14967 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12022), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11889) );
  AOI22_X1 U14968 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11939), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11888) );
  AOI22_X1 U14969 ( .A1(n11922), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11892), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11897) );
  AOI22_X1 U14970 ( .A1(n12067), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12066), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11896) );
  AOI22_X1 U14971 ( .A1(n12614), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11895) );
  AOI22_X1 U14972 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11893), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11894) );
  MUX2_X1 U14973 ( .A(n13000), .B(n11899), .S(n20085), .Z(n11920) );
  INV_X2 U14974 ( .A(n11918), .ZN(n20104) );
  AOI22_X1 U14975 ( .A1(n11922), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12067), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11903) );
  AOI22_X1 U14976 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12396), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11902) );
  AOI22_X1 U14977 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12644), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11901) );
  AOI22_X1 U14978 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11900) );
  AOI22_X1 U14979 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11907) );
  AOI22_X1 U14980 ( .A1(n12641), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11906) );
  AOI22_X1 U14981 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12066), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U14982 ( .A1(n12614), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12022), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11904) );
  NAND2_X2 U14983 ( .A1(n10015), .A2(n9616), .ZN(n12759) );
  AOI22_X1 U14984 ( .A1(n12641), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12396), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11911) );
  AOI22_X1 U14985 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11910) );
  AOI22_X1 U14986 ( .A1(n12469), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12066), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U14987 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12644), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11908) );
  NAND4_X1 U14988 ( .A1(n11911), .A2(n11910), .A3(n11909), .A4(n11908), .ZN(
        n11917) );
  AOI22_X1 U14989 ( .A1(n12067), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12634), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11915) );
  AOI22_X1 U14990 ( .A1(n12614), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11939), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11914) );
  AOI22_X1 U14991 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11913) );
  AOI22_X1 U14992 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12022), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11912) );
  NAND4_X1 U14993 ( .A1(n11915), .A2(n11914), .A3(n11913), .A4(n11912), .ZN(
        n11916) );
  OR2_X2 U14994 ( .A1(n11917), .A2(n11916), .ZN(n13381) );
  NAND2_X1 U14995 ( .A1(n11972), .A2(n13381), .ZN(n11962) );
  NAND3_X1 U14996 ( .A1(n11920), .A2(n11989), .A3(n11919), .ZN(n11970) );
  NOR2_X2 U14997 ( .A1(n12759), .A2(n13437), .ZN(n13577) );
  INV_X1 U14998 ( .A(n13577), .ZN(n12999) );
  AOI22_X1 U14999 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11926) );
  AOI22_X1 U15000 ( .A1(n12641), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11925) );
  AOI22_X1 U15001 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12644), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U15002 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11939), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11923) );
  NAND4_X1 U15003 ( .A1(n11926), .A2(n11925), .A3(n11924), .A4(n11923), .ZN(
        n11934) );
  AOI22_X1 U15004 ( .A1(n12067), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11927), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11932) );
  BUF_X4 U15005 ( .A(n11928), .Z(n12645) );
  AOI22_X1 U15006 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12066), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11931) );
  AOI22_X1 U15007 ( .A1(n12614), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11930) );
  AOI22_X1 U15008 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12022), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11929) );
  NAND4_X1 U15009 ( .A1(n11932), .A2(n11931), .A3(n11930), .A4(n11929), .ZN(
        n11933) );
  OR2_X4 U15010 ( .A1(n11934), .A2(n11933), .ZN(n13325) );
  NAND2_X1 U15011 ( .A1(n12999), .A2(n11957), .ZN(n11956) );
  NAND2_X1 U15012 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11938) );
  NAND2_X1 U15013 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11937) );
  NAND2_X1 U15014 ( .A1(n12633), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11936) );
  NAND2_X1 U15015 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11935) );
  NAND2_X1 U15016 ( .A1(n12067), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11943) );
  BUF_X8 U15017 ( .A(n12614), .Z(n12643) );
  NAND2_X1 U15018 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11942) );
  NAND2_X1 U15019 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11941) );
  NAND2_X1 U15020 ( .A1(n11939), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11940) );
  NAND2_X1 U15021 ( .A1(n12641), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11947) );
  NAND2_X1 U15022 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11946) );
  NAND2_X1 U15023 ( .A1(n12544), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11945) );
  NAND2_X1 U15024 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11944) );
  NAND2_X1 U15025 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11951) );
  NAND2_X1 U15026 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11950) );
  NAND2_X1 U15027 ( .A1(n12296), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11949) );
  NAND2_X1 U15028 ( .A1(n12022), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11948) );
  NAND4_X4 U15029 ( .A1(n11955), .A2(n11954), .A3(n11953), .A4(n11952), .ZN(
        n12697) );
  OAI21_X1 U15030 ( .B1(n11970), .B2(n11956), .A(n20072), .ZN(n11967) );
  INV_X1 U15031 ( .A(n12759), .ZN(n20090) );
  NAND2_X1 U15032 ( .A1(n13437), .A2(n12697), .ZN(n11992) );
  NAND2_X1 U15033 ( .A1(n12901), .A2(n11992), .ZN(n12997) );
  AND2_X2 U15034 ( .A1(n11957), .A2(n12697), .ZN(n13271) );
  NAND2_X1 U15035 ( .A1(n13271), .A2(n11972), .ZN(n11958) );
  NAND2_X1 U15036 ( .A1(n12759), .A2(n13325), .ZN(n12900) );
  NAND2_X1 U15037 ( .A1(n13000), .A2(n14243), .ZN(n13419) );
  NAND2_X1 U15038 ( .A1(n11958), .A2(n13419), .ZN(n11994) );
  NOR2_X1 U15039 ( .A1(n12997), .A2(n11994), .ZN(n11966) );
  NAND2_X1 U15040 ( .A1(n20099), .A2(n12671), .ZN(n11959) );
  NAND2_X1 U15041 ( .A1(n12883), .A2(n20094), .ZN(n11961) );
  AND2_X2 U15042 ( .A1(n11995), .A2(n11961), .ZN(n13004) );
  NAND3_X1 U15043 ( .A1(n11967), .A2(n11966), .A3(n11965), .ZN(n12996) );
  NOR2_X1 U15044 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15796) );
  NAND2_X1 U15045 ( .A1(n15796), .A2(n20071), .ZN(n12860) );
  INV_X1 U15046 ( .A(n12860), .ZN(n12011) );
  NAND2_X1 U15047 ( .A1(n20429), .A2(n20773), .ZN(n11968) );
  NAND2_X1 U15048 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n12009) );
  AND2_X1 U15049 ( .A1(n11968), .A2(n12009), .ZN(n20426) );
  NAND2_X1 U15050 ( .A1(n13584), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20686) );
  AND2_X1 U15051 ( .A1(n20686), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12002) );
  AOI21_X1 U15052 ( .B1(n12011), .B2(n20426), .A(n12002), .ZN(n11979) );
  NOR2_X1 U15053 ( .A1(n11970), .A2(n11969), .ZN(n12882) );
  NAND2_X1 U15054 ( .A1(n12882), .A2(n11957), .ZN(n12674) );
  NOR2_X1 U15055 ( .A1(n11972), .A2(n11971), .ZN(n11974) );
  AND2_X4 U15056 ( .A1(n13325), .A2(n12697), .ZN(n13063) );
  NAND2_X1 U15057 ( .A1(n12692), .A2(n13063), .ZN(n11975) );
  NAND2_X1 U15058 ( .A1(n12674), .A2(n11975), .ZN(n12894) );
  XNOR2_X1 U15059 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12874) );
  NAND2_X1 U15060 ( .A1(n11978), .A2(n11986), .ZN(n11982) );
  INV_X1 U15061 ( .A(n11979), .ZN(n11980) );
  OR2_X1 U15062 ( .A1(n11980), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11981) );
  NAND2_X1 U15063 ( .A1(n11986), .A2(n11985), .ZN(n12005) );
  NAND2_X1 U15064 ( .A1(n12005), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11988) );
  INV_X1 U15065 ( .A(n20686), .ZN(n12115) );
  MUX2_X1 U15066 ( .A(n12115), .B(n12860), .S(n20773), .Z(n11987) );
  INV_X1 U15067 ( .A(n11989), .ZN(n11990) );
  INV_X1 U15068 ( .A(n13126), .ZN(n13140) );
  NAND2_X1 U15069 ( .A1(n11990), .A2(n13140), .ZN(n11991) );
  NAND2_X1 U15070 ( .A1(n11970), .A2(n11991), .ZN(n12000) );
  NAND2_X1 U15071 ( .A1(n20072), .A2(n13325), .ZN(n13438) );
  NAND4_X1 U15072 ( .A1(n13438), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n15796), 
        .A4(n11992), .ZN(n11993) );
  OR2_X1 U15073 ( .A1(n11994), .A2(n11993), .ZN(n11997) );
  NAND2_X1 U15074 ( .A1(n13577), .A2(n20104), .ZN(n13009) );
  OAI21_X1 U15075 ( .B1(n11995), .B2(n20789), .A(n13009), .ZN(n11996) );
  NOR2_X1 U15076 ( .A1(n11997), .A2(n11996), .ZN(n11999) );
  NAND3_X1 U15077 ( .A1(n11964), .A2(n13325), .A3(n15460), .ZN(n11998) );
  NAND3_X1 U15078 ( .A1(n12000), .A2(n11999), .A3(n11998), .ZN(n12031) );
  INV_X1 U15079 ( .A(n12078), .ZN(n12001) );
  INV_X1 U15080 ( .A(n12002), .ZN(n12003) );
  NAND2_X1 U15081 ( .A1(n12003), .A2(n12675), .ZN(n12004) );
  NAND2_X1 U15082 ( .A1(n11983), .A2(n12004), .ZN(n12015) );
  NAND2_X1 U15083 ( .A1(n12077), .A2(n12015), .ZN(n12013) );
  AND2_X1 U15084 ( .A1(n20686), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12007) );
  INV_X1 U15085 ( .A(n12009), .ZN(n12008) );
  INV_X1 U15086 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12676) );
  NAND2_X1 U15087 ( .A1(n12008), .A2(n12676), .ZN(n20197) );
  NAND2_X1 U15088 ( .A1(n12009), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12010) );
  NAND2_X1 U15089 ( .A1(n20197), .A2(n12010), .ZN(n20075) );
  NAND2_X1 U15090 ( .A1(n12011), .A2(n20075), .ZN(n12014) );
  NAND2_X1 U15091 ( .A1(n12016), .A2(n12014), .ZN(n12012) );
  NAND2_X1 U15092 ( .A1(n12013), .A2(n12012), .ZN(n12113) );
  NAND4_X1 U15093 ( .A1(n12077), .A2(n12016), .A3(n12015), .A4(n12014), .ZN(
        n12017) );
  NAND2_X1 U15094 ( .A1(n12113), .A2(n12017), .ZN(n13076) );
  AOI22_X1 U15095 ( .A1(n12641), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12396), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12021) );
  AOI22_X1 U15096 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12020) );
  AOI22_X1 U15097 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12019) );
  AOI22_X1 U15098 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12644), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12018) );
  NAND4_X1 U15099 ( .A1(n12021), .A2(n12020), .A3(n12019), .A4(n12018), .ZN(
        n12028) );
  AOI22_X1 U15100 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12634), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12026) );
  AOI22_X1 U15101 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12025) );
  INV_X1 U15102 ( .A(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n20875) );
  AOI22_X1 U15103 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12024) );
  INV_X1 U15104 ( .A(n12022), .ZN(n13575) );
  AOI22_X1 U15105 ( .A1(n12571), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12023) );
  NAND4_X1 U15106 ( .A1(n12026), .A2(n12025), .A3(n12024), .A4(n12023), .ZN(
        n12027) );
  NOR2_X1 U15107 ( .A1(n12028), .A2(n12027), .ZN(n12774) );
  OAI22_X1 U15108 ( .A1(n13076), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n12774), 
        .B2(n12120), .ZN(n12030) );
  INV_X1 U15109 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n20089) );
  OAI22_X1 U15110 ( .A1(n12774), .A2(n12119), .B1(n12718), .B2(n20089), .ZN(
        n12029) );
  XNOR2_X1 U15111 ( .A(n12030), .B(n12029), .ZN(n12087) );
  INV_X1 U15112 ( .A(n12031), .ZN(n12032) );
  XNOR2_X1 U15113 ( .A(n12033), .B(n12032), .ZN(n12104) );
  AOI22_X1 U15114 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12067), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12037) );
  AOI22_X1 U15115 ( .A1(n12570), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12036) );
  AOI22_X1 U15116 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12035) );
  AOI22_X1 U15117 ( .A1(n12571), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12034) );
  NAND4_X1 U15118 ( .A1(n12037), .A2(n12036), .A3(n12035), .A4(n12034), .ZN(
        n12043) );
  AOI22_X1 U15119 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12048), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12041) );
  AOI22_X1 U15120 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12040) );
  AOI22_X1 U15121 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12644), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12039) );
  AOI22_X1 U15122 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12038) );
  NAND4_X1 U15123 ( .A1(n12041), .A2(n12040), .A3(n12039), .A4(n12038), .ZN(
        n12042) );
  NOR2_X1 U15124 ( .A1(n12120), .A2(n12811), .ZN(n12061) );
  INV_X1 U15125 ( .A(n12811), .ZN(n12817) );
  NOR2_X1 U15126 ( .A1(n12120), .A2(n12817), .ZN(n12060) );
  AOI22_X1 U15127 ( .A1(n12641), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12047) );
  AOI22_X1 U15128 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12046) );
  AOI22_X1 U15129 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12571), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12045) );
  AOI22_X1 U15130 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12044) );
  NAND4_X1 U15131 ( .A1(n12047), .A2(n12046), .A3(n12045), .A4(n12044), .ZN(
        n12054) );
  AOI22_X1 U15132 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12052) );
  AOI22_X1 U15133 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12051) );
  AOI22_X1 U15134 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U15135 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12049) );
  NAND4_X1 U15136 ( .A1(n12052), .A2(n12051), .A3(n12050), .A4(n12049), .ZN(
        n12053) );
  INV_X1 U15137 ( .A(n12760), .ZN(n12055) );
  MUX2_X1 U15138 ( .A(n12061), .B(n12060), .S(n12055), .Z(n12056) );
  INV_X1 U15139 ( .A(n12056), .ZN(n12057) );
  INV_X1 U15140 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20080) );
  AOI21_X1 U15141 ( .B1(n20094), .B2(n12811), .A(n20071), .ZN(n12059) );
  NAND2_X1 U15142 ( .A1(n20072), .A2(n12760), .ZN(n12058) );
  OAI211_X1 U15143 ( .C1(n12718), .C2(n20080), .A(n12059), .B(n12058), .ZN(
        n12102) );
  INV_X1 U15144 ( .A(n12060), .ZN(n12750) );
  NAND2_X1 U15145 ( .A1(n12723), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12076) );
  INV_X1 U15146 ( .A(n12061), .ZN(n12075) );
  AOI22_X1 U15147 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12641), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12065) );
  AOI22_X1 U15148 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12634), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12064) );
  AOI22_X1 U15149 ( .A1(n12633), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12063) );
  AOI22_X1 U15150 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12296), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12062) );
  NAND4_X1 U15151 ( .A1(n12065), .A2(n12064), .A3(n12063), .A4(n12062), .ZN(
        n12073) );
  AOI22_X1 U15152 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12071) );
  AOI22_X1 U15153 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12070) );
  BUF_X1 U15154 ( .A(n12067), .Z(n12331) );
  AOI22_X1 U15155 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U15156 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12068) );
  NAND4_X1 U15157 ( .A1(n12071), .A2(n12070), .A3(n12069), .A4(n12068), .ZN(
        n12072) );
  OR2_X1 U15158 ( .A1(n12073), .A2(n12072), .ZN(n12753) );
  INV_X1 U15159 ( .A(n12753), .ZN(n12079) );
  OR2_X1 U15160 ( .A1(n12119), .A2(n12079), .ZN(n12074) );
  XNOR2_X1 U15161 ( .A(n12081), .B(n12082), .ZN(n12095) );
  NAND2_X1 U15162 ( .A1(n12095), .A2(n12752), .ZN(n12085) );
  INV_X1 U15163 ( .A(n12082), .ZN(n12083) );
  NAND2_X1 U15164 ( .A1(n12087), .A2(n12086), .ZN(n12088) );
  NAND2_X1 U15165 ( .A1(n20104), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12311) );
  NAND2_X1 U15166 ( .A1(n13382), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12107) );
  NOR2_X2 U15167 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13041) );
  XNOR2_X1 U15168 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13514) );
  AND2_X1 U15169 ( .A1(n20074), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12667) );
  AOI21_X1 U15170 ( .B1(n13041), .B2(n13514), .A(n12667), .ZN(n12090) );
  INV_X1 U15171 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20074) );
  NOR2_X1 U15172 ( .A1(n13381), .A2(n20074), .ZN(n12195) );
  NAND2_X1 U15173 ( .A1(n12195), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n12089) );
  OAI211_X1 U15174 ( .C1(n12107), .C2(n12091), .A(n12090), .B(n12089), .ZN(
        n12092) );
  INV_X1 U15175 ( .A(n12092), .ZN(n12093) );
  NAND2_X1 U15176 ( .A1(n12667), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12112) );
  NAND2_X1 U15177 ( .A1(n12094), .A2(n12112), .ZN(n13072) );
  INV_X1 U15178 ( .A(n13072), .ZN(n12111) );
  INV_X1 U15179 ( .A(n12095), .ZN(n12097) );
  INV_X1 U15180 ( .A(n12752), .ZN(n12096) );
  NAND2_X1 U15181 ( .A1(n13595), .A2(n12336), .ZN(n12101) );
  AOI22_X1 U15182 ( .A1(n12195), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20074), .ZN(n12099) );
  INV_X1 U15183 ( .A(n12107), .ZN(n12155) );
  NAND2_X1 U15184 ( .A1(n12155), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12098) );
  AND2_X1 U15185 ( .A1(n12099), .A2(n12098), .ZN(n12100) );
  NAND2_X1 U15186 ( .A1(n12101), .A2(n12100), .ZN(n13038) );
  NAND2_X1 U15187 ( .A1(n12758), .A2(n20104), .ZN(n12103) );
  NAND2_X1 U15188 ( .A1(n12103), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13286) );
  NAND2_X1 U15189 ( .A1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20074), .ZN(
        n12106) );
  NAND2_X1 U15190 ( .A1(n12195), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n12105) );
  OAI211_X1 U15191 ( .C1(n12107), .C2(n11846), .A(n12106), .B(n12105), .ZN(
        n12108) );
  AOI21_X1 U15192 ( .B1(n20195), .B2(n12336), .A(n12108), .ZN(n13287) );
  OR2_X1 U15193 ( .A1(n13286), .A2(n13287), .ZN(n13284) );
  NAND2_X1 U15194 ( .A1(n13287), .A2(n13041), .ZN(n12109) );
  NAND2_X1 U15195 ( .A1(n13284), .A2(n12109), .ZN(n13037) );
  NAND2_X1 U15196 ( .A1(n13038), .A2(n13037), .ZN(n13075) );
  NAND2_X1 U15197 ( .A1(n12111), .A2(n12110), .ZN(n13073) );
  INV_X1 U15198 ( .A(n12135), .ZN(n12133) );
  NAND2_X1 U15199 ( .A1(n12006), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12118) );
  NOR3_X1 U15200 ( .A1(n20507), .A2(n12676), .A3(n20429), .ZN(n20631) );
  INV_X1 U15201 ( .A(n20631), .ZN(n20619) );
  NOR2_X1 U15202 ( .A1(n20773), .A2(n20619), .ZN(n20675) );
  NAND3_X1 U15203 ( .A1(n20507), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20327) );
  NOR2_X1 U15204 ( .A1(n20773), .A2(n20327), .ZN(n20351) );
  NOR2_X1 U15205 ( .A1(n20351), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12114) );
  OR2_X1 U15206 ( .A1(n20675), .A2(n12114), .ZN(n20358) );
  OAI22_X1 U15207 ( .A1(n20358), .A2(n12860), .B1(n12115), .B2(n20507), .ZN(
        n12116) );
  INV_X1 U15208 ( .A(n12116), .ZN(n12117) );
  XNOR2_X2 U15209 ( .A(n13588), .B(n20234), .ZN(n20357) );
  AOI22_X1 U15210 ( .A1(n12641), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12396), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12124) );
  AOI22_X1 U15211 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12123) );
  AOI22_X1 U15212 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12122) );
  AOI22_X1 U15213 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12121) );
  NAND4_X1 U15214 ( .A1(n12124), .A2(n12123), .A3(n12122), .A4(n12121), .ZN(
        n12130) );
  AOI22_X1 U15215 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12634), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12128) );
  AOI22_X1 U15216 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12127) );
  AOI22_X1 U15217 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12126) );
  INV_X1 U15218 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n20897) );
  AOI22_X1 U15219 ( .A1(n12571), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12125) );
  NAND4_X1 U15220 ( .A1(n12128), .A2(n12127), .A3(n12126), .A4(n12125), .ZN(
        n12129) );
  OR2_X1 U15221 ( .A1(n12130), .A2(n12129), .ZN(n12789) );
  AOI22_X1 U15222 ( .A1(n12714), .A2(n12789), .B1(n12723), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12131) );
  NAND2_X1 U15223 ( .A1(n12135), .A2(n13625), .ZN(n12136) );
  INV_X1 U15224 ( .A(n12195), .ZN(n12137) );
  NAND2_X1 U15225 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12138) );
  AOI21_X1 U15226 ( .B1(n19895), .B2(n12138), .A(n12176), .ZN(n19908) );
  INV_X1 U15227 ( .A(n12667), .ZN(n12374) );
  OAI22_X1 U15228 ( .A1(n19908), .A2(n12658), .B1(n12374), .B2(n19895), .ZN(
        n12139) );
  AOI21_X1 U15229 ( .B1(n12668), .B2(P1_EAX_REG_3__SCAN_IN), .A(n12139), .ZN(
        n12141) );
  NAND2_X1 U15230 ( .A1(n12155), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12140) );
  NAND2_X1 U15231 ( .A1(n13535), .A2(n13536), .ZN(n13613) );
  AOI22_X1 U15232 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12643), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12145) );
  AOI22_X1 U15233 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12144) );
  AOI22_X1 U15234 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12143) );
  AOI22_X1 U15235 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12142) );
  NAND4_X1 U15236 ( .A1(n12145), .A2(n12144), .A3(n12143), .A4(n12142), .ZN(
        n12152) );
  AOI22_X1 U15237 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12048), .B1(
        n12634), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12150) );
  AOI22_X1 U15238 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12591), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12149) );
  AOI22_X1 U15239 ( .A1(n12641), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U15240 ( .A1(n12571), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12147) );
  NAND4_X1 U15241 ( .A1(n12150), .A2(n12149), .A3(n12148), .A4(n12147), .ZN(
        n12151) );
  OR2_X1 U15242 ( .A1(n12152), .A2(n12151), .ZN(n12788) );
  NAND2_X1 U15243 ( .A1(n12714), .A2(n12788), .ZN(n12154) );
  NAND2_X1 U15244 ( .A1(n12723), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12153) );
  NAND2_X1 U15245 ( .A1(n12154), .A2(n12153), .ZN(n12162) );
  XNOR2_X1 U15246 ( .A(n12161), .B(n12162), .ZN(n12780) );
  NAND2_X1 U15247 ( .A1(n12155), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12159) );
  INV_X1 U15248 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13757) );
  AOI21_X1 U15249 ( .B1(n13757), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12156) );
  AOI21_X1 U15250 ( .B1(n12668), .B2(P1_EAX_REG_4__SCAN_IN), .A(n12156), .ZN(
        n12158) );
  XNOR2_X1 U15251 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B(n12176), .ZN(
        n19994) );
  NOR2_X1 U15252 ( .A1(n19994), .A2(n12658), .ZN(n12157) );
  AOI21_X1 U15253 ( .B1(n12159), .B2(n12158), .A(n12157), .ZN(n12160) );
  AOI21_X1 U15254 ( .B1(n12780), .B2(n12336), .A(n12160), .ZN(n13614) );
  INV_X1 U15255 ( .A(n12161), .ZN(n12163) );
  AOI22_X1 U15256 ( .A1(n12641), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12396), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12167) );
  AOI22_X1 U15257 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12166) );
  AOI22_X1 U15258 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12165) );
  AOI22_X1 U15259 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12164) );
  NAND4_X1 U15260 ( .A1(n12167), .A2(n12166), .A3(n12165), .A4(n12164), .ZN(
        n12173) );
  AOI22_X1 U15261 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12634), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12171) );
  AOI22_X1 U15262 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12170) );
  AOI22_X1 U15263 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12169) );
  INV_X1 U15264 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20103) );
  AOI22_X1 U15265 ( .A1(n12571), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12168) );
  NAND4_X1 U15266 ( .A1(n12171), .A2(n12170), .A3(n12169), .A4(n12168), .ZN(
        n12172) );
  OR2_X1 U15267 ( .A1(n12173), .A2(n12172), .ZN(n12800) );
  NAND2_X1 U15268 ( .A1(n12714), .A2(n12800), .ZN(n12175) );
  NAND2_X1 U15269 ( .A1(n12723), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12174) );
  NAND2_X1 U15270 ( .A1(n12175), .A2(n12174), .ZN(n12184) );
  XNOR2_X1 U15271 ( .A(n12183), .B(n12184), .ZN(n12787) );
  NAND2_X1 U15272 ( .A1(n12787), .A2(n12336), .ZN(n12182) );
  INV_X1 U15273 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19880) );
  INV_X1 U15274 ( .A(n12196), .ZN(n12198) );
  NAND2_X1 U15275 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n12176), .ZN(
        n12177) );
  NAND2_X1 U15276 ( .A1(n19880), .A2(n12177), .ZN(n12178) );
  NAND2_X1 U15277 ( .A1(n12198), .A2(n12178), .ZN(n19891) );
  NAND2_X1 U15278 ( .A1(n19891), .A2(n13041), .ZN(n12179) );
  OAI21_X1 U15279 ( .B1(n19880), .B2(n12374), .A(n12179), .ZN(n12180) );
  AOI21_X1 U15280 ( .B1(n12668), .B2(P1_EAX_REG_5__SCAN_IN), .A(n12180), .ZN(
        n12181) );
  NAND2_X1 U15281 ( .A1(n13607), .A2(n13608), .ZN(n13606) );
  INV_X1 U15282 ( .A(n13606), .ZN(n12204) );
  AOI22_X1 U15283 ( .A1(n12641), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12634), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12188) );
  AOI22_X1 U15284 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12396), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12187) );
  AOI22_X1 U15285 ( .A1(n12633), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12186) );
  AOI22_X1 U15286 ( .A1(n12571), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12185) );
  NAND4_X1 U15287 ( .A1(n12188), .A2(n12187), .A3(n12186), .A4(n12185), .ZN(
        n12194) );
  AOI22_X1 U15288 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12192) );
  AOI22_X1 U15289 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12191) );
  AOI22_X1 U15290 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12190) );
  AOI22_X1 U15291 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12189) );
  NAND4_X1 U15292 ( .A1(n12192), .A2(n12191), .A3(n12190), .A4(n12189), .ZN(
        n12193) );
  OR2_X1 U15293 ( .A1(n12194), .A2(n12193), .ZN(n12809) );
  AOI22_X1 U15294 ( .A1(n12714), .A2(n12809), .B1(n12723), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12206) );
  NAND2_X1 U15295 ( .A1(n12205), .A2(n12206), .ZN(n12797) );
  INV_X1 U15296 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n19933) );
  INV_X1 U15297 ( .A(n12210), .ZN(n12200) );
  INV_X1 U15298 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12197) );
  NAND2_X1 U15299 ( .A1(n12198), .A2(n12197), .ZN(n12199) );
  NAND2_X1 U15300 ( .A1(n12200), .A2(n12199), .ZN(n19868) );
  AOI22_X1 U15301 ( .A1(n19868), .A2(n13041), .B1(n12667), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12201) );
  OAI21_X1 U15302 ( .B1(n12137), .B2(n19933), .A(n12201), .ZN(n12202) );
  INV_X1 U15303 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n20118) );
  NAND2_X1 U15304 ( .A1(n12714), .A2(n12811), .ZN(n12208) );
  OAI21_X1 U15305 ( .B1(n20118), .B2(n12718), .A(n12208), .ZN(n12209) );
  INV_X1 U15306 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n12212) );
  OAI21_X1 U15307 ( .B1(n12210), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n12214), .ZN(n19855) );
  AOI22_X1 U15308 ( .A1(n19855), .A2(n13041), .B1(n12667), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12211) );
  OAI21_X1 U15309 ( .B1(n12137), .B2(n12212), .A(n12211), .ZN(n12213) );
  AOI21_X1 U15310 ( .B1(n12814), .B2(n12336), .A(n12213), .ZN(n13675) );
  INV_X1 U15311 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12245) );
  XOR2_X1 U15312 ( .A(n12245), .B(n12246), .Z(n19842) );
  INV_X1 U15313 ( .A(n19842), .ZN(n12229) );
  AOI22_X1 U15314 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12218) );
  AOI22_X1 U15315 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12217) );
  AOI22_X1 U15316 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12216) );
  AOI22_X1 U15317 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12215) );
  NAND4_X1 U15318 ( .A1(n12218), .A2(n12217), .A3(n12216), .A4(n12215), .ZN(
        n12224) );
  AOI22_X1 U15319 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12048), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12222) );
  AOI22_X1 U15320 ( .A1(n12570), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12221) );
  AOI22_X1 U15321 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12220) );
  AOI22_X1 U15322 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12219) );
  NAND4_X1 U15323 ( .A1(n12222), .A2(n12221), .A3(n12220), .A4(n12219), .ZN(
        n12223) );
  OAI21_X1 U15324 ( .B1(n12224), .B2(n12223), .A(n12336), .ZN(n12227) );
  NAND2_X1 U15325 ( .A1(n12668), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12226) );
  NAND2_X1 U15326 ( .A1(n12667), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12225) );
  NAND3_X1 U15327 ( .A1(n12227), .A2(n12226), .A3(n12225), .ZN(n12228) );
  AOI21_X1 U15328 ( .B1(n12229), .B2(n13041), .A(n12228), .ZN(n13905) );
  AOI22_X1 U15329 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12233) );
  AOI22_X1 U15330 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12232) );
  AOI22_X1 U15331 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12231) );
  AOI22_X1 U15332 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12230) );
  NAND4_X1 U15333 ( .A1(n12233), .A2(n12232), .A3(n12231), .A4(n12230), .ZN(
        n12239) );
  AOI22_X1 U15334 ( .A1(n12570), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12634), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12237) );
  AOI22_X1 U15335 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12236) );
  AOI22_X1 U15336 ( .A1(n12646), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12235) );
  AOI22_X1 U15337 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12234) );
  NAND4_X1 U15338 ( .A1(n12237), .A2(n12236), .A3(n12235), .A4(n12234), .ZN(
        n12238) );
  OAI21_X1 U15339 ( .B1(n12239), .B2(n12238), .A(n12336), .ZN(n12243) );
  XNOR2_X1 U15340 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n12240), .ZN(
        n13914) );
  AOI22_X1 U15341 ( .A1(n13041), .A2(n13914), .B1(n12667), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12242) );
  NAND2_X1 U15342 ( .A1(n12668), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12241) );
  AND3_X1 U15343 ( .A1(n12243), .A2(n12242), .A3(n12241), .ZN(n13876) );
  NOR2_X1 U15344 ( .A1(n13905), .A2(n13876), .ZN(n12244) );
  INV_X1 U15345 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15606) );
  XNOR2_X1 U15346 ( .A(n12262), .B(n15606), .ZN(n15604) );
  OR2_X1 U15347 ( .A1(n15604), .A2(n12658), .ZN(n12261) );
  AOI22_X1 U15348 ( .A1(n12570), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12250) );
  AOI22_X1 U15349 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12249) );
  AOI22_X1 U15350 ( .A1(n12646), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12248) );
  AOI22_X1 U15351 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12247) );
  NAND4_X1 U15352 ( .A1(n12250), .A2(n12249), .A3(n12248), .A4(n12247), .ZN(
        n12256) );
  AOI22_X1 U15353 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12396), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12254) );
  AOI22_X1 U15354 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12634), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U15355 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U15356 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12251) );
  NAND4_X1 U15357 ( .A1(n12254), .A2(n12253), .A3(n12252), .A4(n12251), .ZN(
        n12255) );
  OAI21_X1 U15358 ( .B1(n12256), .B2(n12255), .A(n12336), .ZN(n12259) );
  NAND2_X1 U15359 ( .A1(n12668), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n12258) );
  NAND2_X1 U15360 ( .A1(n12667), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12257) );
  AND3_X1 U15361 ( .A1(n12259), .A2(n12258), .A3(n12257), .ZN(n12260) );
  NAND2_X1 U15362 ( .A1(n12261), .A2(n12260), .ZN(n13834) );
  INV_X1 U15363 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12265) );
  OAI21_X1 U15364 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12263), .A(
        n12303), .ZN(n15659) );
  NAND2_X1 U15365 ( .A1(n15659), .A2(n13041), .ZN(n12264) );
  OAI21_X1 U15366 ( .B1(n12265), .B2(n12374), .A(n12264), .ZN(n12266) );
  AOI21_X1 U15367 ( .B1(n12668), .B2(P1_EAX_REG_11__SCAN_IN), .A(n12266), .ZN(
        n13967) );
  AOI22_X1 U15368 ( .A1(n12469), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12048), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12270) );
  AOI22_X1 U15369 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12269) );
  AOI22_X1 U15370 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12268) );
  AOI22_X1 U15371 ( .A1(n12571), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12267) );
  NAND4_X1 U15372 ( .A1(n12270), .A2(n12269), .A3(n12268), .A4(n12267), .ZN(
        n12276) );
  AOI22_X1 U15373 ( .A1(n12570), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12396), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U15374 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12273) );
  AOI22_X1 U15375 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U15376 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12271) );
  NAND4_X1 U15377 ( .A1(n12274), .A2(n12273), .A3(n12272), .A4(n12271), .ZN(
        n12275) );
  OR2_X1 U15378 ( .A1(n12276), .A2(n12275), .ZN(n12277) );
  NAND2_X1 U15379 ( .A1(n12336), .A2(n12277), .ZN(n14008) );
  INV_X1 U15380 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n13979) );
  AOI22_X1 U15381 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12331), .B1(
        n12570), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12281) );
  AOI22_X1 U15382 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12280) );
  AOI22_X1 U15383 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12279) );
  AOI22_X1 U15384 ( .A1(n12571), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12278) );
  NAND4_X1 U15385 ( .A1(n12281), .A2(n12280), .A3(n12279), .A4(n12278), .ZN(
        n12287) );
  AOI22_X1 U15386 ( .A1(n12469), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12285) );
  AOI22_X1 U15387 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12284) );
  AOI22_X1 U15388 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12634), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12283) );
  AOI22_X1 U15389 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12048), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12282) );
  NAND4_X1 U15390 ( .A1(n12285), .A2(n12284), .A3(n12283), .A4(n12282), .ZN(
        n12286) );
  OAI21_X1 U15391 ( .B1(n12287), .B2(n12286), .A(n12336), .ZN(n12291) );
  XNOR2_X1 U15392 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12303), .ZN(
        n15646) );
  INV_X1 U15393 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12288) );
  OAI22_X1 U15394 ( .A1(n15646), .A2(n12658), .B1(n12374), .B2(n12288), .ZN(
        n12289) );
  INV_X1 U15395 ( .A(n12289), .ZN(n12290) );
  OAI211_X1 U15396 ( .C1(n12137), .C2(n13979), .A(n12291), .B(n12290), .ZN(
        n13975) );
  AOI22_X1 U15397 ( .A1(n12469), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12643), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12295) );
  AOI22_X1 U15398 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12634), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12294) );
  AOI22_X1 U15399 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12146), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12293) );
  AOI22_X1 U15400 ( .A1(n12633), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12066), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12292) );
  NAND4_X1 U15401 ( .A1(n12295), .A2(n12294), .A3(n12293), .A4(n12292), .ZN(
        n12302) );
  AOI22_X1 U15402 ( .A1(n12570), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12645), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12300) );
  AOI22_X1 U15403 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12299) );
  AOI22_X1 U15404 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U15405 ( .A1(n12401), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12297) );
  NAND4_X1 U15406 ( .A1(n12300), .A2(n12299), .A3(n12298), .A4(n12297), .ZN(
        n12301) );
  NOR2_X1 U15407 ( .A1(n12302), .A2(n12301), .ZN(n12310) );
  INV_X1 U15408 ( .A(n12305), .ZN(n12307) );
  INV_X1 U15409 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n20874) );
  INV_X1 U15410 ( .A(n12339), .ZN(n12306) );
  OAI21_X1 U15411 ( .B1(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n12307), .A(
        n12306), .ZN(n13985) );
  AOI22_X1 U15412 ( .A1(n13041), .A2(n13985), .B1(n12667), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12309) );
  NAND2_X1 U15413 ( .A1(n12668), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12308) );
  OAI211_X1 U15414 ( .C1(n12311), .C2(n12310), .A(n12309), .B(n12308), .ZN(
        n13971) );
  NAND2_X1 U15415 ( .A1(n13975), .A2(n13971), .ZN(n12312) );
  INV_X1 U15416 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14006) );
  AOI22_X1 U15417 ( .A1(n12570), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12396), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12317) );
  AOI22_X1 U15418 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12316) );
  AOI22_X1 U15419 ( .A1(n12571), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12315) );
  AOI22_X1 U15420 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12314) );
  NAND4_X1 U15421 ( .A1(n12317), .A2(n12316), .A3(n12315), .A4(n12314), .ZN(
        n12323) );
  AOI22_X1 U15422 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12634), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12321) );
  AOI22_X1 U15423 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12320) );
  AOI22_X1 U15424 ( .A1(n12469), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12066), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12319) );
  AOI22_X1 U15425 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12022), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12318) );
  NAND4_X1 U15426 ( .A1(n12321), .A2(n12320), .A3(n12319), .A4(n12318), .ZN(
        n12322) );
  OAI21_X1 U15427 ( .B1(n12323), .B2(n12322), .A(n12336), .ZN(n12326) );
  XOR2_X1 U15428 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n12339), .Z(
        n15640) );
  INV_X1 U15429 ( .A(n15640), .ZN(n12324) );
  AOI22_X1 U15430 ( .A1(n12667), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n13041), .B2(n12324), .ZN(n12325) );
  OAI211_X1 U15431 ( .C1(n12137), .C2(n14006), .A(n12326), .B(n12325), .ZN(
        n13999) );
  NAND2_X1 U15432 ( .A1(n13970), .A2(n13999), .ZN(n14000) );
  AOI22_X1 U15433 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12330) );
  AOI22_X1 U15434 ( .A1(n12469), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12329) );
  AOI22_X1 U15435 ( .A1(n12571), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12328) );
  AOI22_X1 U15436 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12327) );
  NAND4_X1 U15437 ( .A1(n12330), .A2(n12329), .A3(n12328), .A4(n12327), .ZN(
        n12338) );
  AOI22_X1 U15438 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12570), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12335) );
  AOI22_X1 U15439 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12634), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12334) );
  AOI22_X1 U15440 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12333) );
  AOI22_X1 U15441 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12066), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12332) );
  NAND4_X1 U15442 ( .A1(n12335), .A2(n12334), .A3(n12333), .A4(n12332), .ZN(
        n12337) );
  OAI21_X1 U15443 ( .B1(n12338), .B2(n12337), .A(n12336), .ZN(n12343) );
  NAND2_X1 U15444 ( .A1(n12339), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12358) );
  INV_X1 U15445 ( .A(n12358), .ZN(n12340) );
  XNOR2_X1 U15446 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n12340), .ZN(
        n14573) );
  AOI22_X1 U15447 ( .A1(n13041), .A2(n14573), .B1(n12667), .B2(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12342) );
  NAND2_X1 U15448 ( .A1(n12668), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12341) );
  AND3_X1 U15449 ( .A1(n12343), .A2(n12342), .A3(n12341), .ZN(n14024) );
  NAND2_X1 U15450 ( .A1(n13427), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12661) );
  AOI22_X1 U15451 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12048), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12347) );
  AOI22_X1 U15452 ( .A1(n12469), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12503), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12346) );
  AOI22_X1 U15453 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12345) );
  AOI22_X1 U15454 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12066), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12344) );
  NAND4_X1 U15455 ( .A1(n12347), .A2(n12346), .A3(n12345), .A4(n12344), .ZN(
        n12353) );
  AOI22_X1 U15456 ( .A1(n12570), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12351) );
  AOI22_X1 U15457 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12350) );
  AOI22_X1 U15458 ( .A1(n12571), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12349) );
  AOI22_X1 U15459 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12348) );
  NAND4_X1 U15460 ( .A1(n12351), .A2(n12350), .A3(n12349), .A4(n12348), .ZN(
        n12352) );
  NOR2_X1 U15461 ( .A1(n12353), .A2(n12352), .ZN(n12357) );
  NAND2_X1 U15462 ( .A1(n20074), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12354) );
  NAND2_X1 U15463 ( .A1(n12658), .A2(n12354), .ZN(n12355) );
  AOI21_X1 U15464 ( .B1(n12668), .B2(P1_EAX_REG_16__SCAN_IN), .A(n12355), .ZN(
        n12356) );
  OAI21_X1 U15465 ( .B1(n12661), .B2(n12357), .A(n12356), .ZN(n12361) );
  INV_X1 U15466 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n14033) );
  OAI21_X1 U15467 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12359), .A(
        n12392), .ZN(n15639) );
  OR2_X1 U15468 ( .A1(n12658), .A2(n15639), .ZN(n12360) );
  NAND2_X1 U15469 ( .A1(n12361), .A2(n12360), .ZN(n14052) );
  AOI22_X1 U15470 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12643), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12366) );
  AOI22_X1 U15471 ( .A1(n12570), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12645), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12365) );
  AOI22_X1 U15472 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12364) );
  AOI22_X1 U15473 ( .A1(n12642), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12066), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12363) );
  NAND4_X1 U15474 ( .A1(n12366), .A2(n12365), .A3(n12364), .A4(n12363), .ZN(
        n12372) );
  AOI22_X1 U15475 ( .A1(n12469), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12370) );
  AOI22_X1 U15476 ( .A1(n12571), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12369) );
  AOI22_X1 U15477 ( .A1(n12634), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12368) );
  AOI22_X1 U15478 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12022), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12367) );
  NAND4_X1 U15479 ( .A1(n12370), .A2(n12369), .A3(n12368), .A4(n12367), .ZN(
        n12371) );
  OR2_X1 U15480 ( .A1(n12372), .A2(n12371), .ZN(n12373) );
  NAND2_X1 U15481 ( .A1(n12626), .A2(n12373), .ZN(n12377) );
  XNOR2_X1 U15482 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12392), .ZN(
        n14564) );
  INV_X1 U15483 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14560) );
  OAI22_X1 U15484 ( .A1(n12658), .A2(n14564), .B1(n12374), .B2(n14560), .ZN(
        n12375) );
  AOI21_X1 U15485 ( .B1(n12668), .B2(P1_EAX_REG_17__SCAN_IN), .A(n12375), .ZN(
        n12376) );
  NAND2_X1 U15486 ( .A1(n12377), .A2(n12376), .ZN(n14349) );
  AOI22_X1 U15487 ( .A1(n12570), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11892), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12381) );
  AOI22_X1 U15488 ( .A1(n12469), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12634), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12380) );
  AOI22_X1 U15489 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12571), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12379) );
  AOI22_X1 U15490 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12378) );
  NAND4_X1 U15491 ( .A1(n12381), .A2(n12380), .A3(n12379), .A4(n12378), .ZN(
        n12387) );
  AOI22_X1 U15492 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12385) );
  AOI22_X1 U15493 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12066), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12384) );
  AOI22_X1 U15494 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12644), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12383) );
  AOI22_X1 U15495 ( .A1(n12646), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12382) );
  NAND4_X1 U15496 ( .A1(n12385), .A2(n12384), .A3(n12383), .A4(n12382), .ZN(
        n12386) );
  NOR2_X1 U15497 ( .A1(n12387), .A2(n12386), .ZN(n12391) );
  NAND2_X1 U15498 ( .A1(n20074), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12388) );
  NAND2_X1 U15499 ( .A1(n12658), .A2(n12388), .ZN(n12389) );
  AOI21_X1 U15500 ( .B1(n12668), .B2(P1_EAX_REG_18__SCAN_IN), .A(n12389), .ZN(
        n12390) );
  OAI21_X1 U15501 ( .B1(n12661), .B2(n12391), .A(n12390), .ZN(n12395) );
  OAI21_X1 U15502 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12393), .A(
        n12465), .ZN(n15556) );
  OR2_X1 U15503 ( .A1(n12658), .A2(n15556), .ZN(n12394) );
  AND2_X1 U15504 ( .A1(n12395), .A2(n12394), .ZN(n14393) );
  AOI22_X1 U15505 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12643), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12400) );
  AOI22_X1 U15506 ( .A1(n12634), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12396), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12399) );
  AOI22_X1 U15507 ( .A1(n12633), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12398) );
  AOI22_X1 U15508 ( .A1(n12571), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12397) );
  NAND4_X1 U15509 ( .A1(n12400), .A2(n12399), .A3(n12398), .A4(n12397), .ZN(
        n12407) );
  AOI22_X1 U15510 ( .A1(n12570), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12405) );
  AOI22_X1 U15511 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12404) );
  AOI22_X1 U15512 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12403) );
  AOI22_X1 U15513 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12402) );
  NAND4_X1 U15514 ( .A1(n12405), .A2(n12404), .A3(n12403), .A4(n12402), .ZN(
        n12406) );
  NOR2_X1 U15515 ( .A1(n12407), .A2(n12406), .ZN(n12411) );
  NAND2_X1 U15516 ( .A1(n20074), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12408) );
  NAND2_X1 U15517 ( .A1(n12658), .A2(n12408), .ZN(n12409) );
  AOI21_X1 U15518 ( .B1(n12668), .B2(P1_EAX_REG_22__SCAN_IN), .A(n12409), .ZN(
        n12410) );
  OAI21_X1 U15519 ( .B1(n12661), .B2(n12411), .A(n12410), .ZN(n12418) );
  INV_X1 U15520 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14528) );
  INV_X1 U15521 ( .A(n12413), .ZN(n12415) );
  INV_X1 U15522 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12414) );
  NAND2_X1 U15523 ( .A1(n12415), .A2(n12414), .ZN(n12416) );
  NAND2_X1 U15524 ( .A1(n12514), .A2(n12416), .ZN(n15630) );
  OR2_X1 U15525 ( .A1(n15630), .A2(n12658), .ZN(n12417) );
  AND2_X1 U15526 ( .A1(n12418), .A2(n12417), .ZN(n14442) );
  AOI22_X1 U15527 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11892), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12422) );
  AOI22_X1 U15528 ( .A1(n12570), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12645), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12421) );
  AOI22_X1 U15529 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12420) );
  AOI22_X1 U15530 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12419) );
  NAND4_X1 U15531 ( .A1(n12422), .A2(n12421), .A3(n12420), .A4(n12419), .ZN(
        n12428) );
  AOI22_X1 U15532 ( .A1(n12469), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12426) );
  AOI22_X1 U15533 ( .A1(n12634), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12066), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12425) );
  AOI22_X1 U15534 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12424) );
  AOI22_X1 U15535 ( .A1(n12571), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12022), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12423) );
  NAND4_X1 U15536 ( .A1(n12426), .A2(n12425), .A3(n12424), .A4(n12423), .ZN(
        n12427) );
  NOR2_X1 U15537 ( .A1(n12428), .A2(n12427), .ZN(n12431) );
  AOI21_X1 U15538 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14528), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12429) );
  AOI21_X1 U15539 ( .B1(n12668), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12429), .ZN(
        n12430) );
  OAI21_X1 U15540 ( .B1(n12661), .B2(n12431), .A(n12430), .ZN(n12433) );
  XNOR2_X1 U15541 ( .A(n12448), .B(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15536) );
  NAND2_X1 U15542 ( .A1(n15536), .A2(n13041), .ZN(n12432) );
  NAND2_X1 U15543 ( .A1(n12433), .A2(n12432), .ZN(n14448) );
  AOI22_X1 U15544 ( .A1(n12469), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12570), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12437) );
  AOI22_X1 U15545 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12643), .B1(
        n12503), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12436) );
  AOI22_X1 U15546 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12048), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12435) );
  AOI22_X1 U15547 ( .A1(n12571), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12022), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12434) );
  NAND4_X1 U15548 ( .A1(n12437), .A2(n12436), .A3(n12435), .A4(n12434), .ZN(
        n12443) );
  AOI22_X1 U15549 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12441) );
  AOI22_X1 U15550 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12440) );
  AOI22_X1 U15551 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12331), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12439) );
  AOI22_X1 U15552 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12438) );
  NAND4_X1 U15553 ( .A1(n12441), .A2(n12440), .A3(n12439), .A4(n12438), .ZN(
        n12442) );
  NOR2_X1 U15554 ( .A1(n12443), .A2(n12442), .ZN(n12447) );
  NAND2_X1 U15555 ( .A1(n20074), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12444) );
  NAND2_X1 U15556 ( .A1(n12658), .A2(n12444), .ZN(n12445) );
  AOI21_X1 U15557 ( .B1(n12668), .B2(P1_EAX_REG_20__SCAN_IN), .A(n12445), .ZN(
        n12446) );
  OAI21_X1 U15558 ( .B1(n12661), .B2(n12447), .A(n12446), .ZN(n12451) );
  OAI21_X1 U15559 ( .B1(n12449), .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n12448), .ZN(n15553) );
  OR2_X1 U15560 ( .A1(n15553), .A2(n12658), .ZN(n12450) );
  NAND2_X1 U15561 ( .A1(n12451), .A2(n12450), .ZN(n14385) );
  AOI22_X1 U15562 ( .A1(n12570), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12645), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12455) );
  AOI22_X1 U15563 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12048), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12454) );
  AOI22_X1 U15564 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12453) );
  AOI22_X1 U15565 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12452) );
  NAND4_X1 U15566 ( .A1(n12455), .A2(n12454), .A3(n12453), .A4(n12452), .ZN(
        n12461) );
  AOI22_X1 U15567 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12571), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12459) );
  AOI22_X1 U15568 ( .A1(n12469), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12458) );
  AOI22_X1 U15569 ( .A1(n12634), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12457) );
  AOI22_X1 U15570 ( .A1(n12066), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12456) );
  NAND4_X1 U15571 ( .A1(n12459), .A2(n12458), .A3(n12457), .A4(n12456), .ZN(
        n12460) );
  NOR2_X1 U15572 ( .A1(n12461), .A2(n12460), .ZN(n12464) );
  INV_X1 U15573 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14540) );
  OAI21_X1 U15574 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14540), .A(n12658), 
        .ZN(n12462) );
  AOI21_X1 U15575 ( .B1(n12668), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12462), .ZN(
        n12463) );
  OAI21_X1 U15576 ( .B1(n12661), .B2(n12464), .A(n12463), .ZN(n12467) );
  XNOR2_X1 U15577 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n12465), .ZN(
        n14544) );
  NAND2_X1 U15578 ( .A1(n13041), .A2(n14544), .ZN(n12466) );
  NAND2_X1 U15579 ( .A1(n12467), .A2(n12466), .ZN(n14384) );
  OR2_X1 U15580 ( .A1(n14385), .A2(n14384), .ZN(n14383) );
  NOR2_X1 U15581 ( .A1(n14448), .A2(n14383), .ZN(n14440) );
  AOI22_X1 U15582 ( .A1(n12570), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12645), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12473) );
  AOI22_X1 U15583 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12634), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12472) );
  AOI22_X1 U15584 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12471) );
  AOI22_X1 U15585 ( .A1(n12469), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12470) );
  NAND4_X1 U15586 ( .A1(n12473), .A2(n12472), .A3(n12471), .A4(n12470), .ZN(
        n12479) );
  AOI22_X1 U15587 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12477) );
  AOI22_X1 U15588 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12476) );
  AOI22_X1 U15589 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12475) );
  AOI22_X1 U15590 ( .A1(n12571), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12474) );
  NAND4_X1 U15591 ( .A1(n12477), .A2(n12476), .A3(n12475), .A4(n12474), .ZN(
        n12478) );
  NOR2_X1 U15592 ( .A1(n12479), .A2(n12478), .ZN(n12497) );
  AOI22_X1 U15593 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12483) );
  AOI22_X1 U15594 ( .A1(n12634), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12482) );
  AOI22_X1 U15595 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12481) );
  AOI22_X1 U15596 ( .A1(n12401), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12480) );
  NAND4_X1 U15597 ( .A1(n12483), .A2(n12482), .A3(n12481), .A4(n12480), .ZN(
        n12490) );
  AOI22_X1 U15598 ( .A1(n12641), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12591), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12488) );
  AOI22_X1 U15599 ( .A1(n12331), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12643), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12487) );
  AOI22_X1 U15600 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12571), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12486) );
  AOI22_X1 U15601 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12485) );
  NAND4_X1 U15602 ( .A1(n12488), .A2(n12487), .A3(n12486), .A4(n12485), .ZN(
        n12489) );
  NOR2_X1 U15603 ( .A1(n12490), .A2(n12489), .ZN(n12498) );
  XOR2_X1 U15604 ( .A(n12497), .B(n12498), .Z(n12491) );
  NAND2_X1 U15605 ( .A1(n12491), .A2(n12626), .ZN(n12494) );
  INV_X1 U15606 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15525) );
  OAI21_X1 U15607 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15525), .A(n12658), 
        .ZN(n12492) );
  AOI21_X1 U15608 ( .B1(n12668), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12492), .ZN(
        n12493) );
  NAND2_X1 U15609 ( .A1(n12494), .A2(n12493), .ZN(n12496) );
  XNOR2_X1 U15610 ( .A(n12514), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15515) );
  NAND2_X1 U15611 ( .A1(n15515), .A2(n13041), .ZN(n12495) );
  NAND2_X1 U15612 ( .A1(n12496), .A2(n12495), .ZN(n14373) );
  NOR2_X1 U15613 ( .A1(n12498), .A2(n12497), .ZN(n12524) );
  AOI22_X1 U15614 ( .A1(n12641), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12396), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12502) );
  AOI22_X1 U15615 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12501) );
  AOI22_X1 U15616 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12500) );
  AOI22_X1 U15617 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12499) );
  NAND4_X1 U15618 ( .A1(n12502), .A2(n12501), .A3(n12500), .A4(n12499), .ZN(
        n12509) );
  AOI22_X1 U15619 ( .A1(n12067), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12503), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12507) );
  INV_X1 U15620 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n20084) );
  AOI22_X1 U15621 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12506) );
  AOI22_X1 U15622 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12505) );
  AOI22_X1 U15623 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12504) );
  NAND4_X1 U15624 ( .A1(n12507), .A2(n12506), .A3(n12505), .A4(n12504), .ZN(
        n12508) );
  OR2_X1 U15625 ( .A1(n12509), .A2(n12508), .ZN(n12523) );
  INV_X1 U15626 ( .A(n12523), .ZN(n12510) );
  XNOR2_X1 U15627 ( .A(n12524), .B(n12510), .ZN(n12513) );
  INV_X1 U15628 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14427) );
  NAND2_X1 U15629 ( .A1(n20074), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12511) );
  OAI211_X1 U15630 ( .C1(n12137), .C2(n14427), .A(n12658), .B(n12511), .ZN(
        n12512) );
  AOI21_X1 U15631 ( .B1(n12513), .B2(n12626), .A(n12512), .ZN(n12521) );
  INV_X1 U15632 ( .A(n12514), .ZN(n12515) );
  INV_X1 U15633 ( .A(n12516), .ZN(n12518) );
  INV_X1 U15634 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12517) );
  NAND2_X1 U15635 ( .A1(n12518), .A2(n12517), .ZN(n12519) );
  NAND2_X1 U15636 ( .A1(n12559), .A2(n12519), .ZN(n14515) );
  NOR2_X1 U15637 ( .A1(n14515), .A2(n12658), .ZN(n12520) );
  NAND2_X1 U15638 ( .A1(n12524), .A2(n12523), .ZN(n12541) );
  AOI22_X1 U15639 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12643), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12528) );
  AOI22_X1 U15640 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12635), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12527) );
  AOI22_X1 U15641 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12526) );
  AOI22_X1 U15642 ( .A1(n12634), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12525) );
  NAND4_X1 U15643 ( .A1(n12528), .A2(n12527), .A3(n12526), .A4(n12525), .ZN(
        n12534) );
  AOI22_X1 U15644 ( .A1(n12067), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12048), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12532) );
  AOI22_X1 U15645 ( .A1(n12641), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12531) );
  AOI22_X1 U15646 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12530) );
  AOI22_X1 U15647 ( .A1(n12633), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12529) );
  NAND4_X1 U15648 ( .A1(n12532), .A2(n12531), .A3(n12530), .A4(n12529), .ZN(
        n12533) );
  NOR2_X1 U15649 ( .A1(n12534), .A2(n12533), .ZN(n12542) );
  XOR2_X1 U15650 ( .A(n12541), .B(n12542), .Z(n12535) );
  NAND2_X1 U15651 ( .A1(n12535), .A2(n12626), .ZN(n12540) );
  NAND2_X1 U15652 ( .A1(n20074), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12536) );
  NAND2_X1 U15653 ( .A1(n12658), .A2(n12536), .ZN(n12537) );
  AOI21_X1 U15654 ( .B1(n12668), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12537), .ZN(
        n12539) );
  XNOR2_X1 U15655 ( .A(n12559), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14508) );
  AND2_X1 U15656 ( .A1(n14508), .A2(n13041), .ZN(n12538) );
  AOI21_X1 U15657 ( .B1(n12540), .B2(n12539), .A(n12538), .ZN(n14311) );
  NOR2_X1 U15658 ( .A1(n12542), .A2(n12541), .ZN(n12569) );
  AOI22_X1 U15659 ( .A1(n12641), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12396), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12548) );
  AOI22_X1 U15660 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12547) );
  AOI22_X1 U15661 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12546) );
  AOI22_X1 U15662 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12544), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12545) );
  NAND4_X1 U15663 ( .A1(n12548), .A2(n12547), .A3(n12546), .A4(n12545), .ZN(
        n12554) );
  AOI22_X1 U15664 ( .A1(n12067), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12634), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12552) );
  AOI22_X1 U15665 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12551) );
  AOI22_X1 U15666 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12550) );
  AOI22_X1 U15667 ( .A1(n12146), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12549) );
  NAND4_X1 U15668 ( .A1(n12552), .A2(n12551), .A3(n12550), .A4(n12549), .ZN(
        n12553) );
  OR2_X1 U15669 ( .A1(n12554), .A2(n12553), .ZN(n12568) );
  INV_X1 U15670 ( .A(n12568), .ZN(n12555) );
  XNOR2_X1 U15671 ( .A(n12569), .B(n12555), .ZN(n12556) );
  NAND2_X1 U15672 ( .A1(n12556), .A2(n12626), .ZN(n12567) );
  NAND2_X1 U15673 ( .A1(n20074), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12557) );
  NAND2_X1 U15674 ( .A1(n12658), .A2(n12557), .ZN(n12558) );
  AOI21_X1 U15675 ( .B1(n12668), .B2(P1_EAX_REG_26__SCAN_IN), .A(n12558), .ZN(
        n12566) );
  INV_X1 U15676 ( .A(n12559), .ZN(n12560) );
  INV_X1 U15677 ( .A(n12561), .ZN(n12563) );
  INV_X1 U15678 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12562) );
  NAND2_X1 U15679 ( .A1(n12563), .A2(n12562), .ZN(n12564) );
  NAND2_X1 U15680 ( .A1(n12606), .A2(n12564), .ZN(n14492) );
  NOR2_X1 U15681 ( .A1(n14492), .A2(n12658), .ZN(n12565) );
  AOI21_X1 U15682 ( .B1(n12567), .B2(n12566), .A(n12565), .ZN(n14292) );
  NAND2_X1 U15683 ( .A1(n12569), .A2(n12568), .ZN(n12589) );
  AOI22_X1 U15684 ( .A1(n12067), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12570), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12575) );
  AOI22_X1 U15685 ( .A1(n12634), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12571), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12574) );
  AOI22_X1 U15686 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12644), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12573) );
  AOI22_X1 U15687 ( .A1(n12633), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12572) );
  NAND4_X1 U15688 ( .A1(n12575), .A2(n12574), .A3(n12573), .A4(n12572), .ZN(
        n12581) );
  AOI22_X1 U15689 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12484), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12579) );
  AOI22_X1 U15690 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12578) );
  AOI22_X1 U15691 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12635), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12577) );
  AOI22_X1 U15692 ( .A1(n12614), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12022), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12576) );
  NAND4_X1 U15693 ( .A1(n12579), .A2(n12578), .A3(n12577), .A4(n12576), .ZN(
        n12580) );
  NOR2_X1 U15694 ( .A1(n12581), .A2(n12580), .ZN(n12590) );
  XOR2_X1 U15695 ( .A(n12589), .B(n12590), .Z(n12582) );
  NAND2_X1 U15696 ( .A1(n12582), .A2(n12626), .ZN(n12586) );
  NAND2_X1 U15697 ( .A1(n20074), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12583) );
  NAND2_X1 U15698 ( .A1(n12658), .A2(n12583), .ZN(n12584) );
  AOI21_X1 U15699 ( .B1(n12668), .B2(P1_EAX_REG_27__SCAN_IN), .A(n12584), .ZN(
        n12585) );
  NAND2_X1 U15700 ( .A1(n12586), .A2(n12585), .ZN(n12588) );
  XNOR2_X1 U15701 ( .A(n12606), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14485) );
  NAND2_X1 U15702 ( .A1(n14485), .A2(n13041), .ZN(n12587) );
  NAND2_X1 U15703 ( .A1(n12588), .A2(n12587), .ZN(n14284) );
  NOR2_X1 U15704 ( .A1(n12590), .A2(n12589), .ZN(n12613) );
  AOI22_X1 U15705 ( .A1(n12641), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12396), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12595) );
  AOI22_X1 U15706 ( .A1(n12591), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12594) );
  AOI22_X1 U15707 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12593) );
  AOI22_X1 U15708 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12644), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12592) );
  NAND4_X1 U15709 ( .A1(n12595), .A2(n12594), .A3(n12593), .A4(n12592), .ZN(
        n12601) );
  AOI22_X1 U15710 ( .A1(n12067), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12634), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12599) );
  AOI22_X1 U15711 ( .A1(n12614), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12598) );
  AOI22_X1 U15712 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12597) );
  AOI22_X1 U15713 ( .A1(n12571), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12022), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12596) );
  NAND4_X1 U15714 ( .A1(n12599), .A2(n12598), .A3(n12597), .A4(n12596), .ZN(
        n12600) );
  OR2_X1 U15715 ( .A1(n12601), .A2(n12600), .ZN(n12612) );
  INV_X1 U15716 ( .A(n12612), .ZN(n12602) );
  XNOR2_X1 U15717 ( .A(n12613), .B(n12602), .ZN(n12605) );
  INV_X1 U15718 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n14411) );
  NAND2_X1 U15719 ( .A1(n20074), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12603) );
  OAI211_X1 U15720 ( .C1(n12137), .C2(n14411), .A(n12658), .B(n12603), .ZN(
        n12604) );
  AOI21_X1 U15721 ( .B1(n12605), .B2(n12626), .A(n12604), .ZN(n12610) );
  INV_X1 U15722 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14487) );
  INV_X1 U15723 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14271) );
  NAND2_X1 U15724 ( .A1(n12607), .A2(n14271), .ZN(n12608) );
  NAND2_X1 U15725 ( .A1(n12663), .A2(n12608), .ZN(n14270) );
  NOR2_X1 U15726 ( .A1(n14270), .A2(n12658), .ZN(n12609) );
  AND2_X2 U15727 ( .A1(n12853), .A2(n12611), .ZN(n14213) );
  NAND2_X1 U15728 ( .A1(n12613), .A2(n12612), .ZN(n12653) );
  AOI22_X1 U15729 ( .A1(n12641), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12619) );
  AOI22_X1 U15730 ( .A1(n12067), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12634), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12618) );
  AOI22_X1 U15731 ( .A1(n12614), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12617) );
  AOI22_X1 U15732 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12615), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12616) );
  NAND4_X1 U15733 ( .A1(n12619), .A2(n12618), .A3(n12617), .A4(n12616), .ZN(
        n12625) );
  AOI22_X1 U15734 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12623) );
  AOI22_X1 U15735 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12622) );
  AOI22_X1 U15736 ( .A1(n12571), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12401), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12621) );
  AOI22_X1 U15737 ( .A1(n12635), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12644), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12620) );
  NAND4_X1 U15738 ( .A1(n12623), .A2(n12622), .A3(n12621), .A4(n12620), .ZN(
        n12624) );
  NOR2_X1 U15739 ( .A1(n12625), .A2(n12624), .ZN(n12654) );
  XOR2_X1 U15740 ( .A(n12653), .B(n12654), .Z(n12627) );
  NAND2_X1 U15741 ( .A1(n12627), .A2(n12626), .ZN(n12632) );
  NAND2_X1 U15742 ( .A1(n20074), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12628) );
  NAND2_X1 U15743 ( .A1(n12658), .A2(n12628), .ZN(n12629) );
  AOI21_X1 U15744 ( .B1(n12668), .B2(P1_EAX_REG_29__SCAN_IN), .A(n12629), .ZN(
        n12631) );
  XNOR2_X1 U15745 ( .A(n12663), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14263) );
  AND2_X1 U15746 ( .A1(n14263), .A2(n13041), .ZN(n12630) );
  AOI21_X1 U15747 ( .B1(n12632), .B2(n12631), .A(n12630), .ZN(n14212) );
  NAND2_X2 U15748 ( .A1(n14213), .A2(n14212), .ZN(n14241) );
  AOI22_X1 U15749 ( .A1(n12634), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12633), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12640) );
  AOI22_X1 U15750 ( .A1(n12571), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12639) );
  AOI22_X1 U15751 ( .A1(n12636), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12635), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12638) );
  AOI22_X1 U15752 ( .A1(n12401), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12022), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12637) );
  NAND4_X1 U15753 ( .A1(n12640), .A2(n12639), .A3(n12638), .A4(n12637), .ZN(
        n12652) );
  AOI22_X1 U15754 ( .A1(n12067), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12641), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12650) );
  AOI22_X1 U15755 ( .A1(n12643), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12642), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12649) );
  AOI22_X1 U15756 ( .A1(n12645), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12644), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12648) );
  AOI22_X1 U15757 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12646), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12647) );
  NAND4_X1 U15758 ( .A1(n12650), .A2(n12649), .A3(n12648), .A4(n12647), .ZN(
        n12651) );
  NOR2_X1 U15759 ( .A1(n12652), .A2(n12651), .ZN(n12656) );
  NOR2_X1 U15760 ( .A1(n12654), .A2(n12653), .ZN(n12655) );
  XOR2_X1 U15761 ( .A(n12656), .B(n12655), .Z(n12662) );
  NAND2_X1 U15762 ( .A1(n20074), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12657) );
  NAND2_X1 U15763 ( .A1(n12658), .A2(n12657), .ZN(n12659) );
  AOI21_X1 U15764 ( .B1(n12668), .B2(P1_EAX_REG_30__SCAN_IN), .A(n12659), .ZN(
        n12660) );
  OAI21_X1 U15765 ( .B1(n12662), .B2(n12661), .A(n12660), .ZN(n12666) );
  INV_X1 U15766 ( .A(n12663), .ZN(n12664) );
  NAND2_X1 U15767 ( .A1(n12664), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13045) );
  XNOR2_X1 U15768 ( .A(n13045), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14475) );
  NAND2_X1 U15769 ( .A1(n14475), .A2(n13041), .ZN(n12665) );
  NAND2_X1 U15770 ( .A1(n12666), .A2(n12665), .ZN(n14242) );
  NOR2_X2 U15771 ( .A1(n14241), .A2(n14242), .ZN(n12670) );
  AOI22_X1 U15772 ( .A1(n12668), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12667), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12669) );
  XNOR2_X1 U15773 ( .A(n12670), .B(n12669), .ZN(n14230) );
  AND3_X1 U15774 ( .A1(n20094), .A2(n20109), .A3(n12671), .ZN(n12672) );
  NAND2_X1 U15775 ( .A1(n12673), .A2(n12672), .ZN(n13293) );
  NAND2_X1 U15776 ( .A1(n20773), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12698) );
  MUX2_X1 U15777 ( .A(n20429), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        n12675), .Z(n12687) );
  OAI22_X1 U15778 ( .A1(n12698), .A2(n12687), .B1(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n12675), .ZN(n12689) );
  MUX2_X1 U15779 ( .A(n12676), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n12688) );
  NAND2_X1 U15780 ( .A1(n12689), .A2(n12688), .ZN(n12678) );
  NAND2_X1 U15781 ( .A1(n12676), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12677) );
  NAND2_X1 U15782 ( .A1(n12678), .A2(n12677), .ZN(n12686) );
  MUX2_X1 U15783 ( .A(n20507), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12685) );
  NAND2_X1 U15784 ( .A1(n12686), .A2(n12685), .ZN(n12680) );
  NAND2_X1 U15785 ( .A1(n20507), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12679) );
  NAND2_X1 U15786 ( .A1(n12680), .A2(n12679), .ZN(n12684) );
  INV_X1 U15787 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15799) );
  NOR2_X1 U15788 ( .A1(n15799), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n12681) );
  OR2_X1 U15789 ( .A1(n12684), .A2(n12681), .ZN(n12683) );
  INV_X1 U15790 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20058) );
  OR2_X1 U15791 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20058), .ZN(
        n12682) );
  INV_X1 U15792 ( .A(n12721), .ZN(n12722) );
  XNOR2_X1 U15793 ( .A(n12686), .B(n12685), .ZN(n12719) );
  XNOR2_X1 U15794 ( .A(n12698), .B(n12687), .ZN(n12704) );
  XNOR2_X1 U15795 ( .A(n12689), .B(n12688), .ZN(n12713) );
  NOR4_X1 U15796 ( .A1(n12722), .A2(n12719), .A3(n12704), .A4(n12713), .ZN(
        n12690) );
  NOR2_X1 U15797 ( .A1(n12694), .A2(n12690), .ZN(n13149) );
  NAND2_X1 U15798 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n20786) );
  NAND2_X1 U15799 ( .A1(n13149), .A2(n20786), .ZN(n12877) );
  OR2_X1 U15800 ( .A1(n15793), .A2(n12877), .ZN(n13441) );
  NAND2_X1 U15801 ( .A1(n15460), .A2(n20072), .ZN(n12691) );
  NAND4_X1 U15802 ( .A1(n20085), .A2(n13004), .A3(n12759), .A4(n12691), .ZN(
        n12851) );
  INV_X1 U15803 ( .A(n12851), .ZN(n12892) );
  NAND2_X1 U15804 ( .A1(n12892), .A2(n13126), .ZN(n13560) );
  NAND2_X1 U15805 ( .A1(n12692), .A2(n20786), .ZN(n12878) );
  OR2_X1 U15806 ( .A1(n12878), .A2(n13292), .ZN(n12693) );
  NAND2_X1 U15807 ( .A1(n13560), .A2(n12693), .ZN(n13435) );
  NAND2_X1 U15808 ( .A1(n13325), .A2(n11971), .ZN(n12779) );
  NAND2_X1 U15809 ( .A1(n12694), .A2(n12720), .ZN(n12729) );
  NAND2_X1 U15810 ( .A1(n12694), .A2(n12714), .ZN(n12728) );
  NOR2_X1 U15811 ( .A1(n11971), .A2(n20071), .ZN(n12695) );
  INV_X1 U15812 ( .A(n12706), .ZN(n12696) );
  NOR2_X1 U15813 ( .A1(n12704), .A2(n12696), .ZN(n12703) );
  AOI21_X1 U15814 ( .B1(n20099), .B2(n12697), .A(n13325), .ZN(n12716) );
  OAI21_X1 U15815 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20773), .A(
        n12698), .ZN(n12699) );
  AOI211_X1 U15816 ( .C1(n13000), .C2(n12697), .A(n12716), .B(n12699), .ZN(
        n12702) );
  INV_X1 U15817 ( .A(n12699), .ZN(n12700) );
  AOI21_X1 U15818 ( .B1(n12714), .B2(n12700), .A(n12720), .ZN(n12701) );
  NAND2_X1 U15819 ( .A1(n12703), .A2(n12705), .ZN(n12712) );
  NAND2_X1 U15820 ( .A1(n12706), .A2(n13325), .ZN(n12725) );
  OAI211_X1 U15821 ( .C1(n12706), .C2(n12705), .A(n12704), .B(n12725), .ZN(
        n12711) );
  INV_X1 U15822 ( .A(n12714), .ZN(n12709) );
  NAND2_X1 U15823 ( .A1(n12723), .A2(n12713), .ZN(n12708) );
  INV_X1 U15824 ( .A(n12716), .ZN(n12707) );
  OAI211_X1 U15825 ( .C1(n12709), .C2(n12713), .A(n12708), .B(n12707), .ZN(
        n12710) );
  INV_X1 U15826 ( .A(n12713), .ZN(n12715) );
  NAND3_X1 U15827 ( .A1(n12716), .A2(n12715), .A3(n12714), .ZN(n12717) );
  NAND2_X1 U15828 ( .A1(n12723), .A2(n12722), .ZN(n12724) );
  AOI21_X1 U15829 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20071), .A(
        n12726), .ZN(n12727) );
  NAND2_X1 U15830 ( .A1(n13435), .A2(n13434), .ZN(n12730) );
  OAI211_X1 U15831 ( .C1(n13140), .C2(n13293), .A(n13441), .B(n12730), .ZN(
        n12731) );
  OR2_X1 U15832 ( .A1(n20686), .A2(n20071), .ZN(n19815) );
  INV_X1 U15833 ( .A(n19815), .ZN(n13295) );
  AND2_X1 U15834 ( .A1(n14428), .A2(n20109), .ZN(n12732) );
  NAND2_X1 U15835 ( .A1(n14230), .A2(n12732), .ZN(n12749) );
  NAND2_X1 U15836 ( .A1(n14428), .A2(n13382), .ZN(n13387) );
  NOR4_X1 U15837 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n12736) );
  NOR4_X1 U15838 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_17__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n12735) );
  NOR4_X1 U15839 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12734) );
  NOR4_X1 U15840 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12733) );
  AND4_X1 U15841 ( .A1(n12736), .A2(n12735), .A3(n12734), .A4(n12733), .ZN(
        n12742) );
  NOR4_X1 U15842 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_11__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n12740) );
  NOR4_X1 U15843 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n12739) );
  NOR4_X1 U15844 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n12738) );
  INV_X1 U15845 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n12737) );
  AND4_X1 U15846 ( .A1(n12740), .A2(n12739), .A3(n12738), .A4(n12737), .ZN(
        n12741) );
  NAND2_X1 U15847 ( .A1(n12742), .A2(n12741), .ZN(n12743) );
  AND2_X2 U15848 ( .A1(n12743), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20068)
         );
  NOR2_X2 U15849 ( .A1(n13387), .A2(n20068), .ZN(n14471) );
  INV_X1 U15850 ( .A(n14428), .ZN(n14465) );
  AOI22_X1 U15851 ( .A1(n14471), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14465), .ZN(n12744) );
  INV_X1 U15852 ( .A(n12744), .ZN(n12747) );
  INV_X1 U15853 ( .A(n13387), .ZN(n12745) );
  NAND2_X1 U15854 ( .A1(n12745), .A2(n20068), .ZN(n14469) );
  INV_X1 U15855 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n19084) );
  NOR2_X1 U15856 ( .A1(n14469), .A2(n19084), .ZN(n12746) );
  NAND2_X1 U15857 ( .A1(n12749), .A2(n12748), .ZN(P1_U2873) );
  NOR2_X1 U15858 ( .A1(n12750), .A2(n12779), .ZN(n12751) );
  NAND3_X1 U15859 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14621) );
  INV_X1 U15860 ( .A(n14621), .ZN(n12841) );
  NAND2_X1 U15861 ( .A1(n12752), .A2(n13325), .ZN(n12757) );
  NAND2_X1 U15862 ( .A1(n12760), .A2(n12753), .ZN(n12775) );
  OAI21_X1 U15863 ( .B1(n12753), .B2(n12760), .A(n12775), .ZN(n12754) );
  OAI211_X1 U15864 ( .C1(n12754), .C2(n20789), .A(n20085), .B(n11971), .ZN(
        n12755) );
  INV_X1 U15865 ( .A(n12755), .ZN(n12756) );
  NAND2_X1 U15866 ( .A1(n20072), .A2(n12759), .ZN(n12767) );
  OAI21_X1 U15867 ( .B1(n20789), .B2(n12760), .A(n12767), .ZN(n12761) );
  INV_X1 U15868 ( .A(n12761), .ZN(n12762) );
  INV_X1 U15869 ( .A(n12764), .ZN(n12765) );
  OR2_X1 U15870 ( .A1(n13282), .A2(n12765), .ZN(n12766) );
  INV_X1 U15871 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20029) );
  OR2_X1 U15872 ( .A1(n13600), .A2(n12779), .ZN(n12771) );
  XNOR2_X1 U15873 ( .A(n12775), .B(n12774), .ZN(n12769) );
  INV_X1 U15874 ( .A(n12767), .ZN(n12768) );
  AOI21_X1 U15875 ( .B1(n12769), .B2(n13271), .A(n12768), .ZN(n12770) );
  NAND2_X1 U15876 ( .A1(n12771), .A2(n12770), .ZN(n13516) );
  NAND2_X1 U15877 ( .A1(n12772), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12773) );
  INV_X1 U15878 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20016) );
  XNOR2_X1 U15879 ( .A(n12777), .B(n20016), .ZN(n13632) );
  NAND2_X1 U15880 ( .A1(n12775), .A2(n12774), .ZN(n12791) );
  XNOR2_X1 U15881 ( .A(n12791), .B(n12789), .ZN(n12776) );
  OAI22_X1 U15882 ( .A1(n20060), .A2(n12779), .B1(n20789), .B2(n12776), .ZN(
        n13631) );
  NAND2_X1 U15883 ( .A1(n13632), .A2(n13631), .ZN(n13634) );
  NAND2_X1 U15884 ( .A1(n12777), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12778) );
  NAND2_X1 U15885 ( .A1(n12780), .A2(n9895), .ZN(n12784) );
  NAND2_X1 U15886 ( .A1(n12791), .A2(n12789), .ZN(n12781) );
  XNOR2_X1 U15887 ( .A(n12781), .B(n12788), .ZN(n12782) );
  NAND2_X1 U15888 ( .A1(n12782), .A2(n13271), .ZN(n12783) );
  NAND2_X1 U15889 ( .A1(n12784), .A2(n12783), .ZN(n12785) );
  INV_X1 U15890 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20009) );
  NAND2_X1 U15891 ( .A1(n12785), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12786) );
  NAND2_X1 U15892 ( .A1(n12787), .A2(n9895), .ZN(n12794) );
  AND2_X1 U15893 ( .A1(n12789), .A2(n12788), .ZN(n12790) );
  NAND2_X1 U15894 ( .A1(n12791), .A2(n12790), .ZN(n12799) );
  XNOR2_X1 U15895 ( .A(n12799), .B(n12800), .ZN(n12792) );
  NAND2_X1 U15896 ( .A1(n12792), .A2(n13271), .ZN(n12793) );
  NAND2_X1 U15897 ( .A1(n12794), .A2(n12793), .ZN(n12795) );
  INV_X1 U15898 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15759) );
  XNOR2_X1 U15899 ( .A(n12795), .B(n15759), .ZN(n15672) );
  NAND2_X1 U15900 ( .A1(n12795), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12796) );
  NAND3_X1 U15901 ( .A1(n12798), .A2(n12797), .A3(n9895), .ZN(n12804) );
  INV_X1 U15902 ( .A(n12799), .ZN(n12801) );
  NAND2_X1 U15903 ( .A1(n12801), .A2(n12800), .ZN(n12808) );
  XNOR2_X1 U15904 ( .A(n12808), .B(n12809), .ZN(n12802) );
  NAND2_X1 U15905 ( .A1(n12802), .A2(n13271), .ZN(n12803) );
  INV_X1 U15906 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15666) );
  NAND2_X1 U15907 ( .A1(n15667), .A2(n15666), .ZN(n12805) );
  INV_X1 U15908 ( .A(n15667), .ZN(n12806) );
  NAND2_X1 U15909 ( .A1(n12806), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12807) );
  INV_X1 U15910 ( .A(n12808), .ZN(n12810) );
  NAND2_X1 U15911 ( .A1(n12810), .A2(n12809), .ZN(n12818) );
  XNOR2_X1 U15912 ( .A(n12818), .B(n12811), .ZN(n12812) );
  AND2_X1 U15913 ( .A1(n12812), .A2(n13271), .ZN(n12813) );
  AOI21_X1 U15914 ( .B1(n12814), .B2(n9895), .A(n12813), .ZN(n12815) );
  INV_X1 U15915 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15776) );
  NAND2_X1 U15916 ( .A1(n12815), .A2(n15776), .ZN(n15662) );
  INV_X1 U15917 ( .A(n12815), .ZN(n12816) );
  NAND2_X1 U15918 ( .A1(n12816), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15661) );
  OR3_X1 U15919 ( .A1(n12818), .A2(n12817), .A3(n20789), .ZN(n12819) );
  NAND2_X1 U15920 ( .A1(n13911), .A2(n15771), .ZN(n12820) );
  NAND2_X1 U15921 ( .A1(n13910), .A2(n12820), .ZN(n12823) );
  INV_X1 U15922 ( .A(n13911), .ZN(n12821) );
  NAND2_X1 U15923 ( .A1(n12821), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12822) );
  INV_X1 U15924 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12824) );
  NOR2_X1 U15925 ( .A1(n15651), .A2(n12824), .ZN(n13990) );
  OR2_X2 U15926 ( .A1(n13989), .A2(n13990), .ZN(n14589) );
  NAND2_X1 U15927 ( .A1(n15651), .A2(n12824), .ZN(n13988) );
  AND2_X1 U15928 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13014) );
  NAND2_X1 U15929 ( .A1(n15631), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14042) );
  INV_X1 U15930 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12825) );
  NAND2_X1 U15931 ( .A1(n15651), .A2(n12825), .ZN(n12826) );
  INV_X1 U15932 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12941) );
  NAND2_X1 U15933 ( .A1(n15651), .A2(n12941), .ZN(n14680) );
  NAND2_X1 U15934 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12827) );
  NAND2_X1 U15935 ( .A1(n15651), .A2(n12827), .ZN(n14579) );
  INV_X1 U15936 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15718) );
  NAND2_X1 U15937 ( .A1(n15651), .A2(n15718), .ZN(n12828) );
  NAND2_X1 U15938 ( .A1(n14044), .A2(n12828), .ZN(n14567) );
  NAND2_X1 U15939 ( .A1(n15631), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12829) );
  AND2_X1 U15940 ( .A1(n14042), .A2(n12829), .ZN(n14568) );
  NAND2_X1 U15941 ( .A1(n15631), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12830) );
  INV_X1 U15942 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15716) );
  XNOR2_X1 U15943 ( .A(n15651), .B(n15716), .ZN(n15635) );
  AOI21_X1 U15944 ( .B1(n14567), .B2(n12831), .A(n15635), .ZN(n14553) );
  NAND2_X1 U15945 ( .A1(n15631), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14580) );
  INV_X1 U15946 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15752) );
  INV_X1 U15947 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15741) );
  NAND2_X1 U15948 ( .A1(n15752), .A2(n15741), .ZN(n12832) );
  NAND2_X1 U15949 ( .A1(n15631), .A2(n12832), .ZN(n14577) );
  OAI21_X1 U15950 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n15631), .ZN(n12833) );
  NAND2_X1 U15951 ( .A1(n14566), .A2(n12833), .ZN(n12834) );
  INV_X1 U15952 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12837) );
  INV_X1 U15953 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12836) );
  NAND3_X1 U15954 ( .A1(n9612), .A2(n12837), .A3(n12836), .ZN(n12838) );
  XNOR2_X1 U15955 ( .A(n15651), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14548) );
  NAND2_X1 U15956 ( .A1(n14546), .A2(n14548), .ZN(n14524) );
  NAND2_X1 U15957 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n13026) );
  INV_X1 U15958 ( .A(n13026), .ZN(n12839) );
  OAI21_X2 U15959 ( .B1(n14524), .B2(n12840), .A(n15651), .ZN(n15625) );
  INV_X1 U15960 ( .A(n12842), .ZN(n12845) );
  INV_X1 U15961 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14643) );
  INV_X1 U15962 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12843) );
  NAND2_X1 U15963 ( .A1(n14643), .A2(n12843), .ZN(n12865) );
  NOR4_X1 U15964 ( .A1(n12865), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12844) );
  NAND2_X1 U15965 ( .A1(n12842), .A2(n12844), .ZN(n12847) );
  NAND3_X1 U15966 ( .A1(n12845), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12846) );
  INV_X1 U15967 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12848) );
  NAND2_X1 U15968 ( .A1(n13000), .A2(n13295), .ZN(n12850) );
  NOR2_X1 U15969 ( .A1(n12851), .A2(n12850), .ZN(n12852) );
  INV_X1 U15970 ( .A(n12853), .ZN(n14283) );
  AOI21_X1 U15971 ( .B1(n12854), .B2(n14283), .A(n14213), .ZN(n14365) );
  NAND3_X1 U15972 ( .A1(n20071), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15801) );
  INV_X1 U15973 ( .A(n15801), .ZN(n12855) );
  NOR2_X1 U15974 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20632) );
  AND2_X1 U15975 ( .A1(n12855), .A2(n20618), .ZN(n13319) );
  INV_X1 U15976 ( .A(n20632), .ZN(n20769) );
  NAND2_X1 U15977 ( .A1(n20769), .A2(n12860), .ZN(n20785) );
  AND2_X1 U15978 ( .A1(n20785), .A2(n20071), .ZN(n12856) );
  NAND2_X1 U15979 ( .A1(n20071), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12858) );
  INV_X1 U15980 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20578) );
  NAND2_X1 U15981 ( .A1(n20578), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12857) );
  AND2_X1 U15982 ( .A1(n12858), .A2(n12857), .ZN(n13288) );
  INV_X1 U15983 ( .A(n13288), .ZN(n12859) );
  OR2_X1 U15984 ( .A1(n12860), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20035) );
  NAND2_X1 U15985 ( .A1(n20053), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14071) );
  NAND2_X1 U15986 ( .A1(n19984), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12861) );
  OAI211_X1 U15987 ( .C1(n19995), .C2(n14270), .A(n14071), .B(n12861), .ZN(
        n12862) );
  AOI21_X1 U15988 ( .B1(n14365), .B2(n13319), .A(n12862), .ZN(n12863) );
  INV_X1 U15989 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12866) );
  NAND2_X1 U15990 ( .A1(n12868), .A2(n15651), .ZN(n14500) );
  NAND2_X1 U15991 ( .A1(n14482), .A2(n14500), .ZN(n12869) );
  NOR2_X1 U15992 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12870) );
  INV_X1 U15993 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14607) );
  NAND2_X1 U15994 ( .A1(n14205), .A2(n14607), .ZN(n14473) );
  AND2_X1 U15995 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13028) );
  NAND2_X1 U15996 ( .A1(n15651), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12872) );
  XNOR2_X1 U15997 ( .A(n12873), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14091) );
  INV_X1 U15998 ( .A(n12874), .ZN(n12875) );
  INV_X1 U15999 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n19812) );
  NAND2_X1 U16000 ( .A1(n12875), .A2(n19812), .ZN(n15505) );
  AND2_X1 U16001 ( .A1(n13325), .A2(n15505), .ZN(n12876) );
  OR2_X1 U16002 ( .A1(n12877), .A2(n12876), .ZN(n12881) );
  AOI22_X1 U16003 ( .A1(n12878), .A2(n12697), .B1(n13271), .B2(n15505), .ZN(
        n12879) );
  MUX2_X1 U16004 ( .A(n12881), .B(n12880), .S(n20085), .Z(n12890) );
  OR2_X1 U16005 ( .A1(n13142), .A2(n12892), .ZN(n12886) );
  NAND2_X1 U16006 ( .A1(n12883), .A2(n13325), .ZN(n12995) );
  NAND2_X1 U16007 ( .A1(n12995), .A2(n12697), .ZN(n12884) );
  OR2_X1 U16008 ( .A1(n12885), .A2(n12884), .ZN(n13008) );
  NAND2_X1 U16009 ( .A1(n12886), .A2(n13008), .ZN(n13440) );
  INV_X1 U16010 ( .A(n13440), .ZN(n12889) );
  INV_X1 U16011 ( .A(n12995), .ZN(n12887) );
  NAND2_X1 U16012 ( .A1(n15484), .A2(n12887), .ZN(n12888) );
  NAND3_X1 U16013 ( .A1(n12890), .A2(n12889), .A3(n12888), .ZN(n12891) );
  NAND2_X1 U16014 ( .A1(n12892), .A2(n13000), .ZN(n15475) );
  NAND2_X1 U16015 ( .A1(n13560), .A2(n15475), .ZN(n13143) );
  NOR2_X1 U16016 ( .A1(n12897), .A2(n20094), .ZN(n12893) );
  OR2_X1 U16017 ( .A1(n13143), .A2(n12893), .ZN(n12895) );
  NOR2_X1 U16018 ( .A1(n12895), .A2(n12894), .ZN(n12896) );
  NOR2_X1 U16019 ( .A1(n13138), .A2(n13325), .ZN(n15480) );
  NOR2_X1 U16020 ( .A1(n12897), .A2(n11972), .ZN(n12898) );
  NOR2_X1 U16021 ( .A1(n15480), .A2(n12898), .ZN(n12899) );
  AOI22_X1 U16022 ( .A1(n13315), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n13292), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12994) );
  AOI22_X1 U16023 ( .A1(n13315), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n13292), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14250) );
  AND2_X2 U16024 ( .A1(n14243), .A2(n13063), .ZN(n12973) );
  INV_X1 U16025 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13297) );
  NAND2_X1 U16026 ( .A1(n12973), .A2(n13297), .ZN(n12905) );
  INV_X1 U16027 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20044) );
  NAND2_X1 U16028 ( .A1(n12901), .A2(n20044), .ZN(n12903) );
  NAND2_X1 U16029 ( .A1(n13063), .A2(n13297), .ZN(n12902) );
  NAND3_X1 U16030 ( .A1(n12903), .A2(n12993), .A3(n12902), .ZN(n12904) );
  NAND2_X1 U16031 ( .A1(n12905), .A2(n12904), .ZN(n12908) );
  NAND2_X1 U16032 ( .A1(n12901), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12907) );
  INV_X1 U16033 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13318) );
  NAND2_X1 U16034 ( .A1(n12993), .A2(n13318), .ZN(n12906) );
  NAND2_X1 U16035 ( .A1(n12907), .A2(n12906), .ZN(n13316) );
  XNOR2_X1 U16036 ( .A(n12908), .B(n13316), .ZN(n13064) );
  NAND2_X1 U16037 ( .A1(n13064), .A2(n13063), .ZN(n13066) );
  NAND2_X1 U16038 ( .A1(n13066), .A2(n12908), .ZN(n13081) );
  INV_X1 U16039 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13510) );
  NAND2_X1 U16040 ( .A1(n12973), .A2(n13510), .ZN(n12912) );
  NAND2_X1 U16041 ( .A1(n12901), .A2(n20029), .ZN(n12910) );
  NAND2_X1 U16042 ( .A1(n13063), .A2(n13510), .ZN(n12909) );
  NAND3_X1 U16043 ( .A1(n12910), .A2(n12993), .A3(n12909), .ZN(n12911) );
  AND2_X1 U16044 ( .A1(n12912), .A2(n12911), .ZN(n13080) );
  MUX2_X1 U16045 ( .A(n12986), .B(n12993), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12915) );
  NAND2_X1 U16046 ( .A1(n9993), .A2(n12915), .ZN(n13538) );
  NAND2_X1 U16047 ( .A1(n12901), .A2(n20009), .ZN(n12917) );
  INV_X1 U16048 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13756) );
  NAND2_X1 U16049 ( .A1(n13063), .A2(n13756), .ZN(n12916) );
  NAND3_X1 U16050 ( .A1(n12917), .A2(n12993), .A3(n12916), .ZN(n12918) );
  OAI21_X1 U16051 ( .B1(n12992), .B2(P1_EBX_REG_4__SCAN_IN), .A(n12918), .ZN(
        n13615) );
  MUX2_X1 U16052 ( .A(n12986), .B(n12993), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n12919) );
  NAND2_X1 U16053 ( .A1(n9992), .A2(n12919), .ZN(n13610) );
  MUX2_X1 U16054 ( .A(n12986), .B(n12993), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n12920) );
  INV_X1 U16055 ( .A(n12920), .ZN(n12922) );
  NOR2_X1 U16056 ( .A1(n13315), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12921) );
  NOR2_X1 U16057 ( .A1(n12922), .A2(n12921), .ZN(n13678) );
  INV_X1 U16058 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n19917) );
  NAND2_X1 U16059 ( .A1(n12973), .A2(n19917), .ZN(n12926) );
  NAND2_X1 U16060 ( .A1(n12901), .A2(n15666), .ZN(n12924) );
  NAND2_X1 U16061 ( .A1(n13063), .A2(n19917), .ZN(n12923) );
  NAND3_X1 U16062 ( .A1(n12924), .A2(n12993), .A3(n12923), .ZN(n12925) );
  NAND2_X1 U16063 ( .A1(n12926), .A2(n12925), .ZN(n15778) );
  INV_X1 U16064 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13882) );
  NAND2_X1 U16065 ( .A1(n12973), .A2(n13882), .ZN(n12931) );
  NAND2_X1 U16066 ( .A1(n12901), .A2(n15771), .ZN(n12929) );
  NAND2_X1 U16067 ( .A1(n13063), .A2(n13882), .ZN(n12928) );
  NAND3_X1 U16068 ( .A1(n12929), .A2(n12993), .A3(n12928), .ZN(n12930) );
  AND2_X1 U16069 ( .A1(n12931), .A2(n12930), .ZN(n13877) );
  MUX2_X1 U16070 ( .A(n12986), .B(n12993), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n12932) );
  INV_X1 U16071 ( .A(n12932), .ZN(n12934) );
  NOR2_X1 U16072 ( .A1(n13315), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12933) );
  NOR2_X1 U16073 ( .A1(n12934), .A2(n12933), .ZN(n13919) );
  NAND2_X1 U16074 ( .A1(n13920), .A2(n13919), .ZN(n13918) );
  MUX2_X1 U16075 ( .A(n12992), .B(n12901), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n12937) );
  INV_X1 U16076 ( .A(n12901), .ZN(n12935) );
  NAND2_X1 U16077 ( .A1(n12935), .A2(n13292), .ZN(n12962) );
  NAND2_X1 U16078 ( .A1(n13292), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12936) );
  INV_X1 U16079 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15623) );
  NAND2_X1 U16080 ( .A1(n13063), .A2(n15623), .ZN(n12939) );
  NAND2_X1 U16081 ( .A1(n12993), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12938) );
  NAND3_X1 U16082 ( .A1(n12939), .A2(n12901), .A3(n12938), .ZN(n12940) );
  OAI21_X1 U16083 ( .B1(n12986), .B2(P1_EBX_REG_11__SCAN_IN), .A(n12940), .ZN(
        n15595) );
  NAND2_X1 U16084 ( .A1(n12901), .A2(n12941), .ZN(n12943) );
  INV_X1 U16085 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15585) );
  NAND2_X1 U16086 ( .A1(n13063), .A2(n15585), .ZN(n12942) );
  NAND3_X1 U16087 ( .A1(n12943), .A2(n12993), .A3(n12942), .ZN(n12944) );
  OAI21_X1 U16088 ( .B1(n12992), .B2(P1_EBX_REG_12__SCAN_IN), .A(n12944), .ZN(
        n14013) );
  INV_X1 U16089 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n12945) );
  NAND2_X1 U16090 ( .A1(n13063), .A2(n12945), .ZN(n12947) );
  NAND2_X1 U16091 ( .A1(n12993), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12946) );
  NAND3_X1 U16092 ( .A1(n12947), .A2(n12901), .A3(n12946), .ZN(n12948) );
  OAI21_X1 U16093 ( .B1(n12986), .B2(P1_EBX_REG_13__SCAN_IN), .A(n12948), .ZN(
        n13973) );
  MUX2_X1 U16094 ( .A(n12992), .B(n12901), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n12950) );
  NAND2_X1 U16095 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n13292), .ZN(
        n12949) );
  AND3_X1 U16096 ( .A1(n12950), .A2(n12962), .A3(n12949), .ZN(n14018) );
  MUX2_X1 U16097 ( .A(n12986), .B(n12993), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12951) );
  NAND2_X1 U16098 ( .A1(n9999), .A2(n12951), .ZN(n14026) );
  MUX2_X1 U16099 ( .A(n12992), .B(n12901), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n12953) );
  NAND2_X1 U16100 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n13292), .ZN(
        n12952) );
  AND3_X1 U16101 ( .A1(n12953), .A2(n12962), .A3(n12952), .ZN(n14350) );
  MUX2_X1 U16102 ( .A(n12986), .B(n12993), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n12954) );
  OAI21_X1 U16103 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n13315), .A(
        n12954), .ZN(n14353) );
  NOR2_X1 U16104 ( .A1(n14350), .A2(n14353), .ZN(n12955) );
  INV_X1 U16105 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14400) );
  NAND2_X1 U16106 ( .A1(n12973), .A2(n14400), .ZN(n12959) );
  INV_X1 U16107 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15701) );
  NAND2_X1 U16108 ( .A1(n12901), .A2(n15701), .ZN(n12957) );
  NAND2_X1 U16109 ( .A1(n13063), .A2(n14400), .ZN(n12956) );
  NAND3_X1 U16110 ( .A1(n12957), .A2(n12993), .A3(n12956), .ZN(n12958) );
  AND2_X1 U16111 ( .A1(n12959), .A2(n12958), .ZN(n14396) );
  OR2_X2 U16112 ( .A1(n14397), .A2(n14396), .ZN(n14399) );
  MUX2_X1 U16113 ( .A(n12986), .B(n12993), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12960) );
  OAI21_X1 U16114 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n13315), .A(
        n12960), .ZN(n14335) );
  MUX2_X1 U16115 ( .A(n12992), .B(n12901), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n12964) );
  NAND2_X1 U16116 ( .A1(n13292), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12961) );
  AND2_X1 U16117 ( .A1(n12962), .A2(n12961), .ZN(n12963) );
  NAND2_X1 U16118 ( .A1(n12964), .A2(n12963), .ZN(n14389) );
  INV_X1 U16119 ( .A(n12986), .ZN(n12965) );
  INV_X1 U16120 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15621) );
  NAND2_X1 U16121 ( .A1(n12965), .A2(n15621), .ZN(n12969) );
  NAND2_X1 U16122 ( .A1(n13063), .A2(n15621), .ZN(n12967) );
  NAND2_X1 U16123 ( .A1(n12993), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12966) );
  NAND3_X1 U16124 ( .A1(n12967), .A2(n12901), .A3(n12966), .ZN(n12968) );
  AND2_X1 U16125 ( .A1(n12969), .A2(n12968), .ZN(n14654) );
  MUX2_X1 U16126 ( .A(n12986), .B(n12993), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n12970) );
  INV_X1 U16127 ( .A(n12970), .ZN(n12972) );
  NOR2_X1 U16128 ( .A1(n13315), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12971) );
  NOR2_X1 U16129 ( .A1(n12972), .A2(n12971), .ZN(n14377) );
  INV_X1 U16130 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15617) );
  NAND2_X1 U16131 ( .A1(n12973), .A2(n15617), .ZN(n12978) );
  INV_X1 U16132 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12974) );
  NAND2_X1 U16133 ( .A1(n12901), .A2(n12974), .ZN(n12976) );
  NAND2_X1 U16134 ( .A1(n13063), .A2(n15617), .ZN(n12975) );
  NAND3_X1 U16135 ( .A1(n12976), .A2(n12993), .A3(n12975), .ZN(n12977) );
  NAND2_X1 U16136 ( .A1(n12978), .A2(n12977), .ZN(n15529) );
  NAND2_X1 U16137 ( .A1(n14377), .A2(n15529), .ZN(n12979) );
  MUX2_X1 U16138 ( .A(n12992), .B(n12901), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n12981) );
  NAND2_X1 U16139 ( .A1(n13292), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12980) );
  AND2_X1 U16140 ( .A1(n12981), .A2(n12980), .ZN(n14322) );
  MUX2_X1 U16141 ( .A(n12986), .B(n12993), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n12982) );
  OAI21_X1 U16142 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n13315), .A(
        n12982), .ZN(n12983) );
  INV_X1 U16143 ( .A(n12983), .ZN(n14305) );
  MUX2_X1 U16144 ( .A(n12992), .B(n12901), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n12985) );
  NAND2_X1 U16145 ( .A1(n13292), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12984) );
  NAND2_X1 U16146 ( .A1(n12985), .A2(n12984), .ZN(n14298) );
  MUX2_X1 U16147 ( .A(n12986), .B(n12993), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12987) );
  OAI21_X1 U16148 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n13315), .A(
        n12987), .ZN(n14280) );
  MUX2_X1 U16149 ( .A(n12992), .B(n12901), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n12989) );
  NAND2_X1 U16150 ( .A1(n13292), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12988) );
  AND2_X1 U16151 ( .A1(n12989), .A2(n12988), .ZN(n14069) );
  OR2_X1 U16152 ( .A1(n13315), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12991) );
  INV_X1 U16153 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14229) );
  NAND2_X1 U16154 ( .A1(n13063), .A2(n14229), .ZN(n12990) );
  NAND2_X1 U16155 ( .A1(n12991), .A2(n12990), .ZN(n14245) );
  OAI22_X1 U16156 ( .A1(n14245), .A2(n14243), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n12992), .ZN(n14225) );
  INV_X1 U16157 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20747) );
  NOR2_X1 U16158 ( .A1(n20035), .A2(n20747), .ZN(n14086) );
  INV_X1 U16159 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20034) );
  OAI21_X1 U16160 ( .B1(n20034), .B2(n20044), .A(n20029), .ZN(n20020) );
  NOR2_X1 U16161 ( .A1(n20009), .A2(n20016), .ZN(n19998) );
  NAND3_X1 U16162 ( .A1(n20020), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n19998), .ZN(n14665) );
  INV_X1 U16163 ( .A(n14665), .ZN(n15744) );
  NOR2_X1 U16164 ( .A1(n12996), .A2(n12995), .ZN(n13562) );
  INV_X1 U16165 ( .A(n13562), .ZN(n13145) );
  NOR2_X1 U16166 ( .A1(n15744), .A2(n13023), .ZN(n15763) );
  INV_X1 U16167 ( .A(n12997), .ZN(n13003) );
  NAND2_X1 U16168 ( .A1(n11976), .A2(n13437), .ZN(n12998) );
  OAI211_X1 U16169 ( .C1(n13000), .C2(n12697), .A(n12999), .B(n12998), .ZN(
        n13001) );
  NAND2_X1 U16170 ( .A1(n13001), .A2(n13325), .ZN(n13002) );
  OAI211_X1 U16171 ( .C1(n13004), .C2(n12993), .A(n13003), .B(n13002), .ZN(
        n13005) );
  INV_X1 U16172 ( .A(n13005), .ZN(n13007) );
  NAND2_X1 U16173 ( .A1(n11970), .A2(n13126), .ZN(n13006) );
  NAND3_X1 U16174 ( .A1(n13008), .A2(n13007), .A3(n13006), .ZN(n13422) );
  OAI21_X1 U16175 ( .B1(n13419), .B2(n12697), .A(n13009), .ZN(n13010) );
  NOR2_X1 U16176 ( .A1(n13422), .A2(n13010), .ZN(n13011) );
  AOI22_X1 U16177 ( .A1(n20035), .A2(n13012), .B1(n20034), .B2(n20046), .ZN(
        n15760) );
  INV_X1 U16178 ( .A(n15760), .ZN(n20033) );
  NOR2_X1 U16179 ( .A1(n15763), .A2(n20033), .ZN(n14685) );
  NAND3_X1 U16180 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15748) );
  NAND2_X1 U16181 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15749) );
  NOR2_X1 U16182 ( .A1(n15748), .A2(n15749), .ZN(n14686) );
  NAND2_X1 U16183 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14686), .ZN(
        n14688) );
  NOR2_X1 U16184 ( .A1(n12941), .A2(n14688), .ZN(n14661) );
  NAND2_X1 U16185 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14661), .ZN(
        n13024) );
  NAND2_X1 U16186 ( .A1(n13142), .A2(n13325), .ZN(n15462) );
  INV_X1 U16187 ( .A(n19998), .ZN(n15764) );
  NOR4_X1 U16188 ( .A1(n15759), .A2(n20029), .A3(n20044), .A4(n15764), .ZN(
        n15743) );
  INV_X1 U16189 ( .A(n15743), .ZN(n14662) );
  AOI222_X1 U16190 ( .A1(n13024), .A2(n20018), .B1(n13024), .B2(n20047), .C1(
        n20018), .C2(n14662), .ZN(n13013) );
  NAND3_X1 U16191 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n13014), .ZN(n15694) );
  NOR2_X1 U16192 ( .A1(n15701), .A2(n15694), .ZN(n13025) );
  INV_X1 U16193 ( .A(n13025), .ZN(n13015) );
  NAND2_X1 U16194 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15682) );
  AND2_X1 U16195 ( .A1(n20031), .A2(n15682), .ZN(n13016) );
  NOR2_X1 U16196 ( .A1(n15679), .A2(n13016), .ZN(n14649) );
  NAND2_X1 U16197 ( .A1(n20047), .A2(n12864), .ZN(n13017) );
  NAND2_X1 U16198 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14625) );
  AND2_X1 U16199 ( .A1(n20046), .A2(n14625), .ZN(n13018) );
  INV_X1 U16200 ( .A(n20031), .ZN(n13022) );
  INV_X1 U16201 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n20891) );
  INV_X1 U16202 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13021) );
  OAI22_X1 U16203 ( .A1(n12841), .A2(n20055), .B1(n13023), .B2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n13019) );
  NAND2_X1 U16204 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13020) );
  NAND2_X1 U16205 ( .A1(n20034), .A2(n20055), .ZN(n20032) );
  NAND2_X1 U16206 ( .A1(n20018), .A2(n20032), .ZN(n14689) );
  NAND2_X1 U16207 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14638), .ZN(
        n20030) );
  NAND2_X1 U16208 ( .A1(n15702), .A2(n13025), .ZN(n15693) );
  AND2_X1 U16209 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13027) );
  NAND3_X1 U16210 ( .A1(n14651), .A2(n12841), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14613) );
  NOR2_X1 U16211 ( .A1(n14613), .A2(n9855), .ZN(n14608) );
  NAND4_X1 U16212 ( .A1(n14608), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n20891), .ZN(n13029) );
  AND2_X1 U16213 ( .A1(n13030), .A2(n13029), .ZN(n13031) );
  OAI21_X1 U16214 ( .B1(n14091), .B2(n20050), .A(n13031), .ZN(P1_U3000) );
  INV_X1 U16215 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20783) );
  NOR3_X1 U16216 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n20783), .ZN(n13033) );
  NOR4_X1 U16217 ( .A1(P1_BE_N_REG_1__SCAN_IN), .A2(P1_BE_N_REG_2__SCAN_IN), 
        .A3(P1_BE_N_REG_3__SCAN_IN), .A4(P1_D_C_N_REG_SCAN_IN), .ZN(n13032) );
  NAND4_X1 U16218 ( .A1(n20068), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13033), .A4(
        n13032), .ZN(U214) );
  INV_X1 U16219 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19798) );
  NOR2_X1 U16220 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(n19798), .ZN(n13035) );
  NOR4_X1 U16221 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13034) );
  INV_X1 U16222 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n20925) );
  NAND4_X1 U16223 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(n13035), .A3(n13034), .A4(
        n20925), .ZN(n13036) );
  NOR2_X1 U16224 ( .A1(n15407), .A2(n13036), .ZN(n16150) );
  NAND2_X1 U16225 ( .A1(n16150), .A2(U214), .ZN(U212) );
  NOR2_X1 U16226 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13036), .ZN(n16226)
         );
  OAI21_X1 U16227 ( .B1(n13038), .B2(n13037), .A(n13075), .ZN(n13534) );
  NAND2_X1 U16228 ( .A1(n13142), .A2(n13149), .ZN(n13139) );
  NOR2_X1 U16229 ( .A1(n13138), .A2(n19815), .ZN(n13039) );
  AND2_X1 U16230 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20071), .ZN(n13040) );
  NOR2_X1 U16231 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20790) );
  NAND2_X1 U16232 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20790), .ZN(n15805) );
  INV_X1 U16233 ( .A(n15805), .ZN(n15488) );
  AOI22_X1 U16234 ( .A1(n13041), .A2(n13040), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n15488), .ZN(n13042) );
  AND2_X1 U16235 ( .A1(n20035), .A2(n13042), .ZN(n13043) );
  NOR2_X1 U16236 ( .A1(n13053), .A2(n13140), .ZN(n13050) );
  INV_X1 U16237 ( .A(n13045), .ZN(n13046) );
  NAND2_X1 U16238 ( .A1(n13046), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13048) );
  INV_X1 U16239 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13047) );
  XNOR2_X1 U16240 ( .A(n13048), .B(n13047), .ZN(n14088) );
  NOR2_X1 U16241 ( .A1(n14088), .A2(n13584), .ZN(n13049) );
  OR2_X1 U16242 ( .A1(n13050), .A2(n19870), .ZN(n19886) );
  INV_X1 U16243 ( .A(n19886), .ZN(n19904) );
  NOR2_X1 U16244 ( .A1(n13534), .A2(n19904), .ZN(n13071) );
  OR2_X1 U16245 ( .A1(n13053), .A2(n13438), .ZN(n19898) );
  NOR2_X1 U16246 ( .A1(n20571), .A2(n19898), .ZN(n13070) );
  AND2_X1 U16247 ( .A1(n14088), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13052) );
  OR2_X1 U16248 ( .A1(n13053), .A2(n20072), .ZN(n13062) );
  AND2_X1 U16249 ( .A1(n13325), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13060) );
  AND2_X1 U16250 ( .A1(n20786), .A2(n20578), .ZN(n15482) );
  INV_X1 U16251 ( .A(n15482), .ZN(n13059) );
  AOI21_X1 U16252 ( .B1(n11957), .B2(n15505), .A(n13059), .ZN(n13057) );
  OR2_X1 U16253 ( .A1(n13060), .A2(n13057), .ZN(n13054) );
  NAND2_X1 U16254 ( .A1(n19876), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n13056) );
  INV_X1 U16255 ( .A(n15531), .ZN(n19850) );
  AOI22_X1 U16256 ( .A1(n19866), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19850), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n13055) );
  OAI211_X1 U16257 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n19890), .A(
        n13056), .B(n13055), .ZN(n13069) );
  INV_X1 U16258 ( .A(n13062), .ZN(n13058) );
  OR2_X1 U16259 ( .A1(n19852), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n13078) );
  NAND2_X1 U16260 ( .A1(n13060), .A2(n13059), .ZN(n13061) );
  OR2_X1 U16261 ( .A1(n13064), .A2(n13063), .ZN(n13065) );
  AND2_X1 U16262 ( .A1(n13066), .A2(n13065), .ZN(n13298) );
  INV_X1 U16263 ( .A(n13298), .ZN(n20041) );
  NAND2_X1 U16264 ( .A1(n9561), .A2(n20041), .ZN(n13067) );
  NAND2_X1 U16265 ( .A1(n13078), .A2(n13067), .ZN(n13068) );
  OR4_X1 U16266 ( .A1(n13071), .A2(n13070), .A3(n13069), .A4(n13068), .ZN(
        P1_U2839) );
  INV_X1 U16267 ( .A(n13073), .ZN(n13074) );
  AOI21_X1 U16268 ( .B1(n13072), .B2(n13075), .A(n13074), .ZN(n13521) );
  INV_X1 U16269 ( .A(n13521), .ZN(n13532) );
  NOR2_X1 U16270 ( .A1(n13532), .A2(n19904), .ZN(n13091) );
  NOR2_X1 U16271 ( .A1(n20512), .A2(n19898), .ZN(n13090) );
  INV_X1 U16272 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n13077) );
  AOI21_X1 U16273 ( .B1(n13078), .B2(n15531), .A(n13077), .ZN(n13089) );
  INV_X1 U16274 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20775) );
  NOR2_X1 U16275 ( .A1(n19852), .A2(n20775), .ZN(n19893) );
  NAND2_X1 U16276 ( .A1(n19893), .A2(n13077), .ZN(n13087) );
  INV_X1 U16277 ( .A(n13514), .ZN(n13079) );
  AOI22_X1 U16278 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19866), .B1(
        n19907), .B2(n13079), .ZN(n13086) );
  NAND2_X1 U16279 ( .A1(n13081), .A2(n13080), .ZN(n13082) );
  NAND2_X1 U16280 ( .A1(n13539), .A2(n13082), .ZN(n20024) );
  INV_X1 U16281 ( .A(n20024), .ZN(n13083) );
  NAND2_X1 U16282 ( .A1(n9561), .A2(n13083), .ZN(n13085) );
  NAND2_X1 U16283 ( .A1(n19876), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n13084) );
  NAND4_X1 U16284 ( .A1(n13087), .A2(n13086), .A3(n13085), .A4(n13084), .ZN(
        n13088) );
  OR4_X1 U16285 ( .A1(n13091), .A2(n13090), .A3(n13089), .A4(n13088), .ZN(
        P1_U2838) );
  NAND2_X1 U16286 ( .A1(n18705), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18564) );
  INV_X1 U16287 ( .A(n18564), .ZN(n17369) );
  NAND2_X1 U16288 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17369), .ZN(n17233) );
  NAND2_X1 U16289 ( .A1(n18700), .A2(n18488), .ZN(n17270) );
  INV_X1 U16290 ( .A(n17270), .ZN(n17268) );
  INV_X1 U16291 ( .A(n17271), .ZN(n17269) );
  NAND2_X1 U16292 ( .A1(n18046), .A2(n17269), .ZN(n18548) );
  INV_X1 U16293 ( .A(n18701), .ZN(n18571) );
  AOI21_X1 U16294 ( .B1(n13092), .B2(n18548), .A(n18571), .ZN(n14062) );
  AND2_X1 U16295 ( .A1(n17263), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  OR3_X1 U16296 ( .A1(n16047), .A2(n16076), .A3(n16035), .ZN(n14199) );
  INV_X1 U16297 ( .A(n14199), .ZN(n18876) );
  INV_X1 U16298 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13095) );
  INV_X1 U16299 ( .A(n14200), .ZN(n13093) );
  OAI211_X1 U16300 ( .C1(n18876), .C2(n13095), .A(n13094), .B(n13093), .ZN(
        P2_U2814) );
  INV_X1 U16301 ( .A(n19682), .ZN(n14706) );
  NAND2_X1 U16302 ( .A1(n11404), .A2(n14706), .ZN(n14710) );
  AND2_X1 U16303 ( .A1(n14710), .A2(n19669), .ZN(n13096) );
  OR2_X1 U16304 ( .A1(n13097), .A2(n13096), .ZN(n16051) );
  AND2_X1 U16305 ( .A1(n16051), .A2(n13133), .ZN(n19807) );
  NAND2_X1 U16306 ( .A1(n19048), .A2(n13133), .ZN(n13098) );
  OR2_X1 U16307 ( .A1(n13099), .A2(n13098), .ZN(n13174) );
  OAI21_X1 U16308 ( .B1(n11350), .B2(n19807), .A(n13174), .ZN(P2_U2819) );
  INV_X1 U16309 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14874) );
  OR2_X1 U16310 ( .A1(n16047), .A2(n16076), .ZN(n13102) );
  OR2_X1 U16311 ( .A1(n13101), .A2(n13100), .ZN(n13269) );
  OAI21_X1 U16312 ( .B1(n13372), .B2(n13102), .A(n13269), .ZN(n13103) );
  OR2_X1 U16313 ( .A1(n19028), .A2(n13104), .ZN(n18992) );
  NOR2_X1 U16314 ( .A1(n19668), .A2(n19665), .ZN(n13365) );
  NAND2_X1 U16315 ( .A1(n13365), .A2(n16078), .ZN(n14713) );
  NAND2_X1 U16316 ( .A1(n19028), .A2(n14713), .ZN(n18995) );
  INV_X2 U16317 ( .A(n18995), .ZN(n19025) );
  AOI22_X1 U16318 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n19025), .B1(n19026), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13105) );
  OAI21_X1 U16319 ( .B1(n14874), .B2(n18992), .A(n13105), .ZN(P2_U2926) );
  INV_X1 U16320 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13107) );
  AOI22_X1 U16321 ( .A1(n19026), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13106) );
  OAI21_X1 U16322 ( .B1(n13107), .B2(n18992), .A(n13106), .ZN(P2_U2931) );
  INV_X1 U16323 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13109) );
  AOI22_X1 U16324 ( .A1(n19026), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13108) );
  OAI21_X1 U16325 ( .B1(n13109), .B2(n18992), .A(n13108), .ZN(P2_U2933) );
  INV_X1 U16326 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n14171) );
  AOI22_X1 U16327 ( .A1(n19026), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13110) );
  OAI21_X1 U16328 ( .B1(n14171), .B2(n18992), .A(n13110), .ZN(P2_U2928) );
  AOI22_X1 U16329 ( .A1(n19026), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13111) );
  OAI21_X1 U16330 ( .B1(n14899), .B2(n18992), .A(n13111), .ZN(P2_U2930) );
  INV_X1 U16331 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n14907) );
  AOI22_X1 U16332 ( .A1(n19026), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13112) );
  OAI21_X1 U16333 ( .B1(n14907), .B2(n18992), .A(n13112), .ZN(P2_U2932) );
  INV_X1 U16334 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14859) );
  AOI22_X1 U16335 ( .A1(n19026), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13113) );
  OAI21_X1 U16336 ( .B1(n14859), .B2(n18992), .A(n13113), .ZN(P2_U2924) );
  INV_X1 U16337 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n14850) );
  AOI22_X1 U16338 ( .A1(n19026), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13114) );
  OAI21_X1 U16339 ( .B1(n14850), .B2(n18992), .A(n13114), .ZN(P2_U2923) );
  INV_X1 U16340 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n14883) );
  AOI22_X1 U16341 ( .A1(n19026), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13115) );
  OAI21_X1 U16342 ( .B1(n14883), .B2(n18992), .A(n13115), .ZN(P2_U2927) );
  INV_X1 U16343 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13961) );
  AOI22_X1 U16344 ( .A1(n19026), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13116) );
  OAI21_X1 U16345 ( .B1(n13961), .B2(n18992), .A(n13116), .ZN(P2_U2934) );
  INV_X1 U16346 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14893) );
  AOI22_X1 U16347 ( .A1(n19026), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13117) );
  OAI21_X1 U16348 ( .B1(n14893), .B2(n18992), .A(n13117), .ZN(P2_U2929) );
  INV_X1 U16349 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13270) );
  AOI22_X1 U16350 ( .A1(n19026), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13118) );
  OAI21_X1 U16351 ( .B1(n13270), .B2(n18992), .A(n13118), .ZN(P2_U2925) );
  INV_X1 U16352 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n13120) );
  AOI22_X1 U16353 ( .A1(n19026), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13119) );
  OAI21_X1 U16354 ( .B1(n13120), .B2(n18992), .A(n13119), .ZN(P2_U2922) );
  INV_X1 U16355 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13122) );
  AOI22_X1 U16356 ( .A1(n19026), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13121) );
  OAI21_X1 U16357 ( .B1(n13122), .B2(n18992), .A(n13121), .ZN(P2_U2935) );
  NAND2_X1 U16358 ( .A1(n20618), .A2(n13584), .ZN(n19818) );
  NAND2_X1 U16359 ( .A1(n13326), .A2(n19818), .ZN(n13124) );
  AOI21_X1 U16360 ( .B1(n13125), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n13124), 
        .ZN(n13123) );
  INV_X1 U16361 ( .A(n13123), .ZN(P1_U2801) );
  OR2_X1 U16362 ( .A1(n13124), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n13127) );
  INV_X1 U16363 ( .A(n13127), .ZN(n13130) );
  INV_X1 U16364 ( .A(n13125), .ZN(n13128) );
  OAI22_X1 U16365 ( .A1(n13128), .A2(n13127), .B1(n13126), .B2(n14243), .ZN(
        n13129) );
  OAI21_X1 U16366 ( .B1(n13130), .B2(n20784), .A(n13129), .ZN(P1_U3487) );
  NAND2_X1 U16367 ( .A1(n15373), .A2(n10511), .ZN(n13353) );
  OR2_X1 U16368 ( .A1(n16037), .A2(n16041), .ZN(n13367) );
  NAND2_X1 U16369 ( .A1(n13353), .A2(n13367), .ZN(n13134) );
  AND2_X2 U16370 ( .A1(n13134), .A2(n13133), .ZN(n20956) );
  NAND2_X1 U16371 ( .A1(n20956), .A2(n9586), .ZN(n18919) );
  MUX2_X1 U16372 ( .A(n13135), .B(n11070), .S(n20956), .Z(n13136) );
  OAI21_X1 U16373 ( .B1(n15396), .B2(n18919), .A(n13136), .ZN(P2_U2886) );
  INV_X1 U16374 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13153) );
  AND2_X1 U16375 ( .A1(n15484), .A2(n13140), .ZN(n13137) );
  AOI21_X1 U16376 ( .B1(n13139), .B2(n13138), .A(n13137), .ZN(n19814) );
  NAND3_X1 U16377 ( .A1(n13140), .A2(n13292), .A3(n15505), .ZN(n13141) );
  NAND2_X1 U16378 ( .A1(n13141), .A2(n20786), .ZN(n20787) );
  AND2_X1 U16379 ( .A1(n19814), .A2(n20787), .ZN(n15472) );
  NOR2_X1 U16380 ( .A1(n15472), .A2(n19815), .ZN(n19824) );
  INV_X1 U16381 ( .A(n13142), .ZN(n13148) );
  AOI21_X1 U16382 ( .B1(n13144), .B2(n12697), .A(n13143), .ZN(n13146) );
  MUX2_X1 U16383 ( .A(n13146), .B(n13145), .S(n13434), .Z(n13147) );
  OAI21_X1 U16384 ( .B1(n13149), .B2(n13148), .A(n13147), .ZN(n13150) );
  NAND2_X1 U16385 ( .A1(n13150), .A2(n13381), .ZN(n15474) );
  INV_X1 U16386 ( .A(n15474), .ZN(n13151) );
  NAND2_X1 U16387 ( .A1(n13151), .A2(n19824), .ZN(n13152) );
  OAI21_X1 U16388 ( .B1(n13153), .B2(n19824), .A(n13152), .ZN(P1_U3484) );
  INV_X1 U16389 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13158) );
  NAND2_X1 U16390 ( .A1(n13154), .A2(n19669), .ZN(n13155) );
  NAND2_X1 U16391 ( .A1(n13155), .A2(n13269), .ZN(n13232) );
  NOR2_X2 U16392 ( .A1(n13155), .A2(n16044), .ZN(n19031) );
  INV_X1 U16393 ( .A(n19031), .ZN(n13157) );
  AOI22_X1 U16394 ( .A1(n15405), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n15407), .ZN(n18936) );
  INV_X1 U16395 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13156) );
  OAI222_X1 U16396 ( .A1(n13158), .A2(n13232), .B1(n13157), .B2(n18936), .C1(
        n13156), .C2(n13269), .ZN(P2_U2982) );
  NAND2_X1 U16397 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n16078), .ZN(n13377) );
  OR2_X1 U16398 ( .A1(n13159), .A2(n13377), .ZN(n13163) );
  OAI21_X1 U16399 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(
        P2_STATE2_REG_2__SCAN_IN), .A(n16078), .ZN(n16070) );
  INV_X1 U16400 ( .A(n16070), .ZN(n13161) );
  INV_X1 U16401 ( .A(n13365), .ZN(n13160) );
  NAND2_X1 U16402 ( .A1(n13161), .A2(n13160), .ZN(n13162) );
  NAND3_X1 U16403 ( .A1(n19759), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19609), 
        .ZN(n15406) );
  INV_X1 U16404 ( .A(n15406), .ZN(n19042) );
  AOI21_X1 U16405 ( .B1(n13167), .B2(n13166), .A(n13165), .ZN(n13403) );
  NOR2_X1 U16406 ( .A1(n19701), .A2(n18765), .ZN(n13402) );
  NAND2_X1 U16407 ( .A1(n13169), .A2(n13168), .ZN(n13170) );
  NAND2_X1 U16408 ( .A1(n13171), .A2(n13170), .ZN(n13406) );
  INV_X1 U16409 ( .A(n13174), .ZN(n13172) );
  NAND2_X1 U16410 ( .A1(n13172), .A2(n19054), .ZN(n15976) );
  NAND2_X1 U16411 ( .A1(n19668), .A2(n19611), .ZN(n19666) );
  INV_X1 U16412 ( .A(n19666), .ZN(n19758) );
  OR2_X1 U16413 ( .A1(n19759), .A2(n19758), .ZN(n19780) );
  NAND2_X1 U16414 ( .A1(n19780), .A2(n16078), .ZN(n13173) );
  NAND2_X1 U16415 ( .A1(n13174), .A2(n13173), .ZN(n19047) );
  OAI22_X1 U16416 ( .A1(n13406), .A2(n15976), .B1(n13734), .B2(n19047), .ZN(
        n13175) );
  AOI211_X1 U16417 ( .C1(n13164), .C2(n13403), .A(n13402), .B(n13175), .ZN(
        n13179) );
  NAND2_X1 U16418 ( .A1(n19544), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13176) );
  NAND2_X1 U16419 ( .A1(n13177), .A2(n13176), .ZN(n14133) );
  NAND2_X1 U16420 ( .A1(n19037), .A2(n13731), .ZN(n13178) );
  OAI211_X1 U16421 ( .C1(n15406), .C2(n11040), .A(n13179), .B(n13178), .ZN(
        P2_U3012) );
  INV_X1 U16422 ( .A(n13164), .ZN(n15977) );
  AOI21_X1 U16423 ( .B1(n15366), .B2(n13181), .A(n13180), .ZN(n13182) );
  INV_X1 U16424 ( .A(n13182), .ZN(n13305) );
  INV_X1 U16425 ( .A(n15976), .ZN(n19040) );
  OAI21_X1 U16426 ( .B1(n13843), .B2(n13345), .A(n13183), .ZN(n13184) );
  XOR2_X1 U16427 ( .A(n13184), .B(n15366), .Z(n13308) );
  INV_X1 U16428 ( .A(n19047), .ZN(n15984) );
  AOI22_X1 U16429 ( .A1(n19040), .A2(n13308), .B1(n15984), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13185) );
  NAND2_X1 U16430 ( .A1(n19038), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n13304) );
  OAI211_X1 U16431 ( .C1(n15977), .C2(n13305), .A(n13185), .B(n13304), .ZN(
        n13186) );
  AOI21_X1 U16432 ( .B1(n19037), .B2(n13187), .A(n13186), .ZN(n13188) );
  OAI21_X1 U16433 ( .B1(n11070), .B2(n15406), .A(n13188), .ZN(P2_U3013) );
  NAND2_X1 U16434 ( .A1(n13189), .A2(n9589), .ZN(n13190) );
  NAND2_X1 U16435 ( .A1(n14908), .A2(n13190), .ZN(n18958) );
  OAI22_X1 U16436 ( .A1(n13263), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n15405), .ZN(n19050) );
  INV_X1 U16437 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19053) );
  AND2_X1 U16438 ( .A1(n19611), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13191) );
  OAI211_X1 U16439 ( .C1(n16044), .C2(n19053), .A(n13192), .B(n13191), .ZN(
        n13193) );
  INV_X1 U16440 ( .A(n13193), .ZN(n13194) );
  INV_X1 U16441 ( .A(n13195), .ZN(n13201) );
  INV_X1 U16442 ( .A(n13196), .ZN(n13199) );
  INV_X1 U16443 ( .A(n13197), .ZN(n13198) );
  NAND2_X1 U16444 ( .A1(n13199), .A2(n13198), .ZN(n13200) );
  NAND2_X1 U16445 ( .A1(n13201), .A2(n13200), .ZN(n13202) );
  INV_X1 U16446 ( .A(n13202), .ZN(n18868) );
  NOR2_X1 U16447 ( .A1(n19792), .A2(n13202), .ZN(n18985) );
  INV_X1 U16448 ( .A(n18985), .ZN(n13203) );
  INV_X1 U16449 ( .A(n18986), .ZN(n18970) );
  OAI211_X1 U16450 ( .C1(n19334), .C2(n18868), .A(n13203), .B(n18970), .ZN(
        n13205) );
  INV_X1 U16451 ( .A(n18935), .ZN(n18982) );
  INV_X1 U16452 ( .A(n18956), .ZN(n18981) );
  AOI22_X1 U16453 ( .A1(n18982), .A2(n18868), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n18981), .ZN(n13204) );
  OAI211_X1 U16454 ( .C1(n18990), .C2(n19050), .A(n13205), .B(n13204), .ZN(
        P2_U2919) );
  INV_X2 U16455 ( .A(n13269), .ZN(n19033) );
  AOI22_X1 U16456 ( .A1(n9582), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_12__SCAN_IN), .B2(n19033), .ZN(n13209) );
  INV_X1 U16457 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n13332) );
  OR2_X1 U16458 ( .A1(n13263), .A2(n13332), .ZN(n13207) );
  NAND2_X1 U16459 ( .A1(n13263), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13206) );
  AND2_X1 U16460 ( .A1(n13207), .A2(n13206), .ZN(n18943) );
  INV_X1 U16461 ( .A(n18943), .ZN(n13208) );
  NAND2_X1 U16462 ( .A1(n19031), .A2(n13208), .ZN(n13239) );
  NAND2_X1 U16463 ( .A1(n13209), .A2(n13239), .ZN(P2_U2979) );
  AOI22_X1 U16464 ( .A1(n9582), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_8__SCAN_IN), .B2(n19033), .ZN(n13211) );
  AOI22_X1 U16465 ( .A1(n15405), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n13263), .ZN(n18953) );
  INV_X1 U16466 ( .A(n18953), .ZN(n13210) );
  NAND2_X1 U16467 ( .A1(n19031), .A2(n13210), .ZN(n13249) );
  NAND2_X1 U16468 ( .A1(n13211), .A2(n13249), .ZN(P2_U2975) );
  AOI22_X1 U16469 ( .A1(n9582), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19033), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13213) );
  AOI22_X1 U16470 ( .A1(n15405), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13263), .ZN(n19088) );
  INV_X1 U16471 ( .A(n19088), .ZN(n13212) );
  NAND2_X1 U16472 ( .A1(n19031), .A2(n13212), .ZN(n13251) );
  NAND2_X1 U16473 ( .A1(n13213), .A2(n13251), .ZN(P2_U2974) );
  AOI22_X1 U16474 ( .A1(n9582), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19033), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n13215) );
  AOI22_X1 U16475 ( .A1(n15405), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n15407), .ZN(n19077) );
  INV_X1 U16476 ( .A(n19077), .ZN(n13214) );
  NAND2_X1 U16477 ( .A1(n19031), .A2(n13214), .ZN(n13253) );
  NAND2_X1 U16478 ( .A1(n13215), .A2(n13253), .ZN(P2_U2973) );
  AOI22_X1 U16479 ( .A1(n9582), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19033), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n13216) );
  AOI22_X1 U16480 ( .A1(n15405), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n15407), .ZN(n19072) );
  INV_X1 U16481 ( .A(n19072), .ZN(n18959) );
  NAND2_X1 U16482 ( .A1(n19031), .A2(n18959), .ZN(n13243) );
  NAND2_X1 U16483 ( .A1(n13216), .A2(n13243), .ZN(P2_U2972) );
  AOI22_X1 U16484 ( .A1(n9582), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19033), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n13220) );
  INV_X1 U16485 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n14009) );
  OR2_X1 U16486 ( .A1(n13263), .A2(n14009), .ZN(n13218) );
  NAND2_X1 U16487 ( .A1(n13263), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13217) );
  AND2_X1 U16488 ( .A1(n13218), .A2(n13217), .ZN(n18945) );
  INV_X1 U16489 ( .A(n18945), .ZN(n13219) );
  NAND2_X1 U16490 ( .A1(n19031), .A2(n13219), .ZN(n13241) );
  NAND2_X1 U16491 ( .A1(n13220), .A2(n13241), .ZN(P2_U2978) );
  AOI22_X1 U16492 ( .A1(n9582), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_9__SCAN_IN), .B2(n19033), .ZN(n13225) );
  INV_X1 U16493 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n13221) );
  OR2_X1 U16494 ( .A1(n13263), .A2(n13221), .ZN(n13223) );
  NAND2_X1 U16495 ( .A1(n13263), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13222) );
  AND2_X1 U16496 ( .A1(n13223), .A2(n13222), .ZN(n18950) );
  INV_X1 U16497 ( .A(n18950), .ZN(n13224) );
  NAND2_X1 U16498 ( .A1(n19031), .A2(n13224), .ZN(n13247) );
  NAND2_X1 U16499 ( .A1(n13225), .A2(n13247), .ZN(P2_U2976) );
  AOI22_X1 U16500 ( .A1(n9582), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n19033), .ZN(n13226) );
  INV_X1 U16501 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16191) );
  INV_X1 U16502 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18058) );
  AOI22_X1 U16503 ( .A1(n15405), .A2(n16191), .B1(n18058), .B2(n15407), .ZN(
        n15895) );
  NAND2_X1 U16504 ( .A1(n19031), .A2(n15895), .ZN(n13257) );
  NAND2_X1 U16505 ( .A1(n13226), .A2(n13257), .ZN(P2_U2971) );
  AOI22_X1 U16506 ( .A1(n9582), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n19033), .ZN(n13228) );
  AOI22_X1 U16507 ( .A1(n15405), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13263), .ZN(n19066) );
  INV_X1 U16508 ( .A(n19066), .ZN(n13227) );
  NAND2_X1 U16509 ( .A1(n19031), .A2(n13227), .ZN(n13259) );
  NAND2_X1 U16510 ( .A1(n13228), .A2(n13259), .ZN(P2_U2970) );
  AOI22_X1 U16511 ( .A1(n9582), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_2__SCAN_IN), .B2(n19033), .ZN(n13229) );
  OAI22_X1 U16512 ( .A1(n13263), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n15405), .ZN(n19062) );
  INV_X1 U16513 ( .A(n19062), .ZN(n15902) );
  NAND2_X1 U16514 ( .A1(n19031), .A2(n15902), .ZN(n13261) );
  NAND2_X1 U16515 ( .A1(n13229), .A2(n13261), .ZN(P2_U2969) );
  AOI22_X1 U16516 ( .A1(n9582), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19033), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n13231) );
  AOI22_X1 U16517 ( .A1(n15405), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n15407), .ZN(n19056) );
  INV_X1 U16518 ( .A(n19056), .ZN(n13230) );
  NAND2_X1 U16519 ( .A1(n19031), .A2(n13230), .ZN(n13255) );
  NAND2_X1 U16520 ( .A1(n13231), .A2(n13255), .ZN(P2_U2968) );
  AOI22_X1 U16521 ( .A1(n9582), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_0__SCAN_IN), .B2(n19033), .ZN(n13233) );
  INV_X1 U16522 ( .A(n19050), .ZN(n18925) );
  NAND2_X1 U16523 ( .A1(n19031), .A2(n18925), .ZN(n13245) );
  NAND2_X1 U16524 ( .A1(n13233), .A2(n13245), .ZN(P2_U2967) );
  AOI22_X1 U16525 ( .A1(n9582), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n19033), .ZN(n13236) );
  INV_X1 U16526 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n13996) );
  OR2_X1 U16527 ( .A1(n13263), .A2(n13996), .ZN(n13235) );
  NAND2_X1 U16528 ( .A1(n13263), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13234) );
  AND2_X1 U16529 ( .A1(n13235), .A2(n13234), .ZN(n18941) );
  INV_X1 U16530 ( .A(n18941), .ZN(n14845) );
  NAND2_X1 U16531 ( .A1(n19031), .A2(n14845), .ZN(n13237) );
  NAND2_X1 U16532 ( .A1(n13236), .A2(n13237), .ZN(P2_U2980) );
  AOI22_X1 U16533 ( .A1(n9582), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n19033), .ZN(n13238) );
  NAND2_X1 U16534 ( .A1(n13238), .A2(n13237), .ZN(P2_U2965) );
  AOI22_X1 U16535 ( .A1(n9582), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(
        P2_EAX_REG_28__SCAN_IN), .B2(n19033), .ZN(n13240) );
  NAND2_X1 U16536 ( .A1(n13240), .A2(n13239), .ZN(P2_U2964) );
  AOI22_X1 U16537 ( .A1(n9582), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n19033), .ZN(n13242) );
  NAND2_X1 U16538 ( .A1(n13242), .A2(n13241), .ZN(P2_U2963) );
  AOI22_X1 U16539 ( .A1(n9582), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19033), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n13244) );
  NAND2_X1 U16540 ( .A1(n13244), .A2(n13243), .ZN(P2_U2957) );
  AOI22_X1 U16541 ( .A1(n9582), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_16__SCAN_IN), .B2(n19033), .ZN(n13246) );
  NAND2_X1 U16542 ( .A1(n13246), .A2(n13245), .ZN(P2_U2952) );
  AOI22_X1 U16543 ( .A1(n9582), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n19033), .ZN(n13248) );
  NAND2_X1 U16544 ( .A1(n13248), .A2(n13247), .ZN(P2_U2961) );
  AOI22_X1 U16545 ( .A1(n9582), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(
        P2_EAX_REG_24__SCAN_IN), .B2(n19033), .ZN(n13250) );
  NAND2_X1 U16546 ( .A1(n13250), .A2(n13249), .ZN(P2_U2960) );
  AOI22_X1 U16547 ( .A1(n9582), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19033), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n13252) );
  NAND2_X1 U16548 ( .A1(n13252), .A2(n13251), .ZN(P2_U2959) );
  AOI22_X1 U16549 ( .A1(n9582), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n19033), .ZN(n13254) );
  NAND2_X1 U16550 ( .A1(n13254), .A2(n13253), .ZN(P2_U2958) );
  AOI22_X1 U16551 ( .A1(n9582), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19033), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n13256) );
  NAND2_X1 U16552 ( .A1(n13256), .A2(n13255), .ZN(P2_U2953) );
  AOI22_X1 U16553 ( .A1(n9582), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n19033), .ZN(n13258) );
  NAND2_X1 U16554 ( .A1(n13258), .A2(n13257), .ZN(P2_U2956) );
  AOI22_X1 U16555 ( .A1(n9582), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19033), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n13260) );
  NAND2_X1 U16556 ( .A1(n13260), .A2(n13259), .ZN(P2_U2955) );
  AOI22_X1 U16557 ( .A1(n9582), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n19033), .ZN(n13262) );
  NAND2_X1 U16558 ( .A1(n13262), .A2(n13261), .ZN(P2_U2954) );
  INV_X1 U16559 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19006) );
  NAND2_X1 U16560 ( .A1(n13263), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13265) );
  INV_X1 U16561 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16181) );
  OR2_X1 U16562 ( .A1(n13263), .A2(n16181), .ZN(n13264) );
  NAND2_X1 U16563 ( .A1(n13265), .A2(n13264), .ZN(n18947) );
  NAND2_X1 U16564 ( .A1(n19031), .A2(n18947), .ZN(n13268) );
  NAND2_X1 U16565 ( .A1(n9582), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13266) );
  OAI211_X1 U16566 ( .C1(n19006), .C2(n13269), .A(n13268), .B(n13266), .ZN(
        P2_U2977) );
  NAND2_X1 U16567 ( .A1(n9582), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13267) );
  OAI211_X1 U16568 ( .C1(n13270), .C2(n13269), .A(n13268), .B(n13267), .ZN(
        P2_U2962) );
  NOR2_X1 U16569 ( .A1(n13271), .A2(n20786), .ZN(n13272) );
  OR2_X2 U16570 ( .A1(n13326), .A2(n13272), .ZN(n19974) );
  OR2_X1 U16571 ( .A1(n19974), .A2(n13325), .ZN(n13462) );
  INV_X1 U16572 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14039) );
  NAND2_X1 U16573 ( .A1(n13466), .A2(n13325), .ZN(n13331) );
  INV_X1 U16574 ( .A(DATAI_15_), .ZN(n13273) );
  NOR2_X1 U16575 ( .A1(n20068), .A2(n13273), .ZN(n13274) );
  AOI21_X1 U16576 ( .B1(n20068), .B2(BUF1_REG_15__SCAN_IN), .A(n13274), .ZN(
        n14037) );
  INV_X1 U16577 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n19921) );
  OAI222_X1 U16578 ( .A1(n13462), .A2(n14039), .B1(n13331), .B2(n14037), .C1(
        n13466), .C2(n19921), .ZN(P1_U2967) );
  NOR2_X1 U16579 ( .A1(n20956), .A2(n10143), .ZN(n13279) );
  AOI21_X1 U16580 ( .B1(n11061), .B2(n20956), .A(n13279), .ZN(n13280) );
  OAI21_X1 U16581 ( .B1(n19761), .B2(n18919), .A(n13280), .ZN(P2_U2884) );
  INV_X2 U16582 ( .A(n20956), .ZN(n20964) );
  MUX2_X1 U16583 ( .A(n15355), .B(n11161), .S(n20964), .Z(n13281) );
  OAI21_X1 U16584 ( .B1(n19792), .B2(n18919), .A(n13281), .ZN(P2_U2887) );
  OAI21_X1 U16585 ( .B1(n13283), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13282), .ZN(n20051) );
  INV_X1 U16586 ( .A(n13284), .ZN(n13285) );
  AOI21_X1 U16587 ( .B1(n13287), .B2(n13286), .A(n13285), .ZN(n13664) );
  NAND2_X1 U16588 ( .A1(n13664), .A2(n13319), .ZN(n13291) );
  NAND2_X1 U16589 ( .A1(n13288), .A2(n14592), .ZN(n13289) );
  AOI22_X1 U16590 ( .A1(n20053), .A2(P1_REIP_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n13289), .ZN(n13290) );
  OAI211_X1 U16591 ( .C1(n19822), .C2(n20051), .A(n13291), .B(n13290), .ZN(
        P1_U2999) );
  NAND2_X1 U16592 ( .A1(n13562), .A2(n15484), .ZN(n13443) );
  OR2_X1 U16593 ( .A1(n13293), .A2(n13292), .ZN(n13294) );
  NAND2_X1 U16594 ( .A1(n13443), .A2(n13294), .ZN(n13296) );
  AND2_X2 U16595 ( .A1(n13296), .A2(n13295), .ZN(n19918) );
  NAND2_X1 U16596 ( .A1(n19918), .A2(n13381), .ZN(n14406) );
  NAND2_X1 U16597 ( .A1(n19918), .A2(n20109), .ZN(n14401) );
  OAI22_X1 U16598 ( .A1(n14401), .A2(n13298), .B1(n13297), .B2(n19918), .ZN(
        n13299) );
  INV_X1 U16599 ( .A(n13299), .ZN(n13300) );
  OAI21_X1 U16600 ( .B1(n13534), .B2(n14406), .A(n13300), .ZN(P1_U2871) );
  MUX2_X1 U16601 ( .A(n13735), .B(n11040), .S(n20956), .Z(n13303) );
  OAI21_X1 U16602 ( .B1(n19770), .B2(n18919), .A(n13303), .ZN(P2_U2885) );
  INV_X1 U16603 ( .A(n13396), .ZN(n13313) );
  OAI21_X1 U16604 ( .B1(n15352), .B2(n13305), .A(n13304), .ZN(n13312) );
  INV_X1 U16605 ( .A(n15225), .ZN(n15206) );
  OAI211_X1 U16606 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n15206), .B(n13398), .ZN(n13310) );
  XNOR2_X1 U16607 ( .A(n13306), .B(n13307), .ZN(n19786) );
  AOI22_X1 U16608 ( .A1(n16010), .A2(n19786), .B1(n16015), .B2(n13308), .ZN(
        n13309) );
  NAND2_X1 U16609 ( .A1(n13310), .A2(n13309), .ZN(n13311) );
  AOI211_X1 U16610 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n13313), .A(
        n13312), .B(n13311), .ZN(n13314) );
  OAI21_X1 U16611 ( .B1(n11070), .B2(n15343), .A(n13314), .ZN(P2_U3045) );
  OR2_X1 U16612 ( .A1(n13315), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13317) );
  NAND2_X1 U16613 ( .A1(n13317), .A2(n13316), .ZN(n20048) );
  INV_X1 U16614 ( .A(n13664), .ZN(n13389) );
  OAI222_X1 U16615 ( .A1(n20048), .A2(n14401), .B1(n13318), .B2(n19918), .C1(
        n13389), .C2(n14406), .ZN(P1_U2872) );
  INV_X1 U16616 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13321) );
  OAI22_X1 U16617 ( .A1(n14592), .A2(n13321), .B1(n20035), .B2(n20775), .ZN(
        n13320) );
  AOI21_X1 U16618 ( .B1(n15647), .B2(n13321), .A(n13320), .ZN(n13324) );
  OR2_X1 U16619 ( .A1(n13322), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20037) );
  NAND3_X1 U16620 ( .A1(n20037), .A2(n20038), .A3(n19990), .ZN(n13323) );
  OAI211_X1 U16621 ( .C1(n13534), .C2(n20067), .A(n13324), .B(n13323), .ZN(
        P1_U2998) );
  INV_X1 U16622 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13330) );
  OR2_X1 U16623 ( .A1(n15484), .A2(n19815), .ZN(n13327) );
  OAI22_X1 U16624 ( .A1(n15462), .A2(n13327), .B1(n13326), .B2(n13325), .ZN(
        n13328) );
  INV_X1 U16625 ( .A(n15505), .ZN(n15479) );
  NAND2_X1 U16626 ( .A1(n19922), .A2(n12697), .ZN(n13558) );
  NOR2_X1 U16627 ( .A1(n20074), .A2(n13584), .ZN(n15802) );
  NAND2_X1 U16628 ( .A1(n20071), .A2(n15802), .ZN(n19920) );
  AOI22_X1 U16629 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n19934), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n19930), .ZN(n13329) );
  OAI21_X1 U16630 ( .B1(n13330), .B2(n13558), .A(n13329), .ZN(P1_U2907) );
  INV_X1 U16631 ( .A(DATAI_12_), .ZN(n13333) );
  MUX2_X1 U16632 ( .A(n13333), .B(n13332), .S(n20068), .Z(n14412) );
  INV_X1 U16633 ( .A(n14412), .ZN(n13334) );
  NAND2_X1 U16634 ( .A1(n19966), .A2(n13334), .ZN(n19977) );
  NAND2_X1 U16635 ( .A1(n19974), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n13335) );
  OAI211_X1 U16636 ( .C1(n13462), .C2(n14411), .A(n19977), .B(n13335), .ZN(
        P1_U2949) );
  AOI22_X1 U16637 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n19930), .B1(n19934), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13336) );
  OAI21_X1 U16638 ( .B1(n14411), .B2(n13558), .A(n13336), .ZN(P1_U2908) );
  INV_X1 U16639 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13338) );
  AOI22_X1 U16640 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n19930), .B1(n19934), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13337) );
  OAI21_X1 U16641 ( .B1(n13338), .B2(n13558), .A(n13337), .ZN(P1_U2911) );
  AOI22_X1 U16642 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n19930), .B1(n19934), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13339) );
  OAI21_X1 U16643 ( .B1(n14427), .B2(n13558), .A(n13339), .ZN(P1_U2912) );
  INV_X1 U16644 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13341) );
  AOI22_X1 U16645 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n19930), .B1(n19934), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13340) );
  OAI21_X1 U16646 ( .B1(n13341), .B2(n13558), .A(n13340), .ZN(P1_U2909) );
  INV_X1 U16647 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13343) );
  AOI22_X1 U16648 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n19930), .B1(n19934), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13342) );
  OAI21_X1 U16649 ( .B1(n13343), .B2(n13558), .A(n13342), .ZN(P1_U2913) );
  NAND2_X1 U16650 ( .A1(n18872), .A2(n13351), .ZN(n13344) );
  NAND2_X1 U16651 ( .A1(n13345), .A2(n13344), .ZN(n14128) );
  OAI21_X1 U16652 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n13347), .A(
        n13346), .ZN(n14130) );
  OAI22_X1 U16653 ( .A1(n15234), .A2(n14128), .B1(n15352), .B2(n14130), .ZN(
        n13350) );
  INV_X1 U16654 ( .A(n15343), .ZN(n16014) );
  AOI22_X1 U16655 ( .A1(n18875), .A2(n16014), .B1(n16010), .B2(n18868), .ZN(
        n13348) );
  NAND2_X1 U16656 ( .A1(n19038), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n14129) );
  OAI211_X1 U16657 ( .C1(n13351), .C2(n13396), .A(n13348), .B(n14129), .ZN(
        n13349) );
  AOI211_X1 U16658 ( .C1(n13351), .C2(n15206), .A(n13350), .B(n13349), .ZN(
        n13352) );
  INV_X1 U16659 ( .A(n13352), .ZN(P2_U3046) );
  INV_X1 U16660 ( .A(n19761), .ZN(n13364) );
  AND2_X1 U16661 ( .A1(n16041), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16071) );
  INV_X1 U16662 ( .A(n15373), .ZN(n15387) );
  NAND2_X1 U16663 ( .A1(n13278), .A2(n15387), .ZN(n13363) );
  NOR2_X1 U16664 ( .A1(n11616), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13354) );
  NOR2_X1 U16665 ( .A1(n10280), .A2(n13354), .ZN(n13361) );
  AND2_X1 U16666 ( .A1(n16042), .A2(n16037), .ZN(n15384) );
  NOR2_X1 U16667 ( .A1(n13355), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15377) );
  XNOR2_X1 U16668 ( .A(n15377), .B(n10156), .ZN(n13359) );
  INV_X1 U16669 ( .A(n13356), .ZN(n13357) );
  OAI211_X1 U16670 ( .C1(n10092), .C2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n15379), .B(n13357), .ZN(n13358) );
  OAI21_X1 U16671 ( .B1(n15384), .B2(n13359), .A(n13358), .ZN(n13360) );
  AOI21_X1 U16672 ( .B1(n15378), .B2(n13361), .A(n13360), .ZN(n13362) );
  NAND2_X1 U16673 ( .A1(n13363), .A2(n13362), .ZN(n16029) );
  AOI22_X1 U16674 ( .A1(n13364), .A2(n16071), .B1(n19758), .B2(n16029), .ZN(
        n13380) );
  NAND2_X1 U16675 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13365), .ZN(n16079) );
  INV_X1 U16676 ( .A(n16079), .ZN(n16064) );
  NAND2_X1 U16677 ( .A1(n13367), .A2(n13366), .ZN(n13369) );
  NOR2_X1 U16678 ( .A1(n13369), .A2(n13368), .ZN(n13376) );
  INV_X1 U16679 ( .A(n16047), .ZN(n13370) );
  OAI21_X1 U16680 ( .B1(n13372), .B2(n13371), .A(n13370), .ZN(n13374) );
  NAND2_X1 U16681 ( .A1(n13374), .A2(n13373), .ZN(n13375) );
  AND2_X1 U16682 ( .A1(n13376), .A2(n13375), .ZN(n16054) );
  OAI21_X1 U16683 ( .B1(n16054), .B2(n16076), .A(n13377), .ZN(n13378) );
  AOI21_X1 U16684 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16064), .A(n13378), .ZN(
        n15393) );
  NAND2_X1 U16685 ( .A1(n15393), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13379) );
  OAI21_X1 U16686 ( .B1(n13380), .B2(n15393), .A(n13379), .ZN(P2_U3596) );
  AND2_X1 U16687 ( .A1(n20099), .A2(n13381), .ZN(n13386) );
  NOR2_X1 U16688 ( .A1(n13386), .A2(n13382), .ZN(n13383) );
  INV_X1 U16689 ( .A(DATAI_0_), .ZN(n13385) );
  NAND2_X1 U16690 ( .A1(n20068), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13384) );
  OAI21_X1 U16691 ( .B1(n20068), .B2(n13385), .A(n13384), .ZN(n20073) );
  INV_X1 U16692 ( .A(n20073), .ZN(n13388) );
  NAND2_X1 U16693 ( .A1(n14428), .A2(n13386), .ZN(n14429) );
  INV_X1 U16694 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n19948) );
  OAI222_X1 U16695 ( .A1(n14434), .A2(n13389), .B1(n13388), .B2(n14038), .C1(
        n14428), .C2(n19948), .ZN(P1_U2904) );
  NAND2_X1 U16696 ( .A1(n13391), .A2(n13390), .ZN(n13394) );
  INV_X1 U16697 ( .A(n13392), .ZN(n13393) );
  AND2_X1 U16698 ( .A1(n13394), .A2(n13393), .ZN(n19772) );
  INV_X1 U16699 ( .A(n19772), .ZN(n13733) );
  INV_X1 U16700 ( .A(n13398), .ZN(n13395) );
  OR2_X1 U16701 ( .A1(n15221), .A2(n13395), .ZN(n13397) );
  OAI211_X1 U16702 ( .C1(n15223), .C2(n13398), .A(n13397), .B(n13396), .ZN(
        n13401) );
  NOR2_X1 U16703 ( .A1(n15221), .A2(n13398), .ZN(n13400) );
  MUX2_X1 U16704 ( .A(n13401), .B(n13400), .S(n13399), .Z(n13408) );
  AOI21_X1 U16705 ( .B1(n13403), .B2(n16011), .A(n13402), .ZN(n13405) );
  OAI211_X1 U16706 ( .C1(n15234), .C2(n13406), .A(n13405), .B(n13404), .ZN(
        n13407) );
  AOI211_X1 U16707 ( .C1(n13733), .C2(n16010), .A(n13408), .B(n13407), .ZN(
        n13409) );
  OAI21_X1 U16708 ( .B1(n11040), .B2(n15343), .A(n13409), .ZN(P2_U3044) );
  AND2_X1 U16709 ( .A1(n13410), .A2(n13411), .ZN(n18912) );
  INV_X1 U16710 ( .A(n18919), .ZN(n18891) );
  NAND2_X1 U16711 ( .A1(n13410), .A2(n13412), .ZN(n18904) );
  OAI211_X1 U16712 ( .C1(n18912), .C2(n13413), .A(n18891), .B(n18904), .ZN(
        n13417) );
  NOR2_X1 U16713 ( .A1(n13775), .A2(n13414), .ZN(n13415) );
  OR2_X1 U16714 ( .A1(n13787), .A2(n13415), .ZN(n18843) );
  INV_X1 U16715 ( .A(n18843), .ZN(n15980) );
  NAND2_X1 U16716 ( .A1(n15980), .A2(n20956), .ZN(n13416) );
  OAI211_X1 U16717 ( .C1(n20956), .C2(n10611), .A(n13417), .B(n13416), .ZN(
        P2_U2878) );
  INV_X1 U16718 ( .A(n20571), .ZN(n20580) );
  INV_X1 U16719 ( .A(n13418), .ZN(n13420) );
  NAND3_X1 U16720 ( .A1(n13420), .A2(n13433), .A3(n13419), .ZN(n13421) );
  NOR2_X1 U16721 ( .A1(n13422), .A2(n13421), .ZN(n13423) );
  AND2_X1 U16722 ( .A1(n13423), .A2(n15793), .ZN(n15461) );
  INV_X1 U16723 ( .A(n15461), .ZN(n13582) );
  NAND2_X1 U16724 ( .A1(n20580), .A2(n13582), .ZN(n13429) );
  INV_X1 U16725 ( .A(n13424), .ZN(n13587) );
  INV_X1 U16726 ( .A(n13425), .ZN(n13426) );
  NAND3_X1 U16727 ( .A1(n13427), .A2(n13587), .A3(n13426), .ZN(n13428) );
  OAI211_X1 U16728 ( .C1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n15462), .A(
        n13429), .B(n13428), .ZN(n15459) );
  INV_X1 U16729 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20756) );
  NAND2_X1 U16730 ( .A1(n13587), .A2(n14696), .ZN(n13430) );
  AOI22_X1 U16731 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n20044), .B2(n20891), .ZN(
        n14695) );
  NAND2_X1 U16732 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14694) );
  OAI22_X1 U16733 ( .A1(n13430), .A2(n13425), .B1(n14695), .B2(n14694), .ZN(
        n13431) );
  AOI21_X1 U16734 ( .B1(n15459), .B2(n15796), .A(n13431), .ZN(n13446) );
  INV_X1 U16735 ( .A(n20786), .ZN(n20693) );
  OR2_X1 U16736 ( .A1(n15505), .A2(n20693), .ZN(n13432) );
  AOI21_X1 U16737 ( .B1(n15462), .B2(n13433), .A(n13432), .ZN(n13436) );
  OAI21_X1 U16738 ( .B1(n13436), .B2(n13435), .A(n13434), .ZN(n13444) );
  NOR2_X1 U16739 ( .A1(n13438), .A2(n13437), .ZN(n13439) );
  NOR2_X1 U16740 ( .A1(n13440), .A2(n13439), .ZN(n13442) );
  NAND4_X1 U16741 ( .A1(n13444), .A2(n13443), .A3(n13442), .A4(n13441), .ZN(
        n15458) );
  INV_X1 U16742 ( .A(n15458), .ZN(n13590) );
  NAND2_X1 U16743 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15802), .ZN(n15808) );
  INV_X1 U16744 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19823) );
  OAI22_X1 U16745 ( .A1(n13590), .A2(n19815), .B1(n15808), .B2(n19823), .ZN(
        n15794) );
  AOI21_X1 U16746 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20071), .A(n15794), 
        .ZN(n20763) );
  NAND2_X1 U16747 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20763), .ZN(
        n13445) );
  OAI21_X1 U16748 ( .B1(n13446), .B2(n20763), .A(n13445), .ZN(P1_U3473) );
  OR2_X1 U16749 ( .A1(n13447), .A2(n9657), .ZN(n13449) );
  NAND2_X1 U16750 ( .A1(n13449), .A2(n13448), .ZN(n13952) );
  NAND2_X1 U16751 ( .A1(n13410), .A2(n18909), .ZN(n14187) );
  NOR2_X1 U16752 ( .A1(n14187), .A2(n13450), .ZN(n13452) );
  OR2_X1 U16753 ( .A1(n14187), .A2(n13451), .ZN(n13455) );
  OAI211_X1 U16754 ( .C1(n13452), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n18891), .B(n13455), .ZN(n13454) );
  NAND2_X1 U16755 ( .A1(n20964), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n13453) );
  OAI211_X1 U16756 ( .C1(n13952), .C2(n20964), .A(n13454), .B(n13453), .ZN(
        P2_U2881) );
  XOR2_X1 U16757 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n13455), .Z(n13461)
         );
  NAND2_X1 U16758 ( .A1(n13456), .A2(n13448), .ZN(n13459) );
  INV_X1 U16759 ( .A(n13457), .ZN(n13458) );
  NAND2_X1 U16760 ( .A1(n13459), .A2(n13458), .ZN(n18857) );
  MUX2_X1 U16761 ( .A(n10602), .B(n18857), .S(n20956), .Z(n13460) );
  OAI21_X1 U16762 ( .B1(n13461), .B2(n18919), .A(n13460), .ZN(P2_U2880) );
  INV_X2 U16763 ( .A(n13462), .ZN(n19981) );
  AOI22_X1 U16764 ( .A1(n19981), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n19974), .ZN(n13465) );
  INV_X1 U16765 ( .A(DATAI_6_), .ZN(n13464) );
  NAND2_X1 U16766 ( .A1(n20068), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13463) );
  OAI21_X1 U16767 ( .B1(n20068), .B2(n13464), .A(n13463), .ZN(n20105) );
  NAND2_X1 U16768 ( .A1(n19966), .A2(n20105), .ZN(n13470) );
  NAND2_X1 U16769 ( .A1(n13465), .A2(n13470), .ZN(P1_U2958) );
  AOI22_X1 U16770 ( .A1(n19981), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n19974), .ZN(n13469) );
  INV_X1 U16771 ( .A(DATAI_2_), .ZN(n13468) );
  NAND2_X1 U16772 ( .A1(n20068), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13467) );
  OAI21_X1 U16773 ( .B1(n20068), .B2(n13468), .A(n13467), .ZN(n20086) );
  NAND2_X1 U16774 ( .A1(n19966), .A2(n20086), .ZN(n13492) );
  NAND2_X1 U16775 ( .A1(n13469), .A2(n13492), .ZN(P1_U2939) );
  AOI22_X1 U16776 ( .A1(n19981), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n19974), .ZN(n13471) );
  NAND2_X1 U16777 ( .A1(n13471), .A2(n13470), .ZN(P1_U2943) );
  AOI22_X1 U16778 ( .A1(n19981), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n19974), .ZN(n13474) );
  INV_X1 U16779 ( .A(DATAI_7_), .ZN(n13473) );
  NAND2_X1 U16780 ( .A1(n20068), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13472) );
  OAI21_X1 U16781 ( .B1(n20068), .B2(n13473), .A(n13472), .ZN(n20113) );
  NAND2_X1 U16782 ( .A1(n19966), .A2(n20113), .ZN(n13475) );
  NAND2_X1 U16783 ( .A1(n13474), .A2(n13475), .ZN(P1_U2959) );
  AOI22_X1 U16784 ( .A1(n19981), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n19974), .ZN(n13476) );
  NAND2_X1 U16785 ( .A1(n13476), .A2(n13475), .ZN(P1_U2944) );
  AOI22_X1 U16786 ( .A1(n19981), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n19974), .ZN(n13479) );
  INV_X1 U16787 ( .A(DATAI_3_), .ZN(n13478) );
  NAND2_X1 U16788 ( .A1(n20068), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13477) );
  OAI21_X1 U16789 ( .B1(n20068), .B2(n13478), .A(n13477), .ZN(n20091) );
  NAND2_X1 U16790 ( .A1(n19966), .A2(n20091), .ZN(n13494) );
  NAND2_X1 U16791 ( .A1(n13479), .A2(n13494), .ZN(P1_U2940) );
  AOI22_X1 U16792 ( .A1(n19981), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n19974), .ZN(n13482) );
  INV_X1 U16793 ( .A(DATAI_4_), .ZN(n13481) );
  NAND2_X1 U16794 ( .A1(n20068), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13480) );
  OAI21_X1 U16795 ( .B1(n20068), .B2(n13481), .A(n13480), .ZN(n20095) );
  NAND2_X1 U16796 ( .A1(n19966), .A2(n20095), .ZN(n13496) );
  NAND2_X1 U16797 ( .A1(n13482), .A2(n13496), .ZN(P1_U2941) );
  AOI22_X1 U16798 ( .A1(n19981), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n19974), .ZN(n13483) );
  NAND2_X1 U16799 ( .A1(n19966), .A2(n20073), .ZN(n13487) );
  NAND2_X1 U16800 ( .A1(n13483), .A2(n13487), .ZN(P1_U2937) );
  AOI22_X1 U16801 ( .A1(n19981), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n19974), .ZN(n13486) );
  INV_X1 U16802 ( .A(DATAI_5_), .ZN(n13485) );
  NAND2_X1 U16803 ( .A1(n20068), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13484) );
  OAI21_X1 U16804 ( .B1(n20068), .B2(n13485), .A(n13484), .ZN(n20100) );
  NAND2_X1 U16805 ( .A1(n19966), .A2(n20100), .ZN(n13500) );
  NAND2_X1 U16806 ( .A1(n13486), .A2(n13500), .ZN(P1_U2942) );
  AOI22_X1 U16807 ( .A1(n19981), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n19974), .ZN(n13488) );
  NAND2_X1 U16808 ( .A1(n13488), .A2(n13487), .ZN(P1_U2952) );
  AOI22_X1 U16809 ( .A1(n19981), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n19974), .ZN(n13491) );
  INV_X1 U16810 ( .A(DATAI_1_), .ZN(n13490) );
  NAND2_X1 U16811 ( .A1(n20068), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13489) );
  OAI21_X1 U16812 ( .B1(n20068), .B2(n13490), .A(n13489), .ZN(n20081) );
  NAND2_X1 U16813 ( .A1(n19966), .A2(n20081), .ZN(n13498) );
  NAND2_X1 U16814 ( .A1(n13491), .A2(n13498), .ZN(P1_U2953) );
  AOI22_X1 U16815 ( .A1(n19981), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n19974), .ZN(n13493) );
  NAND2_X1 U16816 ( .A1(n13493), .A2(n13492), .ZN(P1_U2954) );
  AOI22_X1 U16817 ( .A1(n19981), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n19974), .ZN(n13495) );
  NAND2_X1 U16818 ( .A1(n13495), .A2(n13494), .ZN(P1_U2955) );
  AOI22_X1 U16819 ( .A1(n19981), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n19974), .ZN(n13497) );
  NAND2_X1 U16820 ( .A1(n13497), .A2(n13496), .ZN(P1_U2956) );
  AOI22_X1 U16821 ( .A1(n19981), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n19974), .ZN(n13499) );
  NAND2_X1 U16822 ( .A1(n13499), .A2(n13498), .ZN(P1_U2938) );
  AOI22_X1 U16823 ( .A1(n19981), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n19974), .ZN(n13501) );
  NAND2_X1 U16824 ( .A1(n13501), .A2(n13500), .ZN(P1_U2957) );
  XNOR2_X1 U16825 ( .A(n19770), .B(n19772), .ZN(n13506) );
  INV_X1 U16826 ( .A(n19786), .ZN(n13502) );
  NAND2_X1 U16827 ( .A1(n15396), .A2(n13502), .ZN(n13503) );
  OAI21_X1 U16828 ( .B1(n15396), .B2(n13502), .A(n13503), .ZN(n18984) );
  NOR2_X1 U16829 ( .A1(n18984), .A2(n18985), .ZN(n18983) );
  INV_X1 U16830 ( .A(n13503), .ZN(n13504) );
  NOR2_X1 U16831 ( .A1(n18983), .A2(n13504), .ZN(n13505) );
  NOR2_X1 U16832 ( .A1(n13505), .A2(n13506), .ZN(n18960) );
  AOI21_X1 U16833 ( .B1(n13506), .B2(n13505), .A(n18960), .ZN(n13509) );
  AOI22_X1 U16834 ( .A1(n18958), .A2(n15902), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n18981), .ZN(n13508) );
  NAND2_X1 U16835 ( .A1(n13733), .A2(n18982), .ZN(n13507) );
  OAI211_X1 U16836 ( .C1(n13509), .C2(n18986), .A(n13508), .B(n13507), .ZN(
        P2_U2917) );
  OAI22_X1 U16837 ( .A1(n14401), .A2(n20024), .B1(n13510), .B2(n19918), .ZN(
        n13511) );
  AOI21_X1 U16838 ( .B1(n13521), .B2(n19914), .A(n13511), .ZN(n13512) );
  INV_X1 U16839 ( .A(n13512), .ZN(P1_U2870) );
  AOI22_X1 U16840 ( .A1(n19984), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20053), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13513) );
  OAI21_X1 U16841 ( .B1(n19995), .B2(n13514), .A(n13513), .ZN(n13520) );
  NOR2_X1 U16842 ( .A1(n13515), .A2(n13516), .ZN(n20019) );
  INV_X1 U16843 ( .A(n13517), .ZN(n13518) );
  NOR3_X1 U16844 ( .A1(n20019), .A2(n13518), .A3(n19822), .ZN(n13519) );
  AOI211_X1 U16845 ( .C1(n13319), .C2(n13521), .A(n13520), .B(n13519), .ZN(
        n13522) );
  INV_X1 U16846 ( .A(n13522), .ZN(P1_U2997) );
  AND2_X1 U16847 ( .A1(n13410), .A2(n13523), .ZN(n18903) );
  XNOR2_X1 U16848 ( .A(n18903), .B(n18897), .ZN(n13530) );
  NAND2_X1 U16849 ( .A1(n13524), .A2(n13785), .ZN(n13527) );
  INV_X1 U16850 ( .A(n13525), .ZN(n13526) );
  AND2_X1 U16851 ( .A1(n13527), .A2(n13526), .ZN(n15965) );
  INV_X1 U16852 ( .A(n15965), .ZN(n18822) );
  MUX2_X1 U16853 ( .A(n13528), .B(n18822), .S(n20956), .Z(n13529) );
  OAI21_X1 U16854 ( .B1(n13530), .B2(n18919), .A(n13529), .ZN(P2_U2876) );
  INV_X1 U16855 ( .A(n20086), .ZN(n13531) );
  INV_X1 U16856 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n19942) );
  OAI222_X1 U16857 ( .A1(n14434), .A2(n13532), .B1(n13531), .B2(n14038), .C1(
        n14428), .C2(n19942), .ZN(P1_U2902) );
  INV_X1 U16858 ( .A(n20081), .ZN(n13533) );
  INV_X1 U16859 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n19944) );
  OAI222_X1 U16860 ( .A1(n14434), .A2(n13534), .B1(n13533), .B2(n14038), .C1(
        n14428), .C2(n19944), .ZN(P1_U2903) );
  XNOR2_X1 U16861 ( .A(n13535), .B(n13536), .ZN(n19905) );
  INV_X1 U16862 ( .A(n20091), .ZN(n13537) );
  INV_X1 U16863 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n19940) );
  OAI222_X1 U16864 ( .A1(n14434), .A2(n19905), .B1(n13537), .B2(n14038), .C1(
        n14428), .C2(n19940), .ZN(P1_U2901) );
  AOI21_X1 U16865 ( .B1(n13539), .B2(n13538), .A(n13616), .ZN(n20010) );
  INV_X1 U16866 ( .A(n20010), .ZN(n13540) );
  INV_X1 U16867 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n19896) );
  OAI222_X1 U16868 ( .A1(n13540), .A2(n14401), .B1(n19896), .B2(n19918), .C1(
        n19905), .C2(n14406), .ZN(P1_U2869) );
  INV_X1 U16869 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13542) );
  AOI22_X1 U16870 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n19930), .B1(n19945), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13541) );
  OAI21_X1 U16871 ( .B1(n13542), .B2(n13558), .A(n13541), .ZN(P1_U2914) );
  INV_X1 U16872 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13544) );
  AOI22_X1 U16873 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n19930), .B1(n19945), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13543) );
  OAI21_X1 U16874 ( .B1(n13544), .B2(n13558), .A(n13543), .ZN(P1_U2906) );
  INV_X1 U16875 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13546) );
  AOI22_X1 U16876 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n19930), .B1(n19945), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13545) );
  OAI21_X1 U16877 ( .B1(n13546), .B2(n13558), .A(n13545), .ZN(P1_U2910) );
  INV_X1 U16878 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13548) );
  AOI22_X1 U16879 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n19930), .B1(n19945), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13547) );
  OAI21_X1 U16880 ( .B1(n13548), .B2(n13558), .A(n13547), .ZN(P1_U2920) );
  INV_X1 U16881 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13550) );
  AOI22_X1 U16882 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n19930), .B1(n19945), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13549) );
  OAI21_X1 U16883 ( .B1(n13550), .B2(n13558), .A(n13549), .ZN(P1_U2918) );
  INV_X1 U16884 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13552) );
  AOI22_X1 U16885 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n19930), .B1(n19945), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13551) );
  OAI21_X1 U16886 ( .B1(n13552), .B2(n13558), .A(n13551), .ZN(P1_U2917) );
  INV_X1 U16887 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13554) );
  AOI22_X1 U16888 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n19930), .B1(n19945), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13553) );
  OAI21_X1 U16889 ( .B1(n13554), .B2(n13558), .A(n13553), .ZN(P1_U2919) );
  INV_X1 U16890 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13556) );
  AOI22_X1 U16891 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n19930), .B1(n19945), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13555) );
  OAI21_X1 U16892 ( .B1(n13556), .B2(n13558), .A(n13555), .ZN(P1_U2915) );
  INV_X1 U16893 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13559) );
  AOI22_X1 U16894 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n19930), .B1(n19945), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13557) );
  OAI21_X1 U16895 ( .B1(n13559), .B2(n13558), .A(n13557), .ZN(P1_U2916) );
  NOR2_X1 U16896 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13584), .ZN(n13591) );
  INV_X1 U16897 ( .A(n20512), .ZN(n20063) );
  XNOR2_X1 U16898 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13566) );
  INV_X1 U16899 ( .A(n13560), .ZN(n13561) );
  OR2_X1 U16900 ( .A1(n13562), .A2(n13561), .ZN(n13573) );
  XNOR2_X1 U16901 ( .A(n13425), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13563) );
  NAND2_X1 U16902 ( .A1(n13573), .A2(n13563), .ZN(n13565) );
  INV_X1 U16903 ( .A(n13563), .ZN(n14697) );
  NAND3_X1 U16904 ( .A1(n15461), .A2(n13577), .A3(n14697), .ZN(n13564) );
  OAI211_X1 U16905 ( .C1(n15462), .C2(n13566), .A(n13565), .B(n13564), .ZN(
        n13567) );
  AOI21_X1 U16906 ( .B1(n20063), .B2(n13582), .A(n13567), .ZN(n14699) );
  INV_X1 U16907 ( .A(n14699), .ZN(n13568) );
  MUX2_X1 U16908 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13568), .S(
        n15458), .Z(n15469) );
  AOI22_X1 U16909 ( .A1(n13591), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15469), .B2(n13584), .ZN(n13586) );
  XNOR2_X1 U16910 ( .A(n13569), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13580) );
  MUX2_X1 U16911 ( .A(n11860), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n13425), .Z(n13571) );
  NOR2_X1 U16912 ( .A1(n13571), .A2(n13570), .ZN(n13572) );
  NAND2_X1 U16913 ( .A1(n13573), .A2(n13572), .ZN(n13579) );
  NOR2_X1 U16914 ( .A1(n13425), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13574) );
  NOR2_X1 U16915 ( .A1(n13574), .A2(n11860), .ZN(n13576) );
  AND2_X1 U16916 ( .A1(n13576), .A2(n13575), .ZN(n14701) );
  NAND3_X1 U16917 ( .A1(n15461), .A2(n13577), .A3(n14701), .ZN(n13578) );
  OAI211_X1 U16918 ( .C1(n15462), .C2(n13580), .A(n13579), .B(n13578), .ZN(
        n13581) );
  AOI21_X1 U16919 ( .B1(n20357), .B2(n13582), .A(n13581), .ZN(n14703) );
  NOR2_X1 U16920 ( .A1(n15458), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13583) );
  AOI21_X1 U16921 ( .B1(n14703), .B2(n15458), .A(n13583), .ZN(n15457) );
  AOI22_X1 U16922 ( .A1(n13591), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n13584), .B2(n15457), .ZN(n13585) );
  NOR2_X1 U16923 ( .A1(n13586), .A2(n13585), .ZN(n15477) );
  NAND2_X1 U16924 ( .A1(n15477), .A2(n13587), .ZN(n15487) );
  INV_X1 U16925 ( .A(n20234), .ZN(n20511) );
  NOR2_X1 U16926 ( .A1(n13588), .A2(n20511), .ZN(n13589) );
  XNOR2_X1 U16927 ( .A(n13589), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n15792) );
  OAI21_X1 U16928 ( .B1(n15792), .B2(n15793), .A(n15458), .ZN(n13593) );
  AOI21_X1 U16929 ( .B1(n13590), .B2(n15799), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n13592) );
  AOI22_X1 U16930 ( .A1(n13593), .A2(n13592), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n13591), .ZN(n15486) );
  AND3_X1 U16931 ( .A1(n15487), .A2(n15486), .A3(n19823), .ZN(n13594) );
  OAI21_X1 U16932 ( .B1(n13594), .B2(n15808), .A(n20242), .ZN(n20774) );
  INV_X1 U16933 ( .A(n20774), .ZN(n13605) );
  NAND2_X1 U16934 ( .A1(n20756), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13622) );
  INV_X1 U16935 ( .A(n9569), .ZN(n13596) );
  NAND2_X1 U16936 ( .A1(n9569), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20627) );
  NAND2_X1 U16937 ( .A1(n20627), .A2(n20632), .ZN(n20193) );
  AOI21_X1 U16938 ( .B1(n13596), .B2(n20578), .A(n20193), .ZN(n13597) );
  AOI21_X1 U16939 ( .B1(n20580), .B2(n13622), .A(n13597), .ZN(n13599) );
  NAND2_X1 U16940 ( .A1(n13605), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13598) );
  OAI21_X1 U16941 ( .B1(n13605), .B2(n13599), .A(n13598), .ZN(P1_U3477) );
  INV_X1 U16942 ( .A(n20193), .ZN(n13601) );
  NOR2_X1 U16943 ( .A1(n20627), .A2(n20769), .ZN(n20475) );
  MUX2_X1 U16944 ( .A(n13601), .B(n20475), .S(n20059), .Z(n13602) );
  AOI21_X1 U16945 ( .B1(n13622), .B2(n20063), .A(n13602), .ZN(n13604) );
  NAND2_X1 U16946 ( .A1(n13605), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13603) );
  OAI21_X1 U16947 ( .B1(n13605), .B2(n13604), .A(n13603), .ZN(P1_U3476) );
  OR2_X1 U16948 ( .A1(n13607), .A2(n13608), .ZN(n13609) );
  NAND2_X1 U16949 ( .A1(n13606), .A2(n13609), .ZN(n19884) );
  AOI21_X1 U16950 ( .B1(n13610), .B2(n13618), .A(n12927), .ZN(n19877) );
  INV_X1 U16951 ( .A(n19918), .ZN(n14404) );
  AOI22_X1 U16952 ( .A1(n19877), .A2(n19913), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n14404), .ZN(n13611) );
  OAI21_X1 U16953 ( .B1(n19884), .B2(n14406), .A(n13611), .ZN(P1_U2867) );
  INV_X1 U16954 ( .A(n20100), .ZN(n13612) );
  INV_X1 U16955 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n19936) );
  OAI222_X1 U16956 ( .A1(n14434), .A2(n19884), .B1(n13612), .B2(n14038), .C1(
        n14428), .C2(n19936), .ZN(P1_U2899) );
  AOI21_X1 U16957 ( .B1(n13614), .B2(n13613), .A(n13607), .ZN(n19989) );
  OR2_X1 U16958 ( .A1(n13616), .A2(n13615), .ZN(n13617) );
  NAND2_X1 U16959 ( .A1(n13618), .A2(n13617), .ZN(n20000) );
  OAI22_X1 U16960 ( .A1(n14401), .A2(n20000), .B1(n13756), .B2(n19918), .ZN(
        n13619) );
  AOI21_X1 U16961 ( .B1(n19989), .B2(n19914), .A(n13619), .ZN(n13620) );
  INV_X1 U16962 ( .A(n13620), .ZN(P1_U2868) );
  INV_X1 U16963 ( .A(n19989), .ZN(n13765) );
  INV_X1 U16964 ( .A(n20095), .ZN(n13621) );
  INV_X1 U16965 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19938) );
  OAI222_X1 U16966 ( .A1(n13765), .A2(n14434), .B1(n13621), .B2(n14038), .C1(
        n19938), .C2(n14428), .ZN(P1_U2900) );
  INV_X1 U16967 ( .A(n20357), .ZN(n19899) );
  INV_X1 U16968 ( .A(n13622), .ZN(n20768) );
  INV_X1 U16969 ( .A(n20060), .ZN(n13623) );
  OAI21_X1 U16970 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n20060), .A(n20480), 
        .ZN(n13624) );
  NOR2_X1 U16971 ( .A1(n20272), .A2(n20627), .ZN(n20331) );
  OAI21_X1 U16972 ( .B1(n13624), .B2(n20331), .A(n20618), .ZN(n13628) );
  OR2_X1 U16973 ( .A1(n9569), .A2(n20578), .ZN(n20399) );
  INV_X1 U16974 ( .A(n20399), .ZN(n13626) );
  AND3_X1 U16975 ( .A1(n20624), .A2(n20632), .A3(n13626), .ZN(n20544) );
  INV_X1 U16976 ( .A(n20544), .ZN(n13627) );
  OAI211_X1 U16977 ( .C1(n19899), .C2(n20768), .A(n13628), .B(n13627), .ZN(
        n13629) );
  NAND2_X1 U16978 ( .A1(n20774), .A2(n13629), .ZN(n13630) );
  OAI21_X1 U16979 ( .B1(n20774), .B2(n20507), .A(n13630), .ZN(P1_U3475) );
  OR2_X1 U16980 ( .A1(n13632), .A2(n13631), .ZN(n13633) );
  NAND2_X1 U16981 ( .A1(n13634), .A2(n13633), .ZN(n20011) );
  INV_X1 U16982 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n13635) );
  OAI22_X1 U16983 ( .A1(n14592), .A2(n19895), .B1(n20035), .B2(n13635), .ZN(
        n13637) );
  NOR2_X1 U16984 ( .A1(n19905), .A2(n20067), .ZN(n13636) );
  AOI211_X1 U16985 ( .C1(n15647), .C2(n19908), .A(n13637), .B(n13636), .ZN(
        n13638) );
  OAI21_X1 U16986 ( .B1(n19822), .B2(n20011), .A(n13638), .ZN(P1_U2996) );
  NAND2_X1 U16987 ( .A1(n13640), .A2(n13639), .ZN(n13642) );
  XNOR2_X1 U16988 ( .A(n13642), .B(n13641), .ZN(n13663) );
  OR2_X1 U16989 ( .A1(n9658), .A2(n13643), .ZN(n13645) );
  NAND2_X1 U16990 ( .A1(n13645), .A2(n13644), .ZN(n18961) );
  OAI22_X1 U16991 ( .A1(n18961), .A2(n15348), .B1(n13657), .B2(n18765), .ZN(
        n13651) );
  INV_X1 U16992 ( .A(n13646), .ZN(n13649) );
  MUX2_X1 U16993 ( .A(n13649), .B(n13648), .S(n13647), .Z(n13650) );
  AOI211_X1 U16994 ( .C1(n16014), .C2(n13278), .A(n13651), .B(n13650), .ZN(
        n13656) );
  NAND2_X1 U16995 ( .A1(n13654), .A2(n13653), .ZN(n13660) );
  NAND3_X1 U16996 ( .A1(n13652), .A2(n13660), .A3(n16011), .ZN(n13655) );
  OAI211_X1 U16997 ( .C1(n13663), .C2(n15234), .A(n13656), .B(n13655), .ZN(
        P2_U3043) );
  NOR2_X1 U16998 ( .A1(n18765), .A2(n13657), .ZN(n13659) );
  INV_X1 U16999 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13689) );
  OAI22_X1 U17000 ( .A1(n13689), .A2(n19047), .B1(n15997), .B2(n13687), .ZN(
        n13658) );
  AOI211_X1 U17001 ( .C1(n19042), .C2(n13278), .A(n13659), .B(n13658), .ZN(
        n13662) );
  NAND3_X1 U17002 ( .A1(n13652), .A2(n13660), .A3(n13164), .ZN(n13661) );
  OAI211_X1 U17003 ( .C1(n13663), .C2(n15976), .A(n13662), .B(n13661), .ZN(
        P2_U3011) );
  INV_X1 U17004 ( .A(n20195), .ZN(n20767) );
  NAND2_X1 U17005 ( .A1(n13664), .A2(n19886), .ZN(n13671) );
  NAND2_X1 U17006 ( .A1(n19852), .A2(n15531), .ZN(n19892) );
  NAND2_X1 U17007 ( .A1(n19892), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13669) );
  INV_X1 U17008 ( .A(n20048), .ZN(n13665) );
  NAND2_X1 U17009 ( .A1(n9561), .A2(n13665), .ZN(n13668) );
  NAND2_X1 U17010 ( .A1(n19876), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13667) );
  OAI21_X1 U17011 ( .B1(n19866), .B2(n19907), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13666) );
  AND4_X1 U17012 ( .A1(n13669), .A2(n13668), .A3(n13667), .A4(n13666), .ZN(
        n13670) );
  OAI211_X1 U17013 ( .C1(n19898), .C2(n20767), .A(n13671), .B(n13670), .ZN(
        P1_U2840) );
  XOR2_X1 U17014 ( .A(n13606), .B(n13672), .Z(n19915) );
  INV_X1 U17015 ( .A(n19915), .ZN(n13674) );
  INV_X1 U17016 ( .A(n20105), .ZN(n13673) );
  OAI222_X1 U17017 ( .A1(n14434), .A2(n13674), .B1(n19933), .B2(n14428), .C1(
        n14038), .C2(n13673), .ZN(P1_U2898) );
  NAND2_X1 U17018 ( .A1(n13676), .A2(n13675), .ZN(n13677) );
  AND2_X1 U17019 ( .A1(n9639), .A2(n13677), .ZN(n19851) );
  INV_X1 U17020 ( .A(n19851), .ZN(n13684) );
  INV_X1 U17021 ( .A(n15778), .ZN(n13680) );
  INV_X1 U17022 ( .A(n13678), .ZN(n13679) );
  OAI21_X1 U17023 ( .B1(n15779), .B2(n13680), .A(n13679), .ZN(n13681) );
  AND2_X1 U17024 ( .A1(n13681), .A2(n13878), .ZN(n19857) );
  AOI22_X1 U17025 ( .A1(n19857), .A2(n19913), .B1(P1_EBX_REG_7__SCAN_IN), .B2(
        n14404), .ZN(n13682) );
  OAI21_X1 U17026 ( .B1(n13684), .B2(n14406), .A(n13682), .ZN(P1_U2865) );
  INV_X1 U17027 ( .A(n20113), .ZN(n13683) );
  OAI222_X1 U17028 ( .A1(n14434), .A2(n13684), .B1(n13683), .B2(n14038), .C1(
        n14428), .C2(n12212), .ZN(P1_U2897) );
  NOR2_X1 U17029 ( .A1(n18849), .A2(n13686), .ZN(n13688) );
  XNOR2_X1 U17030 ( .A(n13688), .B(n13687), .ZN(n13698) );
  INV_X1 U17031 ( .A(n18961), .ZN(n19767) );
  INV_X1 U17032 ( .A(n18858), .ZN(n18869) );
  OAI22_X1 U17033 ( .A1(n18864), .A2(n10143), .B1(n18821), .B2(n13689), .ZN(
        n13690) );
  INV_X1 U17034 ( .A(n13690), .ZN(n13692) );
  NAND2_X1 U17035 ( .A1(n18853), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n13691) );
  OAI211_X1 U17036 ( .C1(n13693), .C2(n18871), .A(n13692), .B(n13691), .ZN(
        n13694) );
  AOI21_X1 U17037 ( .B1(n19767), .B2(n18869), .A(n13694), .ZN(n13696) );
  INV_X1 U17038 ( .A(n18856), .ZN(n18874) );
  NAND2_X1 U17039 ( .A1(n13278), .A2(n18874), .ZN(n13695) );
  OAI211_X1 U17040 ( .C1(n19761), .C2(n14199), .A(n13696), .B(n13695), .ZN(
        n13697) );
  AOI21_X1 U17041 ( .B1(n13698), .B2(n19673), .A(n13697), .ZN(n13699) );
  INV_X1 U17042 ( .A(n13699), .ZN(P2_U2852) );
  OAI21_X1 U17043 ( .B1(n13700), .B2(n13702), .A(n13701), .ZN(n18965) );
  NOR2_X1 U17044 ( .A1(n18849), .A2(n13703), .ZN(n13704) );
  XNOR2_X1 U17045 ( .A(n13704), .B(n13868), .ZN(n13705) );
  NAND2_X1 U17046 ( .A1(n13705), .A2(n19673), .ZN(n13713) );
  AOI21_X1 U17047 ( .B1(n13706), .B2(n13722), .A(n9657), .ZN(n14183) );
  INV_X1 U17048 ( .A(n18864), .ZN(n18818) );
  OAI21_X1 U17049 ( .B1(n18821), .B2(n9711), .A(n18765), .ZN(n13707) );
  AOI21_X1 U17050 ( .B1(n18818), .B2(P2_EBX_REG_5__SCAN_IN), .A(n13707), .ZN(
        n13708) );
  OAI21_X1 U17051 ( .B1(n18866), .B2(n13861), .A(n13708), .ZN(n13711) );
  NOR2_X1 U17052 ( .A1(n13709), .A2(n18871), .ZN(n13710) );
  AOI211_X1 U17053 ( .C1(n14183), .C2(n18874), .A(n13711), .B(n13710), .ZN(
        n13712) );
  OAI211_X1 U17054 ( .C1(n18965), .C2(n18858), .A(n13713), .B(n13712), .ZN(
        P2_U2850) );
  XOR2_X1 U17055 ( .A(n13715), .B(n13714), .Z(n19039) );
  INV_X1 U17056 ( .A(n19039), .ZN(n13729) );
  XNOR2_X1 U17057 ( .A(n13716), .B(n13860), .ZN(n13717) );
  XNOR2_X1 U17058 ( .A(n13718), .B(n13717), .ZN(n19043) );
  NAND2_X1 U17059 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19038), .ZN(n13719) );
  OAI221_X1 U17060 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n13858), .C1(
        n13860), .C2(n13862), .A(n13719), .ZN(n13727) );
  OR2_X1 U17061 ( .A1(n13721), .A2(n13720), .ZN(n13723) );
  AND2_X1 U17062 ( .A1(n13723), .A2(n13722), .ZN(n19041) );
  INV_X1 U17063 ( .A(n19041), .ZN(n18918) );
  AOI21_X1 U17064 ( .B1(n13724), .B2(n13644), .A(n13700), .ZN(n18967) );
  INV_X1 U17065 ( .A(n18967), .ZN(n13725) );
  OAI22_X1 U17066 ( .A1(n18918), .A2(n15343), .B1(n15348), .B2(n13725), .ZN(
        n13726) );
  AOI211_X1 U17067 ( .C1(n19043), .C2(n16011), .A(n13727), .B(n13726), .ZN(
        n13728) );
  OAI21_X1 U17068 ( .B1(n13729), .B2(n15234), .A(n13728), .ZN(P2_U3042) );
  NAND2_X1 U17069 ( .A1(n9567), .A2(n13847), .ZN(n13730) );
  XNOR2_X1 U17070 ( .A(n13731), .B(n13730), .ZN(n13732) );
  NAND2_X1 U17071 ( .A1(n13732), .A2(n19673), .ZN(n13742) );
  NAND2_X1 U17072 ( .A1(n13733), .A2(n18869), .ZN(n13739) );
  OAI22_X1 U17073 ( .A1(n18864), .A2(n13735), .B1(n18821), .B2(n13734), .ZN(
        n13736) );
  AOI21_X1 U17074 ( .B1(n18786), .B2(n13737), .A(n13736), .ZN(n13738) );
  OAI211_X1 U17075 ( .C1(n19701), .C2(n18866), .A(n13739), .B(n13738), .ZN(
        n13740) );
  AOI21_X1 U17076 ( .B1(n15388), .B2(n18874), .A(n13740), .ZN(n13741) );
  OAI211_X1 U17077 ( .C1(n14199), .C2(n19770), .A(n13742), .B(n13741), .ZN(
        P2_U2853) );
  XNOR2_X1 U17078 ( .A(n13744), .B(n13743), .ZN(n18957) );
  NAND2_X1 U17079 ( .A1(n9567), .A2(n13745), .ZN(n13746) );
  XNOR2_X1 U17080 ( .A(n13944), .B(n13746), .ZN(n13747) );
  NAND2_X1 U17081 ( .A1(n13747), .A2(n19673), .ZN(n13755) );
  INV_X1 U17082 ( .A(n13748), .ZN(n13753) );
  NAND2_X1 U17083 ( .A1(n18818), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n13749) );
  OAI211_X1 U17084 ( .C1(n18821), .C2(n13942), .A(n13749), .B(n18765), .ZN(
        n13750) );
  AOI21_X1 U17085 ( .B1(n18853), .B2(P2_REIP_REG_6__SCAN_IN), .A(n13750), .ZN(
        n13751) );
  OAI21_X1 U17086 ( .B1(n13952), .B2(n18856), .A(n13751), .ZN(n13752) );
  AOI21_X1 U17087 ( .B1(n18786), .B2(n13753), .A(n13752), .ZN(n13754) );
  OAI211_X1 U17088 ( .C1(n18957), .C2(n18858), .A(n13755), .B(n13754), .ZN(
        P2_U2849) );
  NOR2_X1 U17089 ( .A1(n19897), .A2(n13756), .ZN(n13761) );
  OAI22_X1 U17090 ( .A1(n13757), .A2(n19894), .B1(n19890), .B2(n19994), .ZN(
        n13760) );
  INV_X1 U17091 ( .A(n19818), .ZN(n13758) );
  NAND2_X1 U17092 ( .A1(n15531), .A2(n13758), .ZN(n19878) );
  INV_X1 U17093 ( .A(n19878), .ZN(n19854) );
  OAI22_X1 U17094 ( .A1(n15586), .A2(n20000), .B1(n15792), .B2(n19898), .ZN(
        n13759) );
  NOR4_X1 U17095 ( .A1(n13761), .A2(n13760), .A3(n19854), .A4(n13759), .ZN(
        n13764) );
  NAND3_X1 U17096 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n13762) );
  NOR2_X1 U17097 ( .A1(n19850), .A2(n13762), .ZN(n19911) );
  INV_X1 U17098 ( .A(n19892), .ZN(n13981) );
  AOI21_X1 U17099 ( .B1(P1_REIP_REG_4__SCAN_IN), .B2(n19911), .A(n13981), .ZN(
        n19885) );
  OAI21_X1 U17100 ( .B1(n19911), .B2(P1_REIP_REG_4__SCAN_IN), .A(n19885), .ZN(
        n13763) );
  OAI211_X1 U17101 ( .C1(n13765), .C2(n19904), .A(n13764), .B(n13763), .ZN(
        P1_U2836) );
  NAND2_X1 U17102 ( .A1(n13685), .A2(n13766), .ZN(n13767) );
  XOR2_X1 U17103 ( .A(n15996), .B(n13767), .Z(n13780) );
  AOI21_X1 U17104 ( .B1(n13769), .B2(n15339), .A(n13768), .ZN(n18952) );
  AOI22_X1 U17105 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18879), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n18853), .ZN(n13770) );
  OAI211_X1 U17106 ( .C1(n18864), .C2(n13771), .A(n13770), .B(n18765), .ZN(
        n13772) );
  AOI21_X1 U17107 ( .B1(n18869), .B2(n18952), .A(n13772), .ZN(n13777) );
  NOR2_X1 U17108 ( .A1(n13773), .A2(n13457), .ZN(n13774) );
  OR2_X1 U17109 ( .A1(n13775), .A2(n13774), .ZN(n18917) );
  INV_X1 U17110 ( .A(n18917), .ZN(n16013) );
  NAND2_X1 U17111 ( .A1(n16013), .A2(n18874), .ZN(n13776) );
  OAI211_X1 U17112 ( .C1(n13778), .C2(n18871), .A(n13777), .B(n13776), .ZN(
        n13779) );
  AOI21_X1 U17113 ( .B1(n13780), .B2(n19673), .A(n13779), .ZN(n13781) );
  INV_X1 U17114 ( .A(n13781), .ZN(P2_U2847) );
  NAND2_X1 U17115 ( .A1(n13685), .A2(n13782), .ZN(n13783) );
  XOR2_X1 U17116 ( .A(n15973), .B(n13783), .Z(n13784) );
  NAND2_X1 U17117 ( .A1(n13784), .A2(n19673), .ZN(n13795) );
  OAI21_X1 U17118 ( .B1(n13787), .B2(n13786), .A(n13785), .ZN(n13788) );
  INV_X1 U17119 ( .A(n13788), .ZN(n18907) );
  NOR2_X1 U17120 ( .A1(n18866), .A2(n10365), .ZN(n13793) );
  XNOR2_X1 U17121 ( .A(n13789), .B(n15332), .ZN(n18949) );
  NOR2_X1 U17122 ( .A1(n18864), .A2(n10614), .ZN(n13790) );
  AOI211_X1 U17123 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n18879), .A(
        n19038), .B(n13790), .ZN(n13791) );
  OAI21_X1 U17124 ( .B1(n18949), .B2(n18858), .A(n13791), .ZN(n13792) );
  AOI211_X1 U17125 ( .C1(n18907), .C2(n18874), .A(n13793), .B(n13792), .ZN(
        n13794) );
  OAI211_X1 U17126 ( .C1(n18871), .C2(n13796), .A(n13795), .B(n13794), .ZN(
        P2_U2845) );
  INV_X1 U17127 ( .A(n13797), .ZN(n13813) );
  NAND2_X1 U17128 ( .A1(n9567), .A2(n13814), .ZN(n13798) );
  XOR2_X1 U17129 ( .A(n15946), .B(n13798), .Z(n13799) );
  NAND2_X1 U17130 ( .A1(n13799), .A2(n19673), .ZN(n13812) );
  OAI21_X1 U17131 ( .B1(n13802), .B2(n13800), .A(n13801), .ZN(n18894) );
  INV_X1 U17132 ( .A(n18894), .ZN(n15999) );
  AOI21_X1 U17133 ( .B1(n13805), .B2(n13803), .A(n13804), .ZN(n18938) );
  AOI21_X1 U17134 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n18879), .A(
        n19038), .ZN(n13806) );
  OAI21_X1 U17135 ( .B1(n18864), .B2(n13807), .A(n13806), .ZN(n13808) );
  AOI21_X1 U17136 ( .B1(n18938), .B2(n18869), .A(n13808), .ZN(n13809) );
  OAI21_X1 U17137 ( .B1(n10423), .B2(n18866), .A(n13809), .ZN(n13810) );
  AOI21_X1 U17138 ( .B1(n15999), .B2(n18874), .A(n13810), .ZN(n13811) );
  OAI211_X1 U17139 ( .C1(n13813), .C2(n18871), .A(n13812), .B(n13811), .ZN(
        P2_U2841) );
  NOR2_X1 U17140 ( .A1(n18863), .A2(n18849), .ZN(n18830) );
  OAI211_X1 U17141 ( .C1(n13815), .C2(n13829), .A(n18830), .B(n13814), .ZN(
        n13827) );
  NAND2_X1 U17142 ( .A1(n13817), .A2(n13816), .ZN(n13819) );
  INV_X1 U17143 ( .A(n13800), .ZN(n13818) );
  OR2_X1 U17144 ( .A1(n13821), .A2(n13820), .ZN(n13822) );
  NAND2_X1 U17145 ( .A1(n13822), .A2(n13803), .ZN(n18942) );
  NAND2_X1 U17146 ( .A1(n18853), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n13824) );
  AOI21_X1 U17147 ( .B1(n18818), .B2(P2_EBX_REG_13__SCAN_IN), .A(n19038), .ZN(
        n13823) );
  OAI211_X1 U17148 ( .C1(n18858), .C2(n18942), .A(n13824), .B(n13823), .ZN(
        n13825) );
  AOI21_X1 U17149 ( .B1(n20957), .B2(n18874), .A(n13825), .ZN(n13826) );
  OAI211_X1 U17150 ( .C1(n13828), .C2(n18871), .A(n13827), .B(n13826), .ZN(
        n13831) );
  NAND2_X1 U17151 ( .A1(n18849), .A2(n19673), .ZN(n18835) );
  OAI22_X1 U17152 ( .A1(n15953), .A2(n18821), .B1(n13829), .B2(n18835), .ZN(
        n13830) );
  OR2_X1 U17153 ( .A1(n13831), .A2(n13830), .ZN(P2_U2842) );
  OR2_X1 U17154 ( .A1(n13833), .A2(n13834), .ZN(n13835) );
  NAND2_X1 U17155 ( .A1(n13832), .A2(n13835), .ZN(n15610) );
  INV_X1 U17156 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13839) );
  NAND2_X1 U17157 ( .A1(n13918), .A2(n13836), .ZN(n13837) );
  AND2_X1 U17158 ( .A1(n9609), .A2(n13837), .ZN(n15746) );
  INV_X1 U17159 ( .A(n15746), .ZN(n13838) );
  OAI222_X1 U17160 ( .A1(n15610), .A2(n14406), .B1(n19918), .B2(n13839), .C1(
        n13838), .C2(n14401), .ZN(P1_U2862) );
  INV_X1 U17161 ( .A(DATAI_10_), .ZN(n13840) );
  MUX2_X1 U17162 ( .A(n13840), .B(n16181), .S(n20068), .Z(n19955) );
  INV_X1 U17163 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n13841) );
  OAI222_X1 U17164 ( .A1(n14434), .A2(n15610), .B1(n19955), .B2(n14038), .C1(
        n13841), .C2(n14428), .ZN(P1_U2894) );
  NOR2_X1 U17165 ( .A1(n18866), .A2(n19699), .ZN(n13845) );
  AOI22_X1 U17166 ( .A1(n18818), .A2(P2_EBX_REG_1__SCAN_IN), .B1(n18879), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13842) );
  OAI21_X1 U17167 ( .B1(n18871), .B2(n13843), .A(n13842), .ZN(n13844) );
  AOI211_X1 U17168 ( .C1(n19786), .C2(n18869), .A(n13845), .B(n13844), .ZN(
        n13846) );
  OAI21_X1 U17169 ( .B1(n11070), .B2(n18856), .A(n13846), .ZN(n13850) );
  OAI211_X1 U17170 ( .C1(n15354), .C2(n13848), .A(n13685), .B(n13847), .ZN(
        n15365) );
  OAI22_X1 U17171 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18835), .B1(
        n15365), .B2(n18863), .ZN(n13849) );
  AOI211_X1 U17172 ( .C1(n18876), .C2(n19782), .A(n13850), .B(n13849), .ZN(
        n13851) );
  INV_X1 U17173 ( .A(n13851), .ZN(P2_U2854) );
  XNOR2_X1 U17174 ( .A(n13852), .B(n13853), .ZN(n13874) );
  NAND2_X1 U17175 ( .A1(n13855), .A2(n13854), .ZN(n13856) );
  XNOR2_X1 U17176 ( .A(n13857), .B(n13856), .ZN(n13871) );
  AOI211_X1 U17177 ( .C1(n11453), .C2(n13860), .A(n13859), .B(n13858), .ZN(
        n13866) );
  NOR2_X1 U17178 ( .A1(n18765), .A2(n13861), .ZN(n13870) );
  NOR2_X1 U17179 ( .A1(n13862), .A2(n11453), .ZN(n13863) );
  AOI211_X1 U17180 ( .C1(n16014), .C2(n14183), .A(n13870), .B(n13863), .ZN(
        n13864) );
  OAI21_X1 U17181 ( .B1(n18965), .B2(n15348), .A(n13864), .ZN(n13865) );
  AOI211_X1 U17182 ( .C1(n13871), .C2(n16011), .A(n13866), .B(n13865), .ZN(
        n13867) );
  OAI21_X1 U17183 ( .B1(n13874), .B2(n15234), .A(n13867), .ZN(P2_U3041) );
  OAI22_X1 U17184 ( .A1(n19047), .A2(n9711), .B1(n15997), .B2(n13868), .ZN(
        n13869) );
  AOI211_X1 U17185 ( .C1(n19042), .C2(n14183), .A(n13870), .B(n13869), .ZN(
        n13873) );
  NAND2_X1 U17186 ( .A1(n13871), .A2(n13164), .ZN(n13872) );
  OAI211_X1 U17187 ( .C1(n13874), .C2(n15976), .A(n13873), .B(n13872), .ZN(
        P2_U3009) );
  INV_X1 U17188 ( .A(n13906), .ZN(n13875) );
  AOI21_X1 U17189 ( .B1(n13876), .B2(n9639), .A(n13875), .ZN(n13916) );
  NAND2_X1 U17190 ( .A1(n13916), .A2(n19914), .ZN(n13881) );
  AND2_X1 U17191 ( .A1(n13878), .A2(n13877), .ZN(n13879) );
  NOR2_X1 U17192 ( .A1(n13920), .A2(n13879), .ZN(n15768) );
  NAND2_X1 U17193 ( .A1(n15768), .A2(n19913), .ZN(n13880) );
  OAI211_X1 U17194 ( .C1(n13882), .C2(n19918), .A(n13881), .B(n13880), .ZN(
        P1_U2864) );
  INV_X1 U17195 ( .A(n13916), .ZN(n13904) );
  INV_X1 U17196 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20710) );
  INV_X1 U17197 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n13883) );
  NAND4_X1 U17198 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n19875)
         );
  NOR2_X1 U17199 ( .A1(n13883), .A2(n19875), .ZN(n19863) );
  NAND2_X1 U17200 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n19863), .ZN(n19864) );
  NOR2_X1 U17201 ( .A1(n20710), .A2(n19864), .ZN(n13888) );
  NAND2_X1 U17202 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n13888), .ZN(n14030) );
  INV_X1 U17203 ( .A(n14030), .ZN(n13886) );
  OR2_X1 U17204 ( .A1(n19852), .A2(n13886), .ZN(n13884) );
  NAND2_X1 U17205 ( .A1(n13884), .A2(n15531), .ZN(n19844) );
  NAND2_X1 U17206 ( .A1(n19876), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n13891) );
  INV_X1 U17207 ( .A(n13914), .ZN(n13885) );
  AOI22_X1 U17208 ( .A1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19866), .B1(
        n19907), .B2(n13885), .ZN(n13890) );
  NOR2_X1 U17209 ( .A1(n13886), .A2(n19852), .ZN(n13887) );
  NAND2_X1 U17210 ( .A1(n13888), .A2(n13887), .ZN(n13889) );
  NAND4_X1 U17211 ( .A1(n13891), .A2(n13890), .A3(n19878), .A4(n13889), .ZN(
        n13892) );
  AOI21_X1 U17212 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(n19844), .A(n13892), .ZN(
        n13894) );
  NAND2_X1 U17213 ( .A1(n15768), .A2(n9561), .ZN(n13893) );
  OAI211_X1 U17214 ( .C1(n13904), .C2(n15609), .A(n13894), .B(n13893), .ZN(
        P1_U2832) );
  OAI21_X1 U17215 ( .B1(n13895), .B2(n13896), .A(n15892), .ZN(n13966) );
  NAND2_X1 U17216 ( .A1(n20964), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13900) );
  OR2_X1 U17217 ( .A1(n13925), .A2(n13897), .ZN(n13898) );
  AND2_X1 U17218 ( .A1(n15057), .A2(n13898), .ZN(n18779) );
  NAND2_X1 U17219 ( .A1(n18779), .A2(n20956), .ZN(n13899) );
  OAI211_X1 U17220 ( .C1(n13966), .C2(n18919), .A(n13900), .B(n13899), .ZN(
        P2_U2870) );
  INV_X1 U17221 ( .A(DATAI_8_), .ZN(n13902) );
  INV_X1 U17222 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n13901) );
  MUX2_X1 U17223 ( .A(n13902), .B(n13901), .S(n20068), .Z(n19949) );
  INV_X1 U17224 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n13903) );
  OAI222_X1 U17225 ( .A1(n13904), .A2(n14434), .B1(n19949), .B2(n14038), .C1(
        n13903), .C2(n14428), .ZN(P1_U2896) );
  AND2_X1 U17226 ( .A1(n13906), .A2(n13905), .ZN(n13907) );
  OR2_X1 U17227 ( .A1(n13907), .A2(n13833), .ZN(n19843) );
  INV_X1 U17228 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n13909) );
  NAND2_X1 U17229 ( .A1(n20068), .A2(n13221), .ZN(n13908) );
  OAI21_X1 U17230 ( .B1(n20068), .B2(DATAI_9_), .A(n13908), .ZN(n19952) );
  OAI222_X1 U17231 ( .A1(n19843), .A2(n14434), .B1(n13909), .B2(n14428), .C1(
        n19952), .C2(n14038), .ZN(P1_U2895) );
  XNOR2_X1 U17232 ( .A(n13911), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13912) );
  XNOR2_X1 U17233 ( .A(n13910), .B(n13912), .ZN(n15766) );
  AOI22_X1 U17234 ( .A1(n19984), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n20053), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13913) );
  OAI21_X1 U17235 ( .B1(n19995), .B2(n13914), .A(n13913), .ZN(n13915) );
  AOI21_X1 U17236 ( .B1(n13916), .B2(n13319), .A(n13915), .ZN(n13917) );
  OAI21_X1 U17237 ( .B1(n15766), .B2(n19822), .A(n13917), .ZN(P1_U2991) );
  OAI21_X1 U17238 ( .B1(n13920), .B2(n13919), .A(n13918), .ZN(n15753) );
  INV_X1 U17239 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n13921) );
  OAI222_X1 U17240 ( .A1(n15753), .A2(n14401), .B1(n13921), .B2(n19918), .C1(
        n19843), .C2(n14406), .ZN(P1_U2863) );
  NAND2_X1 U17241 ( .A1(n13685), .A2(n13922), .ZN(n13923) );
  XOR2_X1 U17242 ( .A(n15925), .B(n13923), .Z(n13924) );
  NAND2_X1 U17243 ( .A1(n13924), .A2(n19673), .ZN(n13937) );
  AOI21_X1 U17244 ( .B1(n13926), .B2(n14083), .A(n13925), .ZN(n15919) );
  INV_X1 U17245 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19719) );
  NOR2_X1 U17246 ( .A1(n18866), .A2(n19719), .ZN(n13935) );
  NAND2_X1 U17247 ( .A1(n13928), .A2(n13927), .ZN(n13931) );
  INV_X1 U17248 ( .A(n13929), .ZN(n13930) );
  NAND2_X1 U17249 ( .A1(n13931), .A2(n13930), .ZN(n18929) );
  NOR2_X1 U17250 ( .A1(n18864), .A2(n18886), .ZN(n13932) );
  AOI211_X1 U17251 ( .C1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n18879), .A(
        n19038), .B(n13932), .ZN(n13933) );
  OAI21_X1 U17252 ( .B1(n18929), .B2(n18858), .A(n13933), .ZN(n13934) );
  AOI211_X1 U17253 ( .C1(n15919), .C2(n18874), .A(n13935), .B(n13934), .ZN(
        n13936) );
  OAI211_X1 U17254 ( .C1(n18871), .C2(n13938), .A(n13937), .B(n13936), .ZN(
        P2_U2839) );
  XNOR2_X1 U17255 ( .A(n13939), .B(n13940), .ZN(n13957) );
  XNOR2_X1 U17256 ( .A(n13941), .B(n13949), .ZN(n13955) );
  OAI22_X1 U17257 ( .A1(n19047), .A2(n13942), .B1(n19707), .B2(n18765), .ZN(
        n13943) );
  AOI21_X1 U17258 ( .B1(n19037), .B2(n13944), .A(n13943), .ZN(n13945) );
  OAI21_X1 U17259 ( .B1(n15406), .B2(n13952), .A(n13945), .ZN(n13946) );
  AOI21_X1 U17260 ( .B1(n13955), .B2(n13164), .A(n13946), .ZN(n13947) );
  OAI21_X1 U17261 ( .B1(n15976), .B2(n13957), .A(n13947), .ZN(P2_U3008) );
  NOR2_X1 U17262 ( .A1(n19707), .A2(n18765), .ZN(n13948) );
  AOI221_X1 U17263 ( .B1(n13950), .B2(n13949), .C1(n15345), .C2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(n13948), .ZN(n13951) );
  INV_X1 U17264 ( .A(n13951), .ZN(n13954) );
  OAI22_X1 U17265 ( .A1(n18957), .A2(n15348), .B1(n15343), .B2(n13952), .ZN(
        n13953) );
  AOI211_X1 U17266 ( .C1(n13955), .C2(n16011), .A(n13954), .B(n13953), .ZN(
        n13956) );
  OAI21_X1 U17267 ( .B1(n15234), .B2(n13957), .A(n13956), .ZN(P2_U3040) );
  OR2_X1 U17268 ( .A1(n13959), .A2(n13929), .ZN(n13960) );
  NAND2_X1 U17269 ( .A1(n13958), .A2(n13960), .ZN(n18792) );
  OAI22_X1 U17270 ( .A1(n18935), .A2(n18792), .B1(n18956), .B2(n13961), .ZN(
        n13964) );
  INV_X1 U17271 ( .A(n18927), .ZN(n14910) );
  INV_X1 U17272 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n13962) );
  OAI22_X1 U17273 ( .A1(n14910), .A2(n13962), .B1(n19056), .B2(n14908), .ZN(
        n13963) );
  AOI211_X1 U17274 ( .C1(n18928), .C2(BUF1_REG_17__SCAN_IN), .A(n13964), .B(
        n13963), .ZN(n13965) );
  OAI21_X1 U17275 ( .B1(n13966), .B2(n18986), .A(n13965), .ZN(P2_U2902) );
  NAND2_X1 U17276 ( .A1(n13832), .A2(n13967), .ZN(n13968) );
  NAND2_X1 U17277 ( .A1(n13969), .A2(n13968), .ZN(n14007) );
  OAI21_X1 U17278 ( .B1(n14007), .B2(n14008), .A(n13969), .ZN(n13976) );
  INV_X1 U17279 ( .A(n13970), .ZN(n14002) );
  INV_X1 U17280 ( .A(n14019), .ZN(n13972) );
  AOI21_X1 U17281 ( .B1(n13973), .B2(n14015), .A(n13972), .ZN(n15730) );
  AOI22_X1 U17282 ( .A1(n15730), .A2(n19913), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14404), .ZN(n13974) );
  OAI21_X1 U17283 ( .B1(n14586), .B2(n14406), .A(n13974), .ZN(P1_U2859) );
  NOR2_X1 U17284 ( .A1(n13976), .A2(n13975), .ZN(n13977) );
  OAI222_X1 U17285 ( .A1(n15593), .A2(n14434), .B1(n14412), .B2(n14038), .C1(
        n13979), .C2(n14428), .ZN(P1_U2892) );
  INV_X1 U17286 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20718) );
  INV_X1 U17287 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n15600) );
  NOR2_X1 U17288 ( .A1(n20718), .A2(n15600), .ZN(n13982) );
  INV_X1 U17289 ( .A(n19852), .ZN(n19882) );
  NAND2_X1 U17290 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n13980) );
  AOI21_X1 U17291 ( .B1(n19882), .B2(n13980), .A(n19844), .ZN(n15615) );
  OAI21_X1 U17292 ( .B1(n13982), .B2(n13981), .A(n15615), .ZN(n15590) );
  INV_X2 U17293 ( .A(n19897), .ZN(n19876) );
  AOI22_X1 U17294 ( .A1(n15730), .A2(n9561), .B1(n19876), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n13983) );
  OAI211_X1 U17295 ( .C1(n19894), .C2(n20874), .A(n13983), .B(n19878), .ZN(
        n13984) );
  AOI21_X1 U17296 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n15590), .A(n13984), 
        .ZN(n13987) );
  INV_X1 U17297 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n15614) );
  INV_X1 U17298 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20713) );
  NOR4_X1 U17299 ( .A1(n15614), .A2(n20713), .A3(n20718), .A4(n15600), .ZN(
        n14028) );
  NOR2_X1 U17300 ( .A1(n19852), .A2(n14030), .ZN(n19840) );
  AND2_X1 U17301 ( .A1(n14028), .A2(n19840), .ZN(n15576) );
  INV_X1 U17302 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20717) );
  INV_X1 U17303 ( .A(n13985), .ZN(n14583) );
  AOI22_X1 U17304 ( .A1(n15576), .A2(n20717), .B1(n14583), .B2(n19907), .ZN(
        n13986) );
  OAI211_X1 U17305 ( .C1(n14586), .C2(n15609), .A(n13987), .B(n13986), .ZN(
        P1_U2827) );
  OAI21_X1 U17306 ( .B1(n9901), .B2(n13990), .A(n13989), .ZN(n13991) );
  OAI21_X1 U17307 ( .B1(n14589), .B2(n9901), .A(n13991), .ZN(n15755) );
  AOI22_X1 U17308 ( .A1(n19984), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n20053), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n13993) );
  NAND2_X1 U17309 ( .A1(n15647), .A2(n19842), .ZN(n13992) );
  OAI211_X1 U17310 ( .C1(n19843), .C2(n20067), .A(n13993), .B(n13992), .ZN(
        n13994) );
  AOI21_X1 U17311 ( .B1(n15755), .B2(n19990), .A(n13994), .ZN(n13995) );
  INV_X1 U17312 ( .A(n13995), .ZN(P1_U2990) );
  INV_X1 U17313 ( .A(DATAI_13_), .ZN(n13997) );
  MUX2_X1 U17314 ( .A(n13997), .B(n13996), .S(n20068), .Z(n19961) );
  INV_X1 U17315 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n13998) );
  OAI222_X1 U17316 ( .A1(n14434), .A2(n14586), .B1(n19961), .B2(n14038), .C1(
        n13998), .C2(n14428), .ZN(P1_U2891) );
  INV_X1 U17317 ( .A(n13999), .ZN(n14003) );
  INV_X1 U17318 ( .A(n14023), .ZN(n14001) );
  INV_X1 U17319 ( .A(n15641), .ZN(n14021) );
  INV_X1 U17320 ( .A(DATAI_14_), .ZN(n14005) );
  INV_X1 U17321 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14004) );
  MUX2_X1 U17322 ( .A(n14005), .B(n14004), .S(n20068), .Z(n19964) );
  OAI222_X1 U17323 ( .A1(n14021), .A2(n14434), .B1(n19964), .B2(n14038), .C1(
        n14006), .C2(n14428), .ZN(P1_U2890) );
  XOR2_X1 U17324 ( .A(n14008), .B(n14007), .Z(n15656) );
  INV_X1 U17325 ( .A(n15656), .ZN(n14012) );
  INV_X1 U17326 ( .A(DATAI_11_), .ZN(n14010) );
  MUX2_X1 U17327 ( .A(n14010), .B(n14009), .S(n20068), .Z(n19958) );
  INV_X1 U17328 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14011) );
  OAI222_X1 U17329 ( .A1(n14012), .A2(n14434), .B1(n19958), .B2(n14038), .C1(
        n14011), .C2(n14428), .ZN(P1_U2893) );
  INV_X1 U17330 ( .A(n15593), .ZN(n15645) );
  OR2_X1 U17331 ( .A1(n15594), .A2(n14013), .ZN(n14014) );
  NAND2_X1 U17332 ( .A1(n14015), .A2(n14014), .ZN(n15587) );
  OAI22_X1 U17333 ( .A1(n15587), .A2(n14401), .B1(n15585), .B2(n19918), .ZN(
        n14016) );
  AOI21_X1 U17334 ( .B1(n15645), .B2(n19914), .A(n14016), .ZN(n14017) );
  INV_X1 U17335 ( .A(n14017), .ZN(P1_U2860) );
  NAND2_X1 U17336 ( .A1(n14019), .A2(n14018), .ZN(n14020) );
  NAND2_X1 U17337 ( .A1(n14025), .A2(n14020), .ZN(n15578) );
  INV_X1 U17338 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n20937) );
  OAI222_X1 U17339 ( .A1(n15578), .A2(n14401), .B1(n19918), .B2(n20937), .C1(
        n14021), .C2(n14406), .ZN(P1_U2858) );
  AOI21_X1 U17340 ( .B1(n14024), .B2(n14023), .A(n14022), .ZN(n14575) );
  INV_X1 U17341 ( .A(n14575), .ZN(n14040) );
  AOI21_X1 U17342 ( .B1(n14026), .B2(n14025), .A(n14352), .ZN(n15719) );
  AOI22_X1 U17343 ( .A1(n15719), .A2(n19913), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n14404), .ZN(n14027) );
  OAI21_X1 U17344 ( .B1(n14040), .B2(n14406), .A(n14027), .ZN(P1_U2857) );
  NAND3_X1 U17345 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(n14028), .ZN(n14029) );
  INV_X1 U17346 ( .A(n19840), .ZN(n15602) );
  NOR2_X1 U17347 ( .A1(n14029), .A2(n15602), .ZN(n15568) );
  INV_X1 U17348 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n15566) );
  NOR2_X1 U17349 ( .A1(n14030), .A2(n14029), .ZN(n14231) );
  OAI21_X1 U17350 ( .B1(n14231), .B2(n19852), .A(n15531), .ZN(n15575) );
  INV_X1 U17351 ( .A(n14573), .ZN(n14031) );
  AOI22_X1 U17352 ( .A1(n19876), .A2(P1_EBX_REG_15__SCAN_IN), .B1(n19907), 
        .B2(n14031), .ZN(n14032) );
  OAI211_X1 U17353 ( .C1(n19894), .C2(n14033), .A(n14032), .B(n19878), .ZN(
        n14034) );
  AOI221_X1 U17354 ( .B1(n15568), .B2(n15566), .C1(n15575), .C2(
        P1_REIP_REG_15__SCAN_IN), .A(n14034), .ZN(n14036) );
  NAND2_X1 U17355 ( .A1(n15719), .A2(n9561), .ZN(n14035) );
  OAI211_X1 U17356 ( .C1(n14040), .C2(n15609), .A(n14036), .B(n14035), .ZN(
        P1_U2825) );
  OAI222_X1 U17357 ( .A1(n14040), .A2(n14434), .B1(n14428), .B2(n14039), .C1(
        n14038), .C2(n14037), .ZN(P1_U2889) );
  NAND2_X1 U17358 ( .A1(n14041), .A2(n14566), .ZN(n14554) );
  INV_X1 U17359 ( .A(n14042), .ZN(n14043) );
  AOI21_X1 U17360 ( .B1(n14554), .B2(n14044), .A(n14043), .ZN(n14046) );
  XNOR2_X1 U17361 ( .A(n15651), .B(n15718), .ZN(n14045) );
  XNOR2_X1 U17362 ( .A(n14046), .B(n14045), .ZN(n15644) );
  INV_X1 U17363 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n14047) );
  INV_X1 U17364 ( .A(n20042), .ZN(n20049) );
  OAI22_X1 U17365 ( .A1(n20035), .A2(n14047), .B1(n20049), .B2(n15578), .ZN(
        n14048) );
  AOI221_X1 U17366 ( .B1(n15702), .B2(n15718), .C1(n15731), .C2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A(n14048), .ZN(n14049) );
  OAI21_X1 U17367 ( .B1(n15644), .B2(n20050), .A(n14049), .ZN(P1_U3017) );
  AOI21_X1 U17368 ( .B1(n14052), .B2(n14051), .A(n14050), .ZN(n15636) );
  INV_X1 U17369 ( .A(n15636), .ZN(n14058) );
  XNOR2_X1 U17370 ( .A(n14352), .B(n14350), .ZN(n15711) );
  AOI22_X1 U17371 ( .A1(n15711), .A2(n19913), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n14404), .ZN(n14053) );
  OAI21_X1 U17372 ( .B1(n14058), .B2(n14406), .A(n14053), .ZN(P1_U2856) );
  INV_X1 U17373 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n14055) );
  INV_X1 U17374 ( .A(n14429), .ZN(n14466) );
  AOI22_X1 U17375 ( .A1(n14466), .A2(n20073), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n14465), .ZN(n14054) );
  OAI21_X1 U17376 ( .B1(n14469), .B2(n14055), .A(n14054), .ZN(n14056) );
  AOI21_X1 U17377 ( .B1(n14471), .B2(DATAI_16_), .A(n14056), .ZN(n14057) );
  OAI21_X1 U17378 ( .B1(n14058), .B2(n14434), .A(n14057), .ZN(P1_U2888) );
  INV_X1 U17379 ( .A(n18716), .ZN(n18666) );
  INV_X1 U17380 ( .A(n18499), .ZN(n18512) );
  INV_X1 U17381 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18496) );
  OAI21_X1 U17382 ( .B1(n18512), .B2(n18661), .A(n18496), .ZN(n15435) );
  NAND2_X1 U17383 ( .A1(n18513), .A2(n15435), .ZN(n18495) );
  NOR2_X1 U17384 ( .A1(n18666), .A2(n18495), .ZN(n14067) );
  INV_X1 U17385 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18653) );
  NOR2_X1 U17386 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18653), .ZN(n18039) );
  INV_X1 U17387 ( .A(n18697), .ZN(n18703) );
  NOR2_X1 U17388 ( .A1(n14060), .A2(n18703), .ZN(n14063) );
  NOR2_X1 U17389 ( .A1(n15430), .A2(n16080), .ZN(n14061) );
  AOI21_X1 U17390 ( .B1(n14063), .B2(n14062), .A(n14061), .ZN(n14064) );
  NAND3_X1 U17391 ( .A1(n14065), .A2(n14064), .A3(n15511), .ZN(n18523) );
  INV_X1 U17392 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n16249) );
  NOR2_X1 U17393 ( .A1(n18705), .A2(n18664), .ZN(n18556) );
  NAND2_X1 U17394 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18556), .ZN(n18651) );
  OAI22_X1 U17395 ( .A1(n18533), .A2(n18552), .B1(n16249), .B2(n18651), .ZN(
        n14066) );
  MUX2_X1 U17396 ( .A(n14067), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18684), .Z(P3_U3284) );
  INV_X1 U17397 ( .A(n14068), .ZN(n14616) );
  NAND2_X1 U17398 ( .A1(n14282), .A2(n14069), .ZN(n14070) );
  NAND2_X1 U17399 ( .A1(n14227), .A2(n14070), .ZN(n14366) );
  OAI21_X1 U17400 ( .B1(n14366), .B2(n20049), .A(n14071), .ZN(n14074) );
  XNOR2_X1 U17401 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14072) );
  NOR2_X1 U17402 ( .A1(n14613), .A2(n14072), .ZN(n14073) );
  AOI211_X1 U17403 ( .C1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n14616), .A(
        n14074), .B(n14073), .ZN(n14075) );
  OAI21_X1 U17404 ( .B1(n14076), .B2(n20050), .A(n14075), .ZN(P1_U3003) );
  OAI21_X1 U17405 ( .B1(n14077), .B2(n14079), .A(n14078), .ZN(n14080) );
  NAND3_X1 U17406 ( .A1(n14080), .A2(n18891), .A3(n18884), .ZN(n14085) );
  NAND2_X1 U17407 ( .A1(n13801), .A2(n14081), .ZN(n14082) );
  AND2_X1 U17408 ( .A1(n14083), .A2(n14082), .ZN(n15930) );
  NAND2_X1 U17409 ( .A1(n15930), .A2(n20956), .ZN(n14084) );
  OAI211_X1 U17410 ( .C1(n20956), .C2(n10632), .A(n14085), .B(n14084), .ZN(
        P2_U2872) );
  AOI21_X1 U17411 ( .B1(n19984), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14086), .ZN(n14087) );
  OAI21_X1 U17412 ( .B1(n19995), .B2(n14088), .A(n14087), .ZN(n14089) );
  AOI21_X1 U17413 ( .B1(n14230), .B2(n13319), .A(n14089), .ZN(n14090) );
  OAI21_X1 U17414 ( .B1(n14091), .B2(n19822), .A(n14090), .ZN(P1_U2968) );
  AOI21_X1 U17415 ( .B1(n14095), .B2(n14094), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14140) );
  NAND3_X1 U17416 ( .A1(n14095), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n14094), .ZN(n14138) );
  OAI21_X1 U17417 ( .B1(n14097), .B2(P2_EBX_REG_30__SCAN_IN), .A(n14096), .ZN(
        n14099) );
  NAND2_X1 U17418 ( .A1(n14099), .A2(n14098), .ZN(n15815) );
  NOR2_X1 U17419 ( .A1(n15815), .A2(n14100), .ZN(n14101) );
  XOR2_X1 U17420 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n14101), .Z(
        n14102) );
  XNOR2_X1 U17421 ( .A(n14103), .B(n14102), .ZN(n14163) );
  NAND2_X1 U17422 ( .A1(n14143), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14104) );
  NAND2_X1 U17423 ( .A1(n14107), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14109) );
  NAND2_X1 U17424 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14108) );
  OAI211_X1 U17425 ( .C1(n15881), .C2(n14110), .A(n14109), .B(n14108), .ZN(
        n14111) );
  AOI21_X1 U17426 ( .B1(n10677), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n14111), .ZN(n14112) );
  NAND2_X1 U17427 ( .A1(n10466), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14115) );
  NAND2_X1 U17428 ( .A1(n14113), .A2(P2_EAX_REG_31__SCAN_IN), .ZN(n14114) );
  OAI211_X1 U17429 ( .C1(n14116), .C2(n19748), .A(n14115), .B(n14114), .ZN(
        n14117) );
  NAND2_X1 U17430 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n14119), .ZN(
        n14123) );
  INV_X1 U17431 ( .A(n14123), .ZN(n14145) );
  NAND4_X1 U17432 ( .A1(n15081), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n14124), .A4(n14145), .ZN(n14120) );
  NAND2_X1 U17433 ( .A1(n19038), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14156) );
  NAND2_X1 U17434 ( .A1(n14120), .A2(n14156), .ZN(n14121) );
  INV_X1 U17435 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14122) );
  AOI211_X1 U17436 ( .C1(n14123), .C2(n15206), .A(n14122), .B(n15101), .ZN(
        n14149) );
  OAI21_X1 U17437 ( .B1(n14163), .B2(n15234), .A(n14127), .ZN(P2_U3015) );
  INV_X1 U17438 ( .A(n14128), .ZN(n14132) );
  OAI21_X1 U17439 ( .B1(n15977), .B2(n14130), .A(n14129), .ZN(n14131) );
  AOI21_X1 U17440 ( .B1(n19040), .B2(n14132), .A(n14131), .ZN(n14135) );
  OAI21_X1 U17441 ( .B1(n15984), .B2(n14133), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14134) );
  OAI211_X1 U17442 ( .C1(n15406), .C2(n15355), .A(n14135), .B(n14134), .ZN(
        P2_U3014) );
  NAND2_X1 U17443 ( .A1(n14137), .A2(n14136), .ZN(n14142) );
  INV_X1 U17444 ( .A(n14138), .ZN(n14139) );
  NOR2_X1 U17445 ( .A1(n14140), .A2(n14139), .ZN(n14141) );
  XNOR2_X1 U17446 ( .A(n14142), .B(n14141), .ZN(n14923) );
  XOR2_X1 U17447 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n14143), .Z(
        n14921) );
  INV_X1 U17448 ( .A(n14919), .ZN(n14151) );
  AOI21_X1 U17449 ( .B1(n15081), .B2(n14145), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14148) );
  NOR2_X1 U17450 ( .A1(n18765), .A2(n14146), .ZN(n14917) );
  INV_X1 U17451 ( .A(n14917), .ZN(n14147) );
  OAI21_X1 U17452 ( .B1(n14923), .B2(n15234), .A(n14154), .ZN(P2_U3016) );
  NAND2_X1 U17453 ( .A1(n15984), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14155) );
  OAI211_X1 U17454 ( .C1(n15997), .C2(n14157), .A(n14156), .B(n14155), .ZN(
        n14158) );
  INV_X1 U17455 ( .A(n14158), .ZN(n14159) );
  OAI21_X1 U17456 ( .B1(n15810), .B2(n15406), .A(n14159), .ZN(n14160) );
  OAI21_X1 U17457 ( .B1(n14163), .B2(n15976), .A(n14162), .ZN(P2_U2983) );
  OAI21_X1 U17458 ( .B1(n14166), .B2(n14165), .A(n14164), .ZN(n14180) );
  OR2_X1 U17459 ( .A1(n14169), .A2(n14168), .ZN(n14170) );
  AND2_X1 U17460 ( .A1(n14167), .A2(n14170), .ZN(n15141) );
  INV_X1 U17461 ( .A(n15141), .ZN(n14736) );
  OAI22_X1 U17462 ( .A1(n18935), .A2(n14736), .B1(n18956), .B2(n14171), .ZN(
        n14174) );
  INV_X1 U17463 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n14172) );
  OAI22_X1 U17464 ( .A1(n14910), .A2(n14172), .B1(n19088), .B2(n14908), .ZN(
        n14173) );
  AOI211_X1 U17465 ( .C1(n18928), .C2(BUF1_REG_23__SCAN_IN), .A(n14174), .B(
        n14173), .ZN(n14175) );
  OAI21_X1 U17466 ( .B1(n14180), .B2(n18986), .A(n14175), .ZN(P2_U2896) );
  NAND2_X1 U17467 ( .A1(n14751), .A2(n14176), .ZN(n14177) );
  NAND2_X1 U17468 ( .A1(n14827), .A2(n14177), .ZN(n15144) );
  NOR2_X1 U17469 ( .A1(n15144), .A2(n20964), .ZN(n14178) );
  AOI21_X1 U17470 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n20964), .A(n14178), .ZN(
        n14179) );
  OAI21_X1 U17471 ( .B1(n14180), .B2(n18919), .A(n14179), .ZN(P2_U2864) );
  XOR2_X1 U17472 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n14187), .Z(n14185)
         );
  NOR2_X1 U17473 ( .A1(n20956), .A2(n14181), .ZN(n14182) );
  AOI21_X1 U17474 ( .B1(n14183), .B2(n20956), .A(n14182), .ZN(n14184) );
  OAI21_X1 U17475 ( .B1(n14185), .B2(n18919), .A(n14184), .ZN(P2_U2882) );
  OR2_X1 U17476 ( .A1(n13410), .A2(n18909), .ZN(n14186) );
  NAND2_X1 U17477 ( .A1(n14187), .A2(n14186), .ZN(n18969) );
  AND2_X1 U17478 ( .A1(n13685), .A2(n14188), .ZN(n14190) );
  AOI21_X1 U17479 ( .B1(n19036), .B2(n14190), .A(n18863), .ZN(n14189) );
  OAI21_X1 U17480 ( .B1(n19036), .B2(n14190), .A(n14189), .ZN(n14198) );
  NAND2_X1 U17481 ( .A1(n18818), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n14191) );
  OAI211_X1 U17482 ( .C1(n18821), .C2(n19046), .A(n14191), .B(n18765), .ZN(
        n14192) );
  AOI21_X1 U17483 ( .B1(n18869), .B2(n18967), .A(n14192), .ZN(n14194) );
  NAND2_X1 U17484 ( .A1(n18853), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n14193) );
  OAI211_X1 U17485 ( .C1(n14195), .C2(n18871), .A(n14194), .B(n14193), .ZN(
        n14196) );
  AOI21_X1 U17486 ( .B1(n19041), .B2(n18874), .A(n14196), .ZN(n14197) );
  OAI211_X1 U17487 ( .C1(n18969), .C2(n14199), .A(n14198), .B(n14197), .ZN(
        P2_U2851) );
  OAI21_X1 U17488 ( .B1(n14200), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n18725), 
        .ZN(n14201) );
  OAI21_X1 U17489 ( .B1(n11404), .B2(n18725), .A(n14201), .ZN(P2_U3612) );
  NOR2_X1 U17490 ( .A1(n14919), .A2(n20964), .ZN(n14202) );
  AOI21_X1 U17491 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n20964), .A(n14202), .ZN(
        n14203) );
  OAI21_X1 U17492 ( .B1(n14204), .B2(n18919), .A(n14203), .ZN(P2_U2857) );
  INV_X1 U17493 ( .A(n14205), .ZN(n14208) );
  INV_X1 U17494 ( .A(n14263), .ZN(n14218) );
  INV_X1 U17495 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14210) );
  NAND2_X1 U17496 ( .A1(n20053), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14603) );
  OAI21_X1 U17497 ( .B1(n14592), .B2(n14210), .A(n14603), .ZN(n14211) );
  INV_X1 U17498 ( .A(n14211), .ZN(n14217) );
  NAND2_X2 U17499 ( .A1(n14241), .A2(n14214), .ZN(n14221) );
  NOR2_X1 U17500 ( .A1(n14221), .A2(n20067), .ZN(n14215) );
  INV_X1 U17501 ( .A(n14215), .ZN(n14216) );
  INV_X1 U17502 ( .A(n14219), .ZN(n14220) );
  OAI21_X1 U17503 ( .B1(n14610), .B2(n19822), .A(n14220), .ZN(P1_U2970) );
  INV_X1 U17504 ( .A(n14221), .ZN(n14260) );
  INV_X1 U17505 ( .A(n14469), .ZN(n14431) );
  OAI22_X1 U17506 ( .A1(n14429), .A2(n19961), .B1(n14428), .B2(n13330), .ZN(
        n14222) );
  AOI21_X1 U17507 ( .B1(n14431), .B2(BUF1_REG_29__SCAN_IN), .A(n14222), .ZN(
        n14224) );
  NAND2_X1 U17508 ( .A1(n14471), .A2(DATAI_29_), .ZN(n14223) );
  OAI211_X1 U17509 ( .C1(n14221), .C2(n14434), .A(n14224), .B(n14223), .ZN(
        P1_U2875) );
  INV_X1 U17510 ( .A(n14225), .ZN(n14226) );
  NAND2_X1 U17511 ( .A1(n14227), .A2(n14226), .ZN(n14228) );
  NAND2_X1 U17512 ( .A1(n14244), .A2(n14228), .ZN(n14605) );
  OAI222_X1 U17513 ( .A1(n14406), .A2(n14221), .B1(n14229), .B2(n19918), .C1(
        n14605), .C2(n14401), .ZN(P1_U2843) );
  INV_X1 U17514 ( .A(n14230), .ZN(n14240) );
  INV_X1 U17515 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n15544) );
  AND4_X1 U17516 ( .A1(n14231), .A2(P1_REIP_REG_17__SCAN_IN), .A3(
        P1_REIP_REG_16__SCAN_IN), .A4(P1_REIP_REG_15__SCAN_IN), .ZN(n14339) );
  NAND3_X1 U17517 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .A3(n14339), .ZN(n15545) );
  NOR2_X1 U17518 ( .A1(n15544), .A2(n15545), .ZN(n15537) );
  AND2_X1 U17519 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n15537), .ZN(n15516) );
  NAND3_X1 U17520 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .A3(n15516), .ZN(n14314) );
  NAND2_X1 U17521 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n14232) );
  NOR2_X1 U17522 ( .A1(n14314), .A2(n14232), .ZN(n14294) );
  NAND2_X1 U17523 ( .A1(n14294), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14293) );
  NAND2_X1 U17524 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n14233) );
  OR2_X1 U17525 ( .A1(n14293), .A2(n14233), .ZN(n14235) );
  INV_X1 U17526 ( .A(n14235), .ZN(n14262) );
  NAND4_X1 U17527 ( .A1(n15531), .A2(P1_REIP_REG_30__SCAN_IN), .A3(
        P1_REIP_REG_29__SCAN_IN), .A4(n14262), .ZN(n14234) );
  NAND2_X1 U17528 ( .A1(n19892), .A2(n14234), .ZN(n14253) );
  NOR3_X1 U17529 ( .A1(n19852), .A2(n20743), .A3(n14235), .ZN(n14255) );
  NAND3_X1 U17530 ( .A1(n14255), .A2(P1_REIP_REG_30__SCAN_IN), .A3(n20747), 
        .ZN(n14237) );
  AOI22_X1 U17531 ( .A1(n19876), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19866), .ZN(n14236) );
  OAI211_X1 U17532 ( .C1(n14253), .C2(n20747), .A(n14237), .B(n14236), .ZN(
        n14238) );
  AOI21_X1 U17533 ( .B1(n14360), .B2(n9561), .A(n14238), .ZN(n14239) );
  OAI21_X1 U17534 ( .B1(n14240), .B2(n15609), .A(n14239), .ZN(P1_U2809) );
  XOR2_X1 U17535 ( .A(n14242), .B(n14241), .Z(n14479) );
  NAND2_X1 U17536 ( .A1(n14244), .A2(n14243), .ZN(n14249) );
  INV_X1 U17537 ( .A(n14245), .ZN(n14246) );
  NAND2_X1 U17538 ( .A1(n14247), .A2(n14246), .ZN(n14248) );
  NAND2_X1 U17539 ( .A1(n14249), .A2(n14248), .ZN(n14252) );
  INV_X1 U17540 ( .A(n14250), .ZN(n14251) );
  XNOR2_X1 U17541 ( .A(n14252), .B(n14251), .ZN(n14363) );
  INV_X1 U17542 ( .A(n14363), .ZN(n14599) );
  INV_X1 U17543 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14364) );
  INV_X1 U17544 ( .A(n14253), .ZN(n14254) );
  OAI21_X1 U17545 ( .B1(n14255), .B2(P1_REIP_REG_30__SCAN_IN), .A(n14254), 
        .ZN(n14257) );
  AOI22_X1 U17546 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19866), .B1(
        n19907), .B2(n14475), .ZN(n14256) );
  OAI211_X1 U17547 ( .C1(n19897), .C2(n14364), .A(n14257), .B(n14256), .ZN(
        n14258) );
  AOI21_X1 U17548 ( .B1(n14599), .B2(n9561), .A(n14258), .ZN(n14259) );
  OAI21_X1 U17549 ( .B1(n14410), .B2(n15609), .A(n14259), .ZN(P1_U2810) );
  NAND2_X1 U17550 ( .A1(n14260), .A2(n19870), .ZN(n14269) );
  OR2_X1 U17551 ( .A1(n19852), .A2(n14262), .ZN(n14261) );
  NAND2_X1 U17552 ( .A1(n14261), .A2(n15531), .ZN(n14272) );
  INV_X1 U17553 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20743) );
  NAND2_X1 U17554 ( .A1(n14262), .A2(n20743), .ZN(n14266) );
  NAND2_X1 U17555 ( .A1(n19876), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14265) );
  AOI22_X1 U17556 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19866), .B1(
        n19907), .B2(n14263), .ZN(n14264) );
  OAI211_X1 U17557 ( .C1(n19852), .C2(n14266), .A(n14265), .B(n14264), .ZN(
        n14267) );
  AOI21_X1 U17558 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(n14272), .A(n14267), 
        .ZN(n14268) );
  OAI211_X1 U17559 ( .C1(n15586), .C2(n14605), .A(n14269), .B(n14268), .ZN(
        P1_U2811) );
  NAND2_X1 U17560 ( .A1(n14365), .A2(n19870), .ZN(n14279) );
  OAI22_X1 U17561 ( .A1(n14271), .A2(n19894), .B1(n19890), .B2(n14270), .ZN(
        n14277) );
  INV_X1 U17562 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14275) );
  INV_X1 U17563 ( .A(n14293), .ZN(n14285) );
  NAND3_X1 U17564 ( .A1(n19882), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14285), 
        .ZN(n14274) );
  INV_X1 U17565 ( .A(n14272), .ZN(n14273) );
  AOI21_X1 U17566 ( .B1(n14275), .B2(n14274), .A(n14273), .ZN(n14276) );
  AOI211_X1 U17567 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n19876), .A(n14277), .B(
        n14276), .ZN(n14278) );
  OAI211_X1 U17568 ( .C1(n15586), .C2(n14366), .A(n14279), .B(n14278), .ZN(
        P1_U2812) );
  NAND2_X1 U17569 ( .A1(n14300), .A2(n14280), .ZN(n14281) );
  NAND2_X1 U17570 ( .A1(n14282), .A2(n14281), .ZN(n14612) );
  AOI21_X1 U17571 ( .B1(n14284), .B2(n14291), .A(n12853), .ZN(n14489) );
  NAND2_X1 U17572 ( .A1(n14489), .A2(n19870), .ZN(n14290) );
  OAI21_X1 U17573 ( .B1(n19852), .B2(n14285), .A(n15531), .ZN(n14303) );
  NOR3_X1 U17574 ( .A1(n19852), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14293), 
        .ZN(n14288) );
  INV_X1 U17575 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14368) );
  AOI22_X1 U17576 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19866), .B1(
        n19907), .B2(n14485), .ZN(n14286) );
  OAI21_X1 U17577 ( .B1(n19897), .B2(n14368), .A(n14286), .ZN(n14287) );
  AOI211_X1 U17578 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n14303), .A(n14288), 
        .B(n14287), .ZN(n14289) );
  OAI211_X1 U17579 ( .C1(n15586), .C2(n14612), .A(n14290), .B(n14289), .ZN(
        P1_U2813) );
  OAI21_X1 U17580 ( .B1(n14309), .B2(n14292), .A(n14291), .ZN(n14499) );
  INV_X1 U17581 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14369) );
  NAND3_X1 U17582 ( .A1(n19882), .A2(n14294), .A3(n14293), .ZN(n14297) );
  INV_X1 U17583 ( .A(n14492), .ZN(n14295) );
  AOI22_X1 U17584 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19866), .B1(
        n19907), .B2(n14295), .ZN(n14296) );
  OAI211_X1 U17585 ( .C1(n19897), .C2(n14369), .A(n14297), .B(n14296), .ZN(
        n14302) );
  OR2_X1 U17586 ( .A1(n14307), .A2(n14298), .ZN(n14299) );
  NAND2_X1 U17587 ( .A1(n14300), .A2(n14299), .ZN(n14620) );
  NOR2_X1 U17588 ( .A1(n14620), .A2(n15586), .ZN(n14301) );
  AOI211_X1 U17589 ( .C1(P1_REIP_REG_26__SCAN_IN), .C2(n14303), .A(n14302), 
        .B(n14301), .ZN(n14304) );
  OAI21_X1 U17590 ( .B1(n14499), .B2(n15609), .A(n14304), .ZN(P1_U2814) );
  NOR2_X1 U17591 ( .A1(n14323), .A2(n14305), .ZN(n14306) );
  OR2_X1 U17592 ( .A1(n14307), .A2(n14306), .ZN(n14631) );
  INV_X1 U17593 ( .A(n14309), .ZN(n14310) );
  OAI21_X1 U17594 ( .B1(n14311), .B2(n14308), .A(n14310), .ZN(n14505) );
  INV_X1 U17595 ( .A(n14505), .ZN(n14312) );
  NAND2_X1 U17596 ( .A1(n14312), .A2(n19870), .ZN(n14321) );
  INV_X1 U17597 ( .A(n14314), .ZN(n14327) );
  NAND2_X1 U17598 ( .A1(n15531), .A2(n14327), .ZN(n14313) );
  AND2_X1 U17599 ( .A1(n19892), .A2(n14313), .ZN(n15517) );
  OAI21_X1 U17600 ( .B1(n14314), .B2(P1_REIP_REG_25__SCAN_IN), .A(
        P1_REIP_REG_24__SCAN_IN), .ZN(n14315) );
  OAI21_X1 U17601 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(P1_REIP_REG_24__SCAN_IN), 
        .A(n14315), .ZN(n14318) );
  NAND2_X1 U17602 ( .A1(n19876), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n14317) );
  AOI22_X1 U17603 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19866), .B1(
        n19907), .B2(n14508), .ZN(n14316) );
  OAI211_X1 U17604 ( .C1(n19852), .C2(n14318), .A(n14317), .B(n14316), .ZN(
        n14319) );
  AOI21_X1 U17605 ( .B1(n15517), .B2(P1_REIP_REG_25__SCAN_IN), .A(n14319), 
        .ZN(n14320) );
  OAI211_X1 U17606 ( .C1(n15586), .C2(n14631), .A(n14321), .B(n14320), .ZN(
        P1_U2815) );
  AND2_X1 U17607 ( .A1(n14380), .A2(n14322), .ZN(n14324) );
  OR2_X1 U17608 ( .A1(n14324), .A2(n14323), .ZN(n14636) );
  INV_X1 U17609 ( .A(n14325), .ZN(n14374) );
  AOI21_X1 U17610 ( .B1(n14326), .B2(n14374), .A(n14308), .ZN(n14517) );
  NAND2_X1 U17611 ( .A1(n14517), .A2(n19870), .ZN(n14334) );
  INV_X1 U17612 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20733) );
  NAND2_X1 U17613 ( .A1(n14327), .A2(n20733), .ZN(n14331) );
  NAND2_X1 U17614 ( .A1(n19876), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n14330) );
  INV_X1 U17615 ( .A(n14515), .ZN(n14328) );
  AOI22_X1 U17616 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19866), .B1(
        n19907), .B2(n14328), .ZN(n14329) );
  OAI211_X1 U17617 ( .C1(n19852), .C2(n14331), .A(n14330), .B(n14329), .ZN(
        n14332) );
  AOI21_X1 U17618 ( .B1(n15517), .B2(P1_REIP_REG_24__SCAN_IN), .A(n14332), 
        .ZN(n14333) );
  OAI211_X1 U17619 ( .C1(n15586), .C2(n14636), .A(n14334), .B(n14333), .ZN(
        P1_U2816) );
  INV_X1 U17620 ( .A(n14441), .ZN(n14395) );
  XNOR2_X1 U17621 ( .A(n14395), .B(n14384), .ZN(n14541) );
  AND2_X1 U17622 ( .A1(n14399), .A2(n14335), .ZN(n14336) );
  NOR2_X1 U17623 ( .A1(n14390), .A2(n14336), .ZN(n15689) );
  AOI22_X1 U17624 ( .A1(P1_EBX_REG_19__SCAN_IN), .A2(n19876), .B1(n19907), 
        .B2(n14544), .ZN(n14337) );
  OAI211_X1 U17625 ( .C1(n19894), .C2(n14540), .A(n14337), .B(n19878), .ZN(
        n14338) );
  INV_X1 U17626 ( .A(n14338), .ZN(n14342) );
  OR2_X1 U17627 ( .A1(n19852), .A2(n14339), .ZN(n14340) );
  NAND2_X1 U17628 ( .A1(n14340), .A2(n15531), .ZN(n15558) );
  NAND4_X1 U17629 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .A4(n15568), .ZN(n14344) );
  NOR2_X1 U17630 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n14344), .ZN(n15559) );
  OAI21_X1 U17631 ( .B1(n15558), .B2(n15559), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n14341) );
  NAND2_X1 U17632 ( .A1(n14342), .A2(n14341), .ZN(n14343) );
  AOI21_X1 U17633 ( .B1(n15689), .B2(n9561), .A(n14343), .ZN(n14346) );
  INV_X1 U17634 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20725) );
  OR3_X1 U17635 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n20725), .A3(n14344), .ZN(
        n14345) );
  OAI211_X1 U17636 ( .C1(n14541), .C2(n15609), .A(n14346), .B(n14345), .ZN(
        P1_U2821) );
  INV_X1 U17637 ( .A(n14347), .ZN(n14348) );
  OAI21_X1 U17638 ( .B1(n14050), .B2(n14349), .A(n14348), .ZN(n14561) );
  INV_X1 U17639 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20723) );
  NOR2_X1 U17640 ( .A1(n20723), .A2(n15566), .ZN(n15565) );
  OAI221_X1 U17641 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n15565), .C1(
        P1_REIP_REG_17__SCAN_IN), .C2(n15568), .A(n15558), .ZN(n14359) );
  INV_X1 U17642 ( .A(n14350), .ZN(n14351) );
  NAND2_X1 U17643 ( .A1(n14352), .A2(n14351), .ZN(n14354) );
  NAND2_X1 U17644 ( .A1(n14354), .A2(n14353), .ZN(n14355) );
  AND2_X1 U17645 ( .A1(n14355), .A2(n14397), .ZN(n15704) );
  AOI22_X1 U17646 ( .A1(P1_EBX_REG_17__SCAN_IN), .A2(n19876), .B1(n19907), 
        .B2(n14564), .ZN(n14356) );
  OAI211_X1 U17647 ( .C1(n19894), .C2(n14560), .A(n14356), .B(n19878), .ZN(
        n14357) );
  AOI21_X1 U17648 ( .B1(n15704), .B2(n9561), .A(n14357), .ZN(n14358) );
  OAI211_X1 U17649 ( .C1(n14561), .C2(n15609), .A(n14359), .B(n14358), .ZN(
        P1_U2823) );
  INV_X1 U17650 ( .A(n14360), .ZN(n14362) );
  INV_X1 U17651 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14361) );
  OAI22_X1 U17652 ( .A1(n14362), .A2(n14401), .B1(n19918), .B2(n14361), .ZN(
        P1_U2841) );
  OAI222_X1 U17653 ( .A1(n14406), .A2(n14410), .B1(n14364), .B2(n19918), .C1(
        n14363), .C2(n14401), .ZN(P1_U2842) );
  INV_X1 U17654 ( .A(n14365), .ZN(n14416) );
  INV_X1 U17655 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14367) );
  OAI222_X1 U17656 ( .A1(n14406), .A2(n14416), .B1(n14367), .B2(n19918), .C1(
        n14366), .C2(n14401), .ZN(P1_U2844) );
  INV_X1 U17657 ( .A(n14489), .ZN(n14420) );
  OAI222_X1 U17658 ( .A1(n14406), .A2(n14420), .B1(n14368), .B2(n19918), .C1(
        n14612), .C2(n14401), .ZN(P1_U2845) );
  OAI222_X1 U17659 ( .A1(n14406), .A2(n14499), .B1(n14369), .B2(n19918), .C1(
        n14620), .C2(n14401), .ZN(P1_U2846) );
  INV_X1 U17660 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14370) );
  OAI222_X1 U17661 ( .A1(n14406), .A2(n14505), .B1(n14370), .B2(n19918), .C1(
        n14631), .C2(n14401), .ZN(P1_U2847) );
  INV_X1 U17662 ( .A(n14517), .ZN(n14435) );
  INV_X1 U17663 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14371) );
  OAI222_X1 U17664 ( .A1(n14406), .A2(n14435), .B1(n19918), .B2(n14371), .C1(
        n14636), .C2(n14401), .ZN(P1_U2848) );
  INV_X1 U17665 ( .A(n14372), .ZN(n14376) );
  INV_X1 U17666 ( .A(n14373), .ZN(n14375) );
  OAI21_X1 U17667 ( .B1(n14376), .B2(n14375), .A(n14374), .ZN(n15520) );
  INV_X1 U17668 ( .A(n15529), .ZN(n14379) );
  INV_X1 U17669 ( .A(n14377), .ZN(n14378) );
  OAI21_X1 U17670 ( .B1(n15530), .B2(n14379), .A(n14378), .ZN(n14381) );
  AND2_X1 U17671 ( .A1(n14381), .A2(n14380), .ZN(n15522) );
  AOI22_X1 U17672 ( .A1(n15522), .A2(n19913), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n14404), .ZN(n14382) );
  OAI21_X1 U17673 ( .B1(n15520), .B2(n14406), .A(n14382), .ZN(P1_U2849) );
  OR2_X1 U17674 ( .A1(n14395), .A2(n14384), .ZN(n14386) );
  NAND2_X1 U17675 ( .A1(n14386), .A2(n14385), .ZN(n14387) );
  NAND2_X1 U17676 ( .A1(n14447), .A2(n14387), .ZN(n15547) );
  INV_X1 U17677 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14391) );
  INV_X1 U17678 ( .A(n14655), .ZN(n14388) );
  OAI21_X1 U17679 ( .B1(n14390), .B2(n14389), .A(n14388), .ZN(n15546) );
  OAI222_X1 U17680 ( .A1(n15547), .A2(n14406), .B1(n19918), .B2(n14391), .C1(
        n15546), .C2(n14401), .ZN(P1_U2852) );
  AOI22_X1 U17681 ( .A1(n15689), .A2(n19913), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n14404), .ZN(n14392) );
  OAI21_X1 U17682 ( .B1(n14541), .B2(n14406), .A(n14392), .ZN(P1_U2853) );
  OR2_X1 U17683 ( .A1(n14347), .A2(n14393), .ZN(n14394) );
  NAND2_X1 U17684 ( .A1(n14395), .A2(n14394), .ZN(n15562) );
  INV_X1 U17685 ( .A(n15562), .ZN(n14551) );
  NAND2_X1 U17686 ( .A1(n14397), .A2(n14396), .ZN(n14398) );
  NAND2_X1 U17687 ( .A1(n14399), .A2(n14398), .ZN(n15695) );
  OAI22_X1 U17688 ( .A1(n15695), .A2(n14401), .B1(n14400), .B2(n19918), .ZN(
        n14402) );
  AOI21_X1 U17689 ( .B1(n14551), .B2(n19914), .A(n14402), .ZN(n14403) );
  INV_X1 U17690 ( .A(n14403), .ZN(P1_U2854) );
  AOI22_X1 U17691 ( .A1(n15704), .A2(n19913), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n14404), .ZN(n14405) );
  OAI21_X1 U17692 ( .B1(n14561), .B2(n14406), .A(n14405), .ZN(P1_U2855) );
  OAI22_X1 U17693 ( .A1(n14429), .A2(n19964), .B1(n14428), .B2(n13544), .ZN(
        n14407) );
  AOI21_X1 U17694 ( .B1(n14431), .B2(BUF1_REG_30__SCAN_IN), .A(n14407), .ZN(
        n14409) );
  NAND2_X1 U17695 ( .A1(n14471), .A2(DATAI_30_), .ZN(n14408) );
  OAI211_X1 U17696 ( .C1(n14410), .C2(n14434), .A(n14409), .B(n14408), .ZN(
        P1_U2874) );
  OAI22_X1 U17697 ( .A1(n14429), .A2(n14412), .B1(n14428), .B2(n14411), .ZN(
        n14414) );
  INV_X1 U17698 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16156) );
  NOR2_X1 U17699 ( .A1(n14469), .A2(n16156), .ZN(n14413) );
  AOI211_X1 U17700 ( .C1(DATAI_28_), .C2(n14471), .A(n14414), .B(n14413), .ZN(
        n14415) );
  OAI21_X1 U17701 ( .B1(n14416), .B2(n14434), .A(n14415), .ZN(P1_U2876) );
  OAI22_X1 U17702 ( .A1(n14429), .A2(n19958), .B1(n14428), .B2(n13341), .ZN(
        n14417) );
  AOI21_X1 U17703 ( .B1(n14431), .B2(BUF1_REG_27__SCAN_IN), .A(n14417), .ZN(
        n14419) );
  NAND2_X1 U17704 ( .A1(n14471), .A2(DATAI_27_), .ZN(n14418) );
  OAI211_X1 U17705 ( .C1(n14420), .C2(n14434), .A(n14419), .B(n14418), .ZN(
        P1_U2877) );
  OAI22_X1 U17706 ( .A1(n14429), .A2(n19955), .B1(n14428), .B2(n13546), .ZN(
        n14421) );
  AOI21_X1 U17707 ( .B1(n14431), .B2(BUF1_REG_26__SCAN_IN), .A(n14421), .ZN(
        n14423) );
  NAND2_X1 U17708 ( .A1(n14471), .A2(DATAI_26_), .ZN(n14422) );
  OAI211_X1 U17709 ( .C1(n14499), .C2(n14434), .A(n14423), .B(n14422), .ZN(
        P1_U2878) );
  OAI22_X1 U17710 ( .A1(n14429), .A2(n19952), .B1(n14428), .B2(n13338), .ZN(
        n14424) );
  AOI21_X1 U17711 ( .B1(n14431), .B2(BUF1_REG_25__SCAN_IN), .A(n14424), .ZN(
        n14426) );
  NAND2_X1 U17712 ( .A1(n14471), .A2(DATAI_25_), .ZN(n14425) );
  OAI211_X1 U17713 ( .C1(n14505), .C2(n14434), .A(n14426), .B(n14425), .ZN(
        P1_U2879) );
  OAI22_X1 U17714 ( .A1(n14429), .A2(n19949), .B1(n14428), .B2(n14427), .ZN(
        n14430) );
  AOI21_X1 U17715 ( .B1(n14431), .B2(BUF1_REG_24__SCAN_IN), .A(n14430), .ZN(
        n14433) );
  NAND2_X1 U17716 ( .A1(n14471), .A2(DATAI_24_), .ZN(n14432) );
  OAI211_X1 U17717 ( .C1(n14435), .C2(n14434), .A(n14433), .B(n14432), .ZN(
        P1_U2880) );
  INV_X1 U17718 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n14437) );
  AOI22_X1 U17719 ( .A1(n14466), .A2(n20113), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n14465), .ZN(n14436) );
  OAI21_X1 U17720 ( .B1(n14469), .B2(n14437), .A(n14436), .ZN(n14438) );
  AOI21_X1 U17721 ( .B1(n14471), .B2(DATAI_23_), .A(n14438), .ZN(n14439) );
  OAI21_X1 U17722 ( .B1(n15520), .B2(n14434), .A(n14439), .ZN(P1_U2881) );
  AND2_X1 U17723 ( .A1(n14441), .A2(n14440), .ZN(n14443) );
  OAI21_X1 U17724 ( .B1(n14443), .B2(n14442), .A(n14372), .ZN(n15528) );
  INV_X1 U17725 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16166) );
  AOI22_X1 U17726 ( .A1(n14466), .A2(n20105), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n14465), .ZN(n14444) );
  OAI21_X1 U17727 ( .B1(n16166), .B2(n14469), .A(n14444), .ZN(n14445) );
  AOI21_X1 U17728 ( .B1(n14471), .B2(DATAI_22_), .A(n14445), .ZN(n14446) );
  OAI21_X1 U17729 ( .B1(n15528), .B2(n14434), .A(n14446), .ZN(P1_U2882) );
  INV_X1 U17730 ( .A(n15619), .ZN(n14452) );
  INV_X1 U17731 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16168) );
  AOI22_X1 U17732 ( .A1(n14466), .A2(n20100), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n14465), .ZN(n14449) );
  OAI21_X1 U17733 ( .B1(n16168), .B2(n14469), .A(n14449), .ZN(n14450) );
  AOI21_X1 U17734 ( .B1(n14471), .B2(DATAI_21_), .A(n14450), .ZN(n14451) );
  OAI21_X1 U17735 ( .B1(n14452), .B2(n14434), .A(n14451), .ZN(P1_U2883) );
  INV_X1 U17736 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n14454) );
  AOI22_X1 U17737 ( .A1(n14466), .A2(n20095), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n14465), .ZN(n14453) );
  OAI21_X1 U17738 ( .B1(n14469), .B2(n14454), .A(n14453), .ZN(n14455) );
  AOI21_X1 U17739 ( .B1(n14471), .B2(DATAI_20_), .A(n14455), .ZN(n14456) );
  OAI21_X1 U17740 ( .B1(n15547), .B2(n14434), .A(n14456), .ZN(P1_U2884) );
  INV_X1 U17741 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n14458) );
  AOI22_X1 U17742 ( .A1(n14466), .A2(n20091), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n14465), .ZN(n14457) );
  OAI21_X1 U17743 ( .B1(n14469), .B2(n14458), .A(n14457), .ZN(n14459) );
  AOI21_X1 U17744 ( .B1(n14471), .B2(DATAI_19_), .A(n14459), .ZN(n14460) );
  OAI21_X1 U17745 ( .B1(n14541), .B2(n14434), .A(n14460), .ZN(P1_U2885) );
  INV_X1 U17746 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n14462) );
  AOI22_X1 U17747 ( .A1(n14466), .A2(n20086), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n14465), .ZN(n14461) );
  OAI21_X1 U17748 ( .B1(n14469), .B2(n14462), .A(n14461), .ZN(n14463) );
  AOI21_X1 U17749 ( .B1(n14471), .B2(DATAI_18_), .A(n14463), .ZN(n14464) );
  OAI21_X1 U17750 ( .B1(n15562), .B2(n14434), .A(n14464), .ZN(P1_U2886) );
  INV_X1 U17751 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n14468) );
  AOI22_X1 U17752 ( .A1(n14466), .A2(n20081), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n14465), .ZN(n14467) );
  OAI21_X1 U17753 ( .B1(n14469), .B2(n14468), .A(n14467), .ZN(n14470) );
  AOI21_X1 U17754 ( .B1(n14471), .B2(DATAI_17_), .A(n14470), .ZN(n14472) );
  OAI21_X1 U17755 ( .B1(n14561), .B2(n14434), .A(n14472), .ZN(P1_U2887) );
  NAND2_X1 U17756 ( .A1(n14473), .A2(n9627), .ZN(n14474) );
  XNOR2_X1 U17757 ( .A(n14474), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14601) );
  INV_X1 U17758 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14477) );
  NAND2_X1 U17759 ( .A1(n15647), .A2(n14475), .ZN(n14476) );
  NAND2_X1 U17760 ( .A1(n20053), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14596) );
  OAI211_X1 U17761 ( .C1(n14477), .C2(n14592), .A(n14476), .B(n14596), .ZN(
        n14478) );
  AOI21_X1 U17762 ( .B1(n14479), .B2(n13319), .A(n14478), .ZN(n14480) );
  OAI21_X1 U17763 ( .B1(n14601), .B2(n19822), .A(n14480), .ZN(P1_U2969) );
  INV_X1 U17764 ( .A(n12868), .ZN(n14481) );
  NAND2_X1 U17765 ( .A1(n14482), .A2(n14481), .ZN(n14483) );
  NAND2_X1 U17766 ( .A1(n15647), .A2(n14485), .ZN(n14486) );
  NAND2_X1 U17767 ( .A1(n20053), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14611) );
  OAI211_X1 U17768 ( .C1(n14592), .C2(n14487), .A(n14486), .B(n14611), .ZN(
        n14488) );
  AOI21_X1 U17769 ( .B1(n14489), .B2(n13319), .A(n14488), .ZN(n14490) );
  OAI21_X1 U17770 ( .B1(n19822), .B2(n14618), .A(n14490), .ZN(P1_U2972) );
  INV_X1 U17771 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n14491) );
  NOR2_X1 U17772 ( .A1(n20035), .A2(n14491), .ZN(n14623) );
  NOR2_X1 U17773 ( .A1(n19995), .A2(n14492), .ZN(n14493) );
  AOI211_X1 U17774 ( .C1(n19984), .C2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n14623), .B(n14493), .ZN(n14498) );
  INV_X1 U17775 ( .A(n14520), .ZN(n14510) );
  OAI21_X1 U17776 ( .B1(n14510), .B2(n14621), .A(n15651), .ZN(n14494) );
  NAND2_X1 U17777 ( .A1(n14495), .A2(n14494), .ZN(n14496) );
  XNOR2_X1 U17778 ( .A(n14496), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14619) );
  NAND2_X1 U17779 ( .A1(n14619), .A2(n19990), .ZN(n14497) );
  OAI211_X1 U17780 ( .C1(n14499), .C2(n20067), .A(n14498), .B(n14497), .ZN(
        P1_U2973) );
  NAND2_X1 U17781 ( .A1(n14500), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14511) );
  MUX2_X1 U17782 ( .A(n14643), .B(n14501), .S(n15631), .Z(n14502) );
  AOI21_X1 U17783 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14511), .A(
        n14502), .ZN(n14503) );
  XNOR2_X1 U17784 ( .A(n14503), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14635) );
  INV_X1 U17785 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14504) );
  NAND2_X1 U17786 ( .A1(n20053), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14630) );
  OAI21_X1 U17787 ( .B1(n14592), .B2(n14504), .A(n14630), .ZN(n14507) );
  NOR2_X1 U17788 ( .A1(n14505), .A2(n20067), .ZN(n14506) );
  AOI211_X1 U17789 ( .C1(n15647), .C2(n14508), .A(n14507), .B(n14506), .ZN(
        n14509) );
  OAI21_X1 U17790 ( .B1(n19822), .B2(n14635), .A(n14509), .ZN(P1_U2974) );
  NAND2_X1 U17791 ( .A1(n14510), .A2(n14511), .ZN(n14512) );
  MUX2_X1 U17792 ( .A(n14512), .B(n14511), .S(n15651), .Z(n14513) );
  XNOR2_X1 U17793 ( .A(n14513), .B(n14643), .ZN(n14646) );
  NOR2_X1 U17794 ( .A1(n20035), .A2(n20733), .ZN(n14641) );
  AOI21_X1 U17795 ( .B1(n19984), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n14641), .ZN(n14514) );
  OAI21_X1 U17796 ( .B1(n19995), .B2(n14515), .A(n14514), .ZN(n14516) );
  AOI21_X1 U17797 ( .B1(n14517), .B2(n13319), .A(n14516), .ZN(n14518) );
  OAI21_X1 U17798 ( .B1(n19822), .B2(n14646), .A(n14518), .ZN(P1_U2975) );
  XNOR2_X1 U17799 ( .A(n15651), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14519) );
  XNOR2_X1 U17800 ( .A(n14520), .B(n14519), .ZN(n14653) );
  NAND2_X1 U17801 ( .A1(n20053), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14648) );
  OAI21_X1 U17802 ( .B1(n14592), .B2(n15525), .A(n14648), .ZN(n14522) );
  NOR2_X1 U17803 ( .A1(n15520), .A2(n20067), .ZN(n14521) );
  AOI211_X1 U17804 ( .C1(n15647), .C2(n15515), .A(n14522), .B(n14521), .ZN(
        n14523) );
  OAI21_X1 U17805 ( .B1(n14653), .B2(n19822), .A(n14523), .ZN(P1_U2976) );
  INV_X1 U17806 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14675) );
  NOR3_X1 U17807 ( .A1(n14547), .A2(n15631), .A3(n14675), .ZN(n14525) );
  AOI21_X1 U17808 ( .B1(n9612), .B2(n15631), .A(n14525), .ZN(n14532) );
  NOR2_X1 U17809 ( .A1(n14532), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14531) );
  AOI22_X1 U17810 ( .A1(n14531), .A2(n15631), .B1(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n14525), .ZN(n14526) );
  XOR2_X1 U17811 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n14526), .Z(
        n14660) );
  NAND2_X1 U17812 ( .A1(n15647), .A2(n15536), .ZN(n14527) );
  NAND2_X1 U17813 ( .A1(n20053), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14656) );
  OAI211_X1 U17814 ( .C1(n14592), .C2(n14528), .A(n14527), .B(n14656), .ZN(
        n14529) );
  AOI21_X1 U17815 ( .B1(n15619), .B2(n13319), .A(n14529), .ZN(n14530) );
  OAI21_X1 U17816 ( .B1(n14660), .B2(n19822), .A(n14530), .ZN(P1_U2978) );
  AOI21_X1 U17817 ( .B1(n14532), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n14531), .ZN(n14678) );
  INV_X1 U17818 ( .A(n15547), .ZN(n14535) );
  NOR2_X1 U17819 ( .A1(n20035), .A2(n15544), .ZN(n14673) );
  AOI21_X1 U17820 ( .B1(n19984), .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n14673), .ZN(n14533) );
  OAI21_X1 U17821 ( .B1(n19995), .B2(n15553), .A(n14533), .ZN(n14534) );
  AOI21_X1 U17822 ( .B1(n14535), .B2(n13319), .A(n14534), .ZN(n14536) );
  OAI21_X1 U17823 ( .B1(n14678), .B2(n19822), .A(n14536), .ZN(P1_U2979) );
  NAND2_X1 U17824 ( .A1(n14547), .A2(n15701), .ZN(n14537) );
  MUX2_X1 U17825 ( .A(n14547), .B(n14537), .S(n15631), .Z(n14538) );
  XOR2_X1 U17826 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n14538), .Z(
        n15688) );
  INV_X1 U17827 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n14539) );
  OAI22_X1 U17828 ( .A1(n14592), .A2(n14540), .B1(n20035), .B2(n14539), .ZN(
        n14543) );
  NOR2_X1 U17829 ( .A1(n14541), .A2(n20067), .ZN(n14542) );
  AOI211_X1 U17830 ( .C1(n15647), .C2(n14544), .A(n14543), .B(n14542), .ZN(
        n14545) );
  OAI21_X1 U17831 ( .B1(n19822), .B2(n15688), .A(n14545), .ZN(P1_U2980) );
  OAI21_X1 U17832 ( .B1(n14546), .B2(n14548), .A(n14547), .ZN(n15696) );
  AOI22_X1 U17833 ( .A1(n19984), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n20053), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14549) );
  OAI21_X1 U17834 ( .B1(n19995), .B2(n15556), .A(n14549), .ZN(n14550) );
  AOI21_X1 U17835 ( .B1(n14551), .B2(n13319), .A(n14550), .ZN(n14552) );
  OAI21_X1 U17836 ( .B1(n19822), .B2(n15696), .A(n14552), .ZN(P1_U2981) );
  INV_X1 U17837 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15725) );
  NOR2_X1 U17838 ( .A1(n15631), .A2(n15725), .ZN(n14557) );
  NOR2_X1 U17839 ( .A1(n15651), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14556) );
  OAI21_X1 U17840 ( .B1(n14554), .B2(n15632), .A(n14553), .ZN(n14555) );
  MUX2_X1 U17841 ( .A(n14557), .B(n14556), .S(n14555), .Z(n14558) );
  XNOR2_X1 U17842 ( .A(n14558), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15703) );
  INV_X1 U17843 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n14559) );
  OAI22_X1 U17844 ( .A1(n14592), .A2(n14560), .B1(n20035), .B2(n14559), .ZN(
        n14563) );
  NOR2_X1 U17845 ( .A1(n14561), .A2(n20067), .ZN(n14562) );
  AOI211_X1 U17846 ( .C1(n15647), .C2(n14564), .A(n14563), .B(n14562), .ZN(
        n14565) );
  OAI21_X1 U17847 ( .B1(n15703), .B2(n19822), .A(n14565), .ZN(P1_U2982) );
  OAI21_X1 U17848 ( .B1(n14041), .B2(n14567), .A(n14566), .ZN(n15633) );
  INV_X1 U17849 ( .A(n14568), .ZN(n14569) );
  NOR2_X1 U17850 ( .A1(n15633), .A2(n14569), .ZN(n14571) );
  XNOR2_X1 U17851 ( .A(n15631), .B(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14570) );
  XNOR2_X1 U17852 ( .A(n14571), .B(n14570), .ZN(n15720) );
  AOI22_X1 U17853 ( .A1(n19984), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20053), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n14572) );
  OAI21_X1 U17854 ( .B1(n19995), .B2(n14573), .A(n14572), .ZN(n14574) );
  AOI21_X1 U17855 ( .B1(n14575), .B2(n13319), .A(n14574), .ZN(n14576) );
  OAI21_X1 U17856 ( .B1(n15720), .B2(n19822), .A(n14576), .ZN(P1_U2984) );
  INV_X1 U17857 ( .A(n14041), .ZN(n15652) );
  INV_X1 U17858 ( .A(n14577), .ZN(n14578) );
  AOI21_X1 U17859 ( .B1(n15652), .B2(n14579), .A(n14578), .ZN(n14679) );
  NAND3_X1 U17860 ( .A1(n14679), .A2(n14680), .A3(n14580), .ZN(n14681) );
  NAND2_X1 U17861 ( .A1(n14681), .A2(n14680), .ZN(n14581) );
  NAND2_X1 U17862 ( .A1(n15732), .A2(n19990), .ZN(n14585) );
  OAI22_X1 U17863 ( .A1(n14592), .A2(n20874), .B1(n20035), .B2(n20717), .ZN(
        n14582) );
  AOI21_X1 U17864 ( .B1(n14583), .B2(n15647), .A(n14582), .ZN(n14584) );
  OAI211_X1 U17865 ( .C1(n20067), .C2(n14586), .A(n14585), .B(n14584), .ZN(
        P1_U2986) );
  NAND2_X1 U17866 ( .A1(n14589), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14588) );
  XNOR2_X1 U17867 ( .A(n14041), .B(n15752), .ZN(n14587) );
  MUX2_X1 U17868 ( .A(n14588), .B(n14587), .S(n15651), .Z(n14591) );
  INV_X1 U17869 ( .A(n14589), .ZN(n14590) );
  NAND3_X1 U17870 ( .A1(n14590), .A2(n15631), .A3(n15752), .ZN(n15653) );
  NAND2_X1 U17871 ( .A1(n14591), .A2(n15653), .ZN(n15747) );
  NAND2_X1 U17872 ( .A1(n15747), .A2(n19990), .ZN(n14595) );
  OAI22_X1 U17873 ( .A1(n14592), .A2(n15606), .B1(n20035), .B2(n15614), .ZN(
        n14593) );
  AOI21_X1 U17874 ( .B1(n15604), .B2(n15647), .A(n14593), .ZN(n14594) );
  OAI211_X1 U17875 ( .C1(n20067), .C2(n15610), .A(n14595), .B(n14594), .ZN(
        P1_U2989) );
  INV_X1 U17876 ( .A(n14596), .ZN(n14598) );
  AOI21_X1 U17877 ( .B1(n14608), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14597) );
  OAI21_X1 U17878 ( .B1(n14601), .B2(n20050), .A(n14600), .ZN(P1_U3001) );
  NAND2_X1 U17879 ( .A1(n14602), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14604) );
  OAI211_X1 U17880 ( .C1(n14605), .C2(n20049), .A(n14604), .B(n14603), .ZN(
        n14606) );
  AOI21_X1 U17881 ( .B1(n14608), .B2(n14607), .A(n14606), .ZN(n14609) );
  OAI21_X1 U17882 ( .B1(n14610), .B2(n20050), .A(n14609), .ZN(P1_U3002) );
  OAI21_X1 U17883 ( .B1(n14612), .B2(n20049), .A(n14611), .ZN(n14615) );
  NOR2_X1 U17884 ( .A1(n14613), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14614) );
  AOI211_X1 U17885 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14616), .A(
        n14615), .B(n14614), .ZN(n14617) );
  OAI21_X1 U17886 ( .B1(n14618), .B2(n20050), .A(n14617), .ZN(P1_U3004) );
  INV_X1 U17887 ( .A(n14619), .ZN(n14629) );
  INV_X1 U17888 ( .A(n14620), .ZN(n14624) );
  INV_X1 U17889 ( .A(n14651), .ZN(n14626) );
  NOR3_X1 U17890 ( .A1(n14626), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14621), .ZN(n14622) );
  AOI211_X1 U17891 ( .C1(n20001), .C2(n14624), .A(n14623), .B(n14622), .ZN(
        n14628) );
  NOR3_X1 U17892 ( .A1(n14626), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n14625), .ZN(n14632) );
  OAI21_X1 U17893 ( .B1(n14632), .B2(n9681), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14627) );
  OAI211_X1 U17894 ( .C1(n14629), .C2(n20050), .A(n14628), .B(n14627), .ZN(
        P1_U3005) );
  OAI21_X1 U17895 ( .B1(n14631), .B2(n20049), .A(n14630), .ZN(n14633) );
  AOI211_X1 U17896 ( .C1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n9681), .A(
        n14633), .B(n14632), .ZN(n14634) );
  OAI21_X1 U17897 ( .B1(n14635), .B2(n20050), .A(n14634), .ZN(P1_U3006) );
  INV_X1 U17898 ( .A(n14636), .ZN(n14642) );
  AOI21_X1 U17899 ( .B1(n12864), .B2(n14638), .A(n14637), .ZN(n14639) );
  NOR2_X1 U17900 ( .A1(n14639), .A2(n14643), .ZN(n14640) );
  AOI211_X1 U17901 ( .C1(n20042), .C2(n14642), .A(n14641), .B(n14640), .ZN(
        n14645) );
  NAND3_X1 U17902 ( .A1(n14651), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n14643), .ZN(n14644) );
  OAI211_X1 U17903 ( .C1(n14646), .C2(n20050), .A(n14645), .B(n14644), .ZN(
        P1_U3007) );
  NAND2_X1 U17904 ( .A1(n15522), .A2(n20042), .ZN(n14647) );
  OAI211_X1 U17905 ( .C1(n14649), .C2(n12864), .A(n14648), .B(n14647), .ZN(
        n14650) );
  AOI21_X1 U17906 ( .B1(n14651), .B2(n12864), .A(n14650), .ZN(n14652) );
  OAI21_X1 U17907 ( .B1(n14653), .B2(n20050), .A(n14652), .ZN(P1_U3008) );
  OAI21_X1 U17908 ( .B1(n14655), .B2(n14654), .A(n15530), .ZN(n15539) );
  NAND2_X1 U17909 ( .A1(n15679), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14657) );
  OAI211_X1 U17910 ( .C1(n20049), .C2(n15539), .A(n14657), .B(n14656), .ZN(
        n14658) );
  AOI21_X1 U17911 ( .B1(n15683), .B2(n12837), .A(n14658), .ZN(n14659) );
  OAI21_X1 U17912 ( .B1(n14660), .B2(n20050), .A(n14659), .ZN(P1_U3010) );
  INV_X1 U17913 ( .A(n15546), .ZN(n14674) );
  INV_X1 U17914 ( .A(n15687), .ZN(n14671) );
  INV_X1 U17915 ( .A(n14661), .ZN(n14666) );
  NOR2_X1 U17916 ( .A1(n14666), .A2(n14662), .ZN(n15728) );
  INV_X1 U17917 ( .A(n15728), .ZN(n14663) );
  NOR2_X1 U17918 ( .A1(n14663), .A2(n20034), .ZN(n14664) );
  NAND2_X1 U17919 ( .A1(n20046), .A2(n14664), .ZN(n14669) );
  NOR2_X1 U17920 ( .A1(n14666), .A2(n14665), .ZN(n14667) );
  NAND2_X1 U17921 ( .A1(n20047), .A2(n14667), .ZN(n14668) );
  NAND2_X1 U17922 ( .A1(n14669), .A2(n14668), .ZN(n15727) );
  OAI21_X1 U17923 ( .B1(n15727), .B2(n15729), .A(n14675), .ZN(n14670) );
  AOI21_X1 U17924 ( .B1(n14671), .B2(n14670), .A(n12836), .ZN(n14672) );
  AOI211_X1 U17925 ( .C1(n20001), .C2(n14674), .A(n14673), .B(n14672), .ZN(
        n14677) );
  OR3_X1 U17926 ( .A1(n15693), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n14675), .ZN(n14676) );
  OAI211_X1 U17927 ( .C1(n14678), .C2(n20050), .A(n14677), .B(n14676), .ZN(
        P1_U3011) );
  INV_X1 U17928 ( .A(n14679), .ZN(n14684) );
  OAI21_X1 U17929 ( .B1(n12941), .B2(n15651), .A(n14680), .ZN(n14683) );
  INV_X1 U17930 ( .A(n14681), .ZN(n14682) );
  AOI21_X1 U17931 ( .B1(n14684), .B2(n14683), .A(n14682), .ZN(n15650) );
  NOR2_X1 U17932 ( .A1(n15784), .A2(n14688), .ZN(n14692) );
  OAI221_X1 U17933 ( .B1(n15762), .B2(n14686), .C1(n15762), .C2(n15743), .A(
        n14685), .ZN(n14687) );
  AOI21_X1 U17934 ( .B1(n20047), .B2(n14688), .A(n14687), .ZN(n15742) );
  OAI21_X1 U17935 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n14689), .A(
        n15742), .ZN(n14691) );
  OAI22_X1 U17936 ( .A1(n20035), .A2(n20718), .B1(n20049), .B2(n15587), .ZN(
        n14690) );
  AOI221_X1 U17937 ( .B1(n14692), .B2(n12941), .C1(n14691), .C2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n14690), .ZN(n14693) );
  OAI21_X1 U17938 ( .B1(n15650), .B2(n20050), .A(n14693), .ZN(P1_U3019) );
  INV_X1 U17939 ( .A(n15796), .ZN(n20766) );
  INV_X1 U17940 ( .A(n14694), .ZN(n20760) );
  AOI22_X1 U17941 ( .A1(n14697), .A2(n14696), .B1(n14695), .B2(n20760), .ZN(
        n14698) );
  OAI21_X1 U17942 ( .B1(n14699), .B2(n20766), .A(n14698), .ZN(n14700) );
  MUX2_X1 U17943 ( .A(n14700), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n20763), .Z(P1_U3472) );
  INV_X1 U17944 ( .A(n14701), .ZN(n14702) );
  OAI22_X1 U17945 ( .A1(n14703), .A2(n20766), .B1(n14702), .B2(n20758), .ZN(
        n14704) );
  MUX2_X1 U17946 ( .A(n14704), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n20763), .Z(P1_U3469) );
  INV_X1 U17947 ( .A(n14705), .ZN(n14709) );
  OAI21_X1 U17948 ( .B1(n19690), .B2(n19665), .A(n16070), .ZN(n14708) );
  OAI211_X1 U17949 ( .C1(n14706), .C2(n19544), .A(n19801), .B(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n14707) );
  OAI211_X1 U17950 ( .C1(n14710), .C2(n14709), .A(n14708), .B(n14707), .ZN(
        n14715) );
  OAI21_X1 U17951 ( .B1(n14711), .B2(n19665), .A(n19611), .ZN(n14712) );
  OAI211_X1 U17952 ( .C1(n19690), .C2(n14713), .A(n18725), .B(n14712), .ZN(
        n14714) );
  MUX2_X1 U17953 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .B(n14715), .S(n14714), 
        .Z(P2_U3610) );
  NOR2_X1 U17954 ( .A1(n14802), .A2(n14716), .ZN(n14717) );
  OR2_X1 U17955 ( .A1(n14718), .A2(n14717), .ZN(n15087) );
  OAI211_X1 U17956 ( .C1(n14720), .C2(n14942), .A(n19673), .B(n14719), .ZN(
        n14731) );
  NAND2_X1 U17957 ( .A1(n14721), .A2(n14722), .ZN(n14723) );
  NAND2_X1 U17958 ( .A1(n14724), .A2(n14723), .ZN(n15082) );
  OAI22_X1 U17959 ( .A1(n18864), .A2(n14725), .B1(n18821), .B2(n10052), .ZN(
        n14726) );
  AOI21_X1 U17960 ( .B1(n18853), .B2(P2_REIP_REG_28__SCAN_IN), .A(n14726), 
        .ZN(n14727) );
  OAI21_X1 U17961 ( .B1(n15082), .B2(n18858), .A(n14727), .ZN(n14728) );
  AOI21_X1 U17962 ( .B1(n14729), .B2(n18786), .A(n14728), .ZN(n14730) );
  OAI211_X1 U17963 ( .C1(n18856), .C2(n15087), .A(n14731), .B(n14730), .ZN(
        P2_U2827) );
  OAI211_X1 U17964 ( .C1(n14734), .C2(n14733), .A(n19673), .B(n14732), .ZN(
        n14740) );
  AOI22_X1 U17965 ( .A1(n18818), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18879), .ZN(n14735) );
  OAI21_X1 U17966 ( .B1(n18858), .B2(n14736), .A(n14735), .ZN(n14738) );
  NOR2_X1 U17967 ( .A1(n15144), .A2(n18856), .ZN(n14737) );
  AOI211_X1 U17968 ( .C1(n18853), .C2(P2_REIP_REG_23__SCAN_IN), .A(n14738), 
        .B(n14737), .ZN(n14739) );
  OAI211_X1 U17969 ( .C1(n14741), .C2(n18871), .A(n14740), .B(n14739), .ZN(
        P2_U2832) );
  INV_X1 U17970 ( .A(n14742), .ZN(n14756) );
  OAI211_X1 U17971 ( .C1(n15915), .C2(n14744), .A(n19673), .B(n14743), .ZN(
        n14755) );
  XNOR2_X1 U17972 ( .A(n14746), .B(n14745), .ZN(n15158) );
  AOI22_X1 U17973 ( .A1(n18818), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n18879), .ZN(n14747) );
  OAI21_X1 U17974 ( .B1(n18858), .B2(n15158), .A(n14747), .ZN(n14753) );
  NAND2_X1 U17975 ( .A1(n14748), .A2(n14749), .ZN(n14750) );
  NAND2_X1 U17976 ( .A1(n14751), .A2(n14750), .ZN(n15908) );
  NOR2_X1 U17977 ( .A1(n15908), .A2(n18856), .ZN(n14752) );
  AOI211_X1 U17978 ( .C1(n18853), .C2(P2_REIP_REG_22__SCAN_IN), .A(n14753), 
        .B(n14752), .ZN(n14754) );
  OAI211_X1 U17979 ( .C1(n14756), .C2(n18871), .A(n14755), .B(n14754), .ZN(
        P2_U2833) );
  XNOR2_X1 U17980 ( .A(n14780), .B(n15019), .ZN(n14768) );
  OR2_X1 U17981 ( .A1(n14757), .A2(n14758), .ZN(n14759) );
  NAND2_X1 U17982 ( .A1(n14748), .A2(n14759), .ZN(n15176) );
  OAI22_X1 U17983 ( .A1(n14760), .A2(n18821), .B1(n19728), .B2(n18866), .ZN(
        n14763) );
  OAI21_X1 U17984 ( .B1(n14775), .B2(n14761), .A(n14745), .ZN(n15170) );
  NOR2_X1 U17985 ( .A1(n15170), .A2(n18858), .ZN(n14762) );
  AOI211_X1 U17986 ( .C1(n18818), .C2(P2_EBX_REG_21__SCAN_IN), .A(n14763), .B(
        n14762), .ZN(n14764) );
  OAI21_X1 U17987 ( .B1(n15176), .B2(n18856), .A(n14764), .ZN(n14765) );
  AOI21_X1 U17988 ( .B1(n14766), .B2(n18786), .A(n14765), .ZN(n14767) );
  OAI21_X1 U17989 ( .B1(n14768), .B2(n18863), .A(n14767), .ZN(P2_U2834) );
  NOR2_X1 U17990 ( .A1(n14839), .A2(n14769), .ZN(n14770) );
  OR2_X1 U17991 ( .A1(n14757), .A2(n14770), .ZN(n15889) );
  INV_X1 U17992 ( .A(n18835), .ZN(n18878) );
  NAND2_X1 U17993 ( .A1(n15035), .A2(n18878), .ZN(n14779) );
  OAI22_X1 U17994 ( .A1(n18864), .A2(n14771), .B1(n18821), .B2(n9707), .ZN(
        n14777) );
  NOR2_X1 U17995 ( .A1(n14772), .A2(n14773), .ZN(n14774) );
  OR2_X1 U17996 ( .A1(n14775), .A2(n14774), .ZN(n15896) );
  NOR2_X1 U17997 ( .A1(n15896), .A2(n18858), .ZN(n14776) );
  AOI211_X1 U17998 ( .C1(n18853), .C2(P2_REIP_REG_20__SCAN_IN), .A(n14777), 
        .B(n14776), .ZN(n14778) );
  OAI211_X1 U17999 ( .C1(n18856), .C2(n15889), .A(n14779), .B(n14778), .ZN(
        n14783) );
  AOI211_X1 U18000 ( .C1(n15035), .C2(n14781), .A(n18863), .B(n14780), .ZN(
        n14782) );
  AOI211_X1 U18001 ( .C1(n18786), .C2(n14784), .A(n14783), .B(n14782), .ZN(
        n14785) );
  INV_X1 U18002 ( .A(n14785), .ZN(P2_U2835) );
  INV_X1 U18003 ( .A(n14786), .ZN(n14844) );
  NAND2_X1 U18004 ( .A1(n14788), .A2(n14787), .ZN(n14843) );
  NAND3_X1 U18005 ( .A1(n14844), .A2(n18891), .A3(n14843), .ZN(n14790) );
  NAND2_X1 U18006 ( .A1(n20964), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14789) );
  OAI211_X1 U18007 ( .C1(n20964), .C2(n15821), .A(n14790), .B(n14789), .ZN(
        P2_U2858) );
  NAND2_X1 U18008 ( .A1(n14792), .A2(n14791), .ZN(n14794) );
  XNOR2_X1 U18009 ( .A(n14794), .B(n14793), .ZN(n14855) );
  NOR2_X1 U18010 ( .A1(n15087), .A2(n20964), .ZN(n14795) );
  AOI21_X1 U18011 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n20964), .A(n14795), .ZN(
        n14796) );
  OAI21_X1 U18012 ( .B1(n14855), .B2(n18919), .A(n14796), .ZN(P2_U2859) );
  AOI21_X1 U18013 ( .B1(n14799), .B2(n14798), .A(n14797), .ZN(n14800) );
  INV_X1 U18014 ( .A(n14800), .ZN(n14864) );
  AND2_X1 U18015 ( .A1(n14811), .A2(n14801), .ZN(n14803) );
  OR2_X1 U18016 ( .A1(n14803), .A2(n14802), .ZN(n15835) );
  NOR2_X1 U18017 ( .A1(n15835), .A2(n20964), .ZN(n14804) );
  AOI21_X1 U18018 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n20964), .A(n14804), .ZN(
        n14805) );
  OAI21_X1 U18019 ( .B1(n14864), .B2(n18919), .A(n14805), .ZN(P2_U2860) );
  AOI21_X1 U18020 ( .B1(n14808), .B2(n14807), .A(n14806), .ZN(n14809) );
  INV_X1 U18021 ( .A(n14809), .ZN(n14871) );
  NAND2_X1 U18022 ( .A1(n20964), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14815) );
  INV_X1 U18023 ( .A(n14811), .ZN(n14812) );
  AOI21_X1 U18024 ( .B1(n14813), .B2(n14810), .A(n14812), .ZN(n15849) );
  NAND2_X1 U18025 ( .A1(n15849), .A2(n20956), .ZN(n14814) );
  OAI211_X1 U18026 ( .C1(n14871), .C2(n18919), .A(n14815), .B(n14814), .ZN(
        P2_U2861) );
  OAI21_X1 U18027 ( .B1(n14818), .B2(n14817), .A(n14816), .ZN(n14879) );
  OR2_X1 U18028 ( .A1(n14825), .A2(n14819), .ZN(n14820) );
  NAND2_X1 U18029 ( .A1(n14810), .A2(n14820), .ZN(n15117) );
  MUX2_X1 U18030 ( .A(n15117), .B(n14821), .S(n20964), .Z(n14822) );
  OAI21_X1 U18031 ( .B1(n14879), .B2(n18919), .A(n14822), .ZN(P2_U2862) );
  OR2_X1 U18032 ( .A1(n14824), .A2(n14823), .ZN(n14880) );
  NAND3_X1 U18033 ( .A1(n11704), .A2(n14880), .A3(n18891), .ZN(n14831) );
  INV_X1 U18034 ( .A(n14825), .ZN(n14829) );
  NAND2_X1 U18035 ( .A1(n14827), .A2(n14826), .ZN(n14828) );
  NAND2_X1 U18036 ( .A1(n14829), .A2(n14828), .ZN(n15872) );
  INV_X1 U18037 ( .A(n15872), .ZN(n14987) );
  NAND2_X1 U18038 ( .A1(n14987), .A2(n20956), .ZN(n14830) );
  OAI211_X1 U18039 ( .C1(n20956), .C2(n10660), .A(n14831), .B(n14830), .ZN(
        P2_U2863) );
  OAI21_X1 U18040 ( .B1(n15886), .B2(n14832), .A(n14891), .ZN(n14904) );
  NOR2_X1 U18041 ( .A1(n15176), .A2(n20964), .ZN(n14833) );
  AOI21_X1 U18042 ( .B1(P2_EBX_REG_21__SCAN_IN), .B2(n20964), .A(n14833), .ZN(
        n14834) );
  OAI21_X1 U18043 ( .B1(n14904), .B2(n18919), .A(n14834), .ZN(P2_U2866) );
  AOI21_X1 U18044 ( .B1(n14836), .B2(n15890), .A(n14835), .ZN(n14837) );
  INV_X1 U18045 ( .A(n14837), .ZN(n14914) );
  AND2_X1 U18046 ( .A1(n15059), .A2(n14838), .ZN(n14840) );
  OR2_X1 U18047 ( .A1(n14840), .A2(n14839), .ZN(n18758) );
  NOR2_X1 U18048 ( .A1(n18758), .A2(n20964), .ZN(n14841) );
  AOI21_X1 U18049 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n20964), .A(n14841), .ZN(
        n14842) );
  OAI21_X1 U18050 ( .B1(n14914), .B2(n18919), .A(n14842), .ZN(P2_U2868) );
  NAND3_X1 U18051 ( .A1(n14844), .A2(n18970), .A3(n14843), .ZN(n14849) );
  AOI22_X1 U18052 ( .A1(n15822), .A2(n18982), .B1(P2_EAX_REG_29__SCAN_IN), 
        .B2(n18981), .ZN(n14848) );
  AOI22_X1 U18053 ( .A1(n18927), .A2(BUF2_REG_29__SCAN_IN), .B1(n18926), .B2(
        n14845), .ZN(n14847) );
  NAND2_X1 U18054 ( .A1(n18928), .A2(BUF1_REG_29__SCAN_IN), .ZN(n14846) );
  NAND4_X1 U18055 ( .A1(n14849), .A2(n14848), .A3(n14847), .A4(n14846), .ZN(
        P2_U2890) );
  OAI22_X1 U18056 ( .A1(n18935), .A2(n15082), .B1(n18956), .B2(n14850), .ZN(
        n14853) );
  INV_X1 U18057 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n14851) );
  OAI22_X1 U18058 ( .A1(n14910), .A2(n14851), .B1(n18943), .B2(n14908), .ZN(
        n14852) );
  AOI211_X1 U18059 ( .C1(n18928), .C2(BUF1_REG_28__SCAN_IN), .A(n14853), .B(
        n14852), .ZN(n14854) );
  OAI21_X1 U18060 ( .B1(n14855), .B2(n18986), .A(n14854), .ZN(P2_U2891) );
  AND2_X1 U18061 ( .A1(n14856), .A2(n14865), .ZN(n14867) );
  OR2_X1 U18062 ( .A1(n14867), .A2(n14857), .ZN(n14858) );
  NAND2_X1 U18063 ( .A1(n14721), .A2(n14858), .ZN(n15834) );
  OAI22_X1 U18064 ( .A1(n18935), .A2(n15834), .B1(n18956), .B2(n14859), .ZN(
        n14862) );
  INV_X1 U18065 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n14860) );
  OAI22_X1 U18066 ( .A1(n14910), .A2(n14860), .B1(n18945), .B2(n14908), .ZN(
        n14861) );
  AOI211_X1 U18067 ( .C1(n18928), .C2(BUF1_REG_27__SCAN_IN), .A(n14862), .B(
        n14861), .ZN(n14863) );
  OAI21_X1 U18068 ( .B1(n14864), .B2(n18986), .A(n14863), .ZN(P2_U2892) );
  NOR2_X1 U18069 ( .A1(n14856), .A2(n14865), .ZN(n14866) );
  OAI22_X1 U18070 ( .A1(n18935), .A2(n15847), .B1(n18956), .B2(n13270), .ZN(
        n14868) );
  AOI21_X1 U18071 ( .B1(n18928), .B2(BUF1_REG_26__SCAN_IN), .A(n14868), .ZN(
        n14870) );
  AOI22_X1 U18072 ( .A1(n18927), .A2(BUF2_REG_26__SCAN_IN), .B1(n18926), .B2(
        n18947), .ZN(n14869) );
  OAI211_X1 U18073 ( .C1(n14871), .C2(n18986), .A(n14870), .B(n14869), .ZN(
        P2_U2893) );
  AND2_X1 U18074 ( .A1(n9629), .A2(n14872), .ZN(n14873) );
  OR2_X1 U18075 ( .A1(n14873), .A2(n14856), .ZN(n15858) );
  OAI22_X1 U18076 ( .A1(n18935), .A2(n15858), .B1(n18956), .B2(n14874), .ZN(
        n14877) );
  INV_X1 U18077 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n14875) );
  OAI22_X1 U18078 ( .A1(n14910), .A2(n14875), .B1(n18950), .B2(n14908), .ZN(
        n14876) );
  AOI211_X1 U18079 ( .C1(n18928), .C2(BUF1_REG_25__SCAN_IN), .A(n14877), .B(
        n14876), .ZN(n14878) );
  OAI21_X1 U18080 ( .B1(n14879), .B2(n18986), .A(n14878), .ZN(P2_U2894) );
  NAND3_X1 U18081 ( .A1(n11704), .A2(n14880), .A3(n18970), .ZN(n14888) );
  NAND2_X1 U18082 ( .A1(n14167), .A2(n14881), .ZN(n14882) );
  NAND2_X1 U18083 ( .A1(n9629), .A2(n14882), .ZN(n15871) );
  OAI22_X1 U18084 ( .A1(n18935), .A2(n15871), .B1(n18956), .B2(n14883), .ZN(
        n14886) );
  INV_X1 U18085 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n14884) );
  OAI22_X1 U18086 ( .A1(n14910), .A2(n14884), .B1(n18953), .B2(n14908), .ZN(
        n14885) );
  AOI211_X1 U18087 ( .C1(n18928), .C2(BUF1_REG_24__SCAN_IN), .A(n14886), .B(
        n14885), .ZN(n14887) );
  NAND2_X1 U18088 ( .A1(n14888), .A2(n14887), .ZN(P2_U2895) );
  INV_X1 U18089 ( .A(n14889), .ZN(n14890) );
  AOI21_X1 U18090 ( .B1(n14892), .B2(n14891), .A(n14890), .ZN(n15882) );
  INV_X1 U18091 ( .A(n15882), .ZN(n14898) );
  OAI22_X1 U18092 ( .A1(n18935), .A2(n15158), .B1(n18956), .B2(n14893), .ZN(
        n14896) );
  INV_X1 U18093 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n14894) );
  OAI22_X1 U18094 ( .A1(n14910), .A2(n14894), .B1(n19077), .B2(n14908), .ZN(
        n14895) );
  AOI211_X1 U18095 ( .C1(n18928), .C2(BUF1_REG_22__SCAN_IN), .A(n14896), .B(
        n14895), .ZN(n14897) );
  OAI21_X1 U18096 ( .B1(n14898), .B2(n18986), .A(n14897), .ZN(P2_U2897) );
  OAI22_X1 U18097 ( .A1(n18935), .A2(n15170), .B1(n18956), .B2(n14899), .ZN(
        n14902) );
  INV_X1 U18098 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n14900) );
  OAI22_X1 U18099 ( .A1(n14910), .A2(n14900), .B1(n19072), .B2(n14908), .ZN(
        n14901) );
  AOI211_X1 U18100 ( .C1(n18928), .C2(BUF1_REG_21__SCAN_IN), .A(n14902), .B(
        n14901), .ZN(n14903) );
  OAI21_X1 U18101 ( .B1(n14904), .B2(n18986), .A(n14903), .ZN(P2_U2898) );
  AND2_X1 U18102 ( .A1(n15211), .A2(n14905), .ZN(n14906) );
  NOR2_X1 U18103 ( .A1(n14772), .A2(n14906), .ZN(n15198) );
  INV_X1 U18104 ( .A(n15198), .ZN(n18757) );
  OAI22_X1 U18105 ( .A1(n18935), .A2(n18757), .B1(n18956), .B2(n14907), .ZN(
        n14912) );
  INV_X1 U18106 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n14909) );
  OAI22_X1 U18107 ( .A1(n14910), .A2(n14909), .B1(n19066), .B2(n14908), .ZN(
        n14911) );
  AOI211_X1 U18108 ( .C1(n18928), .C2(BUF1_REG_19__SCAN_IN), .A(n14912), .B(
        n14911), .ZN(n14913) );
  OAI21_X1 U18109 ( .B1(n14914), .B2(n18986), .A(n14913), .ZN(P2_U2900) );
  NOR2_X1 U18110 ( .A1(n15997), .A2(n14915), .ZN(n14916) );
  AOI211_X1 U18111 ( .C1(n15984), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14917), .B(n14916), .ZN(n14918) );
  OAI21_X1 U18112 ( .B1(n14919), .B2(n15406), .A(n14918), .ZN(n14920) );
  AOI21_X1 U18113 ( .B1(n14921), .B2(n13164), .A(n14920), .ZN(n14922) );
  OAI21_X1 U18114 ( .B1(n14923), .B2(n15976), .A(n14922), .ZN(P2_U2984) );
  OAI21_X1 U18115 ( .B1(n19047), .B2(n14925), .A(n14924), .ZN(n14926) );
  AOI21_X1 U18116 ( .B1(n19037), .B2(n14927), .A(n14926), .ZN(n14928) );
  OAI21_X1 U18117 ( .B1(n15821), .B2(n15406), .A(n14928), .ZN(n14929) );
  AOI21_X1 U18118 ( .B1(n14930), .B2(n13164), .A(n14929), .ZN(n14931) );
  OAI21_X1 U18119 ( .B1(n14932), .B2(n15976), .A(n14931), .ZN(P2_U2985) );
  NAND2_X1 U18120 ( .A1(n14934), .A2(n14933), .ZN(n14935) );
  INV_X1 U18121 ( .A(n14935), .ZN(n14937) );
  NAND2_X1 U18122 ( .A1(n14951), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14952) );
  OAI21_X1 U18123 ( .B1(n14937), .B2(n14936), .A(n14952), .ZN(n14940) );
  XNOR2_X1 U18124 ( .A(n14938), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14939) );
  XNOR2_X1 U18125 ( .A(n14940), .B(n14939), .ZN(n15093) );
  INV_X1 U18126 ( .A(n15087), .ZN(n14946) );
  NOR2_X1 U18127 ( .A1(n18765), .A2(n19740), .ZN(n15083) );
  AOI21_X1 U18128 ( .B1(n15984), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15083), .ZN(n14941) );
  OAI21_X1 U18129 ( .B1(n15997), .B2(n14942), .A(n14941), .ZN(n14945) );
  AND2_X1 U18130 ( .A1(n14948), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14949) );
  OAI21_X1 U18131 ( .B1(n15093), .B2(n15976), .A(n14947), .ZN(P2_U2986) );
  INV_X1 U18132 ( .A(n14949), .ZN(n14950) );
  OAI21_X1 U18133 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14948), .A(
        n14950), .ZN(n15104) );
  OR2_X1 U18134 ( .A1(n14951), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15094) );
  NAND3_X1 U18135 ( .A1(n15094), .A2(n14952), .A3(n19040), .ZN(n14957) );
  NAND2_X1 U18136 ( .A1(n19038), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15095) );
  OAI21_X1 U18137 ( .B1(n19047), .B2(n15831), .A(n15095), .ZN(n14954) );
  NOR2_X1 U18138 ( .A1(n15835), .A2(n15406), .ZN(n14953) );
  AOI211_X1 U18139 ( .C1(n19037), .C2(n14955), .A(n14954), .B(n14953), .ZN(
        n14956) );
  OAI211_X1 U18140 ( .C1(n15977), .C2(n15104), .A(n14957), .B(n14956), .ZN(
        P2_U2987) );
  NOR2_X1 U18141 ( .A1(n14958), .A2(n14968), .ZN(n14959) );
  XOR2_X1 U18142 ( .A(n14960), .B(n14959), .Z(n15114) );
  NOR2_X1 U18143 ( .A1(n18765), .A2(n14961), .ZN(n15106) );
  AOI21_X1 U18144 ( .B1(n15984), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15106), .ZN(n14962) );
  OAI21_X1 U18145 ( .B1(n15997), .B2(n15852), .A(n14962), .ZN(n14965) );
  NOR2_X1 U18146 ( .A1(n14971), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14963) );
  NOR2_X1 U18147 ( .A1(n15109), .A2(n15977), .ZN(n14964) );
  OAI21_X1 U18148 ( .B1(n15114), .B2(n15976), .A(n14966), .ZN(P2_U2988) );
  NOR2_X1 U18149 ( .A1(n14969), .A2(n14968), .ZN(n14970) );
  XOR2_X1 U18150 ( .A(n14967), .B(n14970), .Z(n15126) );
  AOI21_X1 U18151 ( .B1(n15115), .B2(n14984), .A(n14971), .ZN(n15124) );
  NAND2_X1 U18152 ( .A1(n19038), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15118) );
  OAI21_X1 U18153 ( .B1(n19047), .B2(n14972), .A(n15118), .ZN(n14973) );
  AOI21_X1 U18154 ( .B1(n19037), .B2(n14974), .A(n14973), .ZN(n14975) );
  OAI21_X1 U18155 ( .B1(n15117), .B2(n15406), .A(n14975), .ZN(n14976) );
  AOI21_X1 U18156 ( .B1(n15124), .B2(n13164), .A(n14976), .ZN(n14977) );
  OAI21_X1 U18157 ( .B1(n15126), .B2(n15976), .A(n14977), .ZN(P2_U2989) );
  XOR2_X1 U18158 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n14978), .Z(
        n14979) );
  XNOR2_X1 U18159 ( .A(n14980), .B(n14979), .ZN(n15127) );
  INV_X1 U18160 ( .A(n15127), .ZN(n14989) );
  INV_X1 U18161 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15868) );
  INV_X1 U18162 ( .A(n15876), .ZN(n14981) );
  NAND2_X1 U18163 ( .A1(n19037), .A2(n14981), .ZN(n14982) );
  NAND2_X1 U18164 ( .A1(n19038), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n15129) );
  OAI211_X1 U18165 ( .C1(n19047), .C2(n15868), .A(n14982), .B(n15129), .ZN(
        n14986) );
  INV_X1 U18166 ( .A(n14983), .ZN(n14993) );
  OAI21_X1 U18167 ( .B1(n14993), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n14984), .ZN(n15136) );
  NOR2_X1 U18168 ( .A1(n15136), .A2(n15977), .ZN(n14985) );
  AOI211_X1 U18169 ( .C1(n14987), .C2(n19042), .A(n14986), .B(n14985), .ZN(
        n14988) );
  OAI21_X1 U18170 ( .B1(n14989), .B2(n15976), .A(n14988), .ZN(P2_U2990) );
  XNOR2_X1 U18171 ( .A(n14990), .B(n14991), .ZN(n15149) );
  AOI21_X1 U18172 ( .B1(n15139), .B2(n14992), .A(n14993), .ZN(n15147) );
  OAI22_X1 U18173 ( .A1(n19047), .A2(n14994), .B1(n19731), .B2(n18765), .ZN(
        n14995) );
  AOI21_X1 U18174 ( .B1(n19037), .B2(n14996), .A(n14995), .ZN(n14997) );
  OAI21_X1 U18175 ( .B1(n15144), .B2(n15406), .A(n14997), .ZN(n14998) );
  AOI21_X1 U18176 ( .B1(n15147), .B2(n13164), .A(n14998), .ZN(n14999) );
  OAI21_X1 U18177 ( .B1(n15149), .B2(n15976), .A(n14999), .ZN(P2_U2991) );
  NAND2_X1 U18178 ( .A1(n15001), .A2(n15000), .ZN(n15016) );
  NAND2_X1 U18179 ( .A1(n15937), .A2(n15003), .ZN(n15261) );
  OAI21_X2 U18180 ( .B1(n15939), .B2(n15004), .A(n15941), .ZN(n15249) );
  INV_X1 U18181 ( .A(n15005), .ZN(n15246) );
  INV_X1 U18182 ( .A(n15247), .ZN(n15006) );
  INV_X1 U18183 ( .A(n15007), .ZN(n15236) );
  OAI21_X2 U18184 ( .B1(n15237), .B2(n15236), .A(n15008), .ZN(n15065) );
  INV_X1 U18185 ( .A(n15009), .ZN(n15011) );
  NAND2_X1 U18186 ( .A1(n15011), .A2(n15010), .ZN(n15066) );
  INV_X1 U18187 ( .A(n15012), .ZN(n15014) );
  NAND2_X1 U18188 ( .A1(n15027), .A2(n15031), .ZN(n15015) );
  XOR2_X1 U18189 ( .A(n15016), .B(n15015), .Z(n15181) );
  NAND2_X1 U18190 ( .A1(n15320), .A2(n15017), .ZN(n15025) );
  AND2_X1 U18191 ( .A1(n15320), .A2(n15018), .ZN(n15163) );
  AOI21_X1 U18192 ( .B1(n15168), .B2(n15025), .A(n15163), .ZN(n15179) );
  NOR2_X1 U18193 ( .A1(n18765), .A2(n19728), .ZN(n15173) );
  NOR2_X1 U18194 ( .A1(n15997), .A2(n15019), .ZN(n15020) );
  AOI211_X1 U18195 ( .C1(n15984), .C2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15173), .B(n15020), .ZN(n15021) );
  OAI21_X1 U18196 ( .B1(n15406), .B2(n15176), .A(n15021), .ZN(n15022) );
  AOI21_X1 U18197 ( .B1(n15179), .B2(n13164), .A(n15022), .ZN(n15023) );
  OAI21_X1 U18198 ( .B1(n15181), .B2(n15976), .A(n15023), .ZN(P2_U2993) );
  INV_X1 U18199 ( .A(n15320), .ZN(n15024) );
  NOR2_X1 U18200 ( .A1(n15024), .A2(n15212), .ZN(n15053) );
  NAND2_X1 U18201 ( .A1(n15053), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15054) );
  OAI21_X1 U18202 ( .B1(n15054), .B2(n15200), .A(n15188), .ZN(n15026) );
  NAND2_X1 U18203 ( .A1(n15026), .A2(n15025), .ZN(n15194) );
  INV_X1 U18204 ( .A(n15027), .ZN(n15032) );
  AOI21_X1 U18205 ( .B1(n15029), .B2(n15031), .A(n15028), .ZN(n15030) );
  AOI21_X1 U18206 ( .B1(n15032), .B2(n15031), .A(n15030), .ZN(n15182) );
  NAND2_X1 U18207 ( .A1(n15182), .A2(n19040), .ZN(n15037) );
  NAND2_X1 U18208 ( .A1(n19038), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n15184) );
  NAND2_X1 U18209 ( .A1(n15984), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15033) );
  OAI211_X1 U18210 ( .C1(n15889), .C2(n15406), .A(n15184), .B(n15033), .ZN(
        n15034) );
  AOI21_X1 U18211 ( .B1(n19037), .B2(n15035), .A(n15034), .ZN(n15036) );
  OAI211_X1 U18212 ( .C1(n15977), .C2(n15194), .A(n15037), .B(n15036), .ZN(
        P2_U2994) );
  NAND2_X1 U18213 ( .A1(n15039), .A2(n15038), .ZN(n15042) );
  INV_X1 U18214 ( .A(n15050), .ZN(n15040) );
  AOI21_X1 U18215 ( .B1(n15052), .B2(n15049), .A(n15040), .ZN(n15041) );
  XOR2_X1 U18216 ( .A(n15042), .B(n15041), .Z(n15205) );
  XNOR2_X1 U18217 ( .A(n15054), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15203) );
  NAND2_X1 U18218 ( .A1(n19038), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15196) );
  OAI21_X1 U18219 ( .B1(n19047), .B2(n15043), .A(n15196), .ZN(n15044) );
  AOI21_X1 U18220 ( .B1(n15045), .B2(n19037), .A(n15044), .ZN(n15046) );
  OAI21_X1 U18221 ( .B1(n15406), .B2(n18758), .A(n15046), .ZN(n15047) );
  AOI21_X1 U18222 ( .B1(n15203), .B2(n13164), .A(n15047), .ZN(n15048) );
  OAI21_X1 U18223 ( .B1(n15205), .B2(n15976), .A(n15048), .ZN(P2_U2995) );
  NAND2_X1 U18224 ( .A1(n15050), .A2(n15049), .ZN(n15051) );
  XNOR2_X1 U18225 ( .A(n15052), .B(n15051), .ZN(n15220) );
  INV_X1 U18226 ( .A(n15053), .ZN(n15071) );
  INV_X1 U18227 ( .A(n15054), .ZN(n15055) );
  AOI21_X1 U18228 ( .B1(n15207), .B2(n15071), .A(n15055), .ZN(n15218) );
  NOR2_X1 U18229 ( .A1(n18765), .A2(n19723), .ZN(n15214) );
  NAND2_X1 U18230 ( .A1(n15057), .A2(n15056), .ZN(n15058) );
  NAND2_X1 U18231 ( .A1(n15059), .A2(n15058), .ZN(n18772) );
  NOR2_X1 U18232 ( .A1(n15406), .A2(n18772), .ZN(n15060) );
  AOI211_X1 U18233 ( .C1(n15984), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15214), .B(n15060), .ZN(n15061) );
  OAI21_X1 U18234 ( .B1(n15997), .B2(n15062), .A(n15061), .ZN(n15063) );
  AOI21_X1 U18235 ( .B1(n15218), .B2(n13164), .A(n15063), .ZN(n15064) );
  OAI21_X1 U18236 ( .B1(n15220), .B2(n15976), .A(n15064), .ZN(P2_U2996) );
  XOR2_X1 U18237 ( .A(n15066), .B(n15065), .Z(n15235) );
  NOR2_X1 U18238 ( .A1(n19721), .A2(n18765), .ZN(n15069) );
  OAI22_X1 U18239 ( .A1(n19047), .A2(n15067), .B1(n15997), .B2(n18796), .ZN(
        n15068) );
  AOI211_X1 U18240 ( .C1(n19042), .C2(n18779), .A(n15069), .B(n15068), .ZN(
        n15073) );
  NAND2_X1 U18241 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15070) );
  OAI211_X1 U18242 ( .C1(n15917), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15071), .B(n13164), .ZN(n15072) );
  OAI211_X1 U18243 ( .C1(n15235), .C2(n15976), .A(n15073), .B(n15072), .ZN(
        P2_U2997) );
  XNOR2_X1 U18244 ( .A(n15074), .B(n15075), .ZN(n15353) );
  NAND2_X1 U18245 ( .A1(n11221), .A2(n15986), .ZN(n15077) );
  XNOR2_X1 U18246 ( .A(n15076), .B(n15077), .ZN(n15350) );
  OAI22_X1 U18247 ( .A1(n19047), .A2(n9712), .B1(n15997), .B2(n18851), .ZN(
        n15079) );
  OAI22_X1 U18248 ( .A1(n15406), .A2(n18857), .B1(n18765), .B2(n19709), .ZN(
        n15078) );
  AOI211_X1 U18249 ( .C1(n15350), .C2(n19040), .A(n15079), .B(n15078), .ZN(
        n15080) );
  OAI21_X1 U18250 ( .B1(n15353), .B2(n15977), .A(n15080), .ZN(P2_U3007) );
  NAND3_X1 U18251 ( .A1(n15081), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n9950), .ZN(n15086) );
  INV_X1 U18252 ( .A(n15082), .ZN(n15084) );
  AOI21_X1 U18253 ( .B1(n16010), .B2(n15084), .A(n15083), .ZN(n15085) );
  OAI211_X1 U18254 ( .C1(n15087), .C2(n15343), .A(n15086), .B(n15085), .ZN(
        n15090) );
  NOR2_X1 U18255 ( .A1(n15088), .A2(n15352), .ZN(n15089) );
  OAI21_X1 U18256 ( .B1(n15093), .B2(n15234), .A(n15092), .ZN(P2_U3018) );
  NAND3_X1 U18257 ( .A1(n15094), .A2(n14952), .A3(n16015), .ZN(n15103) );
  INV_X1 U18258 ( .A(n15835), .ZN(n15097) );
  OAI21_X1 U18259 ( .B1(n15348), .B2(n15834), .A(n15095), .ZN(n15096) );
  AOI21_X1 U18260 ( .B1(n15097), .B2(n16014), .A(n15096), .ZN(n15098) );
  OAI21_X1 U18261 ( .B1(n15099), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15098), .ZN(n15100) );
  AOI21_X1 U18262 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15101), .A(
        n15100), .ZN(n15102) );
  OAI211_X1 U18263 ( .C1(n15104), .C2(n15352), .A(n15103), .B(n15102), .ZN(
        P2_U3019) );
  INV_X1 U18264 ( .A(n15116), .ZN(n15112) );
  XNOR2_X1 U18265 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15108) );
  NOR2_X1 U18266 ( .A1(n15348), .A2(n15847), .ZN(n15105) );
  AOI211_X1 U18267 ( .C1(n15849), .C2(n16014), .A(n15106), .B(n15105), .ZN(
        n15107) );
  OAI21_X1 U18268 ( .B1(n15121), .B2(n15108), .A(n15107), .ZN(n15111) );
  NOR2_X1 U18269 ( .A1(n15109), .A2(n15352), .ZN(n15110) );
  OAI21_X1 U18270 ( .B1(n15114), .B2(n15234), .A(n15113), .ZN(P2_U3020) );
  NOR2_X1 U18271 ( .A1(n15116), .A2(n15115), .ZN(n15123) );
  INV_X1 U18272 ( .A(n15117), .ZN(n15860) );
  OAI21_X1 U18273 ( .B1(n15348), .B2(n15858), .A(n15118), .ZN(n15119) );
  AOI21_X1 U18274 ( .B1(n15860), .B2(n16014), .A(n15119), .ZN(n15120) );
  OAI21_X1 U18275 ( .B1(n15121), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15120), .ZN(n15122) );
  AOI211_X1 U18276 ( .C1(n15124), .C2(n16011), .A(n15123), .B(n15122), .ZN(
        n15125) );
  OAI21_X1 U18277 ( .B1(n15126), .B2(n15234), .A(n15125), .ZN(P2_U3021) );
  NAND2_X1 U18278 ( .A1(n15127), .A2(n16015), .ZN(n15135) );
  INV_X1 U18279 ( .A(n15140), .ZN(n15137) );
  OAI21_X1 U18280 ( .B1(n15137), .B2(n15128), .A(n11312), .ZN(n15132) );
  NOR2_X1 U18281 ( .A1(n15872), .A2(n15343), .ZN(n15131) );
  OAI21_X1 U18282 ( .B1(n15348), .B2(n15871), .A(n15129), .ZN(n15130) );
  AOI211_X1 U18283 ( .C1(n15133), .C2(n15132), .A(n15131), .B(n15130), .ZN(
        n15134) );
  OAI211_X1 U18284 ( .C1(n15352), .C2(n15136), .A(n15135), .B(n15134), .ZN(
        P2_U3022) );
  NOR2_X1 U18285 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n15137), .ZN(
        n15155) );
  INV_X1 U18286 ( .A(n15155), .ZN(n15138) );
  AOI21_X1 U18287 ( .B1(n15169), .B2(n15138), .A(n15139), .ZN(n15146) );
  NAND3_X1 U18288 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n15140), .A3(
        n15139), .ZN(n15143) );
  AOI22_X1 U18289 ( .A1(n16010), .A2(n15141), .B1(P2_REIP_REG_23__SCAN_IN), 
        .B2(n19038), .ZN(n15142) );
  OAI211_X1 U18290 ( .C1(n15343), .C2(n15144), .A(n15143), .B(n15142), .ZN(
        n15145) );
  AOI211_X1 U18291 ( .C1(n15147), .C2(n16011), .A(n15146), .B(n15145), .ZN(
        n15148) );
  OAI21_X1 U18292 ( .B1(n15149), .B2(n15234), .A(n15148), .ZN(P2_U3023) );
  INV_X1 U18293 ( .A(n15150), .ZN(n15152) );
  AND2_X1 U18294 ( .A1(n15152), .A2(n15151), .ZN(n15153) );
  XNOR2_X1 U18295 ( .A(n15154), .B(n15153), .ZN(n15907) );
  INV_X1 U18296 ( .A(n15908), .ZN(n15160) );
  INV_X1 U18297 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19729) );
  NOR2_X1 U18298 ( .A1(n19729), .A2(n18765), .ZN(n15156) );
  NOR2_X1 U18299 ( .A1(n15156), .A2(n15155), .ZN(n15157) );
  OAI21_X1 U18300 ( .B1(n15348), .B2(n15158), .A(n15157), .ZN(n15159) );
  AOI21_X1 U18301 ( .B1(n15160), .B2(n16014), .A(n15159), .ZN(n15161) );
  OAI21_X1 U18302 ( .B1(n15169), .B2(n15162), .A(n15161), .ZN(n15166) );
  OR2_X1 U18303 ( .A1(n15163), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15164) );
  NAND2_X1 U18304 ( .A1(n15164), .A2(n14992), .ZN(n15911) );
  NOR2_X1 U18305 ( .A1(n15911), .A2(n15352), .ZN(n15165) );
  AOI211_X1 U18306 ( .C1(n16015), .C2(n15907), .A(n15166), .B(n15165), .ZN(
        n15167) );
  INV_X1 U18307 ( .A(n15167), .ZN(P2_U3024) );
  NOR2_X1 U18308 ( .A1(n15169), .A2(n15168), .ZN(n15178) );
  INV_X1 U18309 ( .A(n15170), .ZN(n15174) );
  NOR2_X1 U18310 ( .A1(n15171), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15172) );
  AOI211_X1 U18311 ( .C1(n16010), .C2(n15174), .A(n15173), .B(n15172), .ZN(
        n15175) );
  OAI21_X1 U18312 ( .B1(n15176), .B2(n15343), .A(n15175), .ZN(n15177) );
  AOI211_X1 U18313 ( .C1(n15179), .C2(n16011), .A(n15178), .B(n15177), .ZN(
        n15180) );
  OAI21_X1 U18314 ( .B1(n15181), .B2(n15234), .A(n15180), .ZN(P2_U3025) );
  NAND2_X1 U18315 ( .A1(n15182), .A2(n16015), .ZN(n15193) );
  INV_X1 U18316 ( .A(n15889), .ZN(n15191) );
  AND2_X1 U18317 ( .A1(n15330), .A2(n15185), .ZN(n15187) );
  NAND3_X1 U18318 ( .A1(n15188), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n15187), .ZN(n15183) );
  OAI211_X1 U18319 ( .C1(n15348), .C2(n15896), .A(n15184), .B(n15183), .ZN(
        n15190) );
  INV_X1 U18320 ( .A(n15185), .ZN(n15186) );
  INV_X1 U18321 ( .A(n16020), .ZN(n15328) );
  AOI21_X1 U18322 ( .B1(n15186), .B2(n15206), .A(n15328), .ZN(n15201) );
  NAND2_X1 U18323 ( .A1(n15200), .A2(n15187), .ZN(n15195) );
  AOI21_X1 U18324 ( .B1(n15201), .B2(n15195), .A(n15188), .ZN(n15189) );
  AOI211_X1 U18325 ( .C1(n15191), .C2(n16014), .A(n15190), .B(n15189), .ZN(
        n15192) );
  OAI211_X1 U18326 ( .C1(n15194), .C2(n15352), .A(n15193), .B(n15192), .ZN(
        P2_U3026) );
  OAI211_X1 U18327 ( .C1(n18758), .C2(n15343), .A(n15196), .B(n15195), .ZN(
        n15197) );
  AOI21_X1 U18328 ( .B1(n16010), .B2(n15198), .A(n15197), .ZN(n15199) );
  OAI21_X1 U18329 ( .B1(n15201), .B2(n15200), .A(n15199), .ZN(n15202) );
  AOI21_X1 U18330 ( .B1(n15203), .B2(n16011), .A(n15202), .ZN(n15204) );
  OAI21_X1 U18331 ( .B1(n15205), .B2(n15234), .A(n15204), .ZN(P2_U3027) );
  AOI21_X1 U18332 ( .B1(n15212), .B2(n15206), .A(n15328), .ZN(n15208) );
  NOR2_X1 U18333 ( .A1(n15208), .A2(n15207), .ZN(n15217) );
  NAND2_X1 U18334 ( .A1(n13958), .A2(n15209), .ZN(n15210) );
  AND2_X1 U18335 ( .A1(n15211), .A2(n15210), .ZN(n18770) );
  NOR3_X1 U18336 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15226), .A3(
        n15212), .ZN(n15213) );
  AOI211_X1 U18337 ( .C1(n16010), .C2(n18770), .A(n15214), .B(n15213), .ZN(
        n15215) );
  OAI21_X1 U18338 ( .B1(n15343), .B2(n18772), .A(n15215), .ZN(n15216) );
  AOI211_X1 U18339 ( .C1(n15218), .C2(n16011), .A(n15217), .B(n15216), .ZN(
        n15219) );
  OAI21_X1 U18340 ( .B1(n15220), .B2(n15234), .A(n15219), .ZN(P2_U3028) );
  INV_X1 U18341 ( .A(n15221), .ZN(n15224) );
  OAI21_X1 U18342 ( .B1(n15225), .B2(n15222), .A(n16020), .ZN(n15251) );
  OAI21_X1 U18343 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15225), .A(
        n15240), .ZN(n15232) );
  NOR2_X1 U18344 ( .A1(n15227), .A2(n15226), .ZN(n16003) );
  INV_X1 U18345 ( .A(n16003), .ZN(n15262) );
  OAI22_X1 U18346 ( .A1(n15916), .A2(n15352), .B1(n15262), .B2(n16002), .ZN(
        n15243) );
  INV_X1 U18347 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15228) );
  NAND4_X1 U18348 ( .A1(n15243), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15228), .A4(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15230) );
  AOI22_X1 U18349 ( .A1(n16014), .A2(n18779), .B1(n19038), .B2(
        P2_REIP_REG_17__SCAN_IN), .ZN(n15229) );
  OAI211_X1 U18350 ( .C1(n15348), .C2(n18792), .A(n15230), .B(n15229), .ZN(
        n15231) );
  AOI21_X1 U18351 ( .B1(n15232), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15231), .ZN(n15233) );
  OAI21_X1 U18352 ( .B1(n15235), .B2(n15234), .A(n15233), .ZN(P2_U3029) );
  XNOR2_X1 U18353 ( .A(n15237), .B(n15236), .ZN(n15920) );
  NOR2_X1 U18354 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n15252), .ZN(
        n15244) );
  AOI22_X1 U18355 ( .A1(n15919), .A2(n16014), .B1(P2_REIP_REG_16__SCAN_IN), 
        .B2(n19038), .ZN(n15238) );
  OAI21_X1 U18356 ( .B1(n15348), .B2(n18929), .A(n15238), .ZN(n15242) );
  NOR2_X1 U18357 ( .A1(n15240), .A2(n15239), .ZN(n15241) );
  AOI211_X1 U18358 ( .C1(n15244), .C2(n15243), .A(n15242), .B(n15241), .ZN(
        n15245) );
  OAI21_X1 U18359 ( .B1(n15234), .B2(n15920), .A(n15245), .ZN(P2_U3030) );
  XNOR2_X1 U18360 ( .A(n15916), .B(n15252), .ZN(n15927) );
  NOR2_X1 U18361 ( .A1(n15247), .A2(n15246), .ZN(n15248) );
  XNOR2_X1 U18362 ( .A(n15249), .B(n15248), .ZN(n15928) );
  INV_X1 U18363 ( .A(n15928), .ZN(n15259) );
  NOR2_X1 U18364 ( .A1(n16002), .A2(n15262), .ZN(n15253) );
  INV_X1 U18365 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19717) );
  NOR2_X1 U18366 ( .A1(n19717), .A2(n18765), .ZN(n15250) );
  AOI221_X1 U18367 ( .B1(n15253), .B2(n15252), .C1(n15251), .C2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(n15250), .ZN(n15254) );
  INV_X1 U18368 ( .A(n15254), .ZN(n15258) );
  INV_X1 U18369 ( .A(n15930), .ZN(n18803) );
  OR2_X1 U18370 ( .A1(n15255), .A2(n13804), .ZN(n15256) );
  NAND2_X1 U18371 ( .A1(n15256), .A2(n13927), .ZN(n18937) );
  OAI22_X1 U18372 ( .A1(n15343), .A2(n18803), .B1(n15348), .B2(n18937), .ZN(
        n15257) );
  AOI211_X1 U18373 ( .C1(n15259), .C2(n16015), .A(n15258), .B(n15257), .ZN(
        n15260) );
  OAI21_X1 U18374 ( .B1(n15352), .B2(n15927), .A(n15260), .ZN(P2_U3031) );
  AOI21_X1 U18375 ( .B1(n15002), .B2(n15261), .A(n15939), .ZN(n15949) );
  NOR2_X1 U18376 ( .A1(n15329), .A2(n15328), .ZN(n15292) );
  AOI21_X1 U18377 ( .B1(n15292), .B2(n15294), .A(n15293), .ZN(n15998) );
  INV_X1 U18378 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n19716) );
  NOR2_X1 U18379 ( .A1(n19716), .A2(n18765), .ZN(n15264) );
  AOI211_X1 U18380 ( .C1(n11268), .C2(n11247), .A(n16004), .B(n15262), .ZN(
        n15263) );
  AOI211_X1 U18381 ( .C1(n15998), .C2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15264), .B(n15263), .ZN(n15269) );
  NOR2_X2 U18382 ( .A1(n11247), .A2(n15283), .ZN(n15954) );
  INV_X1 U18383 ( .A(n15283), .ZN(n15266) );
  NAND2_X1 U18384 ( .A1(n15266), .A2(n16004), .ZN(n15936) );
  OAI21_X1 U18385 ( .B1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15954), .A(
        n15936), .ZN(n15948) );
  OAI22_X1 U18386 ( .A1(n15348), .A2(n18942), .B1(n15352), .B2(n15948), .ZN(
        n15267) );
  AOI21_X1 U18387 ( .B1(n16014), .B2(n20957), .A(n15267), .ZN(n15268) );
  OAI211_X1 U18388 ( .C1(n15949), .C2(n15234), .A(n15269), .B(n15268), .ZN(
        P2_U3033) );
  NAND2_X1 U18389 ( .A1(n15283), .A2(n11247), .ZN(n15958) );
  INV_X1 U18390 ( .A(n15954), .ZN(n15270) );
  NAND3_X1 U18391 ( .A1(n15958), .A2(n16011), .A3(n15270), .ZN(n15282) );
  NOR2_X1 U18392 ( .A1(n10397), .A2(n18765), .ZN(n15271) );
  AOI221_X1 U18393 ( .B1(n15998), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), 
        .C1(n16003), .C2(n11247), .A(n15271), .ZN(n15281) );
  XNOR2_X1 U18394 ( .A(n15298), .B(n15272), .ZN(n18944) );
  OR2_X1 U18395 ( .A1(n15273), .A2(n13525), .ZN(n15274) );
  NAND2_X1 U18396 ( .A1(n15274), .A2(n13816), .ZN(n18902) );
  OAI22_X1 U18397 ( .A1(n18944), .A2(n15348), .B1(n15343), .B2(n18902), .ZN(
        n15275) );
  INV_X1 U18398 ( .A(n15275), .ZN(n15280) );
  NAND2_X1 U18399 ( .A1(n9654), .A2(n15276), .ZN(n15277) );
  XNOR2_X1 U18400 ( .A(n15278), .B(n15277), .ZN(n15955) );
  OR2_X1 U18401 ( .A1(n15955), .A2(n15234), .ZN(n15279) );
  NAND4_X1 U18402 ( .A1(n15282), .A2(n15281), .A3(n15280), .A4(n15279), .ZN(
        P2_U3034) );
  NOR2_X1 U18403 ( .A1(n15319), .A2(n11226), .ZN(n15310) );
  OAI21_X1 U18404 ( .B1(n15310), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15283), .ZN(n15963) );
  AND2_X1 U18405 ( .A1(n15285), .A2(n15284), .ZN(n15324) );
  NAND2_X1 U18406 ( .A1(n15324), .A2(n15321), .ZN(n15326) );
  INV_X1 U18407 ( .A(n15307), .ZN(n15287) );
  OAI21_X1 U18408 ( .B1(n15326), .B2(n15287), .A(n15286), .ZN(n15291) );
  AND2_X1 U18409 ( .A1(n15289), .A2(n15288), .ZN(n15290) );
  XNOR2_X1 U18410 ( .A(n15291), .B(n15290), .ZN(n15962) );
  NOR2_X1 U18411 ( .A1(n15293), .A2(n15292), .ZN(n15314) );
  INV_X1 U18412 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19715) );
  NOR2_X1 U18413 ( .A1(n19715), .A2(n18765), .ZN(n15297) );
  NAND2_X1 U18414 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15330), .ZN(
        n15311) );
  AOI211_X1 U18415 ( .C1(n15295), .C2(n11226), .A(n15294), .B(n15311), .ZN(
        n15296) );
  AOI211_X1 U18416 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15314), .A(
        n15297), .B(n15296), .ZN(n15303) );
  OAI21_X1 U18417 ( .B1(n15300), .B2(n15299), .A(n15298), .ZN(n18946) );
  OAI22_X1 U18418 ( .A1(n18946), .A2(n15348), .B1(n15343), .B2(n18822), .ZN(
        n15301) );
  INV_X1 U18419 ( .A(n15301), .ZN(n15302) );
  OAI211_X1 U18420 ( .C1(n15962), .C2(n15234), .A(n15303), .B(n15302), .ZN(
        n15304) );
  INV_X1 U18421 ( .A(n15304), .ZN(n15305) );
  OAI21_X1 U18422 ( .B1(n15963), .B2(n15352), .A(n15305), .ZN(P2_U3035) );
  NAND2_X1 U18423 ( .A1(n15307), .A2(n15306), .ZN(n15309) );
  NAND2_X1 U18424 ( .A1(n15326), .A2(n15322), .ZN(n15308) );
  XOR2_X1 U18425 ( .A(n15309), .B(n15308), .Z(n15968) );
  AOI21_X1 U18426 ( .B1(n11226), .B2(n15319), .A(n15310), .ZN(n15969) );
  NAND2_X1 U18427 ( .A1(n15969), .A2(n16011), .ZN(n15318) );
  NOR2_X1 U18428 ( .A1(n10365), .A2(n18765), .ZN(n15313) );
  NOR2_X1 U18429 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n15311), .ZN(
        n15312) );
  AOI211_X1 U18430 ( .C1(n15314), .C2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n15313), .B(n15312), .ZN(n15315) );
  OAI21_X1 U18431 ( .B1(n15348), .B2(n18949), .A(n15315), .ZN(n15316) );
  AOI21_X1 U18432 ( .B1(n16014), .B2(n18907), .A(n15316), .ZN(n15317) );
  OAI211_X1 U18433 ( .C1(n15968), .C2(n15234), .A(n15318), .B(n15317), .ZN(
        P2_U3036) );
  OAI21_X1 U18434 ( .B1(n15320), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15319), .ZN(n15978) );
  INV_X1 U18435 ( .A(n15322), .ZN(n15325) );
  AND2_X1 U18436 ( .A1(n15322), .A2(n15321), .ZN(n15323) );
  OAI22_X1 U18437 ( .A1(n15326), .A2(n15325), .B1(n15324), .B2(n15323), .ZN(
        n15975) );
  INV_X1 U18438 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19712) );
  NOR2_X1 U18439 ( .A1(n19712), .A2(n18765), .ZN(n15327) );
  AOI221_X1 U18440 ( .B1(n15330), .B2(n15329), .C1(n15328), .C2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n15327), .ZN(n15336) );
  OR2_X1 U18441 ( .A1(n15331), .A2(n13768), .ZN(n15333) );
  NAND2_X1 U18442 ( .A1(n15333), .A2(n15332), .ZN(n18951) );
  OAI22_X1 U18443 ( .A1(n15343), .A2(n18843), .B1(n15348), .B2(n18951), .ZN(
        n15334) );
  INV_X1 U18444 ( .A(n15334), .ZN(n15335) );
  OAI211_X1 U18445 ( .C1(n15975), .C2(n15234), .A(n15336), .B(n15335), .ZN(
        n15337) );
  INV_X1 U18446 ( .A(n15337), .ZN(n15338) );
  OAI21_X1 U18447 ( .B1(n15978), .B2(n15352), .A(n15338), .ZN(P2_U3037) );
  OAI21_X1 U18448 ( .B1(n15341), .B2(n15340), .A(n15339), .ZN(n18955) );
  NAND2_X1 U18449 ( .A1(n16009), .A2(n15342), .ZN(n15347) );
  OAI22_X1 U18450 ( .A1(n15343), .A2(n18857), .B1(n19709), .B2(n18765), .ZN(
        n15344) );
  AOI21_X1 U18451 ( .B1(n15345), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n15344), .ZN(n15346) );
  OAI211_X1 U18452 ( .C1(n15348), .C2(n18955), .A(n15347), .B(n15346), .ZN(
        n15349) );
  AOI21_X1 U18453 ( .B1(n15350), .B2(n16015), .A(n15349), .ZN(n15351) );
  OAI21_X1 U18454 ( .B1(n15353), .B2(n15352), .A(n15351), .ZN(P2_U3039) );
  INV_X1 U18455 ( .A(n16071), .ZN(n15389) );
  NOR2_X1 U18456 ( .A1(n18849), .A2(n15354), .ZN(n18877) );
  AOI21_X1 U18457 ( .B1(n18849), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18877), .ZN(n15367) );
  NAND2_X1 U18458 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15367), .ZN(n15362) );
  OR2_X1 U18459 ( .A1(n15355), .A2(n15373), .ZN(n15360) );
  NAND2_X1 U18460 ( .A1(n15357), .A2(n15356), .ZN(n15371) );
  MUX2_X1 U18461 ( .A(n15371), .B(n15379), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15358) );
  INV_X1 U18462 ( .A(n15358), .ZN(n15359) );
  NAND2_X1 U18463 ( .A1(n15360), .A2(n15359), .ZN(n16023) );
  NAND2_X1 U18464 ( .A1(n16023), .A2(n19758), .ZN(n15361) );
  OAI211_X1 U18465 ( .C1(n15363), .C2(n15389), .A(n15362), .B(n15361), .ZN(
        n15364) );
  MUX2_X1 U18466 ( .A(n15364), .B(n9587), .S(n15393), .Z(P2_U3601) );
  OAI21_X1 U18467 ( .B1(n9567), .B2(n15366), .A(n15365), .ZN(n15392) );
  NOR2_X1 U18468 ( .A1(n15367), .A2(n19668), .ZN(n15391) );
  INV_X1 U18469 ( .A(n15391), .ZN(n15375) );
  NAND2_X1 U18470 ( .A1(n15379), .A2(n15368), .ZN(n15380) );
  XNOR2_X1 U18471 ( .A(n15369), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15370) );
  NAND2_X1 U18472 ( .A1(n15371), .A2(n15370), .ZN(n15372) );
  OAI211_X1 U18473 ( .C1(n11070), .C2(n15373), .A(n15380), .B(n15372), .ZN(
        n16024) );
  AOI22_X1 U18474 ( .A1(n19782), .A2(n16071), .B1(n19758), .B2(n16024), .ZN(
        n15374) );
  OAI21_X1 U18475 ( .B1(n15392), .B2(n15375), .A(n15374), .ZN(n15376) );
  INV_X1 U18476 ( .A(n15393), .ZN(n15446) );
  MUX2_X1 U18477 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15376), .S(
        n15446), .Z(P2_U3600) );
  NOR2_X1 U18478 ( .A1(n15377), .A2(n11659), .ZN(n15385) );
  NAND2_X1 U18479 ( .A1(n15378), .A2(n15385), .ZN(n15383) );
  NAND2_X1 U18480 ( .A1(n15379), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15381) );
  MUX2_X1 U18481 ( .A(n15381), .B(n15380), .S(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n15382) );
  OAI211_X1 U18482 ( .C1(n15385), .C2(n15384), .A(n15383), .B(n15382), .ZN(
        n15386) );
  AOI21_X1 U18483 ( .B1(n15388), .B2(n15387), .A(n15386), .ZN(n16021) );
  OAI22_X1 U18484 ( .A1(n19770), .A2(n15389), .B1(n19666), .B2(n16021), .ZN(
        n15390) );
  AOI21_X1 U18485 ( .B1(n15392), .B2(n15391), .A(n15390), .ZN(n15394) );
  MUX2_X1 U18486 ( .A(n15394), .B(n16022), .S(n15393), .Z(n15395) );
  INV_X1 U18487 ( .A(n15395), .ZN(P2_U3599) );
  NAND2_X1 U18488 ( .A1(n19335), .A2(n19274), .ZN(n19126) );
  OAI21_X1 U18489 ( .B1(n19659), .B2(n19116), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n15397) );
  NAND2_X1 U18490 ( .A1(n15397), .A2(n19759), .ZN(n15400) );
  NAND2_X1 U18491 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15398), .ZN(
        n19607) );
  NOR2_X1 U18492 ( .A1(n19797), .A2(n19607), .ZN(n19654) );
  NAND2_X1 U18493 ( .A1(n19769), .A2(n19779), .ZN(n19160) );
  NOR2_X1 U18494 ( .A1(n19336), .A2(n19160), .ZN(n19087) );
  NOR2_X1 U18495 ( .A1(n19654), .A2(n19087), .ZN(n15403) );
  OAI21_X1 U18496 ( .B1(n15401), .B2(n19087), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15399) );
  INV_X1 U18497 ( .A(n19091), .ZN(n15413) );
  INV_X1 U18498 ( .A(n15895), .ZN(n18974) );
  NOR2_X2 U18499 ( .A1(n19549), .A2(n18974), .ZN(n19635) );
  INV_X1 U18500 ( .A(n19635), .ZN(n15412) );
  INV_X1 U18501 ( .A(n15400), .ZN(n15404) );
  AOI211_X1 U18502 ( .C1(n15401), .C2(n19611), .A(n19087), .B(n19759), .ZN(
        n15402) );
  AOI211_X2 U18503 ( .C1(n15404), .C2(n15403), .A(n19549), .B(n15402), .ZN(
        n19094) );
  INV_X1 U18504 ( .A(n19094), .ZN(n15410) );
  NOR2_X2 U18505 ( .A1(n15405), .A2(n15406), .ZN(n19078) );
  INV_X1 U18506 ( .A(n19078), .ZN(n19090) );
  NOR2_X2 U18507 ( .A1(n15407), .A2(n15406), .ZN(n19079) );
  INV_X1 U18508 ( .A(n19079), .ZN(n19089) );
  OAI22_X1 U18509 ( .A1(n14851), .A2(n19090), .B1(n16156), .B2(n19089), .ZN(
        n19636) );
  INV_X1 U18510 ( .A(n19636), .ZN(n19533) );
  AOI22_X1 U18511 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19079), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19078), .ZN(n19641) );
  INV_X1 U18512 ( .A(n19641), .ZN(n19530) );
  AND2_X1 U18513 ( .A1(n9590), .A2(n19086), .ZN(n19634) );
  AOI22_X1 U18514 ( .A1(n19530), .A2(n19116), .B1(n19087), .B2(n19634), .ZN(
        n15408) );
  OAI21_X1 U18515 ( .B1(n19640), .B2(n19533), .A(n15408), .ZN(n15409) );
  AOI21_X1 U18516 ( .B1(n15410), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A(
        n15409), .ZN(n15411) );
  OAI21_X1 U18517 ( .B1(n15413), .B2(n15412), .A(n15411), .ZN(P2_U3052) );
  AOI22_X1 U18518 ( .A1(n9577), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15415) );
  OAI21_X1 U18519 ( .B1(n10741), .B2(n20936), .A(n15415), .ZN(n15427) );
  INV_X1 U18520 ( .A(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15425) );
  AOI22_X1 U18521 ( .A1(n17010), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15424) );
  INV_X1 U18522 ( .A(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15417) );
  AOI22_X1 U18523 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16734), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15416) );
  OAI21_X1 U18524 ( .B1(n16962), .B2(n15417), .A(n15416), .ZN(n15422) );
  AOI22_X1 U18525 ( .A1(n10758), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15420) );
  AOI22_X1 U18526 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9585), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15419) );
  OAI211_X1 U18527 ( .C1(n15418), .C2(n18069), .A(n15420), .B(n15419), .ZN(
        n15421) );
  AOI211_X1 U18528 ( .C1(n9571), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n15422), .B(n15421), .ZN(n15423) );
  OAI211_X1 U18529 ( .C1(n17001), .C2(n15425), .A(n15424), .B(n15423), .ZN(
        n15426) );
  AOI211_X1 U18530 ( .C1(n17025), .C2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n15427), .B(n15426), .ZN(n17152) );
  NAND2_X1 U18531 ( .A1(n18077), .A2(n18059), .ZN(n15428) );
  NOR2_X2 U18532 ( .A1(n17049), .A2(n18077), .ZN(n17043) );
  INV_X2 U18533 ( .A(n17043), .ZN(n17054) );
  INV_X1 U18534 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17045) );
  NOR2_X2 U18535 ( .A1(n17044), .A2(n17045), .ZN(n17048) );
  INV_X1 U18536 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n17037) );
  INV_X1 U18537 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16558) );
  INV_X1 U18538 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n20863) );
  AND2_X2 U18539 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n16985), .ZN(n17005) );
  INV_X1 U18540 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16951) );
  NOR2_X1 U18541 ( .A1(n17043), .A2(n16932), .ZN(n15433) );
  OAI21_X1 U18542 ( .B1(n16948), .B2(P3_EBX_REG_13__SCAN_IN), .A(n15433), .ZN(
        n15434) );
  OAI21_X1 U18543 ( .B1(n17152), .B2(n17054), .A(n15434), .ZN(P3_U2690) );
  INV_X1 U18544 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18035) );
  NAND2_X1 U18545 ( .A1(n18035), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18082) );
  NOR2_X1 U18546 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18653), .ZN(
        n18678) );
  NOR2_X1 U18547 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18708) );
  AOI21_X1 U18548 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(
        P3_STATE2_REG_2__SCAN_IN), .A(n18708), .ZN(n18561) );
  OR2_X1 U18549 ( .A1(n18678), .A2(n18561), .ZN(n18038) );
  NAND2_X1 U18550 ( .A1(n18705), .A2(n18038), .ZN(n18084) );
  INV_X1 U18551 ( .A(n18084), .ZN(n18354) );
  NOR2_X1 U18552 ( .A1(n16734), .A2(n15435), .ZN(n18027) );
  AOI21_X1 U18553 ( .B1(n18027), .B2(n16249), .A(n18651), .ZN(n15436) );
  NOR2_X1 U18554 ( .A1(n18354), .A2(n15436), .ZN(n18028) );
  INV_X1 U18555 ( .A(n18028), .ZN(n18034) );
  NAND2_X1 U18556 ( .A1(n18082), .A2(n18034), .ZN(n15439) );
  INV_X1 U18557 ( .A(n15439), .ZN(n15438) );
  NAND3_X1 U18558 ( .A1(n18715), .A2(n18653), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18296) );
  OAI21_X1 U18559 ( .B1(n18715), .B2(n18664), .A(n18653), .ZN(n18699) );
  INV_X1 U18560 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16281) );
  NOR2_X1 U18561 ( .A1(n18664), .A2(n16281), .ZN(n17671) );
  OAI22_X1 U18562 ( .A1(n18699), .A2(n17671), .B1(n18653), .B2(n18035), .ZN(
        n15441) );
  NAND3_X1 U18563 ( .A1(n18530), .A2(n18034), .A3(n15441), .ZN(n15437) );
  OAI221_X1 U18564 ( .B1(n18530), .B2(n15438), .C1(n18530), .C2(n18296), .A(
        n15437), .ZN(P3_U2864) );
  NAND2_X1 U18565 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18258) );
  NOR2_X1 U18566 ( .A1(n18699), .A2(n17671), .ZN(n15440) );
  AOI221_X1 U18567 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18258), .C1(n15440), 
        .C2(n18258), .A(n15439), .ZN(n18033) );
  INV_X1 U18568 ( .A(n18296), .ZN(n18406) );
  OAI221_X1 U18569 ( .B1(n18406), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18406), .C2(n15441), .A(n18034), .ZN(n18031) );
  AOI22_X1 U18570 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18033), .B1(
        n18031), .B2(n18535), .ZN(P3_U2865) );
  INV_X1 U18571 ( .A(n16043), .ZN(n15442) );
  NOR4_X1 U18572 ( .A1(n16047), .A2(n15442), .A3(n19666), .A4(n19054), .ZN(
        n15443) );
  NAND2_X1 U18573 ( .A1(n15446), .A2(n15443), .ZN(n15444) );
  OAI21_X1 U18574 ( .B1(n15446), .B2(n15445), .A(n15444), .ZN(P2_U3595) );
  NOR2_X1 U18575 ( .A1(n15448), .A2(n15447), .ZN(n15449) );
  XOR2_X1 U18576 ( .A(n15449), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(
        n16129) );
  OAI21_X1 U18577 ( .B1(n17907), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15450), .ZN(n16133) );
  NOR2_X1 U18578 ( .A1(n15498), .A2(n17702), .ZN(n16125) );
  INV_X1 U18579 ( .A(n16082), .ZN(n17179) );
  NOR2_X1 U18580 ( .A1(n18023), .A2(n18491), .ZN(n18022) );
  NAND2_X1 U18581 ( .A1(n17179), .A2(n18022), .ZN(n17933) );
  NOR2_X1 U18582 ( .A1(n15498), .A2(n17703), .ZN(n16114) );
  NOR2_X1 U18583 ( .A1(n18023), .A2(n17999), .ZN(n18020) );
  OAI22_X1 U18584 ( .A1(n16125), .A2(n17933), .B1(n16114), .B2(n18015), .ZN(
        n15500) );
  AOI21_X1 U18585 ( .B1(n17909), .B2(n16133), .A(n15500), .ZN(n15452) );
  OAI21_X1 U18586 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17972), .A(
        n15452), .ZN(n15453) );
  AOI22_X1 U18587 ( .A1(n17815), .A2(P3_REIP_REG_29__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15453), .ZN(n15456) );
  OAI222_X1 U18588 ( .A1(n18015), .A2(n17703), .B1(n15454), .B2(n18023), .C1(
        n17702), .C2(n17933), .ZN(n15499) );
  NAND3_X1 U18589 ( .A1(n16113), .A2(n20920), .A3(n15499), .ZN(n15455) );
  OAI211_X1 U18590 ( .C1(n16129), .C2(n17939), .A(n15456), .B(n15455), .ZN(
        P3_U2833) );
  INV_X1 U18591 ( .A(n15457), .ZN(n15471) );
  NAND2_X1 U18592 ( .A1(n15459), .A2(n15458), .ZN(n15467) );
  OAI22_X1 U18593 ( .A1(n20767), .A2(n15461), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15460), .ZN(n20757) );
  OR2_X1 U18594 ( .A1(n15462), .A2(n11846), .ZN(n20765) );
  INV_X1 U18595 ( .A(n20765), .ZN(n15463) );
  NOR2_X1 U18596 ( .A1(n20757), .A2(n15463), .ZN(n15464) );
  AOI22_X1 U18597 ( .A1(n15467), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n15464), .B2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n15465) );
  INV_X1 U18598 ( .A(n15465), .ZN(n15466) );
  OAI21_X1 U18599 ( .B1(n15467), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15466), .ZN(n15468) );
  AOI222_X1 U18600 ( .A1(n15469), .A2(n12676), .B1(n15469), .B2(n15468), .C1(
        n12676), .C2(n15468), .ZN(n15470) );
  AOI222_X1 U18601 ( .A1(n15471), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .B1(n15471), .B2(n15470), .C1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .C2(n15470), .ZN(n15478) );
  OAI21_X1 U18602 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15472), .ZN(n15473) );
  NAND4_X1 U18603 ( .A1(n15486), .A2(n15475), .A3(n15474), .A4(n15473), .ZN(
        n15476) );
  AOI211_X1 U18604 ( .C1(n20058), .C2(n15478), .A(n15477), .B(n15476), .ZN(
        n15493) );
  AND2_X1 U18605 ( .A1(n15480), .A2(n15479), .ZN(n15483) );
  NAND3_X1 U18606 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20693), .A3(n20071), 
        .ZN(n15481) );
  AOI22_X1 U18607 ( .A1(n15483), .A2(n15482), .B1(n20686), .B2(n15481), .ZN(
        n15803) );
  OAI221_X1 U18608 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n15493), 
        .A(n15803), .ZN(n15809) );
  NOR2_X1 U18609 ( .A1(n15484), .A2(n15805), .ZN(n15485) );
  NOR2_X1 U18610 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15485), .ZN(n15491) );
  AND3_X1 U18611 ( .A1(n15487), .A2(n15486), .A3(n15802), .ZN(n20771) );
  AOI211_X1 U18612 ( .C1(n20693), .C2(n20074), .A(n20771), .B(n15488), .ZN(
        n15489) );
  NAND2_X1 U18613 ( .A1(n15809), .A2(n15489), .ZN(n15490) );
  AOI22_X1 U18614 ( .A1(n15809), .A2(n15491), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n15490), .ZN(n15492) );
  OAI21_X1 U18615 ( .B1(n15493), .B2(n19815), .A(n15492), .ZN(P1_U3161) );
  NAND2_X1 U18616 ( .A1(n15495), .A2(n15494), .ZN(n15497) );
  XOR2_X1 U18617 ( .A(n15497), .B(n15496), .Z(n16111) );
  INV_X1 U18618 ( .A(n18017), .ZN(n17821) );
  NOR2_X1 U18619 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15498), .ZN(
        n16107) );
  AOI22_X1 U18620 ( .A1(n17821), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n16107), 
        .B2(n15499), .ZN(n15503) );
  OAI21_X1 U18621 ( .B1(n15501), .B2(n15500), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15502) );
  OAI211_X1 U18622 ( .C1(n16111), .C2(n17939), .A(n15503), .B(n15502), .ZN(
        P3_U2832) );
  INV_X1 U18623 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20702) );
  INV_X1 U18624 ( .A(HOLD), .ZN(n19687) );
  NOR2_X1 U18625 ( .A1(n20702), .A2(n19687), .ZN(n20690) );
  AOI22_X1 U18626 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n15506) );
  NAND2_X1 U18627 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20693), .ZN(n15504) );
  OAI211_X1 U18628 ( .C1(n20690), .C2(n15506), .A(n15505), .B(n15504), .ZN(
        P1_U3195) );
  AND2_X1 U18629 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(n19934), .ZN(P1_U2905)
         );
  NAND2_X1 U18630 ( .A1(n19665), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19670) );
  NOR2_X1 U18631 ( .A1(n19669), .A2(n19670), .ZN(n16062) );
  AOI221_X1 U18632 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(
        P2_STATE2_REG_1__SCAN_IN), .C1(P2_STATEBS16_REG_SCAN_IN), .C2(
        P2_STATE2_REG_1__SCAN_IN), .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n15507)
         );
  NOR3_X1 U18633 ( .A1(n16062), .A2(n16064), .A3(n15507), .ZN(P2_U3178) );
  OAI221_X1 U18634 ( .B1(n11350), .B2(n16079), .C1(n16063), .C2(n16079), .A(
        n19549), .ZN(n19796) );
  NOR2_X1 U18635 ( .A1(n15508), .A2(n19796), .ZN(P2_U3047) );
  NAND3_X1 U18636 ( .A1(n18046), .A2(n18040), .A3(n15509), .ZN(n15510) );
  INV_X1 U18637 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17267) );
  NAND2_X1 U18638 ( .A1(n18077), .A2(n15513), .ZN(n17101) );
  NAND2_X2 U18639 ( .A1(n15513), .A2(n17176), .ZN(n17199) );
  NAND2_X1 U18640 ( .A1(n15512), .A2(n17172), .ZN(n17202) );
  AOI22_X1 U18641 ( .A1(n17205), .A2(BUF2_REG_0__SCAN_IN), .B1(n17204), .B2(
        n17695), .ZN(n15514) );
  OAI221_X1 U18642 ( .B1(n17207), .B2(n17267), .C1(n17207), .C2(n17101), .A(
        n15514), .ZN(P3_U2735) );
  AOI22_X1 U18643 ( .A1(n19876), .A2(P1_EBX_REG_23__SCAN_IN), .B1(n15515), 
        .B2(n19907), .ZN(n15524) );
  AND2_X1 U18644 ( .A1(n19882), .A2(n15516), .ZN(n15526) );
  AOI21_X1 U18645 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(n15526), .A(
        P1_REIP_REG_23__SCAN_IN), .ZN(n15519) );
  INV_X1 U18646 ( .A(n15517), .ZN(n15518) );
  OAI22_X1 U18647 ( .A1(n15520), .A2(n15609), .B1(n15519), .B2(n15518), .ZN(
        n15521) );
  AOI21_X1 U18648 ( .B1(n9561), .B2(n15522), .A(n15521), .ZN(n15523) );
  OAI211_X1 U18649 ( .C1(n15525), .C2(n19894), .A(n15524), .B(n15523), .ZN(
        P1_U2817) );
  AOI22_X1 U18650 ( .A1(n19876), .A2(P1_EBX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n19866), .ZN(n15535) );
  INV_X1 U18651 ( .A(n15630), .ZN(n15527) );
  INV_X1 U18652 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20731) );
  AOI22_X1 U18653 ( .A1(n15527), .A2(n19907), .B1(n15526), .B2(n20731), .ZN(
        n15534) );
  INV_X1 U18654 ( .A(n15528), .ZN(n15627) );
  XNOR2_X1 U18655 ( .A(n15530), .B(n15529), .ZN(n15680) );
  AOI22_X1 U18656 ( .A1(n15627), .A2(n19870), .B1(n9561), .B2(n15680), .ZN(
        n15533) );
  NOR2_X1 U18657 ( .A1(n19852), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15538) );
  OAI21_X1 U18658 ( .B1(n15537), .B2(n19852), .A(n15531), .ZN(n15550) );
  OAI21_X1 U18659 ( .B1(n15538), .B2(n15550), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n15532) );
  NAND4_X1 U18660 ( .A1(n15535), .A2(n15534), .A3(n15533), .A4(n15532), .ZN(
        P1_U2818) );
  AOI22_X1 U18661 ( .A1(n15536), .A2(n19907), .B1(P1_REIP_REG_21__SCAN_IN), 
        .B2(n15550), .ZN(n15543) );
  AOI22_X1 U18662 ( .A1(n15538), .A2(n15537), .B1(n19876), .B2(
        P1_EBX_REG_21__SCAN_IN), .ZN(n15542) );
  INV_X1 U18663 ( .A(n15539), .ZN(n15618) );
  AOI22_X1 U18664 ( .A1(n15619), .A2(n19870), .B1(n15618), .B2(n9561), .ZN(
        n15541) );
  NAND2_X1 U18665 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n19866), .ZN(
        n15540) );
  NAND4_X1 U18666 ( .A1(n15543), .A2(n15542), .A3(n15541), .A4(n15540), .ZN(
        P1_U2819) );
  AOI22_X1 U18667 ( .A1(n19876), .A2(P1_EBX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19866), .ZN(n15552) );
  OAI21_X1 U18668 ( .B1(n19852), .B2(n15545), .A(n15544), .ZN(n15549) );
  OAI22_X1 U18669 ( .A1(n15547), .A2(n15609), .B1(n15586), .B2(n15546), .ZN(
        n15548) );
  AOI21_X1 U18670 ( .B1(n15550), .B2(n15549), .A(n15548), .ZN(n15551) );
  OAI211_X1 U18671 ( .C1(n15553), .C2(n19890), .A(n15552), .B(n15551), .ZN(
        P1_U2820) );
  NAND2_X1 U18672 ( .A1(n19876), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n15555) );
  AOI21_X1 U18673 ( .B1(n19866), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n19854), .ZN(n15554) );
  OAI211_X1 U18674 ( .C1(n19890), .C2(n15556), .A(n15555), .B(n15554), .ZN(
        n15557) );
  AOI21_X1 U18675 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n15558), .A(n15557), 
        .ZN(n15561) );
  INV_X1 U18676 ( .A(n15559), .ZN(n15560) );
  OAI211_X1 U18677 ( .C1(n15562), .C2(n15609), .A(n15561), .B(n15560), .ZN(
        n15563) );
  INV_X1 U18678 ( .A(n15563), .ZN(n15564) );
  OAI21_X1 U18679 ( .B1(n15586), .B2(n15695), .A(n15564), .ZN(P1_U2822) );
  AOI21_X1 U18680 ( .B1(n20723), .B2(n15566), .A(n15565), .ZN(n15567) );
  AOI22_X1 U18681 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n15575), .B1(n15568), 
        .B2(n15567), .ZN(n15574) );
  NOR2_X1 U18682 ( .A1(n19890), .A2(n15639), .ZN(n15571) );
  INV_X1 U18683 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15569) );
  OAI21_X1 U18684 ( .B1(n19894), .B2(n15569), .A(n19878), .ZN(n15570) );
  AOI211_X1 U18685 ( .C1(P1_EBX_REG_16__SCAN_IN), .C2(n19876), .A(n15571), .B(
        n15570), .ZN(n15573) );
  AOI22_X1 U18686 ( .A1(n15636), .A2(n19870), .B1(n9561), .B2(n15711), .ZN(
        n15572) );
  NAND3_X1 U18687 ( .A1(n15574), .A2(n15573), .A3(n15572), .ZN(P1_U2824) );
  INV_X1 U18688 ( .A(n15575), .ZN(n15584) );
  AOI21_X1 U18689 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n15576), .A(
        P1_REIP_REG_14__SCAN_IN), .ZN(n15583) );
  INV_X1 U18690 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15577) );
  OAI21_X1 U18691 ( .B1(n19894), .B2(n15577), .A(n19878), .ZN(n15580) );
  NOR2_X1 U18692 ( .A1(n15578), .A2(n15586), .ZN(n15579) );
  AOI211_X1 U18693 ( .C1(n19876), .C2(P1_EBX_REG_14__SCAN_IN), .A(n15580), .B(
        n15579), .ZN(n15582) );
  AOI22_X1 U18694 ( .A1(n15641), .A2(n19870), .B1(n19907), .B2(n15640), .ZN(
        n15581) );
  OAI211_X1 U18695 ( .C1(n15584), .C2(n15583), .A(n15582), .B(n15581), .ZN(
        P1_U2826) );
  OAI22_X1 U18696 ( .A1(n15587), .A2(n15586), .B1(n15585), .B2(n19897), .ZN(
        n15588) );
  AOI211_X1 U18697 ( .C1(n19866), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n19854), .B(n15588), .ZN(n15592) );
  NAND3_X1 U18698 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .A3(n19840), .ZN(n15601) );
  OAI21_X1 U18699 ( .B1(n15600), .B2(n15601), .A(n20718), .ZN(n15589) );
  AOI22_X1 U18700 ( .A1(n15646), .A2(n19907), .B1(n15590), .B2(n15589), .ZN(
        n15591) );
  OAI211_X1 U18701 ( .C1(n15609), .C2(n15593), .A(n15592), .B(n15591), .ZN(
        P1_U2828) );
  AOI21_X1 U18702 ( .B1(n19866), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n19854), .ZN(n15597) );
  AOI21_X1 U18703 ( .B1(n15595), .B2(n9609), .A(n15594), .ZN(n15736) );
  AOI22_X1 U18704 ( .A1(n15736), .A2(n9561), .B1(n19876), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n15596) );
  OAI211_X1 U18705 ( .C1(n15659), .C2(n19890), .A(n15597), .B(n15596), .ZN(
        n15598) );
  AOI21_X1 U18706 ( .B1(n19870), .B2(n15656), .A(n15598), .ZN(n15599) );
  OAI221_X1 U18707 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n15601), .C1(n15600), 
        .C2(n15615), .A(n15599), .ZN(P1_U2829) );
  NOR2_X1 U18708 ( .A1(n20713), .A2(n15602), .ZN(n15603) );
  AOI22_X1 U18709 ( .A1(n15604), .A2(n19907), .B1(n15603), .B2(n15614), .ZN(
        n15613) );
  NAND2_X1 U18710 ( .A1(n19876), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n15605) );
  OAI211_X1 U18711 ( .C1(n19894), .C2(n15606), .A(n15605), .B(n19878), .ZN(
        n15607) );
  AOI21_X1 U18712 ( .B1(n15746), .B2(n9561), .A(n15607), .ZN(n15608) );
  OAI21_X1 U18713 ( .B1(n15610), .B2(n15609), .A(n15608), .ZN(n15611) );
  INV_X1 U18714 ( .A(n15611), .ZN(n15612) );
  OAI211_X1 U18715 ( .C1(n15615), .C2(n15614), .A(n15613), .B(n15612), .ZN(
        P1_U2830) );
  AOI22_X1 U18716 ( .A1(n15627), .A2(n19914), .B1(n19913), .B2(n15680), .ZN(
        n15616) );
  OAI21_X1 U18717 ( .B1(n19918), .B2(n15617), .A(n15616), .ZN(P1_U2850) );
  AOI22_X1 U18718 ( .A1(n15619), .A2(n19914), .B1(n15618), .B2(n19913), .ZN(
        n15620) );
  OAI21_X1 U18719 ( .B1(n19918), .B2(n15621), .A(n15620), .ZN(P1_U2851) );
  AOI22_X1 U18720 ( .A1(n15656), .A2(n19914), .B1(n19913), .B2(n15736), .ZN(
        n15622) );
  OAI21_X1 U18721 ( .B1(n19918), .B2(n15623), .A(n15622), .ZN(P1_U2861) );
  AOI22_X1 U18722 ( .A1(n19984), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n20053), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15629) );
  NAND2_X1 U18723 ( .A1(n15625), .A2(n15624), .ZN(n15626) );
  XNOR2_X1 U18724 ( .A(n15626), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15681) );
  AOI22_X1 U18725 ( .A1(n15627), .A2(n13319), .B1(n19990), .B2(n15681), .ZN(
        n15628) );
  OAI211_X1 U18726 ( .C1(n19995), .C2(n15630), .A(n15629), .B(n15628), .ZN(
        P1_U2977) );
  AOI22_X1 U18727 ( .A1(n19984), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20053), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15638) );
  OAI22_X1 U18728 ( .A1(n15633), .A2(n15632), .B1(n15631), .B2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15634) );
  XOR2_X1 U18729 ( .A(n15635), .B(n15634), .Z(n15713) );
  AOI22_X1 U18730 ( .A1(n15713), .A2(n19990), .B1(n13319), .B2(n15636), .ZN(
        n15637) );
  OAI211_X1 U18731 ( .C1(n19995), .C2(n15639), .A(n15638), .B(n15637), .ZN(
        P1_U2983) );
  AOI22_X1 U18732 ( .A1(n19984), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20053), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15643) );
  AOI22_X1 U18733 ( .A1(n15641), .A2(n13319), .B1(n15647), .B2(n15640), .ZN(
        n15642) );
  OAI211_X1 U18734 ( .C1(n15644), .C2(n19822), .A(n15643), .B(n15642), .ZN(
        P1_U2985) );
  AOI22_X1 U18735 ( .A1(n19984), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20053), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15649) );
  AOI22_X1 U18736 ( .A1(n15647), .A2(n15646), .B1(n13319), .B2(n15645), .ZN(
        n15648) );
  OAI211_X1 U18737 ( .C1(n15650), .C2(n19822), .A(n15649), .B(n15648), .ZN(
        P1_U2987) );
  AOI22_X1 U18738 ( .A1(n19984), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20053), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15658) );
  NAND3_X1 U18739 ( .A1(n15652), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15651), .ZN(n15654) );
  NAND2_X1 U18740 ( .A1(n15654), .A2(n15653), .ZN(n15655) );
  XNOR2_X1 U18741 ( .A(n15655), .B(n15741), .ZN(n15738) );
  AOI22_X1 U18742 ( .A1(n19990), .A2(n15738), .B1(n13319), .B2(n15656), .ZN(
        n15657) );
  OAI211_X1 U18743 ( .C1(n19995), .C2(n15659), .A(n15658), .B(n15657), .ZN(
        P1_U2988) );
  AOI22_X1 U18744 ( .A1(n19984), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20053), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15665) );
  NAND2_X1 U18745 ( .A1(n15662), .A2(n15661), .ZN(n15663) );
  XNOR2_X1 U18746 ( .A(n15660), .B(n15663), .ZN(n15773) );
  AOI22_X1 U18747 ( .A1(n15773), .A2(n19990), .B1(n13319), .B2(n19851), .ZN(
        n15664) );
  OAI211_X1 U18748 ( .C1(n19995), .C2(n19855), .A(n15665), .B(n15664), .ZN(
        P1_U2992) );
  AOI22_X1 U18749 ( .A1(n19984), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20053), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15671) );
  XNOR2_X1 U18750 ( .A(n15667), .B(n15666), .ZN(n15668) );
  XNOR2_X1 U18751 ( .A(n15669), .B(n15668), .ZN(n15781) );
  AOI22_X1 U18752 ( .A1(n15781), .A2(n19990), .B1(n13319), .B2(n19915), .ZN(
        n15670) );
  OAI211_X1 U18753 ( .C1(n19995), .C2(n19868), .A(n15671), .B(n15670), .ZN(
        P1_U2993) );
  AOI22_X1 U18754 ( .A1(n19984), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20053), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n15678) );
  OR2_X1 U18755 ( .A1(n15673), .A2(n15672), .ZN(n15674) );
  AND2_X1 U18756 ( .A1(n15675), .A2(n15674), .ZN(n15787) );
  NOR2_X1 U18757 ( .A1(n19884), .A2(n20067), .ZN(n15676) );
  AOI21_X1 U18758 ( .B1(n15787), .B2(n19990), .A(n15676), .ZN(n15677) );
  OAI211_X1 U18759 ( .C1(n19995), .C2(n19891), .A(n15678), .B(n15677), .ZN(
        P1_U2994) );
  AOI22_X1 U18760 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n15679), .B1(
        n20053), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15686) );
  AOI22_X1 U18761 ( .A1(n15681), .A2(n20036), .B1(n20042), .B2(n15680), .ZN(
        n15685) );
  OAI211_X1 U18762 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15683), .B(n15682), .ZN(
        n15684) );
  NAND3_X1 U18763 ( .A1(n15686), .A2(n15685), .A3(n15684), .ZN(P1_U3009) );
  AOI22_X1 U18764 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15687), .B1(
        n20053), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15692) );
  INV_X1 U18765 ( .A(n15688), .ZN(n15690) );
  AOI22_X1 U18766 ( .A1(n15690), .A2(n20036), .B1(n20042), .B2(n15689), .ZN(
        n15691) );
  OAI211_X1 U18767 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15693), .A(
        n15692), .B(n15691), .ZN(P1_U3012) );
  AOI21_X1 U18768 ( .B1(n15694), .B2(n20031), .A(n15731), .ZN(n15709) );
  NOR2_X1 U18769 ( .A1(n15694), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15698) );
  OAI22_X1 U18770 ( .A1(n15696), .A2(n20050), .B1(n20049), .B2(n15695), .ZN(
        n15697) );
  AOI21_X1 U18771 ( .B1(n15698), .B2(n15702), .A(n15697), .ZN(n15700) );
  NAND2_X1 U18772 ( .A1(n20053), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15699) );
  OAI211_X1 U18773 ( .C1(n15709), .C2(n15701), .A(n15700), .B(n15699), .ZN(
        P1_U3013) );
  NAND2_X1 U18774 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15702), .ZN(
        n15710) );
  NOR2_X1 U18775 ( .A1(n15725), .A2(n15710), .ZN(n15712) );
  AOI21_X1 U18776 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15712), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15708) );
  INV_X1 U18777 ( .A(n15703), .ZN(n15705) );
  AOI22_X1 U18778 ( .A1(n15705), .A2(n20036), .B1(n20001), .B2(n15704), .ZN(
        n15707) );
  NAND2_X1 U18779 ( .A1(n20053), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15706) );
  OAI211_X1 U18780 ( .C1(n15709), .C2(n15708), .A(n15707), .B(n15706), .ZN(
        P1_U3014) );
  NOR2_X1 U18781 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n15710), .ZN(
        n15721) );
  AOI211_X1 U18782 ( .C1(n15718), .C2(n20031), .A(n15721), .B(n15731), .ZN(
        n15717) );
  AOI22_X1 U18783 ( .A1(n20053), .A2(P1_REIP_REG_16__SCAN_IN), .B1(n20001), 
        .B2(n15711), .ZN(n15715) );
  AOI22_X1 U18784 ( .A1(n15713), .A2(n20036), .B1(n15712), .B2(n15716), .ZN(
        n15714) );
  OAI211_X1 U18785 ( .C1(n15717), .C2(n15716), .A(n15715), .B(n15714), .ZN(
        P1_U3015) );
  AOI21_X1 U18786 ( .B1(n15718), .B2(n20031), .A(n15731), .ZN(n15726) );
  AOI22_X1 U18787 ( .A1(n20053), .A2(P1_REIP_REG_15__SCAN_IN), .B1(n20042), 
        .B2(n15719), .ZN(n15724) );
  INV_X1 U18788 ( .A(n15720), .ZN(n15722) );
  AOI21_X1 U18789 ( .B1(n15722), .B2(n20036), .A(n15721), .ZN(n15723) );
  OAI211_X1 U18790 ( .C1(n15726), .C2(n15725), .A(n15724), .B(n15723), .ZN(
        P1_U3016) );
  AOI21_X1 U18791 ( .B1(n15729), .B2(n15728), .A(n15727), .ZN(n15735) );
  AOI22_X1 U18792 ( .A1(n20053), .A2(P1_REIP_REG_13__SCAN_IN), .B1(n20001), 
        .B2(n15730), .ZN(n15734) );
  AOI22_X1 U18793 ( .A1(n15732), .A2(n20036), .B1(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15731), .ZN(n15733) );
  OAI211_X1 U18794 ( .C1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n15735), .A(
        n15734), .B(n15733), .ZN(P1_U3018) );
  AOI22_X1 U18795 ( .A1(n20053), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n20042), 
        .B2(n15736), .ZN(n15740) );
  NOR4_X1 U18796 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15784), .A3(
        n15748), .A4(n15749), .ZN(n15737) );
  AOI21_X1 U18797 ( .B1(n15738), .B2(n20036), .A(n15737), .ZN(n15739) );
  OAI211_X1 U18798 ( .C1(n15742), .C2(n15741), .A(n15740), .B(n15739), .ZN(
        P1_U3020) );
  AOI21_X1 U18799 ( .B1(n15744), .B2(n15762), .A(n15743), .ZN(n15745) );
  AOI221_X1 U18800 ( .B1(n15745), .B2(n20031), .C1(n15748), .C2(n20031), .A(
        n20033), .ZN(n15758) );
  AOI222_X1 U18801 ( .A1(n15747), .A2(n20036), .B1(n20001), .B2(n15746), .C1(
        P1_REIP_REG_10__SCAN_IN), .C2(n20053), .ZN(n15751) );
  NOR2_X1 U18802 ( .A1(n15784), .A2(n15748), .ZN(n15754) );
  OAI211_X1 U18803 ( .C1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n15754), .B(n15749), .ZN(n15750) );
  OAI211_X1 U18804 ( .C1(n15758), .C2(n15752), .A(n15751), .B(n15750), .ZN(
        P1_U3021) );
  INV_X1 U18805 ( .A(n15753), .ZN(n19841) );
  AOI22_X1 U18806 ( .A1(n20053), .A2(P1_REIP_REG_9__SCAN_IN), .B1(n20001), 
        .B2(n19841), .ZN(n15757) );
  AOI22_X1 U18807 ( .A1(n15755), .A2(n20036), .B1(n12824), .B2(n15754), .ZN(
        n15756) );
  OAI211_X1 U18808 ( .C1(n15758), .C2(n12824), .A(n15757), .B(n15756), .ZN(
        P1_U3022) );
  NAND2_X1 U18809 ( .A1(n19998), .A2(n15759), .ZN(n15791) );
  NOR2_X1 U18810 ( .A1(n20029), .A2(n20044), .ZN(n15761) );
  OAI21_X1 U18811 ( .B1(n15762), .B2(n15761), .A(n15760), .ZN(n19996) );
  AOI211_X1 U18812 ( .C1(n20018), .C2(n15764), .A(n15763), .B(n19996), .ZN(
        n15786) );
  OAI21_X1 U18813 ( .B1(n15765), .B2(n15791), .A(n15786), .ZN(n15780) );
  AOI21_X1 U18814 ( .B1(n15666), .B2(n20031), .A(n15780), .ZN(n15777) );
  INV_X1 U18815 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15771) );
  INV_X1 U18816 ( .A(n15766), .ZN(n15767) );
  AOI222_X1 U18817 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20053), .B1(n20001), 
        .B2(n15768), .C1(n20036), .C2(n15767), .ZN(n15770) );
  NOR2_X1 U18818 ( .A1(n15666), .A2(n15784), .ZN(n15772) );
  OAI221_X1 U18819 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n15771), .C2(n15776), .A(
        n15772), .ZN(n15769) );
  OAI211_X1 U18820 ( .C1(n15777), .C2(n15771), .A(n15770), .B(n15769), .ZN(
        P1_U3023) );
  AOI22_X1 U18821 ( .A1(n20053), .A2(P1_REIP_REG_7__SCAN_IN), .B1(n20042), 
        .B2(n19857), .ZN(n15775) );
  AOI22_X1 U18822 ( .A1(n15773), .A2(n20036), .B1(n15772), .B2(n15776), .ZN(
        n15774) );
  OAI211_X1 U18823 ( .C1(n15777), .C2(n15776), .A(n15775), .B(n15774), .ZN(
        P1_U3024) );
  XNOR2_X1 U18824 ( .A(n15779), .B(n15778), .ZN(n19912) );
  AOI22_X1 U18825 ( .A1(n20053), .A2(P1_REIP_REG_6__SCAN_IN), .B1(n20001), 
        .B2(n19912), .ZN(n15783) );
  AOI22_X1 U18826 ( .A1(n15781), .A2(n20036), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15780), .ZN(n15782) );
  OAI211_X1 U18827 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n15784), .A(
        n15783), .B(n15782), .ZN(P1_U3025) );
  NAND2_X1 U18828 ( .A1(n15785), .A2(n20020), .ZN(n20012) );
  AOI22_X1 U18829 ( .A1(n20053), .A2(P1_REIP_REG_5__SCAN_IN), .B1(n20001), 
        .B2(n19877), .ZN(n15790) );
  INV_X1 U18830 ( .A(n15786), .ZN(n15788) );
  AOI22_X1 U18831 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15788), .B1(
        n15787), .B2(n20036), .ZN(n15789) );
  OAI211_X1 U18832 ( .C1(n15791), .C2(n20012), .A(n15790), .B(n15789), .ZN(
        P1_U3026) );
  INV_X1 U18833 ( .A(n20763), .ZN(n20761) );
  INV_X1 U18834 ( .A(n15792), .ZN(n15797) );
  INV_X1 U18835 ( .A(n15793), .ZN(n15795) );
  NAND4_X1 U18836 ( .A1(n15797), .A2(n15796), .A3(n15795), .A4(n15794), .ZN(
        n15798) );
  OAI21_X1 U18837 ( .B1(n20761), .B2(n15799), .A(n15798), .ZN(P1_U3468) );
  NAND4_X1 U18838 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20074), .A4(n20786), .ZN(n15800) );
  AND2_X1 U18839 ( .A1(n15801), .A2(n15800), .ZN(n20687) );
  INV_X1 U18840 ( .A(n15802), .ZN(n15804) );
  AOI21_X1 U18841 ( .B1(n20687), .B2(n15804), .A(n15803), .ZN(n15807) );
  OAI221_X1 U18842 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n15809), 
        .A(n15805), .ZN(n15806) );
  AOI211_X1 U18843 ( .C1(n20790), .C2(n20693), .A(n15807), .B(n15806), .ZN(
        P1_U3162) );
  OAI221_X1 U18844 ( .B1(n20756), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n20756), 
        .C2(n15809), .A(n15808), .ZN(P1_U3466) );
  INV_X1 U18845 ( .A(n18830), .ZN(n18790) );
  INV_X1 U18846 ( .A(n15810), .ZN(n15817) );
  AOI22_X1 U18847 ( .A1(n18818), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n18879), .ZN(n15812) );
  OAI21_X1 U18848 ( .B1(n18866), .B2(n19748), .A(n15812), .ZN(n15813) );
  AOI21_X1 U18849 ( .B1(n15811), .B2(n18869), .A(n15813), .ZN(n15814) );
  OAI21_X1 U18850 ( .B1(n15815), .B2(n18871), .A(n15814), .ZN(n15816) );
  OAI21_X1 U18851 ( .B1(n18790), .B2(n15819), .A(n15818), .ZN(P2_U2824) );
  AOI22_X1 U18852 ( .A1(n18853), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n18818), .ZN(n15830) );
  AOI22_X1 U18853 ( .A1(n15820), .A2(n18786), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18879), .ZN(n15829) );
  INV_X1 U18854 ( .A(n15821), .ZN(n15823) );
  AOI22_X1 U18855 ( .A1(n15823), .A2(n18874), .B1(n15822), .B2(n18869), .ZN(
        n15828) );
  OAI211_X1 U18856 ( .C1(n15826), .C2(n15825), .A(n19673), .B(n15824), .ZN(
        n15827) );
  NAND4_X1 U18857 ( .A1(n15830), .A2(n15829), .A3(n15828), .A4(n15827), .ZN(
        P2_U2826) );
  AOI22_X1 U18858 ( .A1(n18853), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_EBX_REG_27__SCAN_IN), .B2(n18818), .ZN(n15843) );
  OAI22_X1 U18859 ( .A1(n15832), .A2(n18871), .B1(n18821), .B2(n15831), .ZN(
        n15833) );
  INV_X1 U18860 ( .A(n15833), .ZN(n15842) );
  OAI22_X1 U18861 ( .A1(n15835), .A2(n18856), .B1(n15834), .B2(n18858), .ZN(
        n15836) );
  INV_X1 U18862 ( .A(n15836), .ZN(n15841) );
  OAI211_X1 U18863 ( .C1(n15839), .C2(n15838), .A(n19673), .B(n15837), .ZN(
        n15840) );
  NAND4_X1 U18864 ( .A1(n15843), .A2(n15842), .A3(n15841), .A4(n15840), .ZN(
        P2_U2828) );
  AOI22_X1 U18865 ( .A1(n18853), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n18818), .ZN(n15856) );
  INV_X1 U18866 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15844) );
  OAI22_X1 U18867 ( .A1(n15845), .A2(n18871), .B1(n18821), .B2(n15844), .ZN(
        n15846) );
  INV_X1 U18868 ( .A(n15846), .ZN(n15855) );
  INV_X1 U18869 ( .A(n15847), .ZN(n15848) );
  AOI22_X1 U18870 ( .A1(n15849), .A2(n18874), .B1(n15848), .B2(n18869), .ZN(
        n15854) );
  OAI211_X1 U18871 ( .C1(n15852), .C2(n15851), .A(n19673), .B(n15850), .ZN(
        n15853) );
  NAND4_X1 U18872 ( .A1(n15856), .A2(n15855), .A3(n15854), .A4(n15853), .ZN(
        P2_U2829) );
  AOI22_X1 U18873 ( .A1(n18853), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n18818), .ZN(n15867) );
  AOI22_X1 U18874 ( .A1(n15857), .A2(n18786), .B1(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18879), .ZN(n15866) );
  INV_X1 U18875 ( .A(n15858), .ZN(n15859) );
  AOI22_X1 U18876 ( .A1(n15860), .A2(n18874), .B1(n15859), .B2(n18869), .ZN(
        n15865) );
  OAI211_X1 U18877 ( .C1(n15863), .C2(n15862), .A(n19673), .B(n15861), .ZN(
        n15864) );
  NAND4_X1 U18878 ( .A1(n15867), .A2(n15866), .A3(n15865), .A4(n15864), .ZN(
        P2_U2830) );
  AOI22_X1 U18879 ( .A1(n18853), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_EBX_REG_24__SCAN_IN), .B2(n18818), .ZN(n15880) );
  OAI22_X1 U18880 ( .A1(n15869), .A2(n18871), .B1(n18821), .B2(n15868), .ZN(
        n15870) );
  INV_X1 U18881 ( .A(n15870), .ZN(n15879) );
  OAI22_X1 U18882 ( .A1(n15872), .A2(n18856), .B1(n15871), .B2(n18858), .ZN(
        n15873) );
  INV_X1 U18883 ( .A(n15873), .ZN(n15878) );
  OAI211_X1 U18884 ( .C1(n15876), .C2(n15875), .A(n19673), .B(n15874), .ZN(
        n15877) );
  NAND4_X1 U18885 ( .A1(n15880), .A2(n15879), .A3(n15878), .A4(n15877), .ZN(
        P2_U2831) );
  AOI22_X1 U18886 ( .A1(n20956), .A2(n15810), .B1(n15881), .B2(n20964), .ZN(
        P2_U2856) );
  AOI22_X1 U18887 ( .A1(n15882), .A2(n18891), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n20964), .ZN(n15883) );
  OAI21_X1 U18888 ( .B1(n20964), .B2(n15908), .A(n15883), .ZN(P2_U2865) );
  NOR2_X1 U18889 ( .A1(n14835), .A2(n15884), .ZN(n15885) );
  OR2_X1 U18890 ( .A1(n15886), .A2(n15885), .ZN(n15897) );
  OAI22_X1 U18891 ( .A1(n15897), .A2(n18919), .B1(n20956), .B2(n14771), .ZN(
        n15887) );
  INV_X1 U18892 ( .A(n15887), .ZN(n15888) );
  OAI21_X1 U18893 ( .B1(n20964), .B2(n15889), .A(n15888), .ZN(P2_U2867) );
  INV_X1 U18894 ( .A(n15890), .ZN(n15891) );
  AOI21_X1 U18895 ( .B1(n15893), .B2(n15892), .A(n15891), .ZN(n15903) );
  AOI22_X1 U18896 ( .A1(n15903), .A2(n18891), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n20964), .ZN(n15894) );
  OAI21_X1 U18897 ( .B1(n20964), .B2(n18772), .A(n15894), .ZN(P2_U2869) );
  AOI22_X1 U18898 ( .A1(n18926), .A2(n15895), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n18981), .ZN(n15901) );
  AOI22_X1 U18899 ( .A1(n18928), .A2(BUF1_REG_20__SCAN_IN), .B1(n18927), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n15900) );
  OAI22_X1 U18900 ( .A1(n15897), .A2(n18986), .B1(n18935), .B2(n15896), .ZN(
        n15898) );
  INV_X1 U18901 ( .A(n15898), .ZN(n15899) );
  NAND3_X1 U18902 ( .A1(n15901), .A2(n15900), .A3(n15899), .ZN(P2_U2899) );
  AOI22_X1 U18903 ( .A1(n18926), .A2(n15902), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n18981), .ZN(n15906) );
  AOI22_X1 U18904 ( .A1(n18928), .A2(BUF1_REG_18__SCAN_IN), .B1(n18927), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n15905) );
  AOI22_X1 U18905 ( .A1(n15903), .A2(n18970), .B1(n18982), .B2(n18770), .ZN(
        n15904) );
  NAND3_X1 U18906 ( .A1(n15906), .A2(n15905), .A3(n15904), .ZN(P2_U2901) );
  AOI22_X1 U18907 ( .A1(n15984), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19038), .ZN(n15914) );
  NAND2_X1 U18908 ( .A1(n15907), .A2(n19040), .ZN(n15910) );
  OR2_X1 U18909 ( .A1(n15908), .A2(n15406), .ZN(n15909) );
  OAI211_X1 U18910 ( .C1(n15911), .C2(n15977), .A(n15910), .B(n15909), .ZN(
        n15912) );
  INV_X1 U18911 ( .A(n15912), .ZN(n15913) );
  OAI211_X1 U18912 ( .C1(n15997), .C2(n15915), .A(n15914), .B(n15913), .ZN(
        P2_U2992) );
  AOI22_X1 U18913 ( .A1(n15984), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        P2_REIP_REG_16__SCAN_IN), .B2(n19038), .ZN(n15924) );
  INV_X1 U18914 ( .A(n15916), .ZN(n15934) );
  AOI21_X1 U18915 ( .B1(n15934), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15918) );
  NOR3_X1 U18916 ( .A1(n15918), .A2(n15917), .A3(n15977), .ZN(n15922) );
  INV_X1 U18917 ( .A(n15919), .ZN(n18889) );
  OAI22_X1 U18918 ( .A1(n15920), .A2(n15976), .B1(n15406), .B2(n18889), .ZN(
        n15921) );
  NOR2_X1 U18919 ( .A1(n15922), .A2(n15921), .ZN(n15923) );
  OAI211_X1 U18920 ( .C1(n15997), .C2(n15925), .A(n15924), .B(n15923), .ZN(
        P2_U2998) );
  AOI22_X1 U18921 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19038), .B1(n19037), 
        .B2(n15926), .ZN(n15932) );
  OAI22_X1 U18922 ( .A1(n15928), .A2(n15976), .B1(n15977), .B2(n15927), .ZN(
        n15929) );
  AOI21_X1 U18923 ( .B1(n19042), .B2(n15930), .A(n15929), .ZN(n15931) );
  OAI211_X1 U18924 ( .C1(n19047), .C2(n15933), .A(n15932), .B(n15931), .ZN(
        P2_U2999) );
  AOI22_X1 U18925 ( .A1(n15984), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19038), .ZN(n15945) );
  AOI21_X1 U18926 ( .B1(n15936), .B2(n15935), .A(n15934), .ZN(n16001) );
  INV_X1 U18927 ( .A(n15937), .ZN(n15938) );
  NOR2_X1 U18928 ( .A1(n15939), .A2(n15938), .ZN(n15943) );
  NAND2_X1 U18929 ( .A1(n15941), .A2(n15940), .ZN(n15942) );
  XNOR2_X1 U18930 ( .A(n15943), .B(n15942), .ZN(n16000) );
  AOI222_X1 U18931 ( .A1(n16001), .A2(n13164), .B1(n19040), .B2(n16000), .C1(
        n19042), .C2(n15999), .ZN(n15944) );
  OAI211_X1 U18932 ( .C1(n15997), .C2(n15946), .A(n15945), .B(n15944), .ZN(
        P2_U3000) );
  AOI22_X1 U18933 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19038), .B1(n19037), 
        .B2(n15947), .ZN(n15952) );
  OAI22_X1 U18934 ( .A1(n15949), .A2(n15976), .B1(n15948), .B2(n15977), .ZN(
        n15950) );
  AOI21_X1 U18935 ( .B1(n19042), .B2(n20957), .A(n15950), .ZN(n15951) );
  OAI211_X1 U18936 ( .C1(n19047), .C2(n15953), .A(n15952), .B(n15951), .ZN(
        P2_U3001) );
  AOI22_X1 U18937 ( .A1(n15984), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19038), .ZN(n15960) );
  NOR2_X1 U18938 ( .A1(n15977), .A2(n15954), .ZN(n15957) );
  OAI22_X1 U18939 ( .A1(n15955), .A2(n15976), .B1(n15406), .B2(n18902), .ZN(
        n15956) );
  AOI21_X1 U18940 ( .B1(n15958), .B2(n15957), .A(n15956), .ZN(n15959) );
  OAI211_X1 U18941 ( .C1(n15997), .C2(n18813), .A(n15960), .B(n15959), .ZN(
        P2_U3002) );
  AOI22_X1 U18942 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19038), .B1(n19037), 
        .B2(n15961), .ZN(n15967) );
  OAI22_X1 U18943 ( .A1(n15963), .A2(n15977), .B1(n15962), .B2(n15976), .ZN(
        n15964) );
  AOI21_X1 U18944 ( .B1(n19042), .B2(n15965), .A(n15964), .ZN(n15966) );
  OAI211_X1 U18945 ( .C1(n19047), .C2(n18820), .A(n15967), .B(n15966), .ZN(
        P2_U3003) );
  AOI22_X1 U18946 ( .A1(n15984), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19038), .ZN(n15972) );
  INV_X1 U18947 ( .A(n15968), .ZN(n15970) );
  AOI222_X1 U18948 ( .A1(n15970), .A2(n19040), .B1(n19042), .B2(n18907), .C1(
        n13164), .C2(n15969), .ZN(n15971) );
  OAI211_X1 U18949 ( .C1(n15997), .C2(n15973), .A(n15972), .B(n15971), .ZN(
        P2_U3004) );
  AOI22_X1 U18950 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19038), .B1(n19037), 
        .B2(n15974), .ZN(n15982) );
  OAI22_X1 U18951 ( .A1(n15978), .A2(n15977), .B1(n15976), .B2(n15975), .ZN(
        n15979) );
  AOI21_X1 U18952 ( .B1(n19042), .B2(n15980), .A(n15979), .ZN(n15981) );
  OAI211_X1 U18953 ( .C1(n19047), .C2(n15983), .A(n15982), .B(n15981), .ZN(
        P2_U3005) );
  AOI22_X1 U18954 ( .A1(n15984), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19038), .ZN(n15995) );
  AOI21_X1 U18955 ( .B1(n15076), .B2(n15986), .A(n15985), .ZN(n15991) );
  INV_X1 U18956 ( .A(n15987), .ZN(n15988) );
  NOR2_X1 U18957 ( .A1(n15989), .A2(n15988), .ZN(n15990) );
  XNOR2_X1 U18958 ( .A(n15991), .B(n15990), .ZN(n16016) );
  XOR2_X1 U18959 ( .A(n15992), .B(n15993), .Z(n16012) );
  AOI222_X1 U18960 ( .A1(n16016), .A2(n19040), .B1(n19042), .B2(n16013), .C1(
        n16012), .C2(n13164), .ZN(n15994) );
  OAI211_X1 U18961 ( .C1(n15997), .C2(n15996), .A(n15995), .B(n15994), .ZN(
        P2_U3006) );
  AOI22_X1 U18962 ( .A1(n15998), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n16010), .B2(n18938), .ZN(n16008) );
  AOI222_X1 U18963 ( .A1(n16001), .A2(n16011), .B1(n16015), .B2(n16000), .C1(
        n16014), .C2(n15999), .ZN(n16007) );
  NAND2_X1 U18964 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n19038), .ZN(n16006) );
  OAI211_X1 U18965 ( .C1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n16004), .A(
        n16003), .B(n16002), .ZN(n16005) );
  NAND4_X1 U18966 ( .A1(n16008), .A2(n16007), .A3(n16006), .A4(n16005), .ZN(
        P2_U3032) );
  AOI21_X1 U18967 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16009), .A(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16019) );
  AOI22_X1 U18968 ( .A1(n16010), .A2(n18952), .B1(n19038), .B2(
        P2_REIP_REG_8__SCAN_IN), .ZN(n16018) );
  AOI222_X1 U18969 ( .A1(n16016), .A2(n16015), .B1(n16014), .B2(n16013), .C1(
        n16012), .C2(n16011), .ZN(n16017) );
  OAI211_X1 U18970 ( .C1(n16020), .C2(n16019), .A(n16018), .B(n16017), .ZN(
        P2_U3038) );
  INV_X1 U18971 ( .A(n16054), .ZN(n16028) );
  AOI22_X1 U18972 ( .A1(n16054), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n16029), .B2(n16028), .ZN(n16056) );
  INV_X1 U18973 ( .A(n16056), .ZN(n16033) );
  MUX2_X1 U18974 ( .A(n16022), .B(n16021), .S(n16028), .Z(n16057) );
  OR2_X1 U18975 ( .A1(n16057), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n16031) );
  INV_X1 U18976 ( .A(n16024), .ZN(n16026) );
  OAI22_X1 U18977 ( .A1(n16024), .A2(n19788), .B1(n19797), .B2(n16023), .ZN(
        n16025) );
  OAI21_X1 U18978 ( .B1(n16026), .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n16025), .ZN(n16027) );
  OAI211_X1 U18979 ( .C1(n19769), .C2(n16029), .A(n16028), .B(n16027), .ZN(
        n16030) );
  AOI222_X1 U18980 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n16031), 
        .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16030), .C1(n16031), 
        .C2(n16030), .ZN(n16032) );
  AOI21_X1 U18981 ( .B1(n19769), .B2(n16033), .A(n16032), .ZN(n16034) );
  OR2_X1 U18982 ( .A1(n16034), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n16060) );
  NAND2_X1 U18983 ( .A1(n16036), .A2(n16035), .ZN(n16040) );
  INV_X1 U18984 ( .A(n16037), .ZN(n16038) );
  NAND2_X1 U18985 ( .A1(n16038), .A2(n16041), .ZN(n16039) );
  OAI211_X1 U18986 ( .C1(n16042), .C2(n16041), .A(n16040), .B(n16039), .ZN(
        n19803) );
  NOR2_X1 U18987 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(P2_MORE_REG_SCAN_IN), .ZN(
        n16050) );
  NAND2_X1 U18988 ( .A1(n16044), .A2(n16043), .ZN(n16046) );
  OAI22_X1 U18989 ( .A1(n16047), .A2(n16046), .B1(n16045), .B2(n19805), .ZN(
        n16048) );
  INV_X1 U18990 ( .A(n16048), .ZN(n16049) );
  OAI21_X1 U18991 ( .B1(n16051), .B2(n16050), .A(n16049), .ZN(n16052) );
  OR2_X1 U18992 ( .A1(n19803), .A2(n16052), .ZN(n16053) );
  AOI21_X1 U18993 ( .B1(n16054), .B2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n16053), .ZN(n16055) );
  OAI21_X1 U18994 ( .B1(n16057), .B2(n16056), .A(n16055), .ZN(n16058) );
  INV_X1 U18995 ( .A(n16058), .ZN(n16059) );
  AND2_X1 U18996 ( .A1(n16060), .A2(n16059), .ZN(n16077) );
  AOI211_X1 U18997 ( .C1(n16064), .C2(n16063), .A(n16062), .B(n16061), .ZN(
        n16075) );
  NAND2_X1 U18998 ( .A1(n16077), .A2(n19668), .ZN(n16069) );
  NAND3_X1 U18999 ( .A1(n10538), .A2(n19801), .A3(n16065), .ZN(n16067) );
  NAND3_X1 U19000 ( .A1(n16067), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n16066), 
        .ZN(n16068) );
  AOI21_X1 U19001 ( .B1(n16069), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16068), 
        .ZN(n19667) );
  OAI21_X1 U19002 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16071), .A(n16070), 
        .ZN(n16073) );
  NAND2_X1 U19003 ( .A1(n19667), .A2(n19690), .ZN(n16072) );
  AOI22_X1 U19004 ( .A1(n19667), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n16073), 
        .B2(n16072), .ZN(n16074) );
  OAI211_X1 U19005 ( .C1(n16077), .C2(n16076), .A(n16075), .B(n16074), .ZN(
        P2_U3176) );
  NOR2_X1 U19006 ( .A1(n16078), .A2(n19667), .ZN(n19674) );
  OAI21_X1 U19007 ( .B1(n19674), .B2(n19611), .A(n16079), .ZN(P2_U3593) );
  INV_X1 U19008 ( .A(n18492), .ZN(n16081) );
  INV_X1 U19009 ( .A(n16083), .ZN(n16098) );
  INV_X1 U19010 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16119) );
  INV_X1 U19011 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17683) );
  INV_X1 U19012 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17670) );
  NOR2_X2 U19013 ( .A1(n17683), .A2(n17670), .ZN(n17642) );
  NAND3_X1 U19014 ( .A1(n17642), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17628) );
  INV_X1 U19015 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17617) );
  NAND4_X1 U19016 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16473) );
  INV_X1 U19017 ( .A(n16473), .ZN(n16084) );
  INV_X1 U19018 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17546) );
  INV_X1 U19019 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17532) );
  NOR2_X1 U19020 ( .A1(n17546), .A2(n17532), .ZN(n17528) );
  NAND2_X1 U19021 ( .A1(n17528), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17493) );
  NAND3_X1 U19022 ( .A1(n17489), .A2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17479) );
  INV_X1 U19023 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17478) );
  NAND3_X1 U19024 ( .A1(n16279), .A2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17444) );
  INV_X1 U19025 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17443) );
  NAND2_X1 U19026 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17397) );
  INV_X1 U19027 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16369) );
  NAND2_X1 U19028 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17371) );
  INV_X1 U19029 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16085) );
  NAND2_X1 U19030 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17331), .ZN(
        n16118) );
  INV_X1 U19031 ( .A(n16089), .ZN(n16087) );
  NOR2_X2 U19032 ( .A1(n18084), .A2(n18296), .ZN(n18434) );
  NOR2_X1 U19033 ( .A1(n16087), .A2(n17527), .ZN(n16104) );
  INV_X1 U19034 ( .A(n16104), .ZN(n16088) );
  INV_X1 U19035 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17692) );
  NOR2_X1 U19036 ( .A1(n17692), .A2(n17329), .ZN(n16271) );
  NAND2_X1 U19037 ( .A1(n16271), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16270) );
  INV_X1 U19038 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17330) );
  NOR2_X1 U19039 ( .A1(n16270), .A2(n17330), .ZN(n16269) );
  NOR2_X1 U19040 ( .A1(n16269), .A2(n18564), .ZN(n16086) );
  AOI211_X1 U19041 ( .C1(n18434), .C2(n16087), .A(n17601), .B(n16086), .ZN(
        n16117) );
  NAND2_X1 U19042 ( .A1(n17445), .A2(n16119), .ZN(n16116) );
  OAI211_X1 U19043 ( .C1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .C2(n16088), .A(
        n16117), .B(n16116), .ZN(n16105) );
  NAND2_X1 U19044 ( .A1(n16105), .A2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16095) );
  INV_X1 U19045 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16090) );
  NAND2_X1 U19046 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16089), .ZN(
        n16115) );
  INV_X1 U19047 ( .A(n16115), .ZN(n16102) );
  NAND2_X1 U19048 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16102), .ZN(
        n16101) );
  XOR2_X1 U19049 ( .A(n16090), .B(n16101), .Z(n16268) );
  NAND2_X1 U19050 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n17815), .ZN(n16092) );
  NAND3_X1 U19051 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16104), .A3(
        n16090), .ZN(n16091) );
  OAI211_X1 U19052 ( .C1(n17506), .C2(n16587), .A(n16092), .B(n16091), .ZN(
        n16093) );
  AOI21_X1 U19053 ( .B1(n16098), .B2(n17538), .A(n16097), .ZN(n16099) );
  OAI21_X1 U19054 ( .B1(n16100), .B2(n17568), .A(n16099), .ZN(P3_U2799) );
  INV_X1 U19055 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18642) );
  OAI21_X1 U19056 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16102), .A(
        n16101), .ZN(n16301) );
  OAI22_X1 U19057 ( .A1(n18017), .A2(n18642), .B1(n17506), .B2(n16301), .ZN(
        n16103) );
  AOI221_X1 U19058 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16105), .C1(
        n16104), .C2(n16105), .A(n16103), .ZN(n16110) );
  OAI22_X1 U19059 ( .A1(n16125), .A2(n17568), .B1(n16114), .B2(n17700), .ZN(
        n16108) );
  AOI22_X1 U19060 ( .A1(n17567), .A2(n17685), .B1(n17608), .B2(n10902), .ZN(
        n17566) );
  NOR2_X2 U19061 ( .A1(n16106), .A2(n17566), .ZN(n17483) );
  AND2_X1 U19062 ( .A1(n17708), .A2(n17483), .ZN(n17349) );
  AOI22_X1 U19063 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16108), .B1(
        n16107), .B2(n17349), .ZN(n16109) );
  OAI211_X1 U19064 ( .C1(n16111), .C2(n17611), .A(n16110), .B(n16109), .ZN(
        P3_U2800) );
  INV_X1 U19065 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18637) );
  NOR2_X1 U19066 ( .A1(n17909), .A2(n18637), .ZN(n16123) );
  NAND2_X1 U19067 ( .A1(n16113), .A2(n16112), .ZN(n16134) );
  AOI211_X1 U19068 ( .C1(n20920), .C2(n16134), .A(n16114), .B(n17700), .ZN(
        n16122) );
  OAI21_X1 U19069 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16269), .A(
        n16115), .ZN(n16314) );
  AOI21_X1 U19070 ( .B1(n16116), .B2(n17506), .A(n16314), .ZN(n16121) );
  INV_X2 U19071 ( .A(n18434), .ZN(n18262) );
  AOI221_X1 U19072 ( .B1(n18262), .B2(n16119), .C1(n16118), .C2(n16119), .A(
        n16117), .ZN(n16120) );
  NOR4_X1 U19073 ( .A1(n16123), .A2(n16122), .A3(n16121), .A4(n16120), .ZN(
        n16128) );
  NOR2_X1 U19074 ( .A1(n16124), .A2(n17702), .ZN(n16132) );
  NOR2_X1 U19075 ( .A1(n16125), .A2(n17568), .ZN(n16126) );
  OAI21_X1 U19076 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16132), .A(
        n16126), .ZN(n16127) );
  OAI211_X1 U19077 ( .C1(n16129), .C2(n17611), .A(n16128), .B(n16127), .ZN(
        P3_U2801) );
  INV_X1 U19078 ( .A(n10902), .ZN(n17932) );
  OAI22_X1 U19079 ( .A1(n17999), .A2(n17891), .B1(n17835), .B2(n17932), .ZN(
        n17803) );
  AOI21_X1 U19080 ( .B1(n17803), .B2(n17804), .A(n17722), .ZN(n17701) );
  INV_X1 U19081 ( .A(n17769), .ZN(n17794) );
  NAND2_X1 U19082 ( .A1(n16130), .A2(n10916), .ZN(n17340) );
  INV_X1 U19083 ( .A(n17341), .ZN(n16140) );
  OAI21_X1 U19084 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17557), .A(
        n16131), .ZN(n17325) );
  NOR2_X1 U19085 ( .A1(n17326), .A2(n17325), .ZN(n17324) );
  AOI211_X1 U19086 ( .C1(n16141), .C2(n16140), .A(n17324), .B(n17844), .ZN(
        n16138) );
  OR2_X1 U19087 ( .A1(n16132), .A2(n17835), .ZN(n16136) );
  AOI21_X1 U19088 ( .B1(n16134), .B2(n18486), .A(n16133), .ZN(n16135) );
  NAND2_X1 U19089 ( .A1(n16136), .A2(n16135), .ZN(n16137) );
  AND2_X1 U19090 ( .A1(n17909), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16145) );
  AND3_X1 U19091 ( .A1(n17325), .A2(n16139), .A3(n17878), .ZN(n16143) );
  AND4_X1 U19092 ( .A1(n10916), .A2(n16141), .A3(n16140), .A4(n17878), .ZN(
        n16142) );
  NAND2_X1 U19093 ( .A1(n17821), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17334) );
  OAI211_X1 U19094 ( .C1(n17794), .C2(n17340), .A(n16147), .B(n17334), .ZN(
        P3_U2834) );
  NOR3_X1 U19095 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16149) );
  NOR4_X1 U19096 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16148) );
  NAND4_X1 U19097 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16149), .A3(n16148), .A4(
        U215), .ZN(U213) );
  INV_X1 U19098 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n18991) );
  NOR2_X1 U19099 ( .A1(n16199), .A2(n16150), .ZN(n16151) );
  INV_X1 U19100 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16235) );
  OAI222_X1 U19101 ( .A1(U212), .A2(n18991), .B1(n16201), .B2(n19084), .C1(
        U214), .C2(n16235), .ZN(U216) );
  AOI222_X1 U19102 ( .A1(n16199), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16151), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n16198), .C2(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n16152) );
  INV_X1 U19103 ( .A(n16152), .ZN(U217) );
  INV_X1 U19104 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16154) );
  AOI22_X1 U19105 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16198), .ZN(n16153) );
  OAI21_X1 U19106 ( .B1(n16154), .B2(n16201), .A(n16153), .ZN(U218) );
  AOI22_X1 U19107 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16198), .ZN(n16155) );
  OAI21_X1 U19108 ( .B1(n16156), .B2(n16201), .A(n16155), .ZN(U219) );
  INV_X1 U19109 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16158) );
  AOI22_X1 U19110 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16198), .ZN(n16157) );
  OAI21_X1 U19111 ( .B1(n16158), .B2(n16201), .A(n16157), .ZN(U220) );
  INV_X1 U19112 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20828) );
  AOI22_X1 U19113 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16198), .ZN(n16159) );
  OAI21_X1 U19114 ( .B1(n20828), .B2(n16201), .A(n16159), .ZN(U221) );
  INV_X1 U19115 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16161) );
  AOI22_X1 U19116 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n16198), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n16199), .ZN(n16160) );
  OAI21_X1 U19117 ( .B1(n16161), .B2(n16201), .A(n16160), .ZN(U222) );
  INV_X1 U19118 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16163) );
  AOI22_X1 U19119 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16198), .ZN(n16162) );
  OAI21_X1 U19120 ( .B1(n16163), .B2(n16201), .A(n16162), .ZN(U223) );
  AOI22_X1 U19121 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16198), .ZN(n16164) );
  OAI21_X1 U19122 ( .B1(n14437), .B2(n16201), .A(n16164), .ZN(U224) );
  AOI22_X1 U19123 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16198), .ZN(n16165) );
  OAI21_X1 U19124 ( .B1(n16166), .B2(n16201), .A(n16165), .ZN(U225) );
  AOI22_X1 U19125 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16198), .ZN(n16167) );
  OAI21_X1 U19126 ( .B1(n16168), .B2(n16201), .A(n16167), .ZN(U226) );
  AOI22_X1 U19127 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16198), .ZN(n16169) );
  OAI21_X1 U19128 ( .B1(n14454), .B2(n16201), .A(n16169), .ZN(U227) );
  AOI22_X1 U19129 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16198), .ZN(n16170) );
  OAI21_X1 U19130 ( .B1(n14458), .B2(n16201), .A(n16170), .ZN(U228) );
  AOI22_X1 U19131 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16198), .ZN(n16171) );
  OAI21_X1 U19132 ( .B1(n14462), .B2(n16201), .A(n16171), .ZN(U229) );
  AOI22_X1 U19133 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16198), .ZN(n16172) );
  OAI21_X1 U19134 ( .B1(n14468), .B2(n16201), .A(n16172), .ZN(U230) );
  AOI22_X1 U19135 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16198), .ZN(n16173) );
  OAI21_X1 U19136 ( .B1(n14055), .B2(n16201), .A(n16173), .ZN(U231) );
  INV_X1 U19137 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n16175) );
  AOI22_X1 U19138 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16198), .ZN(n16174) );
  OAI21_X1 U19139 ( .B1(n16175), .B2(n16201), .A(n16174), .ZN(U232) );
  AOI22_X1 U19140 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16198), .ZN(n16176) );
  OAI21_X1 U19141 ( .B1(n14004), .B2(n16201), .A(n16176), .ZN(U233) );
  AOI22_X1 U19142 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16198), .ZN(n16177) );
  OAI21_X1 U19143 ( .B1(n13996), .B2(n16201), .A(n16177), .ZN(U234) );
  AOI22_X1 U19144 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16198), .ZN(n16178) );
  OAI21_X1 U19145 ( .B1(n13332), .B2(n16201), .A(n16178), .ZN(U235) );
  AOI22_X1 U19146 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16198), .ZN(n16179) );
  OAI21_X1 U19147 ( .B1(n14009), .B2(n16201), .A(n16179), .ZN(U236) );
  AOI22_X1 U19148 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16198), .ZN(n16180) );
  OAI21_X1 U19149 ( .B1(n16181), .B2(n16201), .A(n16180), .ZN(U237) );
  AOI22_X1 U19150 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16198), .ZN(n16182) );
  OAI21_X1 U19151 ( .B1(n13221), .B2(n16201), .A(n16182), .ZN(U238) );
  AOI22_X1 U19152 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16198), .ZN(n16183) );
  OAI21_X1 U19153 ( .B1(n13901), .B2(n16201), .A(n16183), .ZN(U239) );
  INV_X1 U19154 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16185) );
  AOI22_X1 U19155 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16198), .ZN(n16184) );
  OAI21_X1 U19156 ( .B1(n16185), .B2(n16201), .A(n16184), .ZN(U240) );
  INV_X1 U19157 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16187) );
  AOI22_X1 U19158 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16198), .ZN(n16186) );
  OAI21_X1 U19159 ( .B1(n16187), .B2(n16201), .A(n16186), .ZN(U241) );
  INV_X1 U19160 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16189) );
  AOI22_X1 U19161 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16198), .ZN(n16188) );
  OAI21_X1 U19162 ( .B1(n16189), .B2(n16201), .A(n16188), .ZN(U242) );
  AOI22_X1 U19163 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16198), .ZN(n16190) );
  OAI21_X1 U19164 ( .B1(n16191), .B2(n16201), .A(n16190), .ZN(U243) );
  INV_X1 U19165 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16193) );
  AOI22_X1 U19166 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16198), .ZN(n16192) );
  OAI21_X1 U19167 ( .B1(n16193), .B2(n16201), .A(n16192), .ZN(U244) );
  INV_X1 U19168 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16195) );
  AOI22_X1 U19169 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16198), .ZN(n16194) );
  OAI21_X1 U19170 ( .B1(n16195), .B2(n16201), .A(n16194), .ZN(U245) );
  INV_X1 U19171 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16197) );
  AOI22_X1 U19172 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16198), .ZN(n16196) );
  OAI21_X1 U19173 ( .B1(n16197), .B2(n16201), .A(n16196), .ZN(U246) );
  INV_X1 U19174 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16202) );
  AOI22_X1 U19175 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16199), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16198), .ZN(n16200) );
  OAI21_X1 U19176 ( .B1(n16202), .B2(n16201), .A(n16200), .ZN(U247) );
  OAI22_X1 U19177 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16234), .ZN(n16203) );
  INV_X1 U19178 ( .A(n16203), .ZN(U251) );
  OAI22_X1 U19179 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16234), .ZN(n16204) );
  INV_X1 U19180 ( .A(n16204), .ZN(U252) );
  OAI22_X1 U19181 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16234), .ZN(n16205) );
  INV_X1 U19182 ( .A(n16205), .ZN(U253) );
  OAI22_X1 U19183 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16234), .ZN(n16206) );
  INV_X1 U19184 ( .A(n16206), .ZN(U254) );
  OAI22_X1 U19185 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16234), .ZN(n16207) );
  INV_X1 U19186 ( .A(n16207), .ZN(U255) );
  OAI22_X1 U19187 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16234), .ZN(n16208) );
  INV_X1 U19188 ( .A(n16208), .ZN(U256) );
  OAI22_X1 U19189 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16234), .ZN(n16209) );
  INV_X1 U19190 ( .A(n16209), .ZN(U257) );
  OAI22_X1 U19191 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16234), .ZN(n16210) );
  INV_X1 U19192 ( .A(n16210), .ZN(U258) );
  OAI22_X1 U19193 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16234), .ZN(n16211) );
  INV_X1 U19194 ( .A(n16211), .ZN(U259) );
  OAI22_X1 U19195 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16226), .ZN(n16212) );
  INV_X1 U19196 ( .A(n16212), .ZN(U260) );
  OAI22_X1 U19197 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16226), .ZN(n16213) );
  INV_X1 U19198 ( .A(n16213), .ZN(U261) );
  OAI22_X1 U19199 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16234), .ZN(n16214) );
  INV_X1 U19200 ( .A(n16214), .ZN(U262) );
  OAI22_X1 U19201 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16226), .ZN(n16215) );
  INV_X1 U19202 ( .A(n16215), .ZN(U263) );
  OAI22_X1 U19203 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16234), .ZN(n16216) );
  INV_X1 U19204 ( .A(n16216), .ZN(U264) );
  OAI22_X1 U19205 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16234), .ZN(n16217) );
  INV_X1 U19206 ( .A(n16217), .ZN(U265) );
  OAI22_X1 U19207 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16226), .ZN(n16218) );
  INV_X1 U19208 ( .A(n16218), .ZN(U266) );
  OAI22_X1 U19209 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16226), .ZN(n16219) );
  INV_X1 U19210 ( .A(n16219), .ZN(U267) );
  OAI22_X1 U19211 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16226), .ZN(n16220) );
  INV_X1 U19212 ( .A(n16220), .ZN(U268) );
  OAI22_X1 U19213 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16226), .ZN(n16221) );
  INV_X1 U19214 ( .A(n16221), .ZN(U269) );
  OAI22_X1 U19215 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16226), .ZN(n16222) );
  INV_X1 U19216 ( .A(n16222), .ZN(U270) );
  OAI22_X1 U19217 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16226), .ZN(n16223) );
  INV_X1 U19218 ( .A(n16223), .ZN(U271) );
  OAI22_X1 U19219 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16234), .ZN(n16224) );
  INV_X1 U19220 ( .A(n16224), .ZN(U272) );
  OAI22_X1 U19221 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16234), .ZN(n16225) );
  INV_X1 U19222 ( .A(n16225), .ZN(U273) );
  OAI22_X1 U19223 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16226), .ZN(n16227) );
  INV_X1 U19224 ( .A(n16227), .ZN(U274) );
  OAI22_X1 U19225 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16234), .ZN(n16228) );
  INV_X1 U19226 ( .A(n16228), .ZN(U275) );
  OAI22_X1 U19227 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16234), .ZN(n16229) );
  INV_X1 U19228 ( .A(n16229), .ZN(U276) );
  OAI22_X1 U19229 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16234), .ZN(n16230) );
  INV_X1 U19230 ( .A(n16230), .ZN(U277) );
  OAI22_X1 U19231 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16234), .ZN(n16231) );
  INV_X1 U19232 ( .A(n16231), .ZN(U278) );
  OAI22_X1 U19233 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16234), .ZN(n16232) );
  INV_X1 U19234 ( .A(n16232), .ZN(U279) );
  OAI22_X1 U19235 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16234), .ZN(n16233) );
  INV_X1 U19236 ( .A(n16233), .ZN(U280) );
  INV_X1 U19237 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n20866) );
  INV_X1 U19238 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18070) );
  AOI22_X1 U19239 ( .A1(n16234), .A2(n20866), .B1(n18070), .B2(U215), .ZN(U281) );
  INV_X1 U19240 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19083) );
  AOI22_X1 U19241 ( .A1(n16234), .A2(n18991), .B1(n19083), .B2(U215), .ZN(U282) );
  INV_X1 U19242 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16236) );
  AOI222_X1 U19243 ( .A1(n16236), .A2(P3_DATAO_REG_30__SCAN_IN), .B1(n18991), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16235), .C2(
        P1_DATAO_REG_30__SCAN_IN), .ZN(n16237) );
  INV_X1 U19244 ( .A(n16239), .ZN(n16238) );
  INV_X1 U19245 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18600) );
  INV_X1 U19246 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19713) );
  AOI22_X1 U19247 ( .A1(n16238), .A2(n18600), .B1(n19713), .B2(n16239), .ZN(
        U347) );
  INV_X1 U19248 ( .A(n16239), .ZN(n16240) );
  INV_X1 U19249 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18597) );
  INV_X1 U19250 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19711) );
  AOI22_X1 U19251 ( .A1(n16240), .A2(n18597), .B1(n19711), .B2(n16239), .ZN(
        U348) );
  INV_X1 U19252 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18596) );
  INV_X1 U19253 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19710) );
  AOI22_X1 U19254 ( .A1(n16238), .A2(n18596), .B1(n19710), .B2(n16239), .ZN(
        U349) );
  INV_X1 U19255 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18594) );
  INV_X1 U19256 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19708) );
  AOI22_X1 U19257 ( .A1(n16238), .A2(n18594), .B1(n19708), .B2(n16239), .ZN(
        U350) );
  INV_X1 U19258 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18592) );
  INV_X1 U19259 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19706) );
  AOI22_X1 U19260 ( .A1(n16238), .A2(n18592), .B1(n19706), .B2(n16239), .ZN(
        U351) );
  INV_X1 U19261 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18589) );
  INV_X1 U19262 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19705) );
  AOI22_X1 U19263 ( .A1(n16238), .A2(n18589), .B1(n19705), .B2(n16239), .ZN(
        U352) );
  INV_X1 U19264 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18588) );
  INV_X1 U19265 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19704) );
  AOI22_X1 U19266 ( .A1(n16240), .A2(n18588), .B1(n19704), .B2(n16239), .ZN(
        U353) );
  INV_X1 U19267 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18585) );
  AOI22_X1 U19268 ( .A1(n16238), .A2(n18585), .B1(n19703), .B2(n16239), .ZN(
        U354) );
  INV_X1 U19269 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18641) );
  INV_X1 U19270 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19747) );
  AOI22_X1 U19271 ( .A1(n16238), .A2(n18641), .B1(n19747), .B2(n16239), .ZN(
        U355) );
  INV_X1 U19272 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18638) );
  INV_X1 U19273 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19745) );
  AOI22_X1 U19274 ( .A1(n16238), .A2(n18638), .B1(n19745), .B2(n16239), .ZN(
        U356) );
  INV_X1 U19275 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18635) );
  INV_X1 U19276 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19741) );
  AOI22_X1 U19277 ( .A1(n16238), .A2(n18635), .B1(n19741), .B2(n16239), .ZN(
        U357) );
  INV_X1 U19278 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18634) );
  INV_X1 U19279 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19738) );
  AOI22_X1 U19280 ( .A1(n16238), .A2(n18634), .B1(n19738), .B2(n16239), .ZN(
        U358) );
  INV_X1 U19281 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18632) );
  INV_X1 U19282 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19737) );
  AOI22_X1 U19283 ( .A1(n16238), .A2(n18632), .B1(n19737), .B2(n16239), .ZN(
        U359) );
  INV_X1 U19284 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18630) );
  INV_X1 U19285 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19736) );
  AOI22_X1 U19286 ( .A1(n16238), .A2(n18630), .B1(n19736), .B2(n16239), .ZN(
        U360) );
  INV_X1 U19287 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18628) );
  INV_X1 U19288 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19734) );
  AOI22_X1 U19289 ( .A1(n16238), .A2(n18628), .B1(n19734), .B2(n16239), .ZN(
        U361) );
  INV_X1 U19290 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18625) );
  INV_X1 U19291 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19732) );
  AOI22_X1 U19292 ( .A1(n16238), .A2(n18625), .B1(n19732), .B2(n16239), .ZN(
        U362) );
  INV_X1 U19293 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18624) );
  INV_X1 U19294 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19730) );
  AOI22_X1 U19295 ( .A1(n16238), .A2(n18624), .B1(n19730), .B2(n16239), .ZN(
        U363) );
  INV_X1 U19296 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18621) );
  INV_X1 U19297 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20924) );
  AOI22_X1 U19298 ( .A1(n16238), .A2(n18621), .B1(n20924), .B2(n16239), .ZN(
        U364) );
  INV_X1 U19299 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18583) );
  INV_X1 U19300 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19702) );
  AOI22_X1 U19301 ( .A1(n16238), .A2(n18583), .B1(n19702), .B2(n16239), .ZN(
        U365) );
  INV_X1 U19302 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18620) );
  INV_X1 U19303 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19727) );
  AOI22_X1 U19304 ( .A1(n16238), .A2(n18620), .B1(n19727), .B2(n16239), .ZN(
        U366) );
  INV_X1 U19305 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18617) );
  INV_X1 U19306 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19726) );
  AOI22_X1 U19307 ( .A1(n16238), .A2(n18617), .B1(n19726), .B2(n16239), .ZN(
        U367) );
  INV_X1 U19308 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18616) );
  INV_X1 U19309 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19724) );
  AOI22_X1 U19310 ( .A1(n16238), .A2(n18616), .B1(n19724), .B2(n16239), .ZN(
        U368) );
  INV_X1 U19311 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18613) );
  INV_X1 U19312 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19722) );
  AOI22_X1 U19313 ( .A1(n16238), .A2(n18613), .B1(n19722), .B2(n16239), .ZN(
        U369) );
  INV_X1 U19314 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18612) );
  INV_X1 U19315 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19720) );
  AOI22_X1 U19316 ( .A1(n16238), .A2(n18612), .B1(n19720), .B2(n16239), .ZN(
        U370) );
  INV_X1 U19317 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18610) );
  INV_X1 U19318 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19718) );
  AOI22_X1 U19319 ( .A1(n16240), .A2(n18610), .B1(n19718), .B2(n16239), .ZN(
        U371) );
  INV_X1 U19320 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18607) );
  INV_X1 U19321 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20832) );
  AOI22_X1 U19322 ( .A1(n16240), .A2(n18607), .B1(n20832), .B2(n16239), .ZN(
        U372) );
  INV_X1 U19323 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18606) );
  INV_X1 U19324 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20921) );
  AOI22_X1 U19325 ( .A1(n16240), .A2(n18606), .B1(n20921), .B2(n16239), .ZN(
        U373) );
  INV_X1 U19326 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18604) );
  INV_X1 U19327 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20831) );
  AOI22_X1 U19328 ( .A1(n16240), .A2(n18604), .B1(n20831), .B2(n16239), .ZN(
        U374) );
  INV_X1 U19329 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18602) );
  INV_X1 U19330 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19714) );
  AOI22_X1 U19331 ( .A1(n16240), .A2(n18602), .B1(n19714), .B2(n16239), .ZN(
        U375) );
  INV_X1 U19332 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18581) );
  INV_X1 U19333 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19700) );
  AOI22_X1 U19334 ( .A1(n16240), .A2(n18581), .B1(n19700), .B2(n16239), .ZN(
        U376) );
  INV_X1 U19335 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18580) );
  NAND2_X1 U19336 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18580), .ZN(n18569) );
  AOI22_X1 U19337 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18569), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18578), .ZN(n18650) );
  AOI21_X1 U19338 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18650), .ZN(n16241) );
  INV_X1 U19339 ( .A(n16241), .ZN(P3_U2633) );
  NAND2_X1 U19340 ( .A1(n18715), .A2(n18653), .ZN(n16244) );
  OAI21_X1 U19341 ( .B1(n16242), .B2(n17270), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16243) );
  OAI21_X1 U19342 ( .B1(n16244), .B2(n16284), .A(n16243), .ZN(P3_U2634) );
  AOI21_X1 U19343 ( .B1(n18578), .B2(n18580), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16245) );
  AOI22_X1 U19344 ( .A1(n18712), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16245), 
        .B2(n18713), .ZN(P3_U2635) );
  OAI21_X1 U19345 ( .B1(n18566), .B2(BS16), .A(n18650), .ZN(n18648) );
  OAI21_X1 U19346 ( .B1(n18650), .B2(n16281), .A(n18648), .ZN(P3_U2636) );
  AND3_X1 U19347 ( .A1(n16247), .A2(n18488), .A3(n16246), .ZN(n18493) );
  NOR2_X1 U19348 ( .A1(n18493), .A2(n18552), .ZN(n18695) );
  OAI21_X1 U19349 ( .B1(n18695), .B2(n16249), .A(n16248), .ZN(P3_U2637) );
  NOR4_X1 U19350 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16253) );
  NOR4_X1 U19351 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16252) );
  NOR4_X1 U19352 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16251) );
  NOR4_X1 U19353 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16250) );
  NAND4_X1 U19354 ( .A1(n16253), .A2(n16252), .A3(n16251), .A4(n16250), .ZN(
        n16259) );
  NOR4_X1 U19355 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16257) );
  AOI211_X1 U19356 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_16__SCAN_IN), .B(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16256) );
  NOR4_X1 U19357 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16255) );
  NOR4_X1 U19358 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16254) );
  NAND4_X1 U19359 ( .A1(n16257), .A2(n16256), .A3(n16255), .A4(n16254), .ZN(
        n16258) );
  NOR2_X1 U19360 ( .A1(n16259), .A2(n16258), .ZN(n18689) );
  INV_X1 U19361 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16261) );
  NOR3_X1 U19362 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16262) );
  OAI21_X1 U19363 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16262), .A(n18689), .ZN(
        n16260) );
  OAI21_X1 U19364 ( .B1(n18689), .B2(n16261), .A(n16260), .ZN(P3_U2638) );
  INV_X1 U19365 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18685) );
  INV_X1 U19366 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18649) );
  AOI21_X1 U19367 ( .B1(n18685), .B2(n18649), .A(n16262), .ZN(n16264) );
  INV_X1 U19368 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16263) );
  INV_X1 U19369 ( .A(n18689), .ZN(n18692) );
  AOI22_X1 U19370 ( .A1(n18689), .A2(n16264), .B1(n16263), .B2(n18692), .ZN(
        P3_U2639) );
  NAND2_X1 U19371 ( .A1(n16266), .A2(n18718), .ZN(n16282) );
  INV_X1 U19372 ( .A(n16282), .ZN(n16287) );
  NAND2_X1 U19373 ( .A1(n18697), .A2(n16281), .ZN(n16267) );
  INV_X1 U19374 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17051) );
  NAND2_X1 U19375 ( .A1(n20934), .A2(n17051), .ZN(n16644) );
  NOR2_X1 U19376 ( .A1(n16644), .A2(P3_EBX_REG_2__SCAN_IN), .ZN(n16628) );
  INV_X1 U19377 ( .A(n16628), .ZN(n16615) );
  NOR2_X1 U19378 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n16615), .ZN(n16614) );
  NAND2_X1 U19379 ( .A1(n16614), .A2(n17037), .ZN(n16599) );
  NOR2_X1 U19380 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n16599), .ZN(n16590) );
  NAND2_X1 U19381 ( .A1(n16590), .A2(n20863), .ZN(n16581) );
  NOR2_X1 U19382 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n16581), .ZN(n16563) );
  INV_X1 U19383 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n16554) );
  NAND2_X1 U19384 ( .A1(n16563), .A2(n16554), .ZN(n16553) );
  NOR2_X1 U19385 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n16553), .ZN(n16531) );
  INV_X1 U19386 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n16527) );
  NAND2_X1 U19387 ( .A1(n16531), .A2(n16527), .ZN(n16526) );
  NOR2_X1 U19388 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n16526), .ZN(n16507) );
  INV_X1 U19389 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n16504) );
  NAND2_X1 U19390 ( .A1(n16507), .A2(n16504), .ZN(n16503) );
  NOR2_X1 U19391 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n16503), .ZN(n16490) );
  INV_X1 U19392 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n16479) );
  NAND2_X1 U19393 ( .A1(n16490), .A2(n16479), .ZN(n16478) );
  NOR2_X1 U19394 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n16478), .ZN(n16461) );
  INV_X1 U19395 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n16453) );
  NAND2_X1 U19396 ( .A1(n16461), .A2(n16453), .ZN(n16451) );
  NOR2_X1 U19397 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n16451), .ZN(n16437) );
  INV_X1 U19398 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n16430) );
  NAND2_X1 U19399 ( .A1(n16437), .A2(n16430), .ZN(n16428) );
  NOR2_X1 U19400 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n16428), .ZN(n16416) );
  INV_X1 U19401 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16845) );
  NAND2_X1 U19402 ( .A1(n16416), .A2(n16845), .ZN(n16404) );
  NOR2_X1 U19403 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16404), .ZN(n16391) );
  INV_X1 U19404 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16771) );
  NAND2_X1 U19405 ( .A1(n16391), .A2(n16771), .ZN(n16386) );
  NOR2_X1 U19406 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n16386), .ZN(n16368) );
  INV_X1 U19407 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n16772) );
  NAND2_X1 U19408 ( .A1(n16368), .A2(n16772), .ZN(n16361) );
  NOR2_X1 U19409 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n16361), .ZN(n16346) );
  INV_X1 U19410 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n16773) );
  NAND2_X1 U19411 ( .A1(n16346), .A2(n16773), .ZN(n16345) );
  NOR2_X1 U19412 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16345), .ZN(n16331) );
  INV_X1 U19413 ( .A(n16331), .ZN(n16320) );
  NOR2_X1 U19414 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16321), .ZN(n16302) );
  NAND2_X1 U19415 ( .A1(n16600), .A2(n16302), .ZN(n16303) );
  INV_X1 U19416 ( .A(n9662), .ZN(n16620) );
  NOR2_X1 U19417 ( .A1(n16587), .A2(n16620), .ZN(n16643) );
  AOI21_X1 U19418 ( .B1(n16270), .B2(n17330), .A(n16269), .ZN(n17337) );
  INV_X1 U19419 ( .A(n17337), .ZN(n16325) );
  OAI21_X1 U19420 ( .B1(n16271), .B2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16270), .ZN(n17344) );
  NOR2_X1 U19421 ( .A1(n17692), .A2(n17370), .ZN(n16276) );
  INV_X1 U19422 ( .A(n16276), .ZN(n16275) );
  NOR2_X1 U19423 ( .A1(n17371), .A2(n16275), .ZN(n17327) );
  INV_X1 U19424 ( .A(n16271), .ZN(n16272) );
  OAI21_X1 U19425 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17327), .A(
        n16272), .ZN(n17353) );
  INV_X1 U19426 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17387) );
  NOR2_X1 U19427 ( .A1(n17387), .A2(n16275), .ZN(n16274) );
  INV_X1 U19428 ( .A(n17327), .ZN(n16273) );
  OAI21_X1 U19429 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16274), .A(
        n16273), .ZN(n17373) );
  AOI22_X1 U19430 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16275), .B1(
        n16276), .B2(n17387), .ZN(n17384) );
  INV_X1 U19431 ( .A(n17397), .ZN(n17412) );
  NAND2_X1 U19432 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17396), .ZN(
        n16280) );
  INV_X1 U19433 ( .A(n16280), .ZN(n16278) );
  NAND2_X1 U19434 ( .A1(n17412), .A2(n16278), .ZN(n17368) );
  AOI21_X1 U19435 ( .B1(n16369), .B2(n17368), .A(n16276), .ZN(n17402) );
  INV_X1 U19436 ( .A(n17402), .ZN(n16374) );
  INV_X1 U19437 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17430) );
  NOR2_X1 U19438 ( .A1(n17430), .A2(n16280), .ZN(n16277) );
  OAI21_X1 U19439 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n16277), .A(
        n17368), .ZN(n17416) );
  OAI22_X1 U19440 ( .A1(n17430), .A2(n16280), .B1(n16278), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17428) );
  NAND2_X1 U19441 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17457) );
  INV_X1 U19442 ( .A(n16279), .ZN(n17456) );
  NOR2_X1 U19443 ( .A1(n17692), .A2(n17456), .ZN(n17455) );
  INV_X1 U19444 ( .A(n17455), .ZN(n16435) );
  NOR2_X1 U19445 ( .A1(n17457), .A2(n16435), .ZN(n17415) );
  INV_X1 U19446 ( .A(n17415), .ZN(n16411) );
  NAND2_X1 U19447 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17489), .ZN(
        n16472) );
  INV_X1 U19448 ( .A(n16472), .ZN(n17491) );
  NAND2_X1 U19449 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17491), .ZN(
        n16460) );
  NOR2_X1 U19450 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16460), .ZN(
        n16413) );
  AOI21_X1 U19451 ( .B1(n16617), .B2(n16411), .A(n16462), .ZN(n16403) );
  OAI21_X1 U19452 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17415), .A(
        n16280), .ZN(n17446) );
  NAND2_X1 U19453 ( .A1(n16403), .A2(n17446), .ZN(n16402) );
  NAND2_X1 U19454 ( .A1(n16617), .A2(n16402), .ZN(n16396) );
  NAND2_X1 U19455 ( .A1(n17428), .A2(n16396), .ZN(n16395) );
  NAND2_X1 U19456 ( .A1(n16617), .A2(n16395), .ZN(n16385) );
  NAND2_X1 U19457 ( .A1(n17416), .A2(n16385), .ZN(n16384) );
  NAND2_X1 U19458 ( .A1(n16617), .A2(n16384), .ZN(n16373) );
  NAND2_X1 U19459 ( .A1(n16374), .A2(n16373), .ZN(n16372) );
  NAND2_X1 U19460 ( .A1(n16617), .A2(n16372), .ZN(n16363) );
  NAND2_X1 U19461 ( .A1(n17384), .A2(n16363), .ZN(n16362) );
  NAND2_X1 U19462 ( .A1(n16617), .A2(n16362), .ZN(n16355) );
  NAND2_X1 U19463 ( .A1(n17373), .A2(n16355), .ZN(n16354) );
  NAND2_X1 U19464 ( .A1(n16617), .A2(n16354), .ZN(n16344) );
  NAND2_X1 U19465 ( .A1(n17353), .A2(n16344), .ZN(n16343) );
  NAND2_X1 U19466 ( .A1(n16617), .A2(n16343), .ZN(n16337) );
  NAND2_X1 U19467 ( .A1(n17344), .A2(n16337), .ZN(n16336) );
  NAND2_X1 U19468 ( .A1(n16617), .A2(n16336), .ZN(n16324) );
  NAND2_X1 U19469 ( .A1(n16325), .A2(n16324), .ZN(n16323) );
  NAND2_X1 U19470 ( .A1(n16617), .A2(n16323), .ZN(n16313) );
  NAND2_X1 U19471 ( .A1(n16314), .A2(n16313), .ZN(n16312) );
  NAND2_X1 U19472 ( .A1(n16617), .A2(n16312), .ZN(n16300) );
  AND2_X1 U19473 ( .A1(n16301), .A2(n16300), .ZN(n16291) );
  INV_X1 U19474 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18636) );
  INV_X1 U19475 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18633) );
  NOR2_X1 U19476 ( .A1(n18636), .A2(n18633), .ZN(n16315) );
  INV_X1 U19477 ( .A(n16315), .ZN(n16326) );
  NOR2_X1 U19478 ( .A1(n18637), .A2(n16326), .ZN(n16297) );
  NAND2_X1 U19479 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .ZN(n16296) );
  NAND3_X1 U19480 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .A3(P3_REIP_REG_22__SCAN_IN), .ZN(n16295) );
  NAND3_X1 U19481 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n16294) );
  OAI211_X1 U19482 ( .C1(n18702), .C2(n18701), .A(n18697), .B(n16281), .ZN(
        n18547) );
  NOR2_X2 U19483 ( .A1(n18547), .A2(n16282), .ZN(n16630) );
  INV_X1 U19484 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18605) );
  INV_X1 U19485 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18587) );
  NAND3_X1 U19486 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16612) );
  NOR2_X1 U19487 ( .A1(n18587), .A2(n16612), .ZN(n16585) );
  NAND2_X1 U19488 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16585), .ZN(n16567) );
  NAND3_X1 U19489 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .A3(P3_REIP_REG_6__SCAN_IN), .ZN(n16518) );
  NAND3_X1 U19490 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(P3_REIP_REG_11__SCAN_IN), 
        .A3(P3_REIP_REG_10__SCAN_IN), .ZN(n16283) );
  NOR3_X1 U19491 ( .A1(n16567), .A2(n16518), .A3(n16283), .ZN(n16485) );
  NAND2_X1 U19492 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16485), .ZN(n16483) );
  OR2_X1 U19493 ( .A1(n18605), .A2(n16483), .ZN(n16293) );
  NAND4_X1 U19494 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_20__SCAN_IN), 
        .A3(P3_REIP_REG_18__SCAN_IN), .A4(n16424), .ZN(n16381) );
  NOR2_X1 U19495 ( .A1(n16295), .A2(n16381), .ZN(n16360) );
  NAND2_X1 U19496 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16360), .ZN(n16358) );
  NAND2_X1 U19497 ( .A1(n16297), .A2(n16335), .ZN(n16292) );
  NOR3_X1 U19498 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18642), .A3(n16292), 
        .ZN(n16290) );
  INV_X1 U19499 ( .A(n16284), .ZN(n18555) );
  NAND2_X1 U19500 ( .A1(n18715), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18554) );
  INV_X1 U19501 ( .A(n18554), .ZN(n18400) );
  NAND2_X1 U19502 ( .A1(n17909), .A2(n16620), .ZN(n16285) );
  NAND2_X1 U19503 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18702), .ZN(n16286) );
  NAND3_X1 U19504 ( .A1(n16287), .A2(n18547), .A3(n16286), .ZN(n16654) );
  AOI22_X1 U19505 ( .A1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n16642), .B1(
        P3_EBX_REG_31__SCAN_IN), .B2(n16613), .ZN(n16288) );
  INV_X1 U19506 ( .A(n16288), .ZN(n16289) );
  AOI211_X1 U19507 ( .C1(n16643), .C2(n16291), .A(n16290), .B(n16289), .ZN(
        n16299) );
  NOR2_X1 U19508 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16292), .ZN(n16304) );
  INV_X1 U19509 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18608) );
  NOR3_X1 U19510 ( .A1(n18608), .A2(n16293), .A3(n16649), .ZN(n16476) );
  INV_X1 U19511 ( .A(n16476), .ZN(n16446) );
  NOR2_X1 U19512 ( .A1(n16446), .A2(n16294), .ZN(n16409) );
  NAND4_X1 U19513 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n16409), .A3(
        P3_REIP_REG_20__SCAN_IN), .A4(P3_REIP_REG_18__SCAN_IN), .ZN(n16380) );
  NAND2_X1 U19514 ( .A1(n16657), .A2(n16646), .ZN(n16655) );
  OAI21_X1 U19515 ( .B1(n16380), .B2(n16295), .A(n16655), .ZN(n16377) );
  NAND2_X1 U19516 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16377), .ZN(n16359) );
  OAI21_X1 U19517 ( .B1(n16359), .B2(n16296), .A(n16655), .ZN(n16340) );
  OAI21_X1 U19518 ( .B1(n16297), .B2(n16646), .A(n16340), .ZN(n16311) );
  OAI21_X1 U19519 ( .B1(n16304), .B2(n16311), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n16298) );
  OAI211_X1 U19520 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16303), .A(n16299), .B(
        n16298), .ZN(P3_U2640) );
  XNOR2_X1 U19521 ( .A(n16301), .B(n16300), .ZN(n16308) );
  AOI22_X1 U19522 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16642), .B1(
        P3_REIP_REG_30__SCAN_IN), .B2(n16311), .ZN(n16307) );
  NOR2_X1 U19523 ( .A1(n16302), .A2(n16653), .ZN(n16310) );
  INV_X1 U19524 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16667) );
  NAND2_X1 U19525 ( .A1(n16654), .A2(n16303), .ZN(n16305) );
  AOI221_X1 U19526 ( .B1(n16310), .B2(n16667), .C1(n16305), .C2(
        P3_EBX_REG_30__SCAN_IN), .A(n16304), .ZN(n16306) );
  OAI211_X1 U19527 ( .C1(n16620), .C2(n16308), .A(n16307), .B(n16306), .ZN(
        P3_U2641) );
  AOI22_X1 U19528 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n16642), .B1(
        P3_EBX_REG_29__SCAN_IN), .B2(n16613), .ZN(n16319) );
  NAND2_X1 U19529 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16321), .ZN(n16309) );
  AOI22_X1 U19530 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16311), .B1(n16310), 
        .B2(n16309), .ZN(n16318) );
  OAI211_X1 U19531 ( .C1(n16314), .C2(n16313), .A(n9662), .B(n16312), .ZN(
        n16317) );
  NAND3_X1 U19532 ( .A1(n16315), .A2(n16335), .A3(n18637), .ZN(n16316) );
  NAND4_X1 U19533 ( .A1(n16319), .A2(n16318), .A3(n16317), .A4(n16316), .ZN(
        P3_U2642) );
  AOI22_X1 U19534 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16642), .B1(
        P3_EBX_REG_28__SCAN_IN), .B2(n16613), .ZN(n16330) );
  INV_X1 U19535 ( .A(n16340), .ZN(n16342) );
  AOI21_X1 U19536 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n16320), .A(n16653), .ZN(
        n16322) );
  AOI22_X1 U19537 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n16342), .B1(n16322), 
        .B2(n16321), .ZN(n16329) );
  OAI211_X1 U19538 ( .C1(n16325), .C2(n16324), .A(n9662), .B(n16323), .ZN(
        n16328) );
  OAI211_X1 U19539 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16335), .B(n16326), .ZN(n16327) );
  NAND4_X1 U19540 ( .A1(n16330), .A2(n16329), .A3(n16328), .A4(n16327), .ZN(
        P3_U2643) );
  AOI211_X1 U19541 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n16345), .A(n16331), .B(
        n16653), .ZN(n16334) );
  AOI22_X1 U19542 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16642), .B1(
        P3_EBX_REG_27__SCAN_IN), .B2(n16613), .ZN(n16332) );
  INV_X1 U19543 ( .A(n16332), .ZN(n16333) );
  AOI211_X1 U19544 ( .C1(n16335), .C2(n18633), .A(n16334), .B(n16333), .ZN(
        n16339) );
  OAI211_X1 U19545 ( .C1(n17344), .C2(n16337), .A(n9662), .B(n16336), .ZN(
        n16338) );
  OAI211_X1 U19546 ( .C1(n16340), .C2(n18633), .A(n16339), .B(n16338), .ZN(
        P3_U2644) );
  AOI22_X1 U19547 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16642), .B1(
        P3_EBX_REG_26__SCAN_IN), .B2(n16613), .ZN(n16350) );
  NOR2_X1 U19548 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16358), .ZN(n16341) );
  AOI22_X1 U19549 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16342), .B1(
        P3_REIP_REG_25__SCAN_IN), .B2(n16341), .ZN(n16349) );
  OAI211_X1 U19550 ( .C1(n17353), .C2(n16344), .A(n9662), .B(n16343), .ZN(
        n16348) );
  OAI211_X1 U19551 ( .C1(n16346), .C2(n16773), .A(n16600), .B(n16345), .ZN(
        n16347) );
  NAND4_X1 U19552 ( .A1(n16350), .A2(n16349), .A3(n16348), .A4(n16347), .ZN(
        P3_U2645) );
  AND3_X1 U19553 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16655), .A3(n16359), 
        .ZN(n16353) );
  XNOR2_X1 U19554 ( .A(P3_EBX_REG_25__SCAN_IN), .B(n16361), .ZN(n16351) );
  INV_X1 U19555 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16662) );
  OAI22_X1 U19556 ( .A1(n16653), .A2(n16351), .B1(n16662), .B2(n16654), .ZN(
        n16352) );
  AOI211_X1 U19557 ( .C1(n16642), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16353), .B(n16352), .ZN(n16357) );
  OAI211_X1 U19558 ( .C1(n17373), .C2(n16355), .A(n9662), .B(n16354), .ZN(
        n16356) );
  OAI211_X1 U19559 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n16358), .A(n16357), 
        .B(n16356), .ZN(P3_U2646) );
  AOI22_X1 U19560 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16642), .B1(
        P3_EBX_REG_24__SCAN_IN), .B2(n16613), .ZN(n16367) );
  OAI21_X1 U19561 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n16360), .A(n16359), 
        .ZN(n16366) );
  OAI211_X1 U19562 ( .C1(n16368), .C2(n16772), .A(n16600), .B(n16361), .ZN(
        n16365) );
  OAI211_X1 U19563 ( .C1(n17384), .C2(n16363), .A(n9662), .B(n16362), .ZN(
        n16364) );
  NAND4_X1 U19564 ( .A1(n16367), .A2(n16366), .A3(n16365), .A4(n16364), .ZN(
        P3_U2647) );
  INV_X1 U19565 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18622) );
  NOR2_X1 U19566 ( .A1(n18622), .A2(n16381), .ZN(n16379) );
  AOI21_X1 U19567 ( .B1(P3_REIP_REG_22__SCAN_IN), .B2(n16379), .A(
        P3_REIP_REG_23__SCAN_IN), .ZN(n16378) );
  AOI211_X1 U19568 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n16386), .A(n16368), .B(
        n16653), .ZN(n16371) );
  NOR2_X1 U19569 ( .A1(n16369), .A2(n16607), .ZN(n16370) );
  AOI211_X1 U19570 ( .C1(n16613), .C2(P3_EBX_REG_23__SCAN_IN), .A(n16371), .B(
        n16370), .ZN(n16376) );
  OAI211_X1 U19571 ( .C1(n16374), .C2(n16373), .A(n9662), .B(n16372), .ZN(
        n16375) );
  OAI211_X1 U19572 ( .C1(n16378), .C2(n16377), .A(n16376), .B(n16375), .ZN(
        P3_U2648) );
  AOI22_X1 U19573 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n16642), .B1(
        P3_EBX_REG_22__SCAN_IN), .B2(n16613), .ZN(n16390) );
  INV_X1 U19574 ( .A(n16379), .ZN(n16383) );
  NAND2_X1 U19575 ( .A1(n16655), .A2(n16380), .ZN(n16399) );
  INV_X1 U19576 ( .A(n16399), .ZN(n16401) );
  NOR2_X1 U19577 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16381), .ZN(n16394) );
  NOR2_X1 U19578 ( .A1(n16401), .A2(n16394), .ZN(n16382) );
  MUX2_X1 U19579 ( .A(n16383), .B(n16382), .S(P3_REIP_REG_22__SCAN_IN), .Z(
        n16389) );
  OAI211_X1 U19580 ( .C1(n17416), .C2(n16385), .A(n9662), .B(n16384), .ZN(
        n16388) );
  OAI211_X1 U19581 ( .C1(n16391), .C2(n16771), .A(n16600), .B(n16386), .ZN(
        n16387) );
  NAND4_X1 U19582 ( .A1(n16390), .A2(n16389), .A3(n16388), .A4(n16387), .ZN(
        P3_U2649) );
  AOI211_X1 U19583 ( .C1(P3_EBX_REG_21__SCAN_IN), .C2(n16404), .A(n16391), .B(
        n16653), .ZN(n16393) );
  INV_X1 U19584 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16831) );
  OAI22_X1 U19585 ( .A1(n17430), .A2(n16607), .B1(n16831), .B2(n16654), .ZN(
        n16392) );
  NOR3_X1 U19586 ( .A1(n16394), .A2(n16393), .A3(n16392), .ZN(n16398) );
  OAI211_X1 U19587 ( .C1(n17428), .C2(n16396), .A(n9662), .B(n16395), .ZN(
        n16397) );
  OAI211_X1 U19588 ( .C1(n16399), .C2(n18622), .A(n16398), .B(n16397), .ZN(
        P3_U2650) );
  AOI22_X1 U19589 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n16642), .B1(
        P3_EBX_REG_20__SCAN_IN), .B2(n16613), .ZN(n16408) );
  NAND2_X1 U19590 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16421) );
  NOR2_X1 U19591 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16421), .ZN(n16400) );
  AOI22_X1 U19592 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16401), .B1(n16424), 
        .B2(n16400), .ZN(n16407) );
  OAI211_X1 U19593 ( .C1(n16403), .C2(n17446), .A(n9662), .B(n16402), .ZN(
        n16406) );
  OAI211_X1 U19594 ( .C1(n16416), .C2(n16845), .A(n16600), .B(n16404), .ZN(
        n16405) );
  NAND4_X1 U19595 ( .A1(n16408), .A2(n16407), .A3(n16406), .A4(n16405), .ZN(
        P3_U2651) );
  INV_X1 U19596 ( .A(n16409), .ZN(n16410) );
  NAND2_X1 U19597 ( .A1(n16655), .A2(n16410), .ZN(n16438) );
  INV_X1 U19598 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18618) );
  INV_X1 U19599 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n20909) );
  NOR2_X1 U19600 ( .A1(n20909), .A2(n16435), .ZN(n16412) );
  OAI21_X1 U19601 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16412), .A(
        n16411), .ZN(n17460) );
  NAND2_X1 U19602 ( .A1(n17455), .A2(n16413), .ZN(n16425) );
  OAI21_X1 U19603 ( .B1(n20909), .B2(n16425), .A(n16617), .ZN(n16415) );
  OAI21_X1 U19604 ( .B1(n17460), .B2(n16415), .A(n9662), .ZN(n16414) );
  AOI21_X1 U19605 ( .B1(n17460), .B2(n16415), .A(n16414), .ZN(n16420) );
  AOI211_X1 U19606 ( .C1(P3_EBX_REG_19__SCAN_IN), .C2(n16428), .A(n16416), .B(
        n16653), .ZN(n16419) );
  AOI22_X1 U19607 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n16642), .B1(
        P3_EBX_REG_19__SCAN_IN), .B2(n16613), .ZN(n16417) );
  INV_X1 U19608 ( .A(n16417), .ZN(n16418) );
  NOR4_X1 U19609 ( .A1(n17815), .A2(n16420), .A3(n16419), .A4(n16418), .ZN(
        n16423) );
  OAI211_X1 U19610 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(P3_REIP_REG_18__SCAN_IN), .A(n16424), .B(n16421), .ZN(n16422) );
  OAI211_X1 U19611 ( .C1(n16438), .C2(n18618), .A(n16423), .B(n16422), .ZN(
        P3_U2652) );
  INV_X1 U19612 ( .A(n16424), .ZN(n16434) );
  INV_X1 U19613 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18615) );
  AOI22_X1 U19614 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16435), .B1(
        n17455), .B2(n20909), .ZN(n17465) );
  NAND2_X1 U19615 ( .A1(n16617), .A2(n16425), .ZN(n16427) );
  OAI21_X1 U19616 ( .B1(n17465), .B2(n16427), .A(n9662), .ZN(n16426) );
  AOI21_X1 U19617 ( .B1(n17465), .B2(n16427), .A(n16426), .ZN(n16432) );
  OAI211_X1 U19618 ( .C1(n16437), .C2(n16430), .A(n16600), .B(n16428), .ZN(
        n16429) );
  OAI211_X1 U19619 ( .C1(n16430), .C2(n16654), .A(n18017), .B(n16429), .ZN(
        n16431) );
  AOI211_X1 U19620 ( .C1(n16642), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16432), .B(n16431), .ZN(n16433) );
  OAI221_X1 U19621 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16434), .C1(n18615), 
        .C2(n16438), .A(n16433), .ZN(P3_U2653) );
  NAND2_X1 U19622 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17494) );
  NOR2_X1 U19623 ( .A1(n17494), .A2(n16472), .ZN(n16447) );
  OAI21_X1 U19624 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16447), .A(
        n16435), .ZN(n17486) );
  NOR2_X1 U19625 ( .A1(n17692), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16638) );
  INV_X1 U19626 ( .A(n16638), .ZN(n16605) );
  OAI21_X1 U19627 ( .B1(n17479), .B2(n16605), .A(n16617), .ZN(n16436) );
  XNOR2_X1 U19628 ( .A(n17486), .B(n16436), .ZN(n16445) );
  AOI211_X1 U19629 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n16451), .A(n16437), .B(
        n16653), .ZN(n16443) );
  INV_X1 U19630 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16875) );
  OAI22_X1 U19631 ( .A1(n17478), .A2(n16607), .B1(n16875), .B2(n16654), .ZN(
        n16442) );
  NAND2_X1 U19632 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16456) );
  NOR2_X1 U19633 ( .A1(n16456), .A2(n16470), .ZN(n16440) );
  INV_X1 U19634 ( .A(n16438), .ZN(n16439) );
  MUX2_X1 U19635 ( .A(n16440), .B(n16439), .S(P3_REIP_REG_17__SCAN_IN), .Z(
        n16441) );
  NOR4_X1 U19636 ( .A1(n17815), .A2(n16443), .A3(n16442), .A4(n16441), .ZN(
        n16444) );
  OAI21_X1 U19637 ( .B1(n16620), .B2(n16445), .A(n16444), .ZN(P3_U2654) );
  INV_X1 U19638 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18611) );
  NAND2_X1 U19639 ( .A1(n16655), .A2(n16446), .ZN(n16469) );
  INV_X1 U19640 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16448) );
  AOI21_X1 U19641 ( .B1(n16448), .B2(n16460), .A(n16447), .ZN(n17492) );
  INV_X1 U19642 ( .A(n16462), .ZN(n16450) );
  INV_X1 U19643 ( .A(n17492), .ZN(n16449) );
  AOI221_X1 U19644 ( .B1(n16462), .B2(n17492), .C1(n16450), .C2(n16449), .A(
        n16620), .ZN(n16455) );
  OAI211_X1 U19645 ( .C1(n16461), .C2(n16453), .A(n16600), .B(n16451), .ZN(
        n16452) );
  OAI211_X1 U19646 ( .C1(n16453), .C2(n16654), .A(n18017), .B(n16452), .ZN(
        n16454) );
  AOI211_X1 U19647 ( .C1(n16642), .C2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16455), .B(n16454), .ZN(n16459) );
  INV_X1 U19648 ( .A(n16470), .ZN(n16457) );
  OAI211_X1 U19649 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(P3_REIP_REG_15__SCAN_IN), .A(n16457), .B(n16456), .ZN(n16458) );
  OAI211_X1 U19650 ( .C1(n18611), .C2(n16469), .A(n16459), .B(n16458), .ZN(
        P3_U2655) );
  INV_X1 U19651 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18609) );
  OAI21_X1 U19652 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17491), .A(
        n16460), .ZN(n17505) );
  INV_X1 U19653 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16635) );
  OAI21_X1 U19654 ( .B1(n16587), .B2(n16635), .A(n9662), .ZN(n16652) );
  AOI211_X1 U19655 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n16617), .A(
        n17505), .B(n16652), .ZN(n16467) );
  AOI211_X1 U19656 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n16478), .A(n16461), .B(
        n16653), .ZN(n16466) );
  NAND3_X1 U19657 ( .A1(n17505), .A2(n16462), .A3(n9662), .ZN(n16464) );
  AOI22_X1 U19658 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n16642), .B1(
        P3_EBX_REG_15__SCAN_IN), .B2(n16613), .ZN(n16463) );
  NAND2_X1 U19659 ( .A1(n16464), .A2(n16463), .ZN(n16465) );
  NOR4_X1 U19660 ( .A1(n17815), .A2(n16467), .A3(n16466), .A4(n16465), .ZN(
        n16468) );
  OAI221_X1 U19661 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16470), .C1(n18609), 
        .C2(n16469), .A(n16468), .ZN(P3_U2656) );
  INV_X1 U19662 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16482) );
  AOI21_X1 U19663 ( .B1(P3_REIP_REG_14__SCAN_IN), .B2(n16655), .A(n16471), 
        .ZN(n16475) );
  NAND2_X1 U19664 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17603), .ZN(
        n16508) );
  NOR2_X1 U19665 ( .A1(n16473), .A2(n16508), .ZN(n17529) );
  AND2_X1 U19666 ( .A1(n17528), .A2(n17529), .ZN(n16486) );
  OAI21_X1 U19667 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16486), .A(
        n16472), .ZN(n17518) );
  NAND2_X1 U19668 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17632), .ZN(
        n16586) );
  INV_X1 U19669 ( .A(n16586), .ZN(n16573) );
  NAND2_X1 U19670 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16573), .ZN(
        n16572) );
  NOR2_X1 U19671 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16572), .ZN(
        n16566) );
  NAND2_X1 U19672 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n16566), .ZN(
        n16546) );
  OAI21_X1 U19673 ( .B1(n16473), .B2(n16546), .A(n16617), .ZN(n16499) );
  OAI21_X1 U19674 ( .B1(n17528), .B2(n16587), .A(n16499), .ZN(n16488) );
  XOR2_X1 U19675 ( .A(n17518), .B(n16488), .Z(n16474) );
  OAI22_X1 U19676 ( .A1(n16476), .A2(n16475), .B1(n16620), .B2(n16474), .ZN(
        n16477) );
  AOI211_X1 U19677 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16613), .A(n17821), .B(
        n16477), .ZN(n16481) );
  OAI211_X1 U19678 ( .C1(n16490), .C2(n16479), .A(n16600), .B(n16478), .ZN(
        n16480) );
  OAI211_X1 U19679 ( .C1(n16607), .C2(n16482), .A(n16481), .B(n16480), .ZN(
        P3_U2657) );
  NOR3_X1 U19680 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16646), .A3(n16483), 
        .ZN(n16484) );
  AOI211_X1 U19681 ( .C1(P3_EBX_REG_13__SCAN_IN), .C2(n16613), .A(n17821), .B(
        n16484), .ZN(n16496) );
  INV_X1 U19682 ( .A(n16485), .ZN(n16498) );
  OAI21_X1 U19683 ( .B1(n16649), .B2(n16498), .A(n16655), .ZN(n16513) );
  INV_X1 U19684 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18603) );
  NAND2_X1 U19685 ( .A1(n16630), .A2(n18603), .ZN(n16497) );
  AOI21_X1 U19686 ( .B1(n16513), .B2(n16497), .A(n18605), .ZN(n16494) );
  NAND2_X1 U19687 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17529), .ZN(
        n16487) );
  AOI21_X1 U19688 ( .B1(n17532), .B2(n16487), .A(n16486), .ZN(n17535) );
  INV_X1 U19689 ( .A(n17535), .ZN(n16489) );
  AND3_X1 U19690 ( .A1(n16489), .A2(n16488), .A3(n9662), .ZN(n16493) );
  AOI211_X1 U19691 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n16617), .A(
        n16489), .B(n16652), .ZN(n16492) );
  AOI211_X1 U19692 ( .C1(P3_EBX_REG_13__SCAN_IN), .C2(n16503), .A(n16490), .B(
        n16653), .ZN(n16491) );
  NOR4_X1 U19693 ( .A1(n16494), .A2(n16493), .A3(n16492), .A4(n16491), .ZN(
        n16495) );
  OAI211_X1 U19694 ( .C1(n17532), .C2(n16607), .A(n16496), .B(n16495), .ZN(
        P3_U2658) );
  OAI22_X1 U19695 ( .A1(n16504), .A2(n16654), .B1(n16498), .B2(n16497), .ZN(
        n16502) );
  INV_X1 U19696 ( .A(n17529), .ZN(n16509) );
  AOI22_X1 U19697 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17529), .B1(
        n16509), .B2(n17546), .ZN(n17553) );
  XOR2_X1 U19698 ( .A(n17553), .B(n16499), .Z(n16500) );
  OAI22_X1 U19699 ( .A1(n16620), .A2(n16500), .B1(n18603), .B2(n16513), .ZN(
        n16501) );
  NOR3_X1 U19700 ( .A1(n17821), .A2(n16502), .A3(n16501), .ZN(n16506) );
  OAI211_X1 U19701 ( .C1(n16507), .C2(n16504), .A(n16600), .B(n16503), .ZN(
        n16505) );
  OAI211_X1 U19702 ( .C1(n16607), .C2(n17546), .A(n16506), .B(n16505), .ZN(
        P3_U2659) );
  AOI211_X1 U19703 ( .C1(P3_EBX_REG_11__SCAN_IN), .C2(n16526), .A(n16507), .B(
        n16653), .ZN(n16516) );
  INV_X1 U19704 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18598) );
  NAND2_X1 U19705 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n16568) );
  NOR3_X1 U19706 ( .A1(n16646), .A2(n16567), .A3(n16568), .ZN(n16552) );
  NAND2_X1 U19707 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16552), .ZN(n16539) );
  NOR2_X1 U19708 ( .A1(n18598), .A2(n16539), .ZN(n16525) );
  AOI21_X1 U19709 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n16525), .A(
        P3_REIP_REG_11__SCAN_IN), .ZN(n16514) );
  INV_X1 U19710 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17577) );
  INV_X1 U19711 ( .A(n16508), .ZN(n16559) );
  NAND2_X1 U19712 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16559), .ZN(
        n16545) );
  INV_X1 U19713 ( .A(n16545), .ZN(n16535) );
  NAND2_X1 U19714 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16535), .ZN(
        n16520) );
  NOR2_X1 U19715 ( .A1(n17577), .A2(n16520), .ZN(n16519) );
  OAI21_X1 U19716 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16519), .A(
        n16509), .ZN(n17561) );
  NAND2_X1 U19717 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16510) );
  OAI21_X1 U19718 ( .B1(n16510), .B2(n16546), .A(n16617), .ZN(n16537) );
  OAI21_X1 U19719 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16587), .A(
        n16537), .ZN(n16511) );
  XOR2_X1 U19720 ( .A(n17561), .B(n16511), .Z(n16512) );
  OAI22_X1 U19721 ( .A1(n16514), .A2(n16513), .B1(n16620), .B2(n16512), .ZN(
        n16515) );
  AOI211_X1 U19722 ( .C1(n16642), .C2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n16516), .B(n16515), .ZN(n16517) );
  OAI211_X1 U19723 ( .C1(n16951), .C2(n16654), .A(n16517), .B(n17909), .ZN(
        P3_U2660) );
  AOI22_X1 U19724 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16642), .B1(
        P3_EBX_REG_10__SCAN_IN), .B2(n16613), .ZN(n16530) );
  INV_X1 U19725 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18599) );
  AOI21_X1 U19726 ( .B1(n16567), .B2(n16630), .A(n16649), .ZN(n16596) );
  INV_X1 U19727 ( .A(n16596), .ZN(n16580) );
  AOI21_X1 U19728 ( .B1(n16630), .B2(n16518), .A(n16580), .ZN(n16544) );
  OAI21_X1 U19729 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(n16539), .A(n16544), .ZN(
        n16524) );
  AOI21_X1 U19730 ( .B1(n17577), .B2(n16520), .A(n16519), .ZN(n17580) );
  INV_X1 U19731 ( .A(n16537), .ZN(n16522) );
  INV_X1 U19732 ( .A(n17580), .ZN(n16521) );
  AOI221_X1 U19733 ( .B1(n17580), .B2(n16522), .C1(n16521), .C2(n16537), .A(
        n16620), .ZN(n16523) );
  AOI221_X1 U19734 ( .B1(n16525), .B2(n18599), .C1(n16524), .C2(
        P3_REIP_REG_10__SCAN_IN), .A(n16523), .ZN(n16529) );
  OAI211_X1 U19735 ( .C1(n16531), .C2(n16527), .A(n16600), .B(n16526), .ZN(
        n16528) );
  NAND4_X1 U19736 ( .A1(n16530), .A2(n16529), .A3(n17909), .A4(n16528), .ZN(
        P3_U2661) );
  AOI211_X1 U19737 ( .C1(P3_EBX_REG_9__SCAN_IN), .C2(n16553), .A(n16531), .B(
        n16653), .ZN(n16533) );
  INV_X1 U19738 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16534) );
  OAI22_X1 U19739 ( .A1(n16534), .A2(n16535), .B1(n16545), .B2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16536) );
  INV_X1 U19740 ( .A(n16536), .ZN(n17592) );
  NOR2_X1 U19741 ( .A1(n16620), .A2(n16617), .ZN(n16604) );
  INV_X1 U19742 ( .A(n16604), .ZN(n16641) );
  OAI22_X1 U19743 ( .A1(n17592), .A2(n16641), .B1(n16534), .B2(n16607), .ZN(
        n16532) );
  AOI211_X1 U19744 ( .C1(n16613), .C2(P3_EBX_REG_9__SCAN_IN), .A(n16533), .B(
        n16532), .ZN(n16543) );
  NAND2_X1 U19745 ( .A1(n16535), .A2(n16534), .ZN(n16538) );
  OAI22_X1 U19746 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16538), .B1(
        n16537), .B2(n16536), .ZN(n16541) );
  NOR2_X1 U19747 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16539), .ZN(n16540) );
  OAI211_X1 U19748 ( .C1(n16544), .C2(n18598), .A(n16543), .B(n16542), .ZN(
        P3_U2662) );
  AOI22_X1 U19749 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16642), .B1(
        P3_EBX_REG_8__SCAN_IN), .B2(n16613), .ZN(n16557) );
  INV_X1 U19750 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18595) );
  INV_X1 U19751 ( .A(n16544), .ZN(n16551) );
  OAI21_X1 U19752 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16559), .A(
        n16545), .ZN(n16548) );
  INV_X1 U19753 ( .A(n16548), .ZN(n17602) );
  NAND2_X1 U19754 ( .A1(n16617), .A2(n16546), .ZN(n16547) );
  INV_X1 U19755 ( .A(n16547), .ZN(n16549) );
  AOI221_X1 U19756 ( .B1(n17602), .B2(n16549), .C1(n16548), .C2(n16547), .A(
        n16620), .ZN(n16550) );
  AOI221_X1 U19757 ( .B1(n16552), .B2(n18595), .C1(n16551), .C2(
        P3_REIP_REG_8__SCAN_IN), .A(n16550), .ZN(n16556) );
  OAI211_X1 U19758 ( .C1(n16563), .C2(n16554), .A(n16600), .B(n16553), .ZN(
        n16555) );
  NAND4_X1 U19759 ( .A1(n16557), .A2(n16556), .A3(n17909), .A4(n16555), .ZN(
        P3_U2663) );
  OAI22_X1 U19760 ( .A1(n17617), .A2(n16607), .B1(n16558), .B2(n16654), .ZN(
        n16565) );
  AOI21_X1 U19761 ( .B1(n17617), .B2(n16572), .A(n16559), .ZN(n17622) );
  INV_X1 U19762 ( .A(n16566), .ZN(n16560) );
  NAND2_X1 U19763 ( .A1(n16643), .A2(n16560), .ZN(n16574) );
  AOI21_X1 U19764 ( .B1(n16581), .B2(P3_EBX_REG_7__SCAN_IN), .A(n16653), .ZN(
        n16561) );
  INV_X1 U19765 ( .A(n16561), .ZN(n16562) );
  OAI22_X1 U19766 ( .A1(n17622), .A2(n16574), .B1(n16563), .B2(n16562), .ZN(
        n16564) );
  AOI211_X1 U19767 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(n16580), .A(n16565), .B(
        n16564), .ZN(n16571) );
  OAI211_X1 U19768 ( .C1(n16566), .C2(n16587), .A(n9662), .B(n17622), .ZN(
        n16570) );
  NOR2_X1 U19769 ( .A1(n16646), .A2(n16567), .ZN(n16575) );
  OAI211_X1 U19770 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(P3_REIP_REG_6__SCAN_IN), 
        .A(n16575), .B(n16568), .ZN(n16569) );
  NAND4_X1 U19771 ( .A1(n16571), .A2(n18017), .A3(n16570), .A4(n16569), .ZN(
        P3_U2664) );
  AOI22_X1 U19772 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16642), .B1(
        P3_EBX_REG_6__SCAN_IN), .B2(n16613), .ZN(n16584) );
  OAI21_X1 U19773 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16573), .A(
        n16572), .ZN(n17635) );
  AOI211_X1 U19774 ( .C1(n16586), .C2(n16641), .A(n17635), .B(n16652), .ZN(
        n16579) );
  INV_X1 U19775 ( .A(n16574), .ZN(n16576) );
  INV_X1 U19776 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18591) );
  AOI22_X1 U19777 ( .A1(n17635), .A2(n16576), .B1(n18591), .B2(n16575), .ZN(
        n16577) );
  INV_X1 U19778 ( .A(n16577), .ZN(n16578) );
  AOI211_X1 U19779 ( .C1(P3_REIP_REG_6__SCAN_IN), .C2(n16580), .A(n16579), .B(
        n16578), .ZN(n16583) );
  OAI211_X1 U19780 ( .C1(n16590), .C2(n20863), .A(n16600), .B(n16581), .ZN(
        n16582) );
  NAND4_X1 U19781 ( .A1(n16584), .A2(n16583), .A3(n17909), .A4(n16582), .ZN(
        P3_U2665) );
  AOI21_X1 U19782 ( .B1(n16630), .B2(n16585), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n16595) );
  AOI21_X1 U19783 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n16613), .A(n17815), .ZN(
        n16594) );
  INV_X1 U19784 ( .A(n17642), .ZN(n16616) );
  INV_X1 U19785 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17661) );
  NOR3_X1 U19786 ( .A1(n17692), .A2(n16616), .A3(n17661), .ZN(n16597) );
  OAI21_X1 U19787 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16597), .A(
        n16586), .ZN(n17648) );
  INV_X1 U19788 ( .A(n17648), .ZN(n16589) );
  AOI21_X1 U19789 ( .B1(n16635), .B2(n16597), .A(n16587), .ZN(n16588) );
  INV_X1 U19790 ( .A(n16588), .ZN(n16606) );
  AOI221_X1 U19791 ( .B1(n16589), .B2(n16588), .C1(n17648), .C2(n16606), .A(
        n16620), .ZN(n16592) );
  AOI211_X1 U19792 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n16599), .A(n16590), .B(
        n16653), .ZN(n16591) );
  AOI211_X1 U19793 ( .C1(n16642), .C2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n16592), .B(n16591), .ZN(n16593) );
  OAI211_X1 U19794 ( .C1(n16596), .C2(n16595), .A(n16594), .B(n16593), .ZN(
        P3_U2666) );
  AOI21_X1 U19795 ( .B1(n16630), .B2(n16612), .A(n16649), .ZN(n16621) );
  NAND2_X1 U19796 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17642), .ZN(
        n16598) );
  AOI21_X1 U19797 ( .B1(n17661), .B2(n16598), .A(n16597), .ZN(n17658) );
  NOR3_X1 U19798 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16646), .A3(n16612), .ZN(
        n16603) );
  NAND2_X1 U19799 ( .A1(n18040), .A2(n18718), .ZN(n16660) );
  OAI211_X1 U19800 ( .C1(n16614), .C2(n17037), .A(n16600), .B(n16599), .ZN(
        n16601) );
  OAI221_X1 U19801 ( .B1(n16660), .B2(n10741), .C1(n16660), .C2(n18496), .A(
        n16601), .ZN(n16602) );
  AOI211_X1 U19802 ( .C1(n16604), .C2(n17658), .A(n16603), .B(n16602), .ZN(
        n16611) );
  NAND2_X1 U19803 ( .A1(n17642), .A2(n17661), .ZN(n17653) );
  OAI22_X1 U19804 ( .A1(n17658), .A2(n16606), .B1(n16605), .B2(n17653), .ZN(
        n16609) );
  OAI22_X1 U19805 ( .A1(n17661), .A2(n16607), .B1(n17037), .B2(n16654), .ZN(
        n16608) );
  OAI211_X1 U19806 ( .C1(n16621), .C2(n18587), .A(n16611), .B(n16610), .ZN(
        P3_U2667) );
  NAND2_X1 U19807 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16629) );
  NAND2_X1 U19808 ( .A1(n16630), .A2(n16612), .ZN(n16626) );
  INV_X1 U19809 ( .A(n16660), .ZN(n18720) );
  NOR2_X1 U19810 ( .A1(n18683), .A2(n18512), .ZN(n18504) );
  OAI21_X1 U19811 ( .B1(n18504), .B2(n18661), .A(n16987), .ZN(n18658) );
  AOI22_X1 U19812 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n16613), .B1(n18720), .B2(
        n18658), .ZN(n16625) );
  AOI211_X1 U19813 ( .C1(P3_EBX_REG_3__SCAN_IN), .C2(n16615), .A(n16614), .B(
        n16653), .ZN(n16623) );
  INV_X1 U19814 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18584) );
  NAND2_X1 U19815 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16627) );
  INV_X1 U19816 ( .A(n16627), .ZN(n16636) );
  OAI22_X1 U19817 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n16636), .B1(
        n17692), .B2(n16616), .ZN(n17668) );
  OAI21_X1 U19818 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16627), .A(
        n16617), .ZN(n16618) );
  XNOR2_X1 U19819 ( .A(n17668), .B(n16618), .ZN(n16619) );
  OAI22_X1 U19820 ( .A1(n16621), .A2(n18584), .B1(n16620), .B2(n16619), .ZN(
        n16622) );
  AOI211_X1 U19821 ( .C1(n16642), .C2(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n16623), .B(n16622), .ZN(n16624) );
  OAI211_X1 U19822 ( .C1(n16629), .C2(n16626), .A(n16625), .B(n16624), .ZN(
        P3_U2668) );
  OAI21_X1 U19823 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16627), .ZN(n17679) );
  AOI211_X1 U19824 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16644), .A(n16628), .B(
        n16653), .ZN(n16634) );
  AOI21_X1 U19825 ( .B1(n18671), .B2(n18509), .A(n18504), .ZN(n18669) );
  AOI22_X1 U19826 ( .A1(n16649), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n18669), 
        .B2(n18720), .ZN(n16632) );
  OAI211_X1 U19827 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16630), .B(n16629), .ZN(n16631) );
  OAI211_X1 U19828 ( .C1(n16654), .C2(n17045), .A(n16632), .B(n16631), .ZN(
        n16633) );
  AOI211_X1 U19829 ( .C1(n16642), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n16634), .B(n16633), .ZN(n16640) );
  NAND2_X1 U19830 ( .A1(n16636), .A2(n16635), .ZN(n16637) );
  OAI211_X1 U19831 ( .C1(n16638), .C2(n17679), .A(n16643), .B(n16637), .ZN(
        n16639) );
  OAI211_X1 U19832 ( .C1(n16641), .C2(n17679), .A(n16640), .B(n16639), .ZN(
        P3_U2669) );
  AOI21_X1 U19833 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16643), .A(
        n16642), .ZN(n16651) );
  OAI21_X1 U19834 ( .B1(n17051), .B2(n20934), .A(n16644), .ZN(n17052) );
  OAI22_X1 U19835 ( .A1(n17051), .A2(n16654), .B1(n16653), .B2(n17052), .ZN(
        n16648) );
  NAND2_X1 U19836 ( .A1(n16645), .A2(n18509), .ZN(n18672) );
  OAI22_X1 U19837 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16646), .B1(n18672), 
        .B2(n16660), .ZN(n16647) );
  AOI211_X1 U19838 ( .C1(n16649), .C2(P3_REIP_REG_1__SCAN_IN), .A(n16648), .B(
        n16647), .ZN(n16650) );
  OAI221_X1 U19839 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16652), .C1(
        n17692), .C2(n16651), .A(n16650), .ZN(P3_U2670) );
  NAND2_X1 U19840 ( .A1(n16654), .A2(n16653), .ZN(n16656) );
  AOI22_X1 U19841 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n16656), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n16655), .ZN(n16659) );
  NAND3_X1 U19842 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18666), .A3(
        n16657), .ZN(n16658) );
  OAI211_X1 U19843 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n16660), .A(
        n16659), .B(n16658), .ZN(P3_U2671) );
  AND2_X2 U19844 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n16917), .ZN(n16891) );
  INV_X1 U19845 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16847) );
  NAND2_X1 U19846 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16861), .ZN(n16818) );
  NAND4_X1 U19847 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(P3_EBX_REG_23__SCAN_IN), .A4(P3_EBX_REG_24__SCAN_IN), .ZN(n16661)
         );
  NOR4_X1 U19848 ( .A1(n16662), .A2(n16773), .A3(n16818), .A4(n16661), .ZN(
        n16663) );
  NAND4_X1 U19849 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(P3_EBX_REG_28__SCAN_IN), 
        .A3(P3_EBX_REG_29__SCAN_IN), .A4(n16663), .ZN(n16666) );
  NAND2_X1 U19850 ( .A1(n17054), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16665) );
  NAND2_X1 U19851 ( .A1(n16770), .A2(n18077), .ZN(n16664) );
  OAI22_X1 U19852 ( .A1(n16770), .A2(n16665), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16664), .ZN(P3_U2672) );
  NAND2_X1 U19853 ( .A1(n16667), .A2(n16666), .ZN(n16668) );
  NAND2_X1 U19854 ( .A1(n16668), .A2(n17054), .ZN(n16769) );
  AOI22_X1 U19855 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16678) );
  INV_X1 U19856 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16921) );
  AOI22_X1 U19857 ( .A1(n17025), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17006), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16670) );
  AOI22_X1 U19858 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17009), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16669) );
  OAI211_X1 U19859 ( .C1(n16962), .C2(n16921), .A(n16670), .B(n16669), .ZN(
        n16676) );
  AOI22_X1 U19860 ( .A1(n9579), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16674) );
  AOI22_X1 U19861 ( .A1(n16991), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16673) );
  AOI22_X1 U19862 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9585), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16672) );
  NAND2_X1 U19863 ( .A1(n16734), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n16671) );
  NAND4_X1 U19864 ( .A1(n16674), .A2(n16673), .A3(n16672), .A4(n16671), .ZN(
        n16675) );
  AOI211_X1 U19865 ( .C1(n16965), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n16676), .B(n16675), .ZN(n16677) );
  OAI211_X1 U19866 ( .C1(n17001), .C2(n18286), .A(n16678), .B(n16677), .ZN(
        n16774) );
  AOI22_X1 U19867 ( .A1(n9577), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16679) );
  OAI21_X1 U19868 ( .B1(n16756), .B2(n18069), .A(n16679), .ZN(n16688) );
  AOI22_X1 U19869 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9571), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16686) );
  OAI22_X1 U19870 ( .A1(n10797), .A2(n20936), .B1(n9575), .B2(n18319), .ZN(
        n16684) );
  AOI22_X1 U19871 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17025), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16682) );
  AOI22_X1 U19872 ( .A1(n17009), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16681) );
  AOI22_X1 U19873 ( .A1(n16893), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16680) );
  NAND3_X1 U19874 ( .A1(n16682), .A2(n16681), .A3(n16680), .ZN(n16683) );
  AOI211_X1 U19875 ( .C1(n17006), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n16684), .B(n16683), .ZN(n16685) );
  OAI211_X1 U19876 ( .C1(n17001), .C2(n18283), .A(n16686), .B(n16685), .ZN(
        n16687) );
  AOI211_X1 U19877 ( .C1(n16992), .C2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n16688), .B(n16687), .ZN(n16777) );
  AOI22_X1 U19878 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(n9579), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16689) );
  OAI21_X1 U19879 ( .B1(n16987), .B2(n16961), .A(n16689), .ZN(n16698) );
  AOI22_X1 U19880 ( .A1(n16955), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16696) );
  AOI22_X1 U19881 ( .A1(n16734), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16690) );
  OAI21_X1 U19882 ( .B1(n16756), .B2(n18057), .A(n16690), .ZN(n16694) );
  AOI22_X1 U19883 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16692) );
  AOI22_X1 U19884 ( .A1(n17025), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10887), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16691) );
  OAI211_X1 U19885 ( .C1(n15418), .C2(n16850), .A(n16692), .B(n16691), .ZN(
        n16693) );
  AOI211_X1 U19886 ( .C1(n9571), .C2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n16694), .B(n16693), .ZN(n16695) );
  OAI211_X1 U19887 ( .C1(n10009), .C2(n16954), .A(n16696), .B(n16695), .ZN(
        n16697) );
  AOI211_X1 U19888 ( .C1(n17009), .C2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n16698), .B(n16697), .ZN(n16787) );
  AOI22_X1 U19889 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n16699) );
  OAI21_X1 U19890 ( .B1(n10740), .B2(n16700), .A(n16699), .ZN(n16711) );
  INV_X1 U19891 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n16989) );
  AOI22_X1 U19892 ( .A1(n17025), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17006), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n16709) );
  OAI22_X1 U19893 ( .A1(n16962), .A2(n16702), .B1(n16935), .B2(n16701), .ZN(
        n16707) );
  AOI22_X1 U19894 ( .A1(n9579), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n16705) );
  AOI22_X1 U19895 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n16704) );
  AOI22_X1 U19896 ( .A1(n16893), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9571), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n16703) );
  NAND3_X1 U19897 ( .A1(n16705), .A2(n16704), .A3(n16703), .ZN(n16706) );
  AOI211_X1 U19898 ( .C1(n16955), .C2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A(
        n16707), .B(n16706), .ZN(n16708) );
  OAI211_X1 U19899 ( .C1(n10797), .C2(n16989), .A(n16709), .B(n16708), .ZN(
        n16710) );
  AOI211_X1 U19900 ( .C1(n16903), .C2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n16711), .B(n16710), .ZN(n16796) );
  AOI22_X1 U19901 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n9585), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16721) );
  AOI22_X1 U19902 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n16991), .B1(
        P3_INSTQUEUE_REG_3__0__SCAN_IN), .B2(n17006), .ZN(n16720) );
  AOI22_X1 U19903 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n16893), .B1(
        P3_INSTQUEUE_REG_13__0__SCAN_IN), .B2(n17014), .ZN(n16719) );
  OAI22_X1 U19904 ( .A1(n18303), .A2(n9575), .B1(n17001), .B2(n18267), .ZN(
        n16717) );
  AOI22_X1 U19905 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__0__SCAN_IN), .B2(n10704), .ZN(n16715) );
  AOI22_X1 U19906 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17025), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16714) );
  AOI22_X1 U19907 ( .A1(n17009), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16734), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16713) );
  NAND2_X1 U19908 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n9571), .ZN(
        n16712) );
  NAND4_X1 U19909 ( .A1(n16715), .A2(n16714), .A3(n16713), .A4(n16712), .ZN(
        n16716) );
  AOI211_X1 U19910 ( .C1(n9579), .C2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n16717), .B(n16716), .ZN(n16718) );
  NAND4_X1 U19911 ( .A1(n16721), .A2(n16720), .A3(n16719), .A4(n16718), .ZN(
        n16801) );
  AOI22_X1 U19912 ( .A1(n16955), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16733) );
  AOI22_X1 U19913 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16722) );
  OAI21_X1 U19914 ( .B1(n9575), .B2(n18293), .A(n16722), .ZN(n16731) );
  INV_X1 U19915 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18081) );
  OAI22_X1 U19916 ( .A1(n10797), .A2(n18081), .B1(n16935), .B2(n16724), .ZN(
        n16725) );
  AOI21_X1 U19917 ( .B1(n17014), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n16725), .ZN(n16729) );
  AOI22_X1 U19918 ( .A1(n17009), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17025), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16728) );
  AOI22_X1 U19919 ( .A1(n9577), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10887), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16727) );
  AOI22_X1 U19920 ( .A1(n16893), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9571), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16726) );
  NAND4_X1 U19921 ( .A1(n16729), .A2(n16728), .A3(n16727), .A4(n16726), .ZN(
        n16730) );
  AOI211_X1 U19922 ( .C1(n16992), .C2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n16731), .B(n16730), .ZN(n16732) );
  OAI211_X1 U19923 ( .C1(n17011), .C2(n20923), .A(n16733), .B(n16732), .ZN(
        n16802) );
  NAND2_X1 U19924 ( .A1(n16801), .A2(n16802), .ZN(n16800) );
  NOR2_X1 U19925 ( .A1(n16796), .A2(n16800), .ZN(n16792) );
  AOI22_X1 U19926 ( .A1(n17006), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16744) );
  AOI22_X1 U19927 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17009), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16743) );
  AOI22_X1 U19928 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9571), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n16742) );
  OAI22_X1 U19929 ( .A1(n17001), .A2(n18274), .B1(n9575), .B2(n18309), .ZN(
        n16740) );
  AOI22_X1 U19930 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16738) );
  AOI22_X1 U19931 ( .A1(n9578), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16737) );
  AOI22_X1 U19932 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17025), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n16736) );
  NAND2_X1 U19933 ( .A1(n16734), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n16735) );
  NAND4_X1 U19934 ( .A1(n16738), .A2(n16737), .A3(n16736), .A4(n16735), .ZN(
        n16739) );
  AOI211_X1 U19935 ( .C1(n16965), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n16740), .B(n16739), .ZN(n16741) );
  NAND4_X1 U19936 ( .A1(n16744), .A2(n16743), .A3(n16742), .A4(n16741), .ZN(
        n16791) );
  NAND2_X1 U19937 ( .A1(n16792), .A2(n16791), .ZN(n16790) );
  NOR2_X1 U19938 ( .A1(n16787), .A2(n16790), .ZN(n16783) );
  AOI22_X1 U19939 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9579), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16754) );
  AOI22_X1 U19940 ( .A1(n17009), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16745) );
  OAI21_X1 U19941 ( .B1(n16756), .B2(n18063), .A(n16745), .ZN(n16752) );
  OAI22_X1 U19942 ( .A1(n17001), .A2(n18280), .B1(n16962), .B2(n16934), .ZN(
        n16746) );
  AOI21_X1 U19943 ( .B1(n17006), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n16746), .ZN(n16750) );
  AOI22_X1 U19944 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16749) );
  AOI22_X1 U19945 ( .A1(n17025), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16748) );
  AOI22_X1 U19946 ( .A1(n16893), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9571), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16747) );
  NAND4_X1 U19947 ( .A1(n16750), .A2(n16749), .A3(n16748), .A4(n16747), .ZN(
        n16751) );
  AOI211_X1 U19948 ( .C1(n16992), .C2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n16752), .B(n16751), .ZN(n16753) );
  OAI211_X1 U19949 ( .C1(n10797), .C2(n16834), .A(n16754), .B(n16753), .ZN(
        n16782) );
  NAND2_X1 U19950 ( .A1(n16783), .A2(n16782), .ZN(n16781) );
  NOR2_X1 U19951 ( .A1(n16777), .A2(n16781), .ZN(n16776) );
  NAND2_X1 U19952 ( .A1(n16774), .A2(n16776), .ZN(n16768) );
  AOI22_X1 U19953 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17009), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16755) );
  OAI21_X1 U19954 ( .B1(n16756), .B2(n18081), .A(n16755), .ZN(n16766) );
  AOI22_X1 U19955 ( .A1(n16734), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16763) );
  OAI22_X1 U19956 ( .A1(n17001), .A2(n18293), .B1(n16987), .B2(n20923), .ZN(
        n16761) );
  AOI22_X1 U19957 ( .A1(n17025), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9577), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16759) );
  AOI22_X1 U19958 ( .A1(n17006), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16758) );
  AOI22_X1 U19959 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9571), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16757) );
  NAND3_X1 U19960 ( .A1(n16759), .A2(n16758), .A3(n16757), .ZN(n16760) );
  AOI211_X1 U19961 ( .C1(n9585), .C2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n16761), .B(n16760), .ZN(n16762) );
  OAI211_X1 U19962 ( .C1(n15418), .C2(n16764), .A(n16763), .B(n16762), .ZN(
        n16765) );
  AOI211_X1 U19963 ( .C1(n16903), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n16766), .B(n16765), .ZN(n16767) );
  XNOR2_X1 U19964 ( .A(n16768), .B(n16767), .ZN(n17066) );
  OAI22_X1 U19965 ( .A1(n16770), .A2(n16769), .B1(n17066), .B2(n17054), .ZN(
        P3_U2673) );
  NAND2_X1 U19966 ( .A1(n18077), .A2(n16861), .ZN(n16844) );
  NOR2_X2 U19967 ( .A1(n16845), .A2(n16844), .ZN(n16829) );
  NAND2_X1 U19968 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16829), .ZN(n16817) );
  NOR2_X2 U19969 ( .A1(n16817), .A2(n16771), .ZN(n16799) );
  NAND2_X1 U19970 ( .A1(n16799), .A2(P3_EBX_REG_23__SCAN_IN), .ZN(n16795) );
  XNOR2_X1 U19971 ( .A(n16776), .B(n16774), .ZN(n17071) );
  NAND3_X1 U19972 ( .A1(n16778), .A2(P3_EBX_REG_29__SCAN_IN), .A3(n17054), 
        .ZN(n16775) );
  OAI221_X1 U19973 ( .B1(n16778), .B2(P3_EBX_REG_29__SCAN_IN), .C1(n17054), 
        .C2(n17071), .A(n16775), .ZN(P3_U2674) );
  NAND2_X1 U19974 ( .A1(n16789), .A2(P3_EBX_REG_27__SCAN_IN), .ZN(n16784) );
  AOI21_X1 U19975 ( .B1(n16777), .B2(n16781), .A(n16776), .ZN(n17072) );
  AND2_X1 U19976 ( .A1(n17054), .A2(n16778), .ZN(n16779) );
  AOI22_X1 U19977 ( .A1(n17043), .A2(n17072), .B1(P3_EBX_REG_28__SCAN_IN), 
        .B2(n16779), .ZN(n16780) );
  OAI21_X1 U19978 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n16784), .A(n16780), .ZN(
        P3_U2675) );
  OAI21_X1 U19979 ( .B1(n16783), .B2(n16782), .A(n16781), .ZN(n17080) );
  OAI211_X1 U19980 ( .C1(n16789), .C2(P3_EBX_REG_27__SCAN_IN), .A(n17054), .B(
        n16784), .ZN(n16785) );
  OAI21_X1 U19981 ( .B1(n17080), .B2(n17054), .A(n16785), .ZN(P3_U2676) );
  INV_X1 U19982 ( .A(n16786), .ZN(n16794) );
  AOI21_X1 U19983 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17054), .A(n16794), .ZN(
        n16788) );
  XNOR2_X1 U19984 ( .A(n16787), .B(n16790), .ZN(n17085) );
  OAI22_X1 U19985 ( .A1(n16789), .A2(n16788), .B1(n17054), .B2(n17085), .ZN(
        P3_U2677) );
  AOI21_X1 U19986 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17054), .A(n16798), .ZN(
        n16793) );
  OAI21_X1 U19987 ( .B1(n16792), .B2(n16791), .A(n16790), .ZN(n17090) );
  OAI22_X1 U19988 ( .A1(n16794), .A2(n16793), .B1(n17054), .B2(n17090), .ZN(
        P3_U2678) );
  INV_X1 U19989 ( .A(n16795), .ZN(n16804) );
  AOI21_X1 U19990 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17054), .A(n16804), .ZN(
        n16797) );
  XNOR2_X1 U19991 ( .A(n16796), .B(n16800), .ZN(n17095) );
  OAI22_X1 U19992 ( .A1(n16798), .A2(n16797), .B1(n17054), .B2(n17095), .ZN(
        P3_U2679) );
  AOI21_X1 U19993 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17054), .A(n16799), .ZN(
        n16803) );
  OAI21_X1 U19994 ( .B1(n16802), .B2(n16801), .A(n16800), .ZN(n17100) );
  OAI22_X1 U19995 ( .A1(n16804), .A2(n16803), .B1(n17054), .B2(n17100), .ZN(
        P3_U2680) );
  AOI22_X1 U19996 ( .A1(n9578), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17006), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16805) );
  OAI21_X1 U19997 ( .B1(n16987), .B2(n18323), .A(n16805), .ZN(n16815) );
  AOI22_X1 U19998 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16813) );
  AOI22_X1 U19999 ( .A1(n16955), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9571), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16806) );
  INV_X1 U20000 ( .A(n16806), .ZN(n16811) );
  AOI22_X1 U20001 ( .A1(n16988), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16809) );
  AOI22_X1 U20002 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17025), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16808) );
  AOI22_X1 U20003 ( .A1(n16893), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16807) );
  NAND3_X1 U20004 ( .A1(n16809), .A2(n16808), .A3(n16807), .ZN(n16810) );
  AOI211_X1 U20005 ( .C1(n9585), .C2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        n16811), .B(n16810), .ZN(n16812) );
  OAI211_X1 U20006 ( .C1(n10797), .C2(n18074), .A(n16813), .B(n16812), .ZN(
        n16814) );
  AOI211_X1 U20007 ( .C1(n17009), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n16815), .B(n16814), .ZN(n17104) );
  NAND3_X1 U20008 ( .A1(n16817), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17054), 
        .ZN(n16816) );
  OAI221_X1 U20009 ( .B1(n16817), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17054), 
        .C2(n17104), .A(n16816), .ZN(P3_U2681) );
  NAND2_X1 U20010 ( .A1(n17054), .A2(n16818), .ZN(n16846) );
  AOI22_X1 U20011 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16828) );
  AOI22_X1 U20012 ( .A1(n9577), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16820) );
  AOI22_X1 U20013 ( .A1(n17009), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17010), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16819) );
  OAI211_X1 U20014 ( .C1(n15418), .C2(n20936), .A(n16820), .B(n16819), .ZN(
        n16826) );
  AOI22_X1 U20015 ( .A1(n17025), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17006), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16824) );
  AOI22_X1 U20016 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16823) );
  AOI22_X1 U20017 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16822) );
  NAND2_X1 U20018 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n16821) );
  NAND4_X1 U20019 ( .A1(n16824), .A2(n16823), .A3(n16822), .A4(n16821), .ZN(
        n16825) );
  AOI211_X1 U20020 ( .C1(n9571), .C2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n16826), .B(n16825), .ZN(n16827) );
  OAI211_X1 U20021 ( .C1(n10797), .C2(n18069), .A(n16828), .B(n16827), .ZN(
        n17109) );
  AOI22_X1 U20022 ( .A1(n17043), .A2(n17109), .B1(n16829), .B2(n16831), .ZN(
        n16830) );
  OAI21_X1 U20023 ( .B1(n16831), .B2(n16846), .A(n16830), .ZN(P3_U2682) );
  AOI22_X1 U20024 ( .A1(n17006), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16842) );
  AOI22_X1 U20025 ( .A1(n9579), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16833) );
  AOI22_X1 U20026 ( .A1(n17010), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16832) );
  OAI211_X1 U20027 ( .C1(n15418), .C2(n16834), .A(n16833), .B(n16832), .ZN(
        n16840) );
  AOI22_X1 U20028 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17012), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16838) );
  AOI22_X1 U20029 ( .A1(n17009), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9585), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16837) );
  AOI22_X1 U20030 ( .A1(n17025), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16836) );
  NAND2_X1 U20031 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n16835) );
  NAND4_X1 U20032 ( .A1(n16838), .A2(n16837), .A3(n16836), .A4(n16835), .ZN(
        n16839) );
  AOI211_X1 U20033 ( .C1(n17014), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n16840), .B(n16839), .ZN(n16841) );
  OAI211_X1 U20034 ( .C1(n10797), .C2(n18063), .A(n16842), .B(n16841), .ZN(
        n17114) );
  NAND2_X1 U20035 ( .A1(n17043), .A2(n17114), .ZN(n16843) );
  OAI221_X1 U20036 ( .B1(n16846), .B2(n16845), .C1(n16846), .C2(n16844), .A(
        n16843), .ZN(P3_U2683) );
  AOI21_X1 U20037 ( .B1(n16873), .B2(n16847), .A(n17043), .ZN(n16848) );
  INV_X1 U20038 ( .A(n16848), .ZN(n16860) );
  AOI22_X1 U20039 ( .A1(n9579), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16849) );
  OAI21_X1 U20040 ( .B1(n10741), .B2(n16850), .A(n16849), .ZN(n16859) );
  INV_X1 U20041 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16957) );
  AOI22_X1 U20042 ( .A1(n16955), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16857) );
  OAI22_X1 U20043 ( .A1(n10797), .A2(n18057), .B1(n16958), .B2(n16954), .ZN(
        n16855) );
  AOI22_X1 U20044 ( .A1(n17009), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16853) );
  AOI22_X1 U20045 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17025), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16852) );
  AOI22_X1 U20046 ( .A1(n16893), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16851) );
  NAND3_X1 U20047 ( .A1(n16853), .A2(n16852), .A3(n16851), .ZN(n16854) );
  AOI211_X1 U20048 ( .C1(n10704), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n16855), .B(n16854), .ZN(n16856) );
  OAI211_X1 U20049 ( .C1(n10009), .C2(n16957), .A(n16857), .B(n16856), .ZN(
        n16858) );
  AOI211_X1 U20050 ( .C1(n16903), .C2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n16859), .B(n16858), .ZN(n17124) );
  OAI22_X1 U20051 ( .A1(n16861), .A2(n16860), .B1(n17124), .B2(n17054), .ZN(
        P3_U2684) );
  OAI22_X1 U20052 ( .A1(n10797), .A2(n20898), .B1(n10741), .B2(n20868), .ZN(
        n16872) );
  AOI22_X1 U20053 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17025), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16870) );
  AOI22_X1 U20054 ( .A1(n9577), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16869) );
  OAI22_X1 U20055 ( .A1(n17001), .A2(n16862), .B1(n9575), .B2(n18274), .ZN(
        n16867) );
  AOI22_X1 U20056 ( .A1(n17013), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n16865) );
  AOI22_X1 U20057 ( .A1(n17009), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9585), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n16864) );
  AOI22_X1 U20058 ( .A1(n16893), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n16863) );
  NAND3_X1 U20059 ( .A1(n16865), .A2(n16864), .A3(n16863), .ZN(n16866) );
  AOI211_X1 U20060 ( .C1(n9571), .C2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n16867), .B(n16866), .ZN(n16868) );
  NAND3_X1 U20061 ( .A1(n16870), .A2(n16869), .A3(n16868), .ZN(n16871) );
  AOI211_X1 U20062 ( .C1(n16992), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n16872), .B(n16871), .ZN(n17128) );
  OAI21_X1 U20063 ( .B1(n16890), .B2(P3_EBX_REG_18__SCAN_IN), .A(n16873), .ZN(
        n16874) );
  AOI22_X1 U20064 ( .A1(n17043), .A2(n17128), .B1(n16874), .B2(n17054), .ZN(
        P3_U2685) );
  AOI21_X1 U20065 ( .B1(n16876), .B2(n16875), .A(n17043), .ZN(n16877) );
  INV_X1 U20066 ( .A(n16877), .ZN(n16889) );
  AOI22_X1 U20067 ( .A1(n9578), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17006), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n16878) );
  OAI21_X1 U20068 ( .B1(n9575), .B2(n18271), .A(n16878), .ZN(n16888) );
  INV_X1 U20069 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18049) );
  AOI22_X1 U20070 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n16886) );
  OAI22_X1 U20071 ( .A1(n15418), .A2(n16989), .B1(n16935), .B2(n16879), .ZN(
        n16884) );
  AOI22_X1 U20072 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16882) );
  AOI22_X1 U20073 ( .A1(n17009), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17025), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n16881) );
  AOI22_X1 U20074 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9571), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n16880) );
  NAND3_X1 U20075 ( .A1(n16882), .A2(n16881), .A3(n16880), .ZN(n16883) );
  AOI211_X1 U20076 ( .C1(n16955), .C2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n16884), .B(n16883), .ZN(n16885) );
  OAI211_X1 U20077 ( .C1(n10797), .C2(n18049), .A(n16886), .B(n16885), .ZN(
        n16887) );
  AOI211_X1 U20078 ( .C1(n16992), .C2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n16888), .B(n16887), .ZN(n17134) );
  OAI22_X1 U20079 ( .A1(n16890), .A2(n16889), .B1(n17134), .B2(n17054), .ZN(
        P3_U2686) );
  NAND2_X1 U20080 ( .A1(n18077), .A2(n16891), .ZN(n16916) );
  AOI22_X1 U20081 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n9577), .B1(
        P3_INSTQUEUE_REG_14__0__SCAN_IN), .B2(n10704), .ZN(n16892) );
  OAI21_X1 U20082 ( .B1(n10740), .B2(n20895), .A(n16892), .ZN(n16902) );
  INV_X1 U20083 ( .A(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17008) );
  AOI22_X1 U20084 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n17006), .B1(
        P3_INSTQUEUE_REG_4__0__SCAN_IN), .B2(n9571), .ZN(n16900) );
  INV_X1 U20085 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18045) );
  OAI22_X1 U20086 ( .A1(n18045), .A2(n10797), .B1(n18303), .B2(n16987), .ZN(
        n16898) );
  AOI22_X1 U20087 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9585), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16896) );
  AOI22_X1 U20088 ( .A1(n17025), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__0__SCAN_IN), .B2(n16988), .ZN(n16895) );
  AOI22_X1 U20089 ( .A1(n16893), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n16894) );
  NAND3_X1 U20090 ( .A1(n16896), .A2(n16895), .A3(n16894), .ZN(n16897) );
  AOI211_X1 U20091 ( .C1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .C2(n17010), .A(
        n16898), .B(n16897), .ZN(n16899) );
  OAI211_X1 U20092 ( .C1(n17008), .C2(n17001), .A(n16900), .B(n16899), .ZN(
        n16901) );
  AOI211_X1 U20093 ( .C1(n16903), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n16902), .B(n16901), .ZN(n17140) );
  NAND3_X1 U20094 ( .A1(n16916), .A2(P3_EBX_REG_16__SCAN_IN), .A3(n17054), 
        .ZN(n16904) );
  OAI221_X1 U20095 ( .B1(n16916), .B2(P3_EBX_REG_16__SCAN_IN), .C1(n17054), 
        .C2(n17140), .A(n16904), .ZN(P3_U2687) );
  AOI22_X1 U20096 ( .A1(n17010), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16905) );
  OAI21_X1 U20097 ( .B1(n16987), .B2(n18293), .A(n16905), .ZN(n16915) );
  INV_X1 U20098 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16913) );
  AOI22_X1 U20099 ( .A1(n16734), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17006), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16912) );
  AOI22_X1 U20100 ( .A1(n10758), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16906) );
  OAI21_X1 U20101 ( .B1(n16962), .B2(n20923), .A(n16906), .ZN(n16910) );
  AOI22_X1 U20102 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9585), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16908) );
  AOI22_X1 U20103 ( .A1(n17025), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16907) );
  OAI211_X1 U20104 ( .C1(n15418), .C2(n18081), .A(n16908), .B(n16907), .ZN(
        n16909) );
  AOI211_X1 U20105 ( .C1(n9571), .C2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n16910), .B(n16909), .ZN(n16911) );
  OAI211_X1 U20106 ( .C1(n17011), .C2(n16913), .A(n16912), .B(n16911), .ZN(
        n16914) );
  AOI211_X1 U20107 ( .C1(n9579), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n16915), .B(n16914), .ZN(n17144) );
  OAI211_X1 U20108 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n16917), .A(n17054), .B(
        n16916), .ZN(n16918) );
  OAI21_X1 U20109 ( .B1(n17144), .B2(n17054), .A(n16918), .ZN(P3_U2688) );
  INV_X1 U20110 ( .A(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16920) );
  AOI22_X1 U20111 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17025), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16919) );
  OAI21_X1 U20112 ( .B1(n9575), .B2(n16920), .A(n16919), .ZN(n16930) );
  AOI22_X1 U20113 ( .A1(n17006), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16928) );
  OAI22_X1 U20114 ( .A1(n16987), .A2(n18286), .B1(n16935), .B2(n16921), .ZN(
        n16926) );
  AOI22_X1 U20115 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16924) );
  AOI22_X1 U20116 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9577), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16923) );
  AOI22_X1 U20117 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9571), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16922) );
  NAND3_X1 U20118 ( .A1(n16924), .A2(n16923), .A3(n16922), .ZN(n16925) );
  AOI211_X1 U20119 ( .C1(n16734), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n16926), .B(n16925), .ZN(n16927) );
  OAI211_X1 U20120 ( .C1(n15418), .C2(n18074), .A(n16928), .B(n16927), .ZN(
        n16929) );
  AOI211_X1 U20121 ( .C1(n17009), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n16930), .B(n16929), .ZN(n17150) );
  OAI22_X1 U20122 ( .A1(n17043), .A2(n16932), .B1(P3_EBX_REG_14__SCAN_IN), 
        .B2(n17176), .ZN(n16931) );
  OAI21_X1 U20123 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n16932), .A(n16931), .ZN(
        n16933) );
  OAI21_X1 U20124 ( .B1(n17150), .B2(n17054), .A(n16933), .ZN(P3_U2689) );
  OAI22_X1 U20125 ( .A1(n17001), .A2(n16936), .B1(n16935), .B2(n16934), .ZN(
        n16947) );
  AOI22_X1 U20126 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17025), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16945) );
  AOI22_X1 U20127 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17009), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16944) );
  INV_X1 U20128 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16938) );
  AOI22_X1 U20129 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16937) );
  OAI21_X1 U20130 ( .B1(n10797), .B2(n16938), .A(n16937), .ZN(n16942) );
  AOI22_X1 U20131 ( .A1(n9579), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16940) );
  AOI22_X1 U20132 ( .A1(n17006), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16939) );
  OAI211_X1 U20133 ( .C1(n15418), .C2(n18063), .A(n16940), .B(n16939), .ZN(
        n16941) );
  AOI211_X1 U20134 ( .C1(n9571), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n16942), .B(n16941), .ZN(n16943) );
  NAND3_X1 U20135 ( .A1(n16945), .A2(n16944), .A3(n16943), .ZN(n16946) );
  AOI211_X1 U20136 ( .C1(n17014), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n16947), .B(n16946), .ZN(n17155) );
  INV_X1 U20137 ( .A(n16948), .ZN(n16949) );
  OAI21_X1 U20138 ( .B1(n16971), .B2(P3_EBX_REG_12__SCAN_IN), .A(n16949), .ZN(
        n16950) );
  AOI22_X1 U20139 ( .A1(n17043), .A2(n17155), .B1(n16950), .B2(n17054), .ZN(
        P3_U2691) );
  AOI21_X1 U20140 ( .B1(n16982), .B2(n16951), .A(n17043), .ZN(n16952) );
  INV_X1 U20141 ( .A(n16952), .ZN(n16970) );
  AOI22_X1 U20142 ( .A1(n16988), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16953) );
  OAI21_X1 U20143 ( .B1(n10740), .B2(n16954), .A(n16953), .ZN(n16969) );
  INV_X1 U20144 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18313) );
  AOI22_X1 U20145 ( .A1(n16734), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17006), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16967) );
  AOI22_X1 U20146 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16956) );
  OAI21_X1 U20147 ( .B1(n16958), .B2(n16957), .A(n16956), .ZN(n16964) );
  AOI22_X1 U20148 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16960) );
  AOI22_X1 U20149 ( .A1(n17025), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16959) );
  OAI211_X1 U20150 ( .C1(n16962), .C2(n16961), .A(n16960), .B(n16959), .ZN(
        n16963) );
  AOI211_X1 U20151 ( .C1(n16965), .C2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A(
        n16964), .B(n16963), .ZN(n16966) );
  OAI211_X1 U20152 ( .C1(n17011), .C2(n18313), .A(n16967), .B(n16966), .ZN(
        n16968) );
  AOI211_X1 U20153 ( .C1(n9578), .C2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n16969), .B(n16968), .ZN(n17159) );
  OAI22_X1 U20154 ( .A1(n16971), .A2(n16970), .B1(n17159), .B2(n17054), .ZN(
        P3_U2692) );
  AOI22_X1 U20155 ( .A1(n16734), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17006), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16981) );
  AOI22_X1 U20156 ( .A1(n17025), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17013), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16973) );
  AOI22_X1 U20157 ( .A1(n16991), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16972) );
  OAI211_X1 U20158 ( .C1(n15418), .C2(n20898), .A(n16973), .B(n16972), .ZN(
        n16979) );
  AOI22_X1 U20159 ( .A1(n16903), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16977) );
  AOI22_X1 U20160 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n9578), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n16976) );
  AOI22_X1 U20161 ( .A1(n17009), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n16975) );
  NAND2_X1 U20162 ( .A1(n9571), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n16974) );
  NAND4_X1 U20163 ( .A1(n16977), .A2(n16976), .A3(n16975), .A4(n16974), .ZN(
        n16978) );
  AOI211_X1 U20164 ( .C1(n17014), .C2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n16979), .B(n16978), .ZN(n16980) );
  OAI211_X1 U20165 ( .C1(n10009), .C2(n20868), .A(n16981), .B(n16980), .ZN(
        n17162) );
  INV_X1 U20166 ( .A(n17162), .ZN(n16984) );
  OAI21_X1 U20167 ( .B1(n17005), .B2(P3_EBX_REG_10__SCAN_IN), .A(n16982), .ZN(
        n16983) );
  AOI22_X1 U20168 ( .A1(n17043), .A2(n16984), .B1(n16983), .B2(n17054), .ZN(
        P3_U2693) );
  OAI21_X1 U20169 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n16985), .A(n17054), .ZN(
        n17004) );
  AOI22_X1 U20170 ( .A1(n9585), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10704), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n16986) );
  OAI21_X1 U20171 ( .B1(n16987), .B2(n18271), .A(n16986), .ZN(n17003) );
  INV_X1 U20172 ( .A(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17000) );
  AOI22_X1 U20173 ( .A1(n17025), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n16988), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n16999) );
  OAI22_X1 U20174 ( .A1(n15418), .A2(n18049), .B1(n10741), .B2(n16989), .ZN(
        n16997) );
  AOI22_X1 U20175 ( .A1(n16990), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9578), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n16995) );
  AOI22_X1 U20176 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n16991), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16994) );
  AOI22_X1 U20177 ( .A1(n17014), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9571), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n16993) );
  NAND3_X1 U20178 ( .A1(n16995), .A2(n16994), .A3(n16993), .ZN(n16996) );
  AOI211_X1 U20179 ( .C1(n16734), .C2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A(
        n16997), .B(n16996), .ZN(n16998) );
  OAI211_X1 U20180 ( .C1(n17001), .C2(n17000), .A(n16999), .B(n16998), .ZN(
        n17002) );
  AOI211_X1 U20181 ( .C1(n17009), .C2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A(
        n17003), .B(n17002), .ZN(n17168) );
  OAI22_X1 U20182 ( .A1(n17005), .A2(n17004), .B1(n17168), .B2(n17054), .ZN(
        P3_U2694) );
  AOI22_X1 U20183 ( .A1(n9578), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17006), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17007) );
  OAI21_X1 U20184 ( .B1(n17008), .B2(n9575), .A(n17007), .ZN(n17024) );
  INV_X1 U20185 ( .A(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17022) );
  AOI22_X1 U20186 ( .A1(n16734), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__0__SCAN_IN), .B2(n17010), .ZN(n17021) );
  OAI22_X1 U20187 ( .A1(n17011), .A2(n18303), .B1(n18045), .B2(n15418), .ZN(
        n17019) );
  AOI22_X1 U20188 ( .A1(n17012), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9585), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17017) );
  AOI22_X1 U20189 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n10704), .B1(
        P3_INSTQUEUE_REG_9__0__SCAN_IN), .B2(n17013), .ZN(n17016) );
  AOI22_X1 U20190 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n9571), .B1(
        n17014), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17015) );
  NAND3_X1 U20191 ( .A1(n17017), .A2(n17016), .A3(n17015), .ZN(n17018) );
  AOI211_X1 U20192 ( .C1(n16955), .C2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n17019), .B(n17018), .ZN(n17020) );
  OAI211_X1 U20193 ( .C1(n10740), .C2(n17022), .A(n17021), .B(n17020), .ZN(
        n17023) );
  AOI211_X1 U20194 ( .C1(n17025), .C2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A(
        n17024), .B(n17023), .ZN(n17175) );
  OR2_X1 U20195 ( .A1(n17043), .A2(n17026), .ZN(n17030) );
  AOI21_X1 U20196 ( .B1(n18077), .B2(n17026), .A(P3_EBX_REG_8__SCAN_IN), .ZN(
        n17027) );
  AOI21_X1 U20197 ( .B1(n17030), .B2(P3_EBX_REG_8__SCAN_IN), .A(n17027), .ZN(
        n17028) );
  INV_X1 U20198 ( .A(n17028), .ZN(n17029) );
  OAI21_X1 U20199 ( .B1(n17175), .B2(n17054), .A(n17029), .ZN(P3_U2695) );
  NOR2_X1 U20200 ( .A1(n17176), .A2(n17032), .ZN(n17033) );
  AOI21_X1 U20201 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17033), .A(
        P3_EBX_REG_7__SCAN_IN), .ZN(n17031) );
  OAI22_X1 U20202 ( .A1(n17031), .A2(n17030), .B1(n18081), .B2(n17054), .ZN(
        P3_U2696) );
  NAND2_X1 U20203 ( .A1(n17054), .A2(n17032), .ZN(n17035) );
  AOI22_X1 U20204 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n17043), .B1(
        n17033), .B2(n20863), .ZN(n17034) );
  OAI21_X1 U20205 ( .B1(n20863), .B2(n17035), .A(n17034), .ZN(P3_U2697) );
  NOR2_X1 U20206 ( .A1(n17040), .A2(P3_EBX_REG_5__SCAN_IN), .ZN(n17036) );
  OAI22_X1 U20207 ( .A1(n17036), .A2(n17035), .B1(n18069), .B2(n17054), .ZN(
        P3_U2698) );
  AOI21_X1 U20208 ( .B1(n17041), .B2(n17037), .A(n17043), .ZN(n17038) );
  INV_X1 U20209 ( .A(n17038), .ZN(n17039) );
  OAI22_X1 U20210 ( .A1(n17040), .A2(n17039), .B1(n18063), .B2(n17054), .ZN(
        P3_U2699) );
  OAI21_X1 U20211 ( .B1(n17048), .B2(P3_EBX_REG_3__SCAN_IN), .A(n17041), .ZN(
        n17042) );
  AOI22_X1 U20212 ( .A1(n17043), .A2(n18057), .B1(n17042), .B2(n17054), .ZN(
        P3_U2700) );
  AOI21_X1 U20213 ( .B1(n17045), .B2(n17044), .A(n17043), .ZN(n17046) );
  INV_X1 U20214 ( .A(n17046), .ZN(n17047) );
  OAI22_X1 U20215 ( .A1(n17048), .A2(n17047), .B1(n20898), .B2(n17054), .ZN(
        P3_U2701) );
  INV_X1 U20216 ( .A(n17049), .ZN(n17050) );
  NAND2_X1 U20217 ( .A1(n18077), .A2(n17050), .ZN(n17053) );
  OAI222_X1 U20218 ( .A1(n17053), .A2(n17052), .B1(n17051), .B2(n17050), .C1(
        n18049), .C2(n17054), .ZN(P3_U2702) );
  AND2_X1 U20219 ( .A1(n20934), .A2(n17053), .ZN(n17055) );
  OAI22_X1 U20220 ( .A1(n17056), .A2(n17055), .B1(n18045), .B2(n17054), .ZN(
        P3_U2703) );
  INV_X1 U20221 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17212) );
  INV_X1 U20222 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17218) );
  INV_X1 U20223 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17323) );
  INV_X1 U20224 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17261) );
  NAND2_X1 U20225 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .ZN(n17178) );
  NOR2_X1 U20226 ( .A1(n17261), .A2(n17178), .ZN(n17057) );
  NAND4_X1 U20227 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_7__SCAN_IN), 
        .A3(P3_EAX_REG_6__SCAN_IN), .A4(n17057), .ZN(n17145) );
  INV_X1 U20228 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17243) );
  INV_X1 U20229 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17245) );
  INV_X1 U20230 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17303) );
  NAND2_X1 U20231 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .ZN(n17146) );
  NOR4_X1 U20232 ( .A1(n17243), .A2(n17245), .A3(n17303), .A4(n17146), .ZN(
        n17058) );
  NOR2_X2 U20233 ( .A1(n17323), .A2(n17147), .ZN(n17141) );
  NAND2_X1 U20234 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_21__SCAN_IN), 
        .ZN(n17102) );
  NAND4_X1 U20235 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n17059)
         );
  NAND2_X1 U20236 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17097), .ZN(n17096) );
  NAND2_X1 U20237 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17092), .ZN(n17091) );
  NOR2_X2 U20238 ( .A1(n17218), .A2(n17086), .ZN(n17081) );
  NAND2_X1 U20239 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17081), .ZN(n17077) );
  NOR2_X2 U20240 ( .A1(n17212), .A2(n17073), .ZN(n17067) );
  NAND2_X1 U20241 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17067), .ZN(n17063) );
  NAND3_X1 U20242 ( .A1(n17199), .A2(P3_EAX_REG_31__SCAN_IN), .A3(n17063), 
        .ZN(n17062) );
  NAND2_X1 U20243 ( .A1(n17060), .A2(n17172), .ZN(n17103) );
  NAND2_X1 U20244 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17135), .ZN(n17061) );
  OAI211_X1 U20245 ( .C1(P3_EAX_REG_31__SCAN_IN), .C2(n17063), .A(n17062), .B(
        n17061), .ZN(P3_U2704) );
  NAND2_X1 U20246 ( .A1(n18066), .A2(n17172), .ZN(n17119) );
  AOI22_X1 U20247 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17136), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17135), .ZN(n17065) );
  OAI211_X1 U20248 ( .C1(n17067), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17199), .B(
        n17063), .ZN(n17064) );
  OAI211_X1 U20249 ( .C1(n17066), .C2(n17190), .A(n17065), .B(n17064), .ZN(
        P3_U2705) );
  AOI22_X1 U20250 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17136), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17135), .ZN(n17070) );
  AOI211_X1 U20251 ( .C1(n17212), .C2(n17073), .A(n17067), .B(n17172), .ZN(
        n17068) );
  INV_X1 U20252 ( .A(n17068), .ZN(n17069) );
  OAI211_X1 U20253 ( .C1(n17190), .C2(n17071), .A(n17070), .B(n17069), .ZN(
        P3_U2706) );
  AOI22_X1 U20254 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17136), .B1(n17072), .B2(
        n17204), .ZN(n17076) );
  OAI211_X1 U20255 ( .C1(n17074), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17199), .B(
        n17073), .ZN(n17075) );
  OAI211_X1 U20256 ( .C1(n17103), .C2(n14851), .A(n17076), .B(n17075), .ZN(
        P3_U2707) );
  AOI22_X1 U20257 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17136), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17135), .ZN(n17079) );
  OAI211_X1 U20258 ( .C1(n17081), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17199), .B(
        n17077), .ZN(n17078) );
  OAI211_X1 U20259 ( .C1(n17190), .C2(n17080), .A(n17079), .B(n17078), .ZN(
        P3_U2708) );
  AOI22_X1 U20260 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17136), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17135), .ZN(n17084) );
  AOI211_X1 U20261 ( .C1(n17218), .C2(n17086), .A(n17081), .B(n17172), .ZN(
        n17082) );
  INV_X1 U20262 ( .A(n17082), .ZN(n17083) );
  OAI211_X1 U20263 ( .C1(n17190), .C2(n17085), .A(n17084), .B(n17083), .ZN(
        P3_U2709) );
  AOI22_X1 U20264 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17136), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17135), .ZN(n17089) );
  OAI211_X1 U20265 ( .C1(n17087), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17199), .B(
        n17086), .ZN(n17088) );
  OAI211_X1 U20266 ( .C1(n17190), .C2(n17090), .A(n17089), .B(n17088), .ZN(
        P3_U2710) );
  AOI22_X1 U20267 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17136), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17135), .ZN(n17094) );
  OAI211_X1 U20268 ( .C1(n17092), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17199), .B(
        n17091), .ZN(n17093) );
  OAI211_X1 U20269 ( .C1(n17190), .C2(n17095), .A(n17094), .B(n17093), .ZN(
        P3_U2711) );
  AOI22_X1 U20270 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17136), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17135), .ZN(n17099) );
  OAI211_X1 U20271 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17097), .A(n17199), .B(
        n17096), .ZN(n17098) );
  OAI211_X1 U20272 ( .C1(n17190), .C2(n17100), .A(n17099), .B(n17098), .ZN(
        P3_U2712) );
  INV_X1 U20273 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n20858) );
  INV_X1 U20274 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17274) );
  NOR3_X1 U20275 ( .A1(n17176), .A2(n17137), .A3(n17274), .ZN(n17129) );
  NAND2_X1 U20276 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17129), .ZN(n17125) );
  NAND2_X1 U20277 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17121), .ZN(n17120) );
  NAND2_X1 U20278 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17116), .ZN(n17115) );
  NAND2_X1 U20279 ( .A1(n17199), .A2(n17115), .ZN(n17110) );
  OAI21_X1 U20280 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17101), .A(n17110), .ZN(
        n17107) );
  NOR3_X1 U20281 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17102), .A3(n17120), .ZN(
        n17106) );
  OAI22_X1 U20282 ( .A1(n17104), .A2(n17190), .B1(n14894), .B2(n17103), .ZN(
        n17105) );
  AOI211_X1 U20283 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n17107), .A(n17106), .B(
        n17105), .ZN(n17108) );
  OAI21_X1 U20284 ( .B1(n20858), .B2(n17119), .A(n17108), .ZN(P3_U2713) );
  AOI22_X1 U20285 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n17135), .B1(n17204), .B2(
        n17109), .ZN(n17113) );
  INV_X1 U20286 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18065) );
  INV_X1 U20287 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17227) );
  OAI22_X1 U20288 ( .A1(n18065), .A2(n17119), .B1(n17227), .B2(n17110), .ZN(
        n17111) );
  INV_X1 U20289 ( .A(n17111), .ZN(n17112) );
  OAI211_X1 U20290 ( .C1(P3_EAX_REG_21__SCAN_IN), .C2(n17115), .A(n17113), .B(
        n17112), .ZN(P3_U2714) );
  AOI22_X1 U20291 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17135), .B1(n17204), .B2(
        n17114), .ZN(n17118) );
  OAI211_X1 U20292 ( .C1(n17116), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17199), .B(
        n17115), .ZN(n17117) );
  OAI211_X1 U20293 ( .C1(n17119), .C2(n18058), .A(n17118), .B(n17117), .ZN(
        P3_U2715) );
  AOI22_X1 U20294 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17136), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17135), .ZN(n17123) );
  OAI211_X1 U20295 ( .C1(n17121), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17199), .B(
        n17120), .ZN(n17122) );
  OAI211_X1 U20296 ( .C1(n17124), .C2(n17190), .A(n17123), .B(n17122), .ZN(
        P3_U2716) );
  AOI22_X1 U20297 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17136), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17135), .ZN(n17127) );
  OAI211_X1 U20298 ( .C1(n17129), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17199), .B(
        n17125), .ZN(n17126) );
  OAI211_X1 U20299 ( .C1(n17128), .C2(n17190), .A(n17127), .B(n17126), .ZN(
        P3_U2717) );
  AOI22_X1 U20300 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17136), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17135), .ZN(n17133) );
  INV_X1 U20301 ( .A(n17137), .ZN(n17131) );
  INV_X1 U20302 ( .A(n17129), .ZN(n17130) );
  OAI211_X1 U20303 ( .C1(n17131), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17199), .B(
        n17130), .ZN(n17132) );
  OAI211_X1 U20304 ( .C1(n17134), .C2(n17190), .A(n17133), .B(n17132), .ZN(
        P3_U2718) );
  AOI22_X1 U20305 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17136), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17135), .ZN(n17139) );
  OAI211_X1 U20306 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17141), .A(n17199), .B(
        n17137), .ZN(n17138) );
  OAI211_X1 U20307 ( .C1(n17140), .C2(n17190), .A(n17139), .B(n17138), .ZN(
        P3_U2719) );
  AOI21_X1 U20308 ( .B1(n17323), .B2(n17147), .A(n17141), .ZN(n17142) );
  AOI22_X1 U20309 ( .A1(n17205), .A2(BUF2_REG_15__SCAN_IN), .B1(n17142), .B2(
        n17199), .ZN(n17143) );
  OAI21_X1 U20310 ( .B1(n17144), .B2(n17190), .A(n17143), .ZN(P3_U2720) );
  INV_X1 U20311 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17241) );
  NOR3_X1 U20312 ( .A1(n17176), .A2(n17206), .A3(n17145), .ZN(n17181) );
  NAND2_X1 U20313 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17181), .ZN(n17166) );
  NOR2_X1 U20314 ( .A1(n17146), .A2(n17166), .ZN(n17158) );
  INV_X1 U20315 ( .A(n17158), .ZN(n17163) );
  NOR2_X1 U20316 ( .A1(n17245), .A2(n17163), .ZN(n17161) );
  NAND2_X1 U20317 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17161), .ZN(n17151) );
  NOR2_X1 U20318 ( .A1(n17241), .A2(n17151), .ZN(n17154) );
  INV_X1 U20319 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17318) );
  AOI22_X1 U20320 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17205), .B1(n17154), .B2(
        n17318), .ZN(n17149) );
  NAND3_X1 U20321 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17199), .A3(n17147), 
        .ZN(n17148) );
  OAI211_X1 U20322 ( .C1(n17150), .C2(n17190), .A(n17149), .B(n17148), .ZN(
        P3_U2721) );
  INV_X1 U20323 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17316) );
  INV_X1 U20324 ( .A(n17151), .ZN(n17157) );
  AOI21_X1 U20325 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17199), .A(n17157), .ZN(
        n17153) );
  OAI222_X1 U20326 ( .A1(n17202), .A2(n17316), .B1(n17154), .B2(n17153), .C1(
        n17190), .C2(n17152), .ZN(P3_U2722) );
  INV_X1 U20327 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17312) );
  AOI21_X1 U20328 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17199), .A(n17161), .ZN(
        n17156) );
  OAI222_X1 U20329 ( .A1(n17202), .A2(n17312), .B1(n17157), .B2(n17156), .C1(
        n17190), .C2(n17155), .ZN(P3_U2723) );
  INV_X1 U20330 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17309) );
  AOI21_X1 U20331 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17199), .A(n17158), .ZN(
        n17160) );
  OAI222_X1 U20332 ( .A1(n17202), .A2(n17309), .B1(n17161), .B2(n17160), .C1(
        n17190), .C2(n17159), .ZN(P3_U2724) );
  AOI22_X1 U20333 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17205), .B1(n17204), .B2(
        n17162), .ZN(n17165) );
  INV_X1 U20334 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17249) );
  NOR2_X1 U20335 ( .A1(n17249), .A2(n17166), .ZN(n17170) );
  OAI211_X1 U20336 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n17170), .A(n17199), .B(
        n17163), .ZN(n17164) );
  NAND2_X1 U20337 ( .A1(n17165), .A2(n17164), .ZN(P3_U2725) );
  INV_X1 U20338 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17305) );
  OAI21_X1 U20339 ( .B1(n17249), .B2(n17172), .A(n17166), .ZN(n17167) );
  INV_X1 U20340 ( .A(n17167), .ZN(n17169) );
  OAI222_X1 U20341 ( .A1(n17202), .A2(n17305), .B1(n17170), .B2(n17169), .C1(
        n17190), .C2(n17168), .ZN(P3_U2726) );
  AOI22_X1 U20342 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17205), .B1(n17181), .B2(
        n17303), .ZN(n17174) );
  OR3_X1 U20343 ( .A1(n17303), .A2(n17172), .A3(n17171), .ZN(n17173) );
  OAI211_X1 U20344 ( .C1(n17175), .C2(n17190), .A(n17174), .B(n17173), .ZN(
        P3_U2727) );
  INV_X1 U20345 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n20860) );
  INV_X1 U20346 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17254) );
  NOR2_X1 U20347 ( .A1(n17176), .A2(n17206), .ZN(n17177) );
  NAND2_X1 U20348 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17177), .ZN(n17196) );
  NOR2_X1 U20349 ( .A1(n17178), .A2(n17196), .ZN(n17192) );
  NAND2_X1 U20350 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17192), .ZN(n17182) );
  NOR2_X1 U20351 ( .A1(n17254), .A2(n17182), .ZN(n17185) );
  AOI21_X1 U20352 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17199), .A(n17185), .ZN(
        n17180) );
  OAI222_X1 U20353 ( .A1(n20860), .A2(n17202), .B1(n17181), .B2(n17180), .C1(
        n17190), .C2(n17179), .ZN(P3_U2728) );
  INV_X1 U20354 ( .A(n17182), .ZN(n17188) );
  AOI21_X1 U20355 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17199), .A(n17188), .ZN(
        n17184) );
  OAI222_X1 U20356 ( .A1(n20858), .A2(n17202), .B1(n17185), .B2(n17184), .C1(
        n17190), .C2(n17183), .ZN(P3_U2729) );
  AOI21_X1 U20357 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17199), .A(n17192), .ZN(
        n17187) );
  OAI222_X1 U20358 ( .A1(n18065), .A2(n17202), .B1(n17188), .B2(n17187), .C1(
        n17190), .C2(n17186), .ZN(P3_U2730) );
  INV_X1 U20359 ( .A(n17196), .ZN(n17197) );
  AOI22_X1 U20360 ( .A1(n17197), .A2(P3_EAX_REG_3__SCAN_IN), .B1(
        P3_EAX_REG_4__SCAN_IN), .B2(n17199), .ZN(n17191) );
  OAI222_X1 U20361 ( .A1(n18058), .A2(n17202), .B1(n17192), .B2(n17191), .C1(
        n17190), .C2(n17189), .ZN(P3_U2731) );
  NAND3_X1 U20362 ( .A1(n17199), .A2(P3_EAX_REG_3__SCAN_IN), .A3(n17196), .ZN(
        n17195) );
  AOI22_X1 U20363 ( .A1(n17205), .A2(BUF2_REG_3__SCAN_IN), .B1(n17204), .B2(
        n17193), .ZN(n17194) );
  OAI211_X1 U20364 ( .C1(P3_EAX_REG_3__SCAN_IN), .C2(n17196), .A(n17195), .B(
        n17194), .ZN(P3_U2732) );
  INV_X1 U20365 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18050) );
  AOI21_X1 U20366 ( .B1(n17206), .B2(n17261), .A(n17197), .ZN(n17200) );
  INV_X1 U20367 ( .A(n10754), .ZN(n17198) );
  AOI22_X1 U20368 ( .A1(n17200), .A2(n17199), .B1(n17204), .B2(n17198), .ZN(
        n17201) );
  OAI21_X1 U20369 ( .B1(n18050), .B2(n17202), .A(n17201), .ZN(P3_U2733) );
  AOI22_X1 U20370 ( .A1(n17205), .A2(BUF2_REG_1__SCAN_IN), .B1(n17204), .B2(
        n17203), .ZN(n17209) );
  OAI211_X1 U20371 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(n17207), .A(n17199), .B(
        n17206), .ZN(n17208) );
  NAND2_X1 U20372 ( .A1(n17209), .A2(n17208), .ZN(P3_U2734) );
  INV_X1 U20373 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17290) );
  NOR2_X1 U20374 ( .A1(n17266), .A2(n18040), .ZN(n17231) );
  AOI22_X1 U20375 ( .A1(n17264), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17210) );
  OAI21_X1 U20376 ( .B1(n17290), .B2(n17236), .A(n17210), .ZN(P3_U2737) );
  AOI22_X1 U20377 ( .A1(P3_UWORD_REG_13__SCAN_IN), .A2(n17264), .B1(n17263), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17211) );
  OAI21_X1 U20378 ( .B1(n17212), .B2(n17236), .A(n17211), .ZN(P3_U2738) );
  INV_X1 U20379 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17214) );
  AOI22_X1 U20380 ( .A1(n17264), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17213) );
  OAI21_X1 U20381 ( .B1(n17214), .B2(n17236), .A(n17213), .ZN(P3_U2739) );
  INV_X1 U20382 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17216) );
  AOI22_X1 U20383 ( .A1(P3_UWORD_REG_11__SCAN_IN), .A2(n17264), .B1(n17263), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17215) );
  OAI21_X1 U20384 ( .B1(n17216), .B2(n17236), .A(n17215), .ZN(P3_U2740) );
  AOI22_X1 U20385 ( .A1(n17264), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17217) );
  OAI21_X1 U20386 ( .B1(n17218), .B2(n17236), .A(n17217), .ZN(P3_U2741) );
  INV_X1 U20387 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17220) );
  AOI22_X1 U20388 ( .A1(n17264), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17219) );
  OAI21_X1 U20389 ( .B1(n17220), .B2(n17236), .A(n17219), .ZN(P3_U2742) );
  INV_X1 U20390 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17283) );
  AOI22_X1 U20391 ( .A1(n17264), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17221) );
  OAI21_X1 U20392 ( .B1(n17283), .B2(n17236), .A(n17221), .ZN(P3_U2743) );
  INV_X1 U20393 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17223) );
  AOI22_X1 U20394 ( .A1(P3_DATAO_REG_23__SCAN_IN), .A2(n17263), .B1(n17264), 
        .B2(P3_UWORD_REG_7__SCAN_IN), .ZN(n17222) );
  OAI21_X1 U20395 ( .B1(n17223), .B2(n17236), .A(n17222), .ZN(P3_U2744) );
  INV_X1 U20396 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17225) );
  AOI22_X1 U20397 ( .A1(n17264), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17224) );
  OAI21_X1 U20398 ( .B1(n17225), .B2(n17236), .A(n17224), .ZN(P3_U2745) );
  AOI22_X1 U20399 ( .A1(n17264), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17226) );
  OAI21_X1 U20400 ( .B1(n17227), .B2(n17236), .A(n17226), .ZN(P3_U2746) );
  INV_X1 U20401 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17229) );
  AOI22_X1 U20402 ( .A1(n17264), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17228) );
  OAI21_X1 U20403 ( .B1(n17229), .B2(n17236), .A(n17228), .ZN(P3_U2747) );
  INV_X1 U20404 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17277) );
  AOI22_X1 U20405 ( .A1(n17264), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17230) );
  OAI21_X1 U20406 ( .B1(n17277), .B2(n17236), .A(n17230), .ZN(P3_U2748) );
  INV_X1 U20407 ( .A(P3_UWORD_REG_2__SCAN_IN), .ZN(n20848) );
  AOI22_X1 U20408 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17231), .B1(n17263), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17232) );
  OAI21_X1 U20409 ( .B1(n20848), .B2(n17233), .A(n17232), .ZN(P3_U2749) );
  AOI22_X1 U20410 ( .A1(n17264), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17234) );
  OAI21_X1 U20411 ( .B1(n17274), .B2(n17236), .A(n17234), .ZN(P3_U2750) );
  INV_X1 U20412 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17237) );
  AOI22_X1 U20413 ( .A1(n17264), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17235) );
  OAI21_X1 U20414 ( .B1(n17237), .B2(n17236), .A(n17235), .ZN(P3_U2751) );
  AOI22_X1 U20415 ( .A1(n17264), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17238) );
  OAI21_X1 U20416 ( .B1(n17323), .B2(n17266), .A(n17238), .ZN(P3_U2752) );
  AOI22_X1 U20417 ( .A1(n17264), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17239) );
  OAI21_X1 U20418 ( .B1(n17318), .B2(n17266), .A(n17239), .ZN(P3_U2753) );
  AOI22_X1 U20419 ( .A1(n17264), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17240) );
  OAI21_X1 U20420 ( .B1(n17241), .B2(n17266), .A(n17240), .ZN(P3_U2754) );
  AOI22_X1 U20421 ( .A1(n17264), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17242) );
  OAI21_X1 U20422 ( .B1(n17243), .B2(n17266), .A(n17242), .ZN(P3_U2755) );
  AOI22_X1 U20423 ( .A1(n17264), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17244) );
  OAI21_X1 U20424 ( .B1(n17245), .B2(n17266), .A(n17244), .ZN(P3_U2756) );
  INV_X1 U20425 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17247) );
  AOI22_X1 U20426 ( .A1(P3_LWORD_REG_10__SCAN_IN), .A2(n17264), .B1(n17263), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17246) );
  OAI21_X1 U20427 ( .B1(n17247), .B2(n17266), .A(n17246), .ZN(P3_U2757) );
  AOI22_X1 U20428 ( .A1(n17264), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17248) );
  OAI21_X1 U20429 ( .B1(n17249), .B2(n17266), .A(n17248), .ZN(P3_U2758) );
  AOI22_X1 U20430 ( .A1(n17264), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17250) );
  OAI21_X1 U20431 ( .B1(n17303), .B2(n17266), .A(n17250), .ZN(P3_U2759) );
  INV_X1 U20432 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17252) );
  AOI22_X1 U20433 ( .A1(n17264), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17251) );
  OAI21_X1 U20434 ( .B1(n17252), .B2(n17266), .A(n17251), .ZN(P3_U2760) );
  AOI22_X1 U20435 ( .A1(n17264), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17253) );
  OAI21_X1 U20436 ( .B1(n17254), .B2(n17266), .A(n17253), .ZN(P3_U2761) );
  INV_X1 U20437 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17256) );
  AOI22_X1 U20438 ( .A1(n17264), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17255) );
  OAI21_X1 U20439 ( .B1(n17256), .B2(n17266), .A(n17255), .ZN(P3_U2762) );
  INV_X1 U20440 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17258) );
  AOI22_X1 U20441 ( .A1(n17264), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17257) );
  OAI21_X1 U20442 ( .B1(n17258), .B2(n17266), .A(n17257), .ZN(P3_U2763) );
  INV_X1 U20443 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17297) );
  AOI22_X1 U20444 ( .A1(n17264), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17259) );
  OAI21_X1 U20445 ( .B1(n17297), .B2(n17266), .A(n17259), .ZN(P3_U2764) );
  AOI22_X1 U20446 ( .A1(n17264), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17260) );
  OAI21_X1 U20447 ( .B1(n17261), .B2(n17266), .A(n17260), .ZN(P3_U2765) );
  INV_X1 U20448 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17293) );
  AOI22_X1 U20449 ( .A1(n17264), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17262) );
  OAI21_X1 U20450 ( .B1(n17293), .B2(n17266), .A(n17262), .ZN(P3_U2766) );
  AOI22_X1 U20451 ( .A1(n17264), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17263), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17265) );
  OAI21_X1 U20452 ( .B1(n17267), .B2(n17266), .A(n17265), .ZN(P3_U2767) );
  INV_X1 U20453 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18037) );
  OAI211_X1 U20454 ( .C1(n18697), .C2(n18046), .A(n17269), .B(n17268), .ZN(
        n17294) );
  NOR2_X1 U20455 ( .A1(n17319), .A2(n18046), .ZN(n17320) );
  NOR3_X1 U20456 ( .A1(n18702), .A2(n17271), .A3(n17270), .ZN(n17313) );
  AOI22_X1 U20457 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17310), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17319), .ZN(n17272) );
  OAI21_X1 U20458 ( .B1(n18037), .B2(n17315), .A(n17272), .ZN(P3_U2768) );
  INV_X1 U20459 ( .A(n17313), .ZN(n17322) );
  AOI22_X1 U20460 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17320), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17294), .ZN(n17273) );
  OAI21_X1 U20461 ( .B1(n17274), .B2(n17322), .A(n17273), .ZN(P3_U2769) );
  AOI22_X1 U20462 ( .A1(P3_UWORD_REG_2__SCAN_IN), .A2(n17319), .B1(
        P3_EAX_REG_18__SCAN_IN), .B2(n17310), .ZN(n17275) );
  OAI21_X1 U20463 ( .B1(n18050), .B2(n17315), .A(n17275), .ZN(P3_U2770) );
  AOI22_X1 U20464 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17320), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17294), .ZN(n17276) );
  OAI21_X1 U20465 ( .B1(n17277), .B2(n17322), .A(n17276), .ZN(P3_U2771) );
  AOI22_X1 U20466 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17310), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17319), .ZN(n17278) );
  OAI21_X1 U20467 ( .B1(n18058), .B2(n17315), .A(n17278), .ZN(P3_U2772) );
  AOI22_X1 U20468 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17310), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17319), .ZN(n17279) );
  OAI21_X1 U20469 ( .B1(n18065), .B2(n17315), .A(n17279), .ZN(P3_U2773) );
  AOI22_X1 U20470 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17310), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17319), .ZN(n17280) );
  OAI21_X1 U20471 ( .B1(n20858), .B2(n17315), .A(n17280), .ZN(P3_U2774) );
  AOI22_X1 U20472 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17310), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17294), .ZN(n17281) );
  OAI21_X1 U20473 ( .B1(n20860), .B2(n17315), .A(n17281), .ZN(P3_U2775) );
  AOI22_X1 U20474 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17320), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17294), .ZN(n17282) );
  OAI21_X1 U20475 ( .B1(n17283), .B2(n17322), .A(n17282), .ZN(P3_U2776) );
  AOI22_X1 U20476 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17313), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17294), .ZN(n17284) );
  OAI21_X1 U20477 ( .B1(n17305), .B2(n17315), .A(n17284), .ZN(P3_U2777) );
  INV_X1 U20478 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17307) );
  AOI22_X1 U20479 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17310), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17294), .ZN(n17285) );
  OAI21_X1 U20480 ( .B1(n17307), .B2(n17315), .A(n17285), .ZN(P3_U2778) );
  AOI22_X1 U20481 ( .A1(P3_UWORD_REG_11__SCAN_IN), .A2(n17319), .B1(
        P3_EAX_REG_27__SCAN_IN), .B2(n17310), .ZN(n17286) );
  OAI21_X1 U20482 ( .B1(n17309), .B2(n17315), .A(n17286), .ZN(P3_U2779) );
  AOI22_X1 U20483 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17313), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17294), .ZN(n17287) );
  OAI21_X1 U20484 ( .B1(n17312), .B2(n17315), .A(n17287), .ZN(P3_U2780) );
  AOI22_X1 U20485 ( .A1(P3_UWORD_REG_13__SCAN_IN), .A2(n17319), .B1(
        P3_EAX_REG_29__SCAN_IN), .B2(n17310), .ZN(n17288) );
  OAI21_X1 U20486 ( .B1(n17316), .B2(n17315), .A(n17288), .ZN(P3_U2781) );
  AOI22_X1 U20487 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17320), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17319), .ZN(n17289) );
  OAI21_X1 U20488 ( .B1(n17290), .B2(n17322), .A(n17289), .ZN(P3_U2782) );
  AOI22_X1 U20489 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17310), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17294), .ZN(n17291) );
  OAI21_X1 U20490 ( .B1(n18037), .B2(n17315), .A(n17291), .ZN(P3_U2783) );
  AOI22_X1 U20491 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17320), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17319), .ZN(n17292) );
  OAI21_X1 U20492 ( .B1(n17293), .B2(n17322), .A(n17292), .ZN(P3_U2784) );
  AOI22_X1 U20493 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17313), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17294), .ZN(n17295) );
  OAI21_X1 U20494 ( .B1(n18050), .B2(n17315), .A(n17295), .ZN(P3_U2785) );
  AOI22_X1 U20495 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17320), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17319), .ZN(n17296) );
  OAI21_X1 U20496 ( .B1(n17297), .B2(n17322), .A(n17296), .ZN(P3_U2786) );
  AOI22_X1 U20497 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17310), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17319), .ZN(n17298) );
  OAI21_X1 U20498 ( .B1(n18058), .B2(n17315), .A(n17298), .ZN(P3_U2787) );
  AOI22_X1 U20499 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17310), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17319), .ZN(n17299) );
  OAI21_X1 U20500 ( .B1(n18065), .B2(n17315), .A(n17299), .ZN(P3_U2788) );
  AOI22_X1 U20501 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17310), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17319), .ZN(n17300) );
  OAI21_X1 U20502 ( .B1(n20858), .B2(n17315), .A(n17300), .ZN(P3_U2789) );
  AOI22_X1 U20503 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17310), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17319), .ZN(n17301) );
  OAI21_X1 U20504 ( .B1(n20860), .B2(n17315), .A(n17301), .ZN(P3_U2790) );
  AOI22_X1 U20505 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17320), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17319), .ZN(n17302) );
  OAI21_X1 U20506 ( .B1(n17303), .B2(n17322), .A(n17302), .ZN(P3_U2791) );
  AOI22_X1 U20507 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17310), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17319), .ZN(n17304) );
  OAI21_X1 U20508 ( .B1(n17305), .B2(n17315), .A(n17304), .ZN(P3_U2792) );
  AOI22_X1 U20509 ( .A1(P3_LWORD_REG_10__SCAN_IN), .A2(n17319), .B1(
        P3_EAX_REG_10__SCAN_IN), .B2(n17310), .ZN(n17306) );
  OAI21_X1 U20510 ( .B1(n17307), .B2(n17315), .A(n17306), .ZN(P3_U2793) );
  AOI22_X1 U20511 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17313), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17319), .ZN(n17308) );
  OAI21_X1 U20512 ( .B1(n17309), .B2(n17315), .A(n17308), .ZN(P3_U2794) );
  AOI22_X1 U20513 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17310), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17319), .ZN(n17311) );
  OAI21_X1 U20514 ( .B1(n17312), .B2(n17315), .A(n17311), .ZN(P3_U2795) );
  AOI22_X1 U20515 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17313), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17319), .ZN(n17314) );
  OAI21_X1 U20516 ( .B1(n17316), .B2(n17315), .A(n17314), .ZN(P3_U2796) );
  AOI22_X1 U20517 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17320), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17319), .ZN(n17317) );
  OAI21_X1 U20518 ( .B1(n17318), .B2(n17322), .A(n17317), .ZN(P3_U2797) );
  AOI22_X1 U20519 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17320), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17319), .ZN(n17321) );
  OAI21_X1 U20520 ( .B1(n17323), .B2(n17322), .A(n17321), .ZN(P3_U2798) );
  INV_X1 U20521 ( .A(n17483), .ZN(n17500) );
  AOI211_X1 U20522 ( .C1(n17326), .C2(n17325), .A(n17324), .B(n17611), .ZN(
        n17336) );
  NOR3_X1 U20523 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17527), .A3(
        n17329), .ZN(n17346) );
  INV_X1 U20524 ( .A(n17445), .ZN(n17354) );
  OAI21_X1 U20525 ( .B1(n17327), .B2(n18564), .A(n9594), .ZN(n17328) );
  AOI21_X1 U20526 ( .B1(n17671), .B2(n17329), .A(n17328), .ZN(n17364) );
  OAI21_X1 U20527 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17354), .A(
        n17364), .ZN(n17347) );
  OAI21_X1 U20528 ( .B1(n17346), .B2(n17347), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17333) );
  INV_X1 U20529 ( .A(n17527), .ZN(n17395) );
  NAND3_X1 U20530 ( .A1(n17331), .A2(n17330), .A3(n17395), .ZN(n17332) );
  NAND3_X1 U20531 ( .A1(n17334), .A2(n17333), .A3(n17332), .ZN(n17335) );
  AOI211_X1 U20532 ( .C1(n17554), .C2(n17337), .A(n17336), .B(n17335), .ZN(
        n17339) );
  NAND2_X1 U20533 ( .A1(n17568), .A2(n17700), .ZN(n17442) );
  AOI22_X1 U20534 ( .A1(n17608), .A2(n17702), .B1(n17685), .B2(n17703), .ZN(
        n17359) );
  NAND2_X1 U20535 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17359), .ZN(
        n17348) );
  NAND3_X1 U20536 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17442), .A3(
        n17348), .ZN(n17338) );
  OAI211_X1 U20537 ( .C1(n17340), .C2(n17500), .A(n17339), .B(n17338), .ZN(
        P3_U2802) );
  NAND2_X1 U20538 ( .A1(n17342), .A2(n17341), .ZN(n17343) );
  XOR2_X1 U20539 ( .A(n17597), .B(n17343), .Z(n17711) );
  OAI22_X1 U20540 ( .A1(n18017), .A2(n18633), .B1(n17506), .B2(n17344), .ZN(
        n17345) );
  AOI211_X1 U20541 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17347), .A(
        n17346), .B(n17345), .ZN(n17351) );
  OAI21_X1 U20542 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17349), .A(
        n17348), .ZN(n17350) );
  OAI211_X1 U20543 ( .C1(n17711), .C2(n17611), .A(n17351), .B(n17350), .ZN(
        P3_U2803) );
  AOI21_X1 U20544 ( .B1(n17352), .B2(n18434), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17363) );
  INV_X1 U20545 ( .A(n17353), .ZN(n17355) );
  NAND2_X2 U20546 ( .A1(n17506), .A2(n17354), .ZN(n17688) );
  AOI22_X1 U20547 ( .A1(n17821), .A2(P3_REIP_REG_26__SCAN_IN), .B1(n17355), 
        .B2(n17688), .ZN(n17362) );
  NOR2_X1 U20548 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17356), .ZN(
        n17716) );
  AOI21_X1 U20549 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17358), .A(
        n17357), .ZN(n17718) );
  OAI22_X1 U20550 ( .A1(n17359), .A2(n17714), .B1(n17718), .B2(n17611), .ZN(
        n17360) );
  AOI21_X1 U20551 ( .B1(n17483), .B2(n17716), .A(n17360), .ZN(n17361) );
  OAI211_X1 U20552 ( .C1(n17364), .C2(n17363), .A(n17362), .B(n17361), .ZN(
        P3_U2804) );
  NOR2_X1 U20553 ( .A1(n17847), .A2(n17389), .ZN(n17736) );
  OAI221_X1 U20554 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n17736), .A(n17365), .ZN(
        n17734) );
  OAI21_X1 U20555 ( .B1(n17366), .B2(n18262), .A(n9594), .ZN(n17367) );
  AOI21_X1 U20556 ( .B1(n17369), .B2(n17368), .A(n17367), .ZN(n17398) );
  OAI21_X1 U20557 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18564), .A(
        n17398), .ZN(n17386) );
  NOR2_X1 U20558 ( .A1(n17527), .A2(n17370), .ZN(n17388) );
  OAI211_X1 U20559 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17388), .B(n17371), .ZN(n17372) );
  NAND2_X1 U20560 ( .A1(n17815), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17726) );
  OAI211_X1 U20561 ( .C1(n17506), .C2(n17373), .A(n17372), .B(n17726), .ZN(
        n17380) );
  OAI21_X1 U20562 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17375), .A(
        n17374), .ZN(n17728) );
  OAI21_X1 U20563 ( .B1(n17597), .B2(n17377), .A(n17376), .ZN(n17378) );
  XOR2_X1 U20564 ( .A(n17378), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17729) );
  OAI22_X1 U20565 ( .A1(n17568), .A2(n17728), .B1(n17611), .B2(n17729), .ZN(
        n17379) );
  AOI211_X1 U20566 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17386), .A(
        n17380), .B(n17379), .ZN(n17381) );
  OAI21_X1 U20567 ( .B1(n17700), .B2(n17734), .A(n17381), .ZN(P3_U2805) );
  AOI21_X1 U20568 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17383), .A(
        n17382), .ZN(n17749) );
  INV_X1 U20569 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18627) );
  OAI22_X1 U20570 ( .A1(n17909), .A2(n18627), .B1(n17506), .B2(n17384), .ZN(
        n17385) );
  AOI221_X1 U20571 ( .B1(n17388), .B2(n17387), .C1(n17386), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17385), .ZN(n17391) );
  NAND2_X1 U20572 ( .A1(n17735), .A2(n17608), .ZN(n17392) );
  OAI21_X1 U20573 ( .B1(n17736), .B2(n17700), .A(n17392), .ZN(n17407) );
  NOR2_X1 U20574 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17389), .ZN(
        n17746) );
  AOI22_X1 U20575 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17407), .B1(
        n17483), .B2(n17746), .ZN(n17390) );
  OAI211_X1 U20576 ( .C1(n17749), .C2(n17611), .A(n17391), .B(n17390), .ZN(
        P3_U2806) );
  NOR2_X1 U20577 ( .A1(n17736), .A2(n17700), .ZN(n17394) );
  INV_X1 U20578 ( .A(n17392), .ZN(n17393) );
  AOI22_X1 U20579 ( .A1(n17758), .A2(n17394), .B1(n17836), .B2(n17393), .ZN(
        n17411) );
  INV_X1 U20580 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18626) );
  NOR2_X1 U20581 ( .A1(n18017), .A2(n18626), .ZN(n17752) );
  NAND2_X1 U20582 ( .A1(n17396), .A2(n17395), .ZN(n17431) );
  NOR2_X1 U20583 ( .A1(n17397), .A2(n17431), .ZN(n17400) );
  INV_X1 U20584 ( .A(n17398), .ZN(n17399) );
  MUX2_X1 U20585 ( .A(n17400), .B(n17399), .S(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .Z(n17401) );
  AOI211_X1 U20586 ( .C1(n17554), .C2(n17402), .A(n17752), .B(n17401), .ZN(
        n17409) );
  AOI22_X1 U20587 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17597), .B1(
        n17422), .B2(n17404), .ZN(n17405) );
  NAND2_X1 U20588 ( .A1(n17403), .A2(n17405), .ZN(n17406) );
  XOR2_X1 U20589 ( .A(n17406), .B(n17756), .Z(n17753) );
  AOI22_X1 U20590 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17407), .B1(
        n17538), .B2(n17753), .ZN(n17408) );
  OAI211_X1 U20591 ( .C1(n17411), .C2(n17410), .A(n17409), .B(n17408), .ZN(
        P3_U2807) );
  OAI22_X1 U20592 ( .A1(n17836), .A2(n17568), .B1(n17758), .B2(n17700), .ZN(
        n17469) );
  AOI21_X1 U20593 ( .B1(n17424), .B2(n17442), .A(n17469), .ZN(n17436) );
  INV_X1 U20594 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17417) );
  AOI211_X1 U20595 ( .C1(n17430), .C2(n17417), .A(n17412), .B(n17431), .ZN(
        n17419) );
  AOI21_X1 U20596 ( .B1(n17671), .B2(n17413), .A(n17601), .ZN(n17414) );
  OAI21_X1 U20597 ( .B1(n17415), .B2(n18564), .A(n17414), .ZN(n17449) );
  AOI21_X1 U20598 ( .B1(n17445), .B2(n17443), .A(n17449), .ZN(n17429) );
  OAI22_X1 U20599 ( .A1(n17429), .A2(n17417), .B1(n17506), .B2(n17416), .ZN(
        n17418) );
  AOI211_X1 U20600 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n17815), .A(n17419), 
        .B(n17418), .ZN(n17426) );
  INV_X1 U20601 ( .A(n17403), .ZN(n17421) );
  AOI221_X1 U20602 ( .B1(n9580), .B2(n17422), .C1(n17424), .C2(n17422), .A(
        n17421), .ZN(n17423) );
  XOR2_X1 U20603 ( .A(n17423), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(
        n17770) );
  NOR2_X1 U20604 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17424), .ZN(
        n17768) );
  AOI22_X1 U20605 ( .A1(n17538), .A2(n17770), .B1(n17483), .B2(n17768), .ZN(
        n17425) );
  OAI211_X1 U20606 ( .C1(n17436), .C2(n17427), .A(n17426), .B(n17425), .ZN(
        P3_U2808) );
  NAND2_X1 U20607 ( .A1(n17778), .A2(n17775), .ZN(n17774) );
  NAND2_X1 U20608 ( .A1(n17441), .A2(n17483), .ZN(n17464) );
  INV_X1 U20609 ( .A(n17428), .ZN(n17439) );
  NAND2_X1 U20610 ( .A1(n17815), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n17781) );
  OAI221_X1 U20611 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17431), .C1(
        n17430), .C2(n17429), .A(n17781), .ZN(n17438) );
  NOR3_X1 U20612 ( .A1(n17812), .A2(n17597), .A3(n17432), .ZN(n17453) );
  INV_X1 U20613 ( .A(n17433), .ZN(n17471) );
  AOI22_X1 U20614 ( .A1(n17778), .A2(n17453), .B1(n17434), .B2(n17471), .ZN(
        n17435) );
  XOR2_X1 U20615 ( .A(n17435), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .Z(
        n17783) );
  OAI22_X1 U20616 ( .A1(n17436), .A2(n17775), .B1(n17783), .B2(n17611), .ZN(
        n17437) );
  AOI211_X1 U20617 ( .C1(n17554), .C2(n17439), .A(n17438), .B(n17437), .ZN(
        n17440) );
  OAI21_X1 U20618 ( .B1(n17774), .B2(n17464), .A(n17440), .ZN(P3_U2809) );
  NAND2_X1 U20619 ( .A1(n17441), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n17785) );
  AOI21_X1 U20620 ( .B1(n17442), .B2(n17785), .A(n17469), .ZN(n17463) );
  OAI21_X1 U20621 ( .B1(n17444), .B2(n18262), .A(n17443), .ZN(n17448) );
  AOI21_X1 U20622 ( .B1(n17506), .B2(n17354), .A(n17446), .ZN(n17447) );
  INV_X1 U20623 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18619) );
  NOR2_X1 U20624 ( .A1(n18017), .A2(n18619), .ZN(n17790) );
  AOI211_X1 U20625 ( .C1(n17449), .C2(n17448), .A(n17447), .B(n17790), .ZN(
        n17452) );
  OAI221_X1 U20626 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17470), 
        .C1(n17800), .C2(n17453), .A(n17403), .ZN(n17450) );
  XOR2_X1 U20627 ( .A(n17787), .B(n17450), .Z(n17791) );
  NOR2_X1 U20628 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17785), .ZN(
        n17784) );
  AOI22_X1 U20629 ( .A1(n17538), .A2(n17791), .B1(n17483), .B2(n17784), .ZN(
        n17451) );
  OAI211_X1 U20630 ( .C1(n17463), .C2(n17787), .A(n17452), .B(n17451), .ZN(
        P3_U2810) );
  AOI21_X1 U20631 ( .B1(n17471), .B2(n17470), .A(n17453), .ZN(n17454) );
  XOR2_X1 U20632 ( .A(n17800), .B(n17454), .Z(n17796) );
  AOI21_X1 U20633 ( .B1(n17671), .B2(n17456), .A(n17601), .ZN(n17477) );
  OAI21_X1 U20634 ( .B1(n17455), .B2(n18564), .A(n17477), .ZN(n17467) );
  AOI22_X1 U20635 ( .A1(n17821), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17467), .ZN(n17459) );
  NOR2_X1 U20636 ( .A1(n17527), .A2(n17456), .ZN(n17468) );
  OAI211_X1 U20637 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17468), .B(n17457), .ZN(n17458) );
  OAI211_X1 U20638 ( .C1(n17506), .C2(n17460), .A(n17459), .B(n17458), .ZN(
        n17461) );
  AOI21_X1 U20639 ( .B1(n17538), .B2(n17796), .A(n17461), .ZN(n17462) );
  OAI221_X1 U20640 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17464), 
        .C1(n17800), .C2(n17463), .A(n17462), .ZN(P3_U2811) );
  NAND2_X1 U20641 ( .A1(n17806), .A2(n17812), .ZN(n17818) );
  OAI22_X1 U20642 ( .A1(n17909), .A2(n18615), .B1(n17506), .B2(n17465), .ZN(
        n17466) );
  AOI221_X1 U20643 ( .B1(n17468), .B2(n20909), .C1(n17467), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17466), .ZN(n17474) );
  INV_X1 U20644 ( .A(n17469), .ZN(n17499) );
  OAI21_X1 U20645 ( .B1(n17806), .B2(n17500), .A(n17499), .ZN(n17482) );
  AOI21_X1 U20646 ( .B1(n17557), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17470), .ZN(n17472) );
  XOR2_X1 U20647 ( .A(n17472), .B(n17471), .Z(n17814) );
  AOI22_X1 U20648 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17482), .B1(
        n17538), .B2(n17814), .ZN(n17473) );
  OAI211_X1 U20649 ( .C1(n17500), .C2(n17818), .A(n17474), .B(n17473), .ZN(
        P3_U2812) );
  OAI21_X1 U20650 ( .B1(n17476), .B2(n17819), .A(n17475), .ZN(n17824) );
  INV_X1 U20651 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18614) );
  NOR2_X1 U20652 ( .A1(n17909), .A2(n18614), .ZN(n17481) );
  AOI221_X1 U20653 ( .B1(n17479), .B2(n17478), .C1(n18262), .C2(n17478), .A(
        n17477), .ZN(n17480) );
  AOI211_X1 U20654 ( .C1(n17538), .C2(n17824), .A(n17481), .B(n17480), .ZN(
        n17485) );
  OAI221_X1 U20655 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n17483), .A(n17482), .ZN(
        n17484) );
  OAI211_X1 U20656 ( .C1(n17680), .C2(n17486), .A(n17485), .B(n17484), .ZN(
        P3_U2813) );
  AOI21_X1 U20657 ( .B1(n17557), .B2(n9580), .A(n17487), .ZN(n17488) );
  XOR2_X1 U20658 ( .A(n17488), .B(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .Z(
        n17831) );
  INV_X1 U20659 ( .A(n17489), .ZN(n17490) );
  AOI21_X1 U20660 ( .B1(n17671), .B2(n17490), .A(n17601), .ZN(n17520) );
  OAI21_X1 U20661 ( .B1(n17491), .B2(n18564), .A(n17520), .ZN(n17508) );
  AOI22_X1 U20662 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17508), .B1(
        n17554), .B2(n17492), .ZN(n17496) );
  NOR3_X1 U20663 ( .A1(n17527), .A2(n17493), .A3(n17531), .ZN(n17510) );
  OAI211_X1 U20664 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17510), .B(n17494), .ZN(n17495) );
  OAI211_X1 U20665 ( .C1(n18611), .C2(n18017), .A(n17496), .B(n17495), .ZN(
        n17497) );
  AOI21_X1 U20666 ( .B1(n17538), .B2(n17831), .A(n17497), .ZN(n17498) );
  OAI221_X1 U20667 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17500), 
        .C1(n10903), .C2(n17499), .A(n17498), .ZN(P3_U2814) );
  NAND3_X1 U20668 ( .A1(n17542), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17502) );
  OAI21_X1 U20669 ( .B1(n17572), .B2(n17502), .A(n17501), .ZN(n17503) );
  OAI221_X1 U20670 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17860), 
        .C1(n9757), .C2(n17557), .A(n17503), .ZN(n17504) );
  XOR2_X1 U20671 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17504), .Z(
        n17843) );
  INV_X1 U20672 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17509) );
  OAI22_X1 U20673 ( .A1(n18017), .A2(n18609), .B1(n17506), .B2(n17505), .ZN(
        n17507) );
  AOI221_X1 U20674 ( .B1(n17510), .B2(n17509), .C1(n17508), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17507), .ZN(n17514) );
  NOR2_X1 U20675 ( .A1(n17836), .A2(n17568), .ZN(n17512) );
  NAND2_X1 U20676 ( .A1(n17850), .A2(n17523), .ZN(n17840) );
  NOR2_X1 U20677 ( .A1(n17758), .A2(n17700), .ZN(n17511) );
  NAND3_X1 U20678 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17851), .A3(
        n17567), .ZN(n17516) );
  NAND2_X1 U20679 ( .A1(n17850), .A2(n17516), .ZN(n17846) );
  AOI22_X1 U20680 ( .A1(n17512), .A2(n17840), .B1(n17511), .B2(n17846), .ZN(
        n17513) );
  OAI211_X1 U20681 ( .C1(n17611), .C2(n17843), .A(n17514), .B(n17513), .ZN(
        P3_U2815) );
  NOR2_X1 U20682 ( .A1(n17891), .A2(n17515), .ZN(n17517) );
  OAI21_X1 U20683 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17517), .A(
        n17516), .ZN(n17867) );
  NOR2_X1 U20684 ( .A1(n17531), .A2(n18262), .ZN(n17563) );
  AOI21_X1 U20685 ( .B1(n17528), .B2(n17563), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17519) );
  OAI22_X1 U20686 ( .A1(n17520), .A2(n17519), .B1(n17680), .B2(n17518), .ZN(
        n17525) );
  NAND2_X1 U20687 ( .A1(n17557), .A2(n10902), .ZN(n17586) );
  INV_X1 U20688 ( .A(n17586), .ZN(n17556) );
  AOI21_X1 U20689 ( .B1(n17556), .B2(n17851), .A(n17521), .ZN(n17522) );
  XOR2_X1 U20690 ( .A(n17522), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n17862) );
  OAI221_X1 U20691 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17851), 
        .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n10902), .A(n17523), .ZN(
        n17861) );
  OAI22_X1 U20692 ( .A1(n17862), .A2(n17611), .B1(n17568), .B2(n17861), .ZN(
        n17524) );
  AOI211_X1 U20693 ( .C1(n17821), .C2(P3_REIP_REG_14__SCAN_IN), .A(n17525), 
        .B(n17524), .ZN(n17526) );
  OAI21_X1 U20694 ( .B1(n17700), .B2(n17867), .A(n17526), .ZN(P3_U2816) );
  INV_X1 U20695 ( .A(n17853), .ZN(n17854) );
  NAND2_X1 U20696 ( .A1(n17854), .A2(n10902), .ZN(n17870) );
  NAND2_X1 U20697 ( .A1(n17854), .A2(n17567), .ZN(n17871) );
  AOI22_X1 U20698 ( .A1(n17608), .A2(n17870), .B1(n17685), .B2(n17871), .ZN(
        n17548) );
  OR2_X1 U20699 ( .A1(n17531), .A2(n17527), .ZN(n17547) );
  AOI211_X1 U20700 ( .C1(n17546), .C2(n17532), .A(n17528), .B(n17547), .ZN(
        n17534) );
  OAI21_X1 U20701 ( .B1(n17529), .B2(n18564), .A(n9594), .ZN(n17530) );
  AOI21_X1 U20702 ( .B1(n17671), .B2(n17531), .A(n17530), .ZN(n17545) );
  OAI22_X1 U20703 ( .A1(n17545), .A2(n17532), .B1(n17909), .B2(n18605), .ZN(
        n17533) );
  AOI211_X1 U20704 ( .C1(n17554), .C2(n17535), .A(n17534), .B(n17533), .ZN(
        n17540) );
  OAI22_X1 U20705 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17557), .B1(
        n17572), .B2(n17853), .ZN(n17536) );
  OAI21_X1 U20706 ( .B1(n17557), .B2(n17541), .A(n17536), .ZN(n17537) );
  XOR2_X1 U20707 ( .A(n17537), .B(n17857), .Z(n17877) );
  NOR2_X1 U20708 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17853), .ZN(
        n17876) );
  INV_X1 U20709 ( .A(n17566), .ZN(n17594) );
  AOI22_X1 U20710 ( .A1(n17538), .A2(n17877), .B1(n17876), .B2(n17594), .ZN(
        n17539) );
  OAI211_X1 U20711 ( .C1(n17548), .C2(n17857), .A(n17540), .B(n17539), .ZN(
        P3_U2817) );
  AOI21_X1 U20712 ( .B1(n17556), .B2(n17542), .A(n17541), .ZN(n17543) );
  XOR2_X1 U20713 ( .A(n17543), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n17888) );
  NAND2_X1 U20714 ( .A1(n17815), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n17544) );
  OAI221_X1 U20715 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17547), .C1(
        n17546), .C2(n17545), .A(n17544), .ZN(n17552) );
  NOR2_X1 U20716 ( .A1(n17566), .A2(n17881), .ZN(n17550) );
  INV_X1 U20717 ( .A(n17548), .ZN(n17549) );
  MUX2_X1 U20718 ( .A(n17550), .B(n17549), .S(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n17551) );
  AOI211_X1 U20719 ( .C1(n17554), .C2(n17553), .A(n17552), .B(n17551), .ZN(
        n17555) );
  OAI21_X1 U20720 ( .B1(n17888), .B2(n17611), .A(n17555), .ZN(P3_U2818) );
  NAND2_X1 U20721 ( .A1(n17895), .A2(n17556), .ZN(n17574) );
  OR2_X1 U20722 ( .A1(n17557), .A2(n17931), .ZN(n17585) );
  OR2_X1 U20723 ( .A1(n17585), .A2(n17581), .ZN(n17558) );
  NAND2_X1 U20724 ( .A1(n17574), .A2(n17558), .ZN(n17559) );
  XNOR2_X1 U20725 ( .A(n17559), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17902) );
  NOR2_X1 U20726 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17560), .ZN(
        n17889) );
  INV_X1 U20727 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18601) );
  NOR2_X1 U20728 ( .A1(n18017), .A2(n18601), .ZN(n17565) );
  INV_X1 U20729 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17606) );
  NOR4_X1 U20730 ( .A1(n17616), .A2(n17617), .A3(n17606), .A4(n18262), .ZN(
        n17589) );
  NAND2_X1 U20731 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17589), .ZN(
        n17588) );
  NOR2_X1 U20732 ( .A1(n17577), .A2(n17588), .ZN(n17576) );
  AOI21_X1 U20733 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17650), .A(
        n17576), .ZN(n17562) );
  OAI22_X1 U20734 ( .A1(n17563), .A2(n17562), .B1(n17680), .B2(n17561), .ZN(
        n17564) );
  AOI211_X1 U20735 ( .C1(n17889), .C2(n17594), .A(n17565), .B(n17564), .ZN(
        n17570) );
  NOR2_X1 U20736 ( .A1(n17895), .A2(n17566), .ZN(n17582) );
  OAI22_X1 U20737 ( .A1(n10902), .A2(n17568), .B1(n17567), .B2(n17700), .ZN(
        n17595) );
  OAI21_X1 U20738 ( .B1(n17582), .B2(n17595), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17569) );
  OAI211_X1 U20739 ( .C1(n17902), .C2(n17611), .A(n17570), .B(n17569), .ZN(
        P3_U2819) );
  OAI221_X1 U20740 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17585), .C1(
        n17913), .C2(n17586), .A(n17571), .ZN(n17575) );
  NAND4_X1 U20741 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17913), .A3(
        n17597), .A4(n17572), .ZN(n17573) );
  NAND3_X1 U20742 ( .A1(n17575), .A2(n17574), .A3(n17573), .ZN(n17912) );
  AOI211_X1 U20743 ( .C1(n17588), .C2(n17577), .A(n17693), .B(n17576), .ZN(
        n17579) );
  NOR2_X1 U20744 ( .A1(n17909), .A2(n18599), .ZN(n17578) );
  AOI211_X1 U20745 ( .C1(n17580), .C2(n17688), .A(n17579), .B(n17578), .ZN(
        n17584) );
  AOI22_X1 U20746 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17595), .B1(
        n17582), .B2(n17581), .ZN(n17583) );
  OAI211_X1 U20747 ( .C1(n17611), .C2(n17912), .A(n17584), .B(n17583), .ZN(
        P3_U2820) );
  NAND2_X1 U20748 ( .A1(n17586), .A2(n17585), .ZN(n17587) );
  XOR2_X1 U20749 ( .A(n17587), .B(n17913), .Z(n17921) );
  OAI211_X1 U20750 ( .C1(n17589), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n17650), .B(n17588), .ZN(n17591) );
  NAND2_X1 U20751 ( .A1(n17815), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n17590) );
  OAI211_X1 U20752 ( .C1(n17680), .C2(n17592), .A(n17591), .B(n17590), .ZN(
        n17593) );
  AOI221_X1 U20753 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17595), .C1(
        n17913), .C2(n17594), .A(n17593), .ZN(n17596) );
  OAI21_X1 U20754 ( .B1(n17921), .B2(n17611), .A(n17596), .ZN(P3_U2821) );
  NAND2_X1 U20755 ( .A1(n17931), .A2(n17932), .ZN(n17598) );
  XOR2_X1 U20756 ( .A(n17598), .B(n17597), .Z(n17940) );
  AOI21_X1 U20757 ( .B1(n17600), .B2(n17929), .A(n17599), .ZN(n17934) );
  AOI21_X1 U20758 ( .B1(n17671), .B2(n17616), .A(n17601), .ZN(n17615) );
  AOI22_X1 U20759 ( .A1(n17821), .A2(P3_REIP_REG_8__SCAN_IN), .B1(n17602), 
        .B2(n17688), .ZN(n17605) );
  OAI221_X1 U20760 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17603), .C1(
        n17606), .C2(n17617), .A(n18434), .ZN(n17604) );
  OAI211_X1 U20761 ( .C1(n17615), .C2(n17606), .A(n17605), .B(n17604), .ZN(
        n17607) );
  AOI21_X1 U20762 ( .B1(n17685), .B2(n17934), .A(n17607), .ZN(n17610) );
  NAND2_X1 U20763 ( .A1(n17940), .A2(n17608), .ZN(n17609) );
  OAI211_X1 U20764 ( .C1(n17940), .C2(n17611), .A(n17610), .B(n17609), .ZN(
        P3_U2822) );
  NAND2_X1 U20765 ( .A1(n17613), .A2(n17612), .ZN(n17614) );
  XOR2_X1 U20766 ( .A(n17614), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n17948) );
  INV_X1 U20767 ( .A(n17615), .ZN(n17619) );
  NOR2_X1 U20768 ( .A1(n17616), .A2(n18262), .ZN(n17618) );
  INV_X1 U20769 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18593) );
  NOR2_X1 U20770 ( .A1(n18017), .A2(n18593), .ZN(n17941) );
  AOI221_X1 U20771 ( .B1(n17619), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C1(
        n17618), .C2(n17617), .A(n17941), .ZN(n17624) );
  AOI21_X1 U20772 ( .B1(n17943), .B2(n17621), .A(n17620), .ZN(n17944) );
  AOI22_X1 U20773 ( .A1(n9596), .A2(n17944), .B1(n17622), .B2(n17688), .ZN(
        n17623) );
  OAI211_X1 U20774 ( .C1(n17700), .C2(n17948), .A(n17624), .B(n17623), .ZN(
        P3_U2823) );
  AOI21_X1 U20775 ( .B1(n17627), .B2(n17626), .A(n17625), .ZN(n17955) );
  NOR2_X1 U20776 ( .A1(n18017), .A2(n18591), .ZN(n17952) );
  NOR3_X1 U20777 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17628), .A3(
        n18262), .ZN(n17629) );
  AOI211_X1 U20778 ( .C1(n9596), .C2(n17955), .A(n17952), .B(n17629), .ZN(
        n17634) );
  AOI21_X1 U20779 ( .B1(n17953), .B2(n17631), .A(n17630), .ZN(n17956) );
  AOI21_X1 U20780 ( .B1(n18434), .B2(n17632), .A(n17693), .ZN(n17645) );
  AOI22_X1 U20781 ( .A1(n17685), .A2(n17956), .B1(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17645), .ZN(n17633) );
  OAI211_X1 U20782 ( .C1(n17680), .C2(n17635), .A(n17634), .B(n17633), .ZN(
        P3_U2824) );
  AOI21_X1 U20783 ( .B1(n17638), .B2(n17637), .A(n17636), .ZN(n17961) );
  AOI22_X1 U20784 ( .A1(n17821), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n17685), 
        .B2(n17961), .ZN(n17647) );
  OAI21_X1 U20785 ( .B1(n17640), .B2(n9650), .A(n17639), .ZN(n17641) );
  XNOR2_X1 U20786 ( .A(n17641), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17960) );
  NAND2_X1 U20787 ( .A1(n17642), .A2(n9594), .ZN(n17649) );
  INV_X1 U20788 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17643) );
  OAI21_X1 U20789 ( .B1(n17661), .B2(n17649), .A(n17643), .ZN(n17644) );
  AOI22_X1 U20790 ( .A1(n9596), .A2(n17960), .B1(n17645), .B2(n17644), .ZN(
        n17646) );
  OAI211_X1 U20791 ( .C1(n17680), .C2(n17648), .A(n17647), .B(n17646), .ZN(
        P3_U2825) );
  NAND2_X1 U20792 ( .A1(n17650), .A2(n17649), .ZN(n17667) );
  AOI21_X1 U20793 ( .B1(n17965), .B2(n17652), .A(n17651), .ZN(n17973) );
  OAI22_X1 U20794 ( .A1(n17909), .A2(n18587), .B1(n18262), .B2(n17653), .ZN(
        n17654) );
  AOI21_X1 U20795 ( .B1(n17685), .B2(n17973), .A(n17654), .ZN(n17660) );
  AOI21_X1 U20796 ( .B1(n17657), .B2(n17656), .A(n17655), .ZN(n17967) );
  AOI22_X1 U20797 ( .A1(n9596), .A2(n17967), .B1(n17658), .B2(n17688), .ZN(
        n17659) );
  OAI211_X1 U20798 ( .C1(n17661), .C2(n17667), .A(n17660), .B(n17659), .ZN(
        P3_U2826) );
  XNOR2_X1 U20799 ( .A(n17663), .B(n17662), .ZN(n17986) );
  AOI21_X1 U20800 ( .B1(n17666), .B2(n17665), .A(n17664), .ZN(n17983) );
  NOR2_X1 U20801 ( .A1(n18017), .A2(n18584), .ZN(n17981) );
  OAI22_X1 U20802 ( .A1(n17680), .A2(n17668), .B1(n17670), .B2(n17667), .ZN(
        n17669) );
  AOI211_X1 U20803 ( .C1(n9596), .C2(n17983), .A(n17981), .B(n17669), .ZN(
        n17673) );
  NAND4_X1 U20804 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n17671), .A3(
        n9594), .A4(n17670), .ZN(n17672) );
  OAI211_X1 U20805 ( .C1(n17700), .C2(n17986), .A(n17673), .B(n17672), .ZN(
        P3_U2827) );
  AOI21_X1 U20806 ( .B1(n17676), .B2(n17675), .A(n17674), .ZN(n17992) );
  INV_X1 U20807 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18582) );
  NOR2_X1 U20808 ( .A1(n18017), .A2(n18582), .ZN(n18001) );
  XNOR2_X1 U20809 ( .A(n17678), .B(n17677), .ZN(n18000) );
  OAI22_X1 U20810 ( .A1(n17680), .A2(n17679), .B1(n17700), .B2(n18000), .ZN(
        n17681) );
  AOI211_X1 U20811 ( .C1(n9596), .C2(n17992), .A(n18001), .B(n17681), .ZN(
        n17682) );
  OAI221_X1 U20812 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18262), .C1(
        n17683), .C2(n9594), .A(n17682), .ZN(P3_U2828) );
  NOR2_X1 U20813 ( .A1(n17695), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17684) );
  XNOR2_X1 U20814 ( .A(n17684), .B(n17687), .ZN(n18004) );
  AOI22_X1 U20815 ( .A1(n17821), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n17685), 
        .B2(n18004), .ZN(n17691) );
  AOI21_X1 U20816 ( .B1(n17687), .B2(n17694), .A(n17686), .ZN(n18010) );
  AOI22_X1 U20817 ( .A1(n9596), .A2(n18010), .B1(n17692), .B2(n17688), .ZN(
        n17690) );
  OAI211_X1 U20818 ( .C1(n17693), .C2(n17692), .A(n17691), .B(n17690), .ZN(
        P3_U2829) );
  OAI21_X1 U20819 ( .B1(n17695), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17694), .ZN(n18019) );
  INV_X1 U20820 ( .A(n18019), .ZN(n18021) );
  OAI21_X1 U20821 ( .B1(n18555), .B2(n18708), .A(n9594), .ZN(n17697) );
  AOI22_X1 U20822 ( .A1(n17821), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17697), .ZN(n17698) );
  OAI221_X1 U20823 ( .B1(n18021), .B2(n17700), .C1(n18019), .C2(n17699), .A(
        n17698), .ZN(P3_U2830) );
  AOI22_X1 U20824 ( .A1(n17821), .A2(P3_REIP_REG_27__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17982), .ZN(n17710) );
  INV_X1 U20825 ( .A(n17701), .ZN(n17750) );
  NOR2_X1 U20826 ( .A1(n18514), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17996) );
  NOR2_X1 U20827 ( .A1(n17996), .A2(n17760), .ZN(n17805) );
  AOI22_X1 U20828 ( .A1(n18486), .A2(n17703), .B1(n17890), .B2(n17702), .ZN(
        n17704) );
  OAI221_X1 U20829 ( .B1(n17994), .B2(n17708), .C1(n17994), .C2(n17805), .A(
        n17704), .ZN(n17705) );
  OAI21_X1 U20830 ( .B1(n17706), .B2(n17705), .A(n18006), .ZN(n17713) );
  OAI21_X1 U20831 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18023), .A(
        n17713), .ZN(n17707) );
  OAI221_X1 U20832 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17708), 
        .C1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n17750), .A(n17707), .ZN(
        n17709) );
  OAI211_X1 U20833 ( .C1(n17711), .C2(n17939), .A(n17710), .B(n17709), .ZN(
        P3_U2835) );
  NAND2_X1 U20834 ( .A1(n17815), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17712) );
  OAI221_X1 U20835 ( .B1(n17714), .B2(n18007), .C1(n17714), .C2(n17713), .A(
        n17712), .ZN(n17715) );
  AOI21_X1 U20836 ( .B1(n17769), .B2(n17716), .A(n17715), .ZN(n17717) );
  OAI21_X1 U20837 ( .B1(n17718), .B2(n17939), .A(n17717), .ZN(P3_U2836) );
  AOI21_X1 U20838 ( .B1(n17751), .B2(n17805), .A(n17994), .ZN(n17739) );
  OAI21_X1 U20839 ( .B1(n17719), .B2(n17773), .A(n18497), .ZN(n17763) );
  OAI21_X1 U20840 ( .B1(n17720), .B2(n18519), .A(n17763), .ZN(n17741) );
  AOI211_X1 U20841 ( .C1(n17926), .C2(n17721), .A(n17739), .B(n17741), .ZN(
        n17725) );
  NAND3_X1 U20842 ( .A1(n17723), .A2(n17722), .A3(n17727), .ZN(n17724) );
  OAI21_X1 U20843 ( .B1(n17725), .B2(n17727), .A(n17724), .ZN(n17732) );
  OAI21_X1 U20844 ( .B1(n17727), .B2(n18007), .A(n17726), .ZN(n17731) );
  OAI22_X1 U20845 ( .A1(n17939), .A2(n17729), .B1(n17933), .B2(n17728), .ZN(
        n17730) );
  AOI211_X1 U20846 ( .C1(n18006), .C2(n17732), .A(n17731), .B(n17730), .ZN(
        n17733) );
  OAI21_X1 U20847 ( .B1(n18015), .B2(n17734), .A(n17733), .ZN(P3_U2837) );
  INV_X1 U20848 ( .A(n17735), .ZN(n17737) );
  OAI22_X1 U20849 ( .A1(n17737), .A2(n17835), .B1(n17736), .B2(n17999), .ZN(
        n17738) );
  NOR3_X1 U20850 ( .A1(n17982), .A2(n17739), .A3(n17738), .ZN(n17743) );
  NAND2_X1 U20851 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17743), .ZN(
        n17740) );
  OAI21_X1 U20852 ( .B1(n17741), .B2(n17740), .A(n18017), .ZN(n17757) );
  AOI211_X1 U20853 ( .C1(n17744), .C2(n17743), .A(n17742), .B(n17757), .ZN(
        n17745) );
  AOI21_X1 U20854 ( .B1(n17746), .B2(n17769), .A(n17745), .ZN(n17748) );
  NAND2_X1 U20855 ( .A1(n17815), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n17747) );
  OAI211_X1 U20856 ( .C1(n17749), .C2(n17939), .A(n17748), .B(n17747), .ZN(
        P3_U2838) );
  NAND3_X1 U20857 ( .A1(n17751), .A2(n18007), .A3(n17750), .ZN(n17755) );
  AOI21_X1 U20858 ( .B1(n17753), .B2(n17878), .A(n17752), .ZN(n17754) );
  OAI221_X1 U20859 ( .B1(n17757), .B2(n17756), .C1(n17757), .C2(n17755), .A(
        n17754), .ZN(P3_U2839) );
  OAI22_X1 U20860 ( .A1(n17758), .A2(n17999), .B1(n17836), .B2(n17835), .ZN(
        n17759) );
  NOR2_X1 U20861 ( .A1(n18023), .A2(n17759), .ZN(n17826) );
  OAI21_X1 U20862 ( .B1(n17773), .B2(n17827), .A(n18524), .ZN(n17762) );
  OAI21_X1 U20863 ( .B1(n17760), .B2(n17785), .A(n18506), .ZN(n17761) );
  NAND4_X1 U20864 ( .A1(n17826), .A2(n17763), .A3(n17762), .A4(n17761), .ZN(
        n17786) );
  NAND2_X1 U20865 ( .A1(n17999), .A2(n17835), .ZN(n17810) );
  INV_X1 U20866 ( .A(n17810), .ZN(n17894) );
  OAI22_X1 U20867 ( .A1(n18526), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n17764), .B2(n17894), .ZN(n17765) );
  NOR2_X1 U20868 ( .A1(n17786), .A2(n17765), .ZN(n17777) );
  INV_X1 U20869 ( .A(n17777), .ZN(n17767) );
  OAI221_X1 U20870 ( .B1(n17767), .B2(n17926), .C1(n17767), .C2(n17766), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17772) );
  INV_X1 U20871 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18623) );
  AOI22_X1 U20872 ( .A1(n17878), .A2(n17770), .B1(n17769), .B2(n17768), .ZN(
        n17771) );
  OAI221_X1 U20873 ( .B1(n17821), .B2(n17772), .C1(n18017), .C2(n18623), .A(
        n17771), .ZN(P3_U2840) );
  NOR2_X1 U20874 ( .A1(n17773), .A2(n17794), .ZN(n17795) );
  INV_X1 U20875 ( .A(n17774), .ZN(n17780) );
  NAND2_X1 U20876 ( .A1(n18519), .A2(n18514), .ZN(n18005) );
  INV_X1 U20877 ( .A(n18005), .ZN(n17776) );
  AOI221_X1 U20878 ( .B1(n17778), .B2(n17777), .C1(n17776), .C2(n17777), .A(
        n17775), .ZN(n17779) );
  AOI22_X1 U20879 ( .A1(n17795), .A2(n17780), .B1(n17779), .B2(n17909), .ZN(
        n17782) );
  OAI211_X1 U20880 ( .C1(n17783), .C2(n17939), .A(n17782), .B(n17781), .ZN(
        P3_U2841) );
  INV_X1 U20881 ( .A(n17784), .ZN(n17793) );
  OAI221_X1 U20882 ( .B1(n17786), .B2(n17785), .C1(n17786), .C2(n17810), .A(
        n18017), .ZN(n17799) );
  NAND3_X1 U20883 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n17800), .A3(n18005), 
        .ZN(n17788) );
  AOI21_X1 U20884 ( .B1(n17799), .B2(n17788), .A(n17787), .ZN(n17789) );
  AOI211_X1 U20885 ( .C1(n17791), .C2(n17878), .A(n17790), .B(n17789), .ZN(
        n17792) );
  OAI21_X1 U20886 ( .B1(n17794), .B2(n17793), .A(n17792), .ZN(P3_U2842) );
  AOI22_X1 U20887 ( .A1(n17878), .A2(n17796), .B1(n17795), .B2(n17800), .ZN(
        n17798) );
  NAND2_X1 U20888 ( .A1(n17815), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17797) );
  OAI211_X1 U20889 ( .C1(n17800), .C2(n17799), .A(n17798), .B(n17797), .ZN(
        P3_U2843) );
  NAND2_X1 U20890 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17971) );
  OAI22_X1 U20891 ( .A1(n17968), .A2(n18519), .B1(n17971), .B2(n17988), .ZN(
        n17966) );
  NAND2_X1 U20892 ( .A1(n17801), .A2(n17966), .ZN(n17949) );
  NOR2_X1 U20893 ( .A1(n17802), .A2(n17949), .ZN(n17837) );
  NOR2_X1 U20894 ( .A1(n17837), .A2(n17803), .ZN(n17882) );
  NAND2_X1 U20895 ( .A1(n17804), .A2(n17914), .ZN(n17834) );
  AOI21_X1 U20896 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17805), .A(
        n17994), .ZN(n17809) );
  OAI221_X1 U20897 ( .B1(n18519), .B2(n17807), .C1(n18519), .C2(n17806), .A(
        n17826), .ZN(n17808) );
  AOI211_X1 U20898 ( .C1(n17811), .C2(n17810), .A(n17809), .B(n17808), .ZN(
        n17820) );
  AOI221_X1 U20899 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17820), 
        .C1(n17994), .C2(n17820), .A(n17812), .ZN(n17813) );
  AOI22_X1 U20900 ( .A1(n17814), .A2(n17878), .B1(n17813), .B2(n17909), .ZN(
        n17817) );
  NAND2_X1 U20901 ( .A1(n17815), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17816) );
  OAI211_X1 U20902 ( .C1(n17818), .C2(n17834), .A(n17817), .B(n17816), .ZN(
        P3_U2844) );
  NOR3_X1 U20903 ( .A1(n17821), .A2(n17820), .A3(n17819), .ZN(n17823) );
  NOR3_X1 U20904 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n10903), .A3(
        n17834), .ZN(n17822) );
  AOI211_X1 U20905 ( .C1(n17878), .C2(n17824), .A(n17823), .B(n17822), .ZN(
        n17825) );
  OAI21_X1 U20906 ( .B1(n17909), .B2(n18614), .A(n17825), .ZN(P3_U2845) );
  INV_X1 U20907 ( .A(n17826), .ZN(n17830) );
  AOI22_X1 U20908 ( .A1(n18497), .A2(n17852), .B1(n18506), .B2(n17904), .ZN(
        n17916) );
  OAI21_X1 U20909 ( .B1(n17850), .B2(n18524), .A(n17827), .ZN(n17828) );
  OAI211_X1 U20910 ( .C1(n17907), .C2(n17829), .A(n17916), .B(n17828), .ZN(
        n17838) );
  OAI221_X1 U20911 ( .B1(n17830), .B2(n17926), .C1(n17830), .C2(n17838), .A(
        n17909), .ZN(n17833) );
  AOI22_X1 U20912 ( .A1(n17815), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n17878), 
        .B2(n17831), .ZN(n17832) );
  OAI221_X1 U20913 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17834), 
        .C1(n10903), .C2(n17833), .A(n17832), .ZN(P3_U2846) );
  NOR2_X1 U20914 ( .A1(n17836), .A2(n17835), .ZN(n17841) );
  NAND2_X1 U20915 ( .A1(n17851), .A2(n17837), .ZN(n17859) );
  OAI21_X1 U20916 ( .B1(n17860), .B2(n17859), .A(n17850), .ZN(n17839) );
  AOI22_X1 U20917 ( .A1(n17841), .A2(n17840), .B1(n17839), .B2(n17838), .ZN(
        n17842) );
  OAI21_X1 U20918 ( .B1(n17844), .B2(n17843), .A(n17842), .ZN(n17845) );
  AOI22_X1 U20919 ( .A1(n17815), .A2(P3_REIP_REG_15__SCAN_IN), .B1(n18006), 
        .B2(n17845), .ZN(n17849) );
  NAND3_X1 U20920 ( .A1(n18020), .A2(n17847), .A3(n17846), .ZN(n17848) );
  OAI211_X1 U20921 ( .C1(n17850), .C2(n18007), .A(n17849), .B(n17848), .ZN(
        P3_U2847) );
  AOI21_X1 U20922 ( .B1(n17851), .B2(n17868), .A(n18526), .ZN(n17856) );
  INV_X1 U20923 ( .A(n17917), .ZN(n17892) );
  AND2_X1 U20924 ( .A1(n18497), .A2(n17852), .ZN(n17897) );
  AOI221_X1 U20925 ( .B1(n17853), .B2(n18524), .C1(n17892), .C2(n18524), .A(
        n17897), .ZN(n17873) );
  OAI211_X1 U20926 ( .C1(n17854), .C2(n18519), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17873), .ZN(n17855) );
  AOI211_X1 U20927 ( .C1(n17857), .C2(n18005), .A(n17856), .B(n17855), .ZN(
        n17858) );
  AOI211_X1 U20928 ( .C1(n17860), .C2(n17859), .A(n17858), .B(n18023), .ZN(
        n17865) );
  OAI22_X1 U20929 ( .A1(n18017), .A2(n18608), .B1(n18007), .B2(n17860), .ZN(
        n17864) );
  OAI22_X1 U20930 ( .A1(n17862), .A2(n17939), .B1(n17933), .B2(n17861), .ZN(
        n17863) );
  NOR3_X1 U20931 ( .A1(n17865), .A2(n17864), .A3(n17863), .ZN(n17866) );
  OAI21_X1 U20932 ( .B1(n18015), .B2(n17867), .A(n17866), .ZN(P3_U2848) );
  AOI21_X1 U20933 ( .B1(n17895), .B2(n17868), .A(n18526), .ZN(n17869) );
  AOI21_X1 U20934 ( .B1(n18497), .B2(n17881), .A(n17869), .ZN(n17898) );
  AOI22_X1 U20935 ( .A1(n18486), .A2(n17871), .B1(n17890), .B2(n17870), .ZN(
        n17872) );
  NAND3_X1 U20936 ( .A1(n17898), .A2(n17873), .A3(n17872), .ZN(n17885) );
  OAI21_X1 U20937 ( .B1(n18526), .B2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17884) );
  INV_X1 U20938 ( .A(n17884), .ZN(n17874) );
  OAI21_X1 U20939 ( .B1(n17907), .B2(n17874), .A(n18006), .ZN(n17875) );
  OAI21_X1 U20940 ( .B1(n17885), .B2(n17875), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17880) );
  AOI22_X1 U20941 ( .A1(n17878), .A2(n17877), .B1(n17914), .B2(n17876), .ZN(
        n17879) );
  OAI221_X1 U20942 ( .B1(n17815), .B2(n17880), .C1(n18017), .C2(n18605), .A(
        n17879), .ZN(P3_U2849) );
  AOI22_X1 U20943 ( .A1(n17821), .A2(P3_REIP_REG_12__SCAN_IN), .B1(n17982), 
        .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17887) );
  OAI21_X1 U20944 ( .B1(n17882), .B2(n17881), .A(n9757), .ZN(n17883) );
  OAI211_X1 U20945 ( .C1(n17885), .C2(n17884), .A(n18006), .B(n17883), .ZN(
        n17886) );
  OAI211_X1 U20946 ( .C1(n17888), .C2(n17939), .A(n17887), .B(n17886), .ZN(
        P3_U2850) );
  AOI22_X1 U20947 ( .A1(n17815), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n17914), 
        .B2(n17889), .ZN(n17901) );
  AOI22_X1 U20948 ( .A1(n18486), .A2(n17891), .B1(n17890), .B2(n17932), .ZN(
        n17915) );
  OAI21_X1 U20949 ( .B1(n17913), .B2(n17892), .A(n18524), .ZN(n17893) );
  OAI211_X1 U20950 ( .C1(n17895), .C2(n17894), .A(n17915), .B(n17893), .ZN(
        n17896) );
  NOR3_X1 U20951 ( .A1(n17897), .A2(n18023), .A3(n17896), .ZN(n17906) );
  OAI211_X1 U20952 ( .C1(n18514), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17898), .B(n17906), .ZN(n17899) );
  NAND3_X1 U20953 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17909), .A3(
        n17899), .ZN(n17900) );
  OAI211_X1 U20954 ( .C1(n17902), .C2(n17939), .A(n17901), .B(n17900), .ZN(
        P3_U2851) );
  NOR2_X1 U20955 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17913), .ZN(
        n17903) );
  AOI22_X1 U20956 ( .A1(n17821), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n17914), 
        .B2(n17903), .ZN(n17911) );
  NAND2_X1 U20957 ( .A1(n18506), .A2(n17904), .ZN(n17905) );
  OAI211_X1 U20958 ( .C1(n17907), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17906), .B(n17905), .ZN(n17908) );
  NAND3_X1 U20959 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17909), .A3(
        n17908), .ZN(n17910) );
  OAI211_X1 U20960 ( .C1(n17912), .C2(n17939), .A(n17911), .B(n17910), .ZN(
        P3_U2852) );
  AOI22_X1 U20961 ( .A1(n17821), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n17914), 
        .B2(n17913), .ZN(n17920) );
  OAI211_X1 U20962 ( .C1(n18514), .C2(n17917), .A(n17916), .B(n17915), .ZN(
        n17918) );
  OAI211_X1 U20963 ( .C1(n18023), .C2(n17918), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n17909), .ZN(n17919) );
  OAI211_X1 U20964 ( .C1(n17921), .C2(n17939), .A(n17920), .B(n17919), .ZN(
        P3_U2853) );
  NOR3_X1 U20965 ( .A1(n18023), .A2(n17925), .A3(n17949), .ZN(n17930) );
  AOI21_X1 U20966 ( .B1(n17922), .B2(n17970), .A(n17996), .ZN(n17923) );
  OAI21_X1 U20967 ( .B1(n17924), .B2(n18519), .A(n17923), .ZN(n17950) );
  AOI21_X1 U20968 ( .B1(n17926), .B2(n17925), .A(n17950), .ZN(n17942) );
  OAI21_X1 U20969 ( .B1(n17942), .B2(n17972), .A(n18007), .ZN(n17928) );
  NOR2_X1 U20970 ( .A1(n18017), .A2(n18595), .ZN(n17927) );
  AOI221_X1 U20971 ( .B1(n17930), .B2(n17929), .C1(n17928), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n17927), .ZN(n17938) );
  AND2_X1 U20972 ( .A1(n17932), .A2(n17931), .ZN(n17936) );
  INV_X1 U20973 ( .A(n17933), .ZN(n17935) );
  AOI22_X1 U20974 ( .A1(n17936), .A2(n17935), .B1(n18020), .B2(n17934), .ZN(
        n17937) );
  OAI211_X1 U20975 ( .C1(n17940), .C2(n17939), .A(n17938), .B(n17937), .ZN(
        P3_U2854) );
  AOI21_X1 U20976 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17982), .A(
        n17941), .ZN(n17947) );
  AOI221_X1 U20977 ( .B1(n17953), .B2(n17943), .C1(n17949), .C2(n17943), .A(
        n17942), .ZN(n17945) );
  AOI22_X1 U20978 ( .A1(n18006), .A2(n17945), .B1(n18022), .B2(n17944), .ZN(
        n17946) );
  OAI211_X1 U20979 ( .C1(n18015), .C2(n17948), .A(n17947), .B(n17946), .ZN(
        P3_U2855) );
  NOR2_X1 U20980 ( .A1(n18023), .A2(n17949), .ZN(n17954) );
  AOI21_X1 U20981 ( .B1(n17950), .B2(n18006), .A(n17982), .ZN(n17951) );
  INV_X1 U20982 ( .A(n17951), .ZN(n17959) );
  AOI221_X1 U20983 ( .B1(n17954), .B2(n17953), .C1(n17959), .C2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(n17952), .ZN(n17958) );
  AOI22_X1 U20984 ( .A1(n18020), .A2(n17956), .B1(n18022), .B2(n17955), .ZN(
        n17957) );
  NAND2_X1 U20985 ( .A1(n17958), .A2(n17957), .ZN(P3_U2856) );
  INV_X1 U20986 ( .A(n17966), .ZN(n17979) );
  OR4_X1 U20987 ( .A1(n10739), .A2(n18023), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A4(n17979), .ZN(n17964) );
  AOI22_X1 U20988 ( .A1(n17821), .A2(P3_REIP_REG_5__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17959), .ZN(n17963) );
  AOI22_X1 U20989 ( .A1(n18020), .A2(n17961), .B1(n18022), .B2(n17960), .ZN(
        n17962) );
  OAI211_X1 U20990 ( .C1(n17965), .C2(n17964), .A(n17963), .B(n17962), .ZN(
        P3_U2857) );
  NAND3_X1 U20991 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18006), .A3(
        n17966), .ZN(n17977) );
  AOI22_X1 U20992 ( .A1(n17821), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18022), 
        .B2(n17967), .ZN(n17976) );
  NAND2_X1 U20993 ( .A1(n18497), .A2(n17968), .ZN(n17987) );
  NAND2_X1 U20994 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17987), .ZN(
        n17969) );
  AOI211_X1 U20995 ( .C1(n17971), .C2(n17970), .A(n17996), .B(n17969), .ZN(
        n17978) );
  OAI21_X1 U20996 ( .B1(n17978), .B2(n17972), .A(n18007), .ZN(n17974) );
  AOI22_X1 U20997 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n17974), .B1(
        n18020), .B2(n17973), .ZN(n17975) );
  OAI211_X1 U20998 ( .C1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n17977), .A(
        n17976), .B(n17975), .ZN(P3_U2858) );
  AOI211_X1 U20999 ( .C1(n17979), .C2(n10739), .A(n17978), .B(n18023), .ZN(
        n17980) );
  AOI211_X1 U21000 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n17982), .A(
        n17981), .B(n17980), .ZN(n17985) );
  NAND2_X1 U21001 ( .A1(n18022), .A2(n17983), .ZN(n17984) );
  OAI211_X1 U21002 ( .C1(n17986), .C2(n18015), .A(n17985), .B(n17984), .ZN(
        P3_U2859) );
  INV_X1 U21003 ( .A(n17987), .ZN(n17990) );
  NOR3_X1 U21004 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18663), .A3(
        n17988), .ZN(n17989) );
  AOI211_X1 U21005 ( .C1(n17992), .C2(n17991), .A(n17990), .B(n17989), .ZN(
        n17998) );
  NAND2_X1 U21006 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17993) );
  OAI22_X1 U21007 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17994), .B1(
        n18519), .B2(n17993), .ZN(n17995) );
  OAI21_X1 U21008 ( .B1(n17996), .B2(n17995), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n17997) );
  OAI211_X1 U21009 ( .C1(n18000), .C2(n17999), .A(n17998), .B(n17997), .ZN(
        n18002) );
  AOI21_X1 U21010 ( .B1(n18006), .B2(n18002), .A(n18001), .ZN(n18003) );
  OAI21_X1 U21011 ( .B1(n18007), .B2(n10723), .A(n18003), .ZN(P3_U2860) );
  INV_X1 U21012 ( .A(n18004), .ZN(n18016) );
  NOR2_X1 U21013 ( .A1(n18017), .A2(n18685), .ZN(n18009) );
  NAND3_X1 U21014 ( .A1(n18006), .A2(n18680), .A3(n18005), .ZN(n18025) );
  AOI21_X1 U21015 ( .B1(n18007), .B2(n18025), .A(n18663), .ZN(n18008) );
  AOI211_X1 U21016 ( .C1(n18010), .C2(n18022), .A(n18009), .B(n18008), .ZN(
        n18014) );
  NAND3_X1 U21017 ( .A1(n18012), .A2(n18663), .A3(n18011), .ZN(n18013) );
  OAI211_X1 U21018 ( .C1(n18016), .C2(n18015), .A(n18014), .B(n18013), .ZN(
        P3_U2861) );
  INV_X1 U21019 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18691) );
  NOR2_X1 U21020 ( .A1(n18017), .A2(n18691), .ZN(n18018) );
  AOI221_X1 U21021 ( .B1(n18022), .B2(n18021), .C1(n18020), .C2(n18019), .A(
        n18018), .ZN(n18026) );
  OAI211_X1 U21022 ( .C1(n18506), .C2(n18023), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n17909), .ZN(n18024) );
  NAND3_X1 U21023 ( .A1(n18026), .A2(n18025), .A3(n18024), .ZN(P3_U2862) );
  OAI211_X1 U21024 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n18027), .A(
        P3_STATE2_REG_1__SCAN_IN), .B(P3_STATE2_REG_2__SCAN_IN), .ZN(n18546)
         );
  AOI21_X1 U21025 ( .B1(n18546), .B2(n18082), .A(n18028), .ZN(n18029) );
  INV_X1 U21026 ( .A(n18029), .ZN(n18030) );
  OAI221_X1 U21027 ( .B1(n18035), .B2(n18699), .C1(n18035), .C2(n18034), .A(
        n18030), .ZN(P3_U2863) );
  INV_X1 U21028 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18538) );
  NAND2_X1 U21029 ( .A1(n18535), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18331) );
  INV_X1 U21030 ( .A(n18331), .ZN(n18352) );
  NAND2_X1 U21031 ( .A1(n18538), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18213) );
  INV_X1 U21032 ( .A(n18213), .ZN(n18215) );
  NOR2_X1 U21033 ( .A1(n18352), .A2(n18215), .ZN(n18032) );
  OAI22_X1 U21034 ( .A1(n18033), .A2(n18538), .B1(n18032), .B2(n18031), .ZN(
        P3_U2866) );
  NOR2_X1 U21035 ( .A1(n18539), .A2(n18034), .ZN(P3_U2867) );
  NAND2_X1 U21036 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18529) );
  NOR2_X1 U21037 ( .A1(n18535), .A2(n18538), .ZN(n18036) );
  INV_X1 U21038 ( .A(n18036), .ZN(n18042) );
  NOR2_X2 U21039 ( .A1(n18529), .A2(n18042), .ZN(n18428) );
  NAND2_X1 U21040 ( .A1(n18530), .A2(n18035), .ZN(n18531) );
  NOR2_X1 U21041 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18125) );
  INV_X1 U21042 ( .A(n18125), .ZN(n18167) );
  NOR2_X1 U21043 ( .A1(n18531), .A2(n18167), .ZN(n18138) );
  CLKBUF_X1 U21044 ( .A(n18138), .Z(n18142) );
  NOR2_X1 U21045 ( .A1(n18428), .A2(n18142), .ZN(n18104) );
  AOI21_X1 U21046 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18084), .ZN(n18404) );
  INV_X1 U21047 ( .A(n18404), .ZN(n18295) );
  NAND2_X1 U21048 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18035), .ZN(
        n18294) );
  NAND2_X1 U21049 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18530), .ZN(
        n18264) );
  NAND2_X1 U21050 ( .A1(n18294), .A2(n18264), .ZN(n18351) );
  NAND2_X1 U21051 ( .A1(n18036), .A2(n18351), .ZN(n18401) );
  OAI22_X1 U21052 ( .A1(n18104), .A2(n18295), .B1(n18262), .B2(n18401), .ZN(
        n18080) );
  NOR2_X1 U21053 ( .A1(n18042), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18433) );
  NAND2_X1 U21054 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18433), .ZN(
        n18398) );
  INV_X1 U21055 ( .A(n18398), .ZN(n18480) );
  AND2_X1 U21056 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18434), .ZN(n18435) );
  NOR2_X2 U21057 ( .A1(n18084), .A2(n18037), .ZN(n18429) );
  NOR2_X1 U21058 ( .A1(n18400), .A2(n18104), .ZN(n18075) );
  AOI22_X1 U21059 ( .A1(n18480), .A2(n18435), .B1(n18429), .B2(n18075), .ZN(
        n18044) );
  NAND2_X1 U21060 ( .A1(n18039), .A2(n18038), .ZN(n18076) );
  NOR2_X1 U21061 ( .A1(n18040), .A2(n18076), .ZN(n18300) );
  INV_X1 U21062 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18041) );
  NOR2_X2 U21063 ( .A1(n18262), .A2(n18041), .ZN(n18430) );
  NOR2_X2 U21064 ( .A1(n18042), .A2(n18294), .ZN(n18399) );
  AOI22_X1 U21065 ( .A1(n18142), .A2(n18300), .B1(n18430), .B2(n18399), .ZN(
        n18043) );
  OAI211_X1 U21066 ( .C1(n18045), .C2(n18080), .A(n18044), .B(n18043), .ZN(
        P3_U2868) );
  AND2_X1 U21067 ( .A1(n18434), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18441) );
  AND2_X1 U21068 ( .A1(n18354), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18439) );
  AOI22_X1 U21069 ( .A1(n18399), .A2(n18441), .B1(n18075), .B2(n18439), .ZN(
        n18048) );
  NOR2_X1 U21070 ( .A1(n18046), .A2(n18076), .ZN(n18268) );
  NOR2_X2 U21071 ( .A1(n14875), .A2(n18262), .ZN(n18440) );
  AOI22_X1 U21072 ( .A1(n18138), .A2(n18268), .B1(n18480), .B2(n18440), .ZN(
        n18047) );
  OAI211_X1 U21073 ( .C1(n18049), .C2(n18080), .A(n18048), .B(n18047), .ZN(
        P3_U2869) );
  AND2_X1 U21074 ( .A1(n18434), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18447) );
  NOR2_X2 U21075 ( .A1(n18084), .A2(n18050), .ZN(n18445) );
  AOI22_X1 U21076 ( .A1(n18399), .A2(n18447), .B1(n18075), .B2(n18445), .ZN(
        n18053) );
  NOR2_X1 U21077 ( .A1(n9671), .A2(n18076), .ZN(n18306) );
  INV_X1 U21078 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n18051) );
  NOR2_X2 U21079 ( .A1(n18051), .A2(n18262), .ZN(n18446) );
  AOI22_X1 U21080 ( .A1(n18142), .A2(n18306), .B1(n18480), .B2(n18446), .ZN(
        n18052) );
  OAI211_X1 U21081 ( .C1(n20898), .C2(n18080), .A(n18053), .B(n18052), .ZN(
        P3_U2870) );
  AND2_X1 U21082 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18434), .ZN(n18453) );
  AND2_X1 U21083 ( .A1(n18354), .A2(BUF2_REG_3__SCAN_IN), .ZN(n18451) );
  AOI22_X1 U21084 ( .A1(n18480), .A2(n18453), .B1(n18075), .B2(n18451), .ZN(
        n18056) );
  NOR2_X1 U21085 ( .A1(n18054), .A2(n18076), .ZN(n18310) );
  NOR2_X2 U21086 ( .A1(n18262), .A2(n14909), .ZN(n18452) );
  AOI22_X1 U21087 ( .A1(n18142), .A2(n18310), .B1(n18399), .B2(n18452), .ZN(
        n18055) );
  OAI211_X1 U21088 ( .C1(n18057), .C2(n18080), .A(n18056), .B(n18055), .ZN(
        P3_U2871) );
  NOR2_X2 U21089 ( .A1(n14851), .A2(n18262), .ZN(n18458) );
  NOR2_X2 U21090 ( .A1(n18084), .A2(n18058), .ZN(n18457) );
  AOI22_X1 U21091 ( .A1(n18480), .A2(n18458), .B1(n18075), .B2(n18457), .ZN(
        n18062) );
  NOR2_X1 U21092 ( .A1(n18059), .A2(n18076), .ZN(n18277) );
  INV_X1 U21093 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n18060) );
  NOR2_X2 U21094 ( .A1(n18262), .A2(n18060), .ZN(n18459) );
  AOI22_X1 U21095 ( .A1(n18142), .A2(n18277), .B1(n18399), .B2(n18459), .ZN(
        n18061) );
  OAI211_X1 U21096 ( .C1(n18063), .C2(n18080), .A(n18062), .B(n18061), .ZN(
        P3_U2872) );
  INV_X1 U21097 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18064) );
  NOR2_X2 U21098 ( .A1(n18064), .A2(n18262), .ZN(n18465) );
  NOR2_X2 U21099 ( .A1(n18084), .A2(n18065), .ZN(n18463) );
  AOI22_X1 U21100 ( .A1(n18480), .A2(n18465), .B1(n18075), .B2(n18463), .ZN(
        n18068) );
  NOR2_X1 U21101 ( .A1(n18066), .A2(n18076), .ZN(n18316) );
  AND2_X1 U21102 ( .A1(n18434), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18464) );
  AOI22_X1 U21103 ( .A1(n18142), .A2(n18316), .B1(n18399), .B2(n18464), .ZN(
        n18067) );
  OAI211_X1 U21104 ( .C1(n18069), .C2(n18080), .A(n18068), .B(n18067), .ZN(
        P3_U2873) );
  NOR2_X2 U21105 ( .A1(n18070), .A2(n18262), .ZN(n18469) );
  NOR2_X2 U21106 ( .A1(n18084), .A2(n20858), .ZN(n18470) );
  AOI22_X1 U21107 ( .A1(n18480), .A2(n18469), .B1(n18075), .B2(n18470), .ZN(
        n18073) );
  NOR2_X1 U21108 ( .A1(n18071), .A2(n18076), .ZN(n18320) );
  NOR2_X2 U21109 ( .A1(n18262), .A2(n14894), .ZN(n18471) );
  AOI22_X1 U21110 ( .A1(n18142), .A2(n18320), .B1(n18399), .B2(n18471), .ZN(
        n18072) );
  OAI211_X1 U21111 ( .C1(n18074), .C2(n18080), .A(n18073), .B(n18072), .ZN(
        P3_U2874) );
  NOR2_X2 U21112 ( .A1(n18262), .A2(n19083), .ZN(n18478) );
  NOR2_X2 U21113 ( .A1(n20860), .A2(n18084), .ZN(n18476) );
  AOI22_X1 U21114 ( .A1(n18480), .A2(n18478), .B1(n18075), .B2(n18476), .ZN(
        n18079) );
  NOR2_X1 U21115 ( .A1(n18077), .A2(n18076), .ZN(n18289) );
  NOR2_X2 U21116 ( .A1(n14172), .A2(n18262), .ZN(n18479) );
  AOI22_X1 U21117 ( .A1(n18142), .A2(n18289), .B1(n18399), .B2(n18479), .ZN(
        n18078) );
  OAI211_X1 U21118 ( .C1(n18081), .C2(n18080), .A(n18079), .B(n18078), .ZN(
        P3_U2875) );
  INV_X1 U21119 ( .A(n18300), .ZN(n18438) );
  NOR2_X2 U21120 ( .A1(n18167), .A2(n18264), .ZN(n18163) );
  INV_X1 U21121 ( .A(n18163), .ZN(n18103) );
  NAND2_X1 U21122 ( .A1(n18530), .A2(n18554), .ZN(n18263) );
  NOR2_X1 U21123 ( .A1(n18167), .A2(n18263), .ZN(n18099) );
  AOI22_X1 U21124 ( .A1(n18428), .A2(n18430), .B1(n18429), .B2(n18099), .ZN(
        n18086) );
  NOR2_X1 U21125 ( .A1(n18538), .A2(n18258), .ZN(n18431) );
  INV_X1 U21126 ( .A(n18082), .ZN(n18083) );
  NOR2_X1 U21127 ( .A1(n18084), .A2(n18083), .ZN(n18432) );
  INV_X1 U21128 ( .A(n18432), .ZN(n18260) );
  NOR2_X1 U21129 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18260), .ZN(
        n18168) );
  AOI22_X1 U21130 ( .A1(n18434), .A2(n18431), .B1(n18125), .B2(n18168), .ZN(
        n18100) );
  AOI22_X1 U21131 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18100), .B1(
        n18399), .B2(n18435), .ZN(n18085) );
  OAI211_X1 U21132 ( .C1(n18438), .C2(n18103), .A(n18086), .B(n18085), .ZN(
        P3_U2876) );
  INV_X1 U21133 ( .A(n18268), .ZN(n18444) );
  AOI22_X1 U21134 ( .A1(n18399), .A2(n18440), .B1(n18439), .B2(n18099), .ZN(
        n18088) );
  AOI22_X1 U21135 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18100), .B1(
        n18428), .B2(n18441), .ZN(n18087) );
  OAI211_X1 U21136 ( .C1(n18444), .C2(n18103), .A(n18088), .B(n18087), .ZN(
        P3_U2877) );
  INV_X1 U21137 ( .A(n18306), .ZN(n18450) );
  AOI22_X1 U21138 ( .A1(n18399), .A2(n18446), .B1(n18445), .B2(n18099), .ZN(
        n18090) );
  AOI22_X1 U21139 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18100), .B1(
        n18428), .B2(n18447), .ZN(n18089) );
  OAI211_X1 U21140 ( .C1(n18450), .C2(n18103), .A(n18090), .B(n18089), .ZN(
        P3_U2878) );
  INV_X1 U21141 ( .A(n18310), .ZN(n18456) );
  AOI22_X1 U21142 ( .A1(n18399), .A2(n18453), .B1(n18451), .B2(n18099), .ZN(
        n18092) );
  AOI22_X1 U21143 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18100), .B1(
        n18428), .B2(n18452), .ZN(n18091) );
  OAI211_X1 U21144 ( .C1(n18456), .C2(n18103), .A(n18092), .B(n18091), .ZN(
        P3_U2879) );
  INV_X1 U21145 ( .A(n18277), .ZN(n18462) );
  AOI22_X1 U21146 ( .A1(n18428), .A2(n18459), .B1(n18457), .B2(n18099), .ZN(
        n18094) );
  AOI22_X1 U21147 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18100), .B1(
        n18399), .B2(n18458), .ZN(n18093) );
  OAI211_X1 U21148 ( .C1(n18462), .C2(n18103), .A(n18094), .B(n18093), .ZN(
        P3_U2880) );
  INV_X1 U21149 ( .A(n18316), .ZN(n18468) );
  AOI22_X1 U21150 ( .A1(n18428), .A2(n18464), .B1(n18463), .B2(n18099), .ZN(
        n18096) );
  AOI22_X1 U21151 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18100), .B1(
        n18399), .B2(n18465), .ZN(n18095) );
  OAI211_X1 U21152 ( .C1(n18468), .C2(n18103), .A(n18096), .B(n18095), .ZN(
        P3_U2881) );
  INV_X1 U21153 ( .A(n18320), .ZN(n18474) );
  AOI22_X1 U21154 ( .A1(n18399), .A2(n18469), .B1(n18470), .B2(n18099), .ZN(
        n18098) );
  AOI22_X1 U21155 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18100), .B1(
        n18428), .B2(n18471), .ZN(n18097) );
  OAI211_X1 U21156 ( .C1(n18474), .C2(n18103), .A(n18098), .B(n18097), .ZN(
        P3_U2882) );
  INV_X1 U21157 ( .A(n18289), .ZN(n18484) );
  AOI22_X1 U21158 ( .A1(n18399), .A2(n18478), .B1(n18476), .B2(n18099), .ZN(
        n18102) );
  AOI22_X1 U21159 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18100), .B1(
        n18428), .B2(n18479), .ZN(n18101) );
  OAI211_X1 U21160 ( .C1(n18484), .C2(n18103), .A(n18102), .B(n18101), .ZN(
        P3_U2883) );
  NOR2_X2 U21161 ( .A1(n18167), .A2(n18294), .ZN(n18185) );
  INV_X1 U21162 ( .A(n18185), .ZN(n18124) );
  NOR2_X1 U21163 ( .A1(n18163), .A2(n18185), .ZN(n18146) );
  NOR2_X1 U21164 ( .A1(n18400), .A2(n18146), .ZN(n18120) );
  AOI22_X1 U21165 ( .A1(n18428), .A2(n18435), .B1(n18429), .B2(n18120), .ZN(
        n18107) );
  AOI221_X1 U21166 ( .B1(n18146), .B2(n18296), .C1(n18146), .C2(n18104), .A(
        n18295), .ZN(n18105) );
  INV_X1 U21167 ( .A(n18105), .ZN(n18121) );
  AOI22_X1 U21168 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18121), .B1(
        n18142), .B2(n18430), .ZN(n18106) );
  OAI211_X1 U21169 ( .C1(n18438), .C2(n18124), .A(n18107), .B(n18106), .ZN(
        P3_U2884) );
  AOI22_X1 U21170 ( .A1(n18142), .A2(n18441), .B1(n18439), .B2(n18120), .ZN(
        n18109) );
  AOI22_X1 U21171 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18121), .B1(
        n18428), .B2(n18440), .ZN(n18108) );
  OAI211_X1 U21172 ( .C1(n18444), .C2(n18124), .A(n18109), .B(n18108), .ZN(
        P3_U2885) );
  AOI22_X1 U21173 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18121), .B1(
        n18445), .B2(n18120), .ZN(n18111) );
  AOI22_X1 U21174 ( .A1(n18428), .A2(n18446), .B1(n18138), .B2(n18447), .ZN(
        n18110) );
  OAI211_X1 U21175 ( .C1(n18450), .C2(n18124), .A(n18111), .B(n18110), .ZN(
        P3_U2886) );
  AOI22_X1 U21176 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18121), .B1(
        n18451), .B2(n18120), .ZN(n18113) );
  AOI22_X1 U21177 ( .A1(n18428), .A2(n18453), .B1(n18142), .B2(n18452), .ZN(
        n18112) );
  OAI211_X1 U21178 ( .C1(n18456), .C2(n18124), .A(n18113), .B(n18112), .ZN(
        P3_U2887) );
  AOI22_X1 U21179 ( .A1(n18428), .A2(n18458), .B1(n18457), .B2(n18120), .ZN(
        n18115) );
  AOI22_X1 U21180 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18121), .B1(
        n18138), .B2(n18459), .ZN(n18114) );
  OAI211_X1 U21181 ( .C1(n18462), .C2(n18124), .A(n18115), .B(n18114), .ZN(
        P3_U2888) );
  AOI22_X1 U21182 ( .A1(n18428), .A2(n18465), .B1(n18463), .B2(n18120), .ZN(
        n18117) );
  AOI22_X1 U21183 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18121), .B1(
        n18138), .B2(n18464), .ZN(n18116) );
  OAI211_X1 U21184 ( .C1(n18468), .C2(n18124), .A(n18117), .B(n18116), .ZN(
        P3_U2889) );
  AOI22_X1 U21185 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18121), .B1(
        n18470), .B2(n18120), .ZN(n18119) );
  AOI22_X1 U21186 ( .A1(n18428), .A2(n18469), .B1(n18138), .B2(n18471), .ZN(
        n18118) );
  OAI211_X1 U21187 ( .C1(n18474), .C2(n18124), .A(n18119), .B(n18118), .ZN(
        P3_U2890) );
  AOI22_X1 U21188 ( .A1(n18428), .A2(n18478), .B1(n18476), .B2(n18120), .ZN(
        n18123) );
  AOI22_X1 U21189 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18121), .B1(
        n18142), .B2(n18479), .ZN(n18122) );
  OAI211_X1 U21190 ( .C1(n18484), .C2(n18124), .A(n18123), .B(n18122), .ZN(
        P3_U2891) );
  NOR2_X2 U21191 ( .A1(n18529), .A2(n18167), .ZN(n18208) );
  INV_X1 U21192 ( .A(n18208), .ZN(n18191) );
  AOI22_X1 U21193 ( .A1(n18430), .A2(n18163), .B1(n18429), .B2(n18141), .ZN(
        n18127) );
  AOI21_X1 U21194 ( .B1(n18530), .B2(n18296), .A(n18260), .ZN(n18214) );
  NAND2_X1 U21195 ( .A1(n18125), .A2(n18214), .ZN(n18143) );
  AOI22_X1 U21196 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18143), .B1(
        n18142), .B2(n18435), .ZN(n18126) );
  OAI211_X1 U21197 ( .C1(n18438), .C2(n18191), .A(n18127), .B(n18126), .ZN(
        P3_U2892) );
  AOI22_X1 U21198 ( .A1(n18142), .A2(n18440), .B1(n18439), .B2(n18141), .ZN(
        n18129) );
  AOI22_X1 U21199 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18143), .B1(
        n18441), .B2(n18163), .ZN(n18128) );
  OAI211_X1 U21200 ( .C1(n18444), .C2(n18191), .A(n18129), .B(n18128), .ZN(
        P3_U2893) );
  AOI22_X1 U21201 ( .A1(n18447), .A2(n18163), .B1(n18445), .B2(n18141), .ZN(
        n18131) );
  AOI22_X1 U21202 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18143), .B1(
        n18138), .B2(n18446), .ZN(n18130) );
  OAI211_X1 U21203 ( .C1(n18450), .C2(n18191), .A(n18131), .B(n18130), .ZN(
        P3_U2894) );
  AOI22_X1 U21204 ( .A1(n18452), .A2(n18163), .B1(n18451), .B2(n18141), .ZN(
        n18133) );
  AOI22_X1 U21205 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18143), .B1(
        n18138), .B2(n18453), .ZN(n18132) );
  OAI211_X1 U21206 ( .C1(n18456), .C2(n18191), .A(n18133), .B(n18132), .ZN(
        P3_U2895) );
  AOI22_X1 U21207 ( .A1(n18142), .A2(n18458), .B1(n18457), .B2(n18141), .ZN(
        n18135) );
  AOI22_X1 U21208 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18143), .B1(
        n18459), .B2(n18163), .ZN(n18134) );
  OAI211_X1 U21209 ( .C1(n18462), .C2(n18191), .A(n18135), .B(n18134), .ZN(
        P3_U2896) );
  AOI22_X1 U21210 ( .A1(n18464), .A2(n18163), .B1(n18463), .B2(n18141), .ZN(
        n18137) );
  AOI22_X1 U21211 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18143), .B1(
        n18138), .B2(n18465), .ZN(n18136) );
  OAI211_X1 U21212 ( .C1(n18468), .C2(n18191), .A(n18137), .B(n18136), .ZN(
        P3_U2897) );
  AOI22_X1 U21213 ( .A1(n18471), .A2(n18163), .B1(n18470), .B2(n18141), .ZN(
        n18140) );
  AOI22_X1 U21214 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18143), .B1(
        n18138), .B2(n18469), .ZN(n18139) );
  OAI211_X1 U21215 ( .C1(n18474), .C2(n18191), .A(n18140), .B(n18139), .ZN(
        P3_U2898) );
  AOI22_X1 U21216 ( .A1(n18142), .A2(n18478), .B1(n18476), .B2(n18141), .ZN(
        n18145) );
  AOI22_X1 U21217 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18143), .B1(
        n18479), .B2(n18163), .ZN(n18144) );
  OAI211_X1 U21218 ( .C1(n18484), .C2(n18191), .A(n18145), .B(n18144), .ZN(
        P3_U2899) );
  NOR2_X2 U21219 ( .A1(n18531), .A2(n18213), .ZN(n18231) );
  INV_X1 U21220 ( .A(n18231), .ZN(n18190) );
  AOI21_X1 U21221 ( .B1(n18191), .B2(n18190), .A(n18400), .ZN(n18162) );
  AOI22_X1 U21222 ( .A1(n18435), .A2(n18163), .B1(n18429), .B2(n18162), .ZN(
        n18149) );
  AOI221_X1 U21223 ( .B1(n18146), .B2(n18191), .C1(n18296), .C2(n18191), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18147) );
  OAI21_X1 U21224 ( .B1(n18231), .B2(n18147), .A(n18354), .ZN(n18164) );
  AOI22_X1 U21225 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18164), .B1(
        n18430), .B2(n18185), .ZN(n18148) );
  OAI211_X1 U21226 ( .C1(n18438), .C2(n18190), .A(n18149), .B(n18148), .ZN(
        P3_U2900) );
  AOI22_X1 U21227 ( .A1(n18441), .A2(n18185), .B1(n18439), .B2(n18162), .ZN(
        n18151) );
  AOI22_X1 U21228 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18164), .B1(
        n18440), .B2(n18163), .ZN(n18150) );
  OAI211_X1 U21229 ( .C1(n18444), .C2(n18190), .A(n18151), .B(n18150), .ZN(
        P3_U2901) );
  AOI22_X1 U21230 ( .A1(n18446), .A2(n18163), .B1(n18445), .B2(n18162), .ZN(
        n18153) );
  AOI22_X1 U21231 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18164), .B1(
        n18447), .B2(n18185), .ZN(n18152) );
  OAI211_X1 U21232 ( .C1(n18450), .C2(n18190), .A(n18153), .B(n18152), .ZN(
        P3_U2902) );
  AOI22_X1 U21233 ( .A1(n18452), .A2(n18185), .B1(n18451), .B2(n18162), .ZN(
        n18155) );
  AOI22_X1 U21234 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18164), .B1(
        n18453), .B2(n18163), .ZN(n18154) );
  OAI211_X1 U21235 ( .C1(n18456), .C2(n18190), .A(n18155), .B(n18154), .ZN(
        P3_U2903) );
  AOI22_X1 U21236 ( .A1(n18458), .A2(n18163), .B1(n18457), .B2(n18162), .ZN(
        n18157) );
  AOI22_X1 U21237 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18164), .B1(
        n18459), .B2(n18185), .ZN(n18156) );
  OAI211_X1 U21238 ( .C1(n18462), .C2(n18190), .A(n18157), .B(n18156), .ZN(
        P3_U2904) );
  AOI22_X1 U21239 ( .A1(n18465), .A2(n18163), .B1(n18463), .B2(n18162), .ZN(
        n18159) );
  AOI22_X1 U21240 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18164), .B1(
        n18464), .B2(n18185), .ZN(n18158) );
  OAI211_X1 U21241 ( .C1(n18468), .C2(n18190), .A(n18159), .B(n18158), .ZN(
        P3_U2905) );
  AOI22_X1 U21242 ( .A1(n18470), .A2(n18162), .B1(n18469), .B2(n18163), .ZN(
        n18161) );
  AOI22_X1 U21243 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18164), .B1(
        n18471), .B2(n18185), .ZN(n18160) );
  OAI211_X1 U21244 ( .C1(n18474), .C2(n18190), .A(n18161), .B(n18160), .ZN(
        P3_U2906) );
  AOI22_X1 U21245 ( .A1(n18479), .A2(n18185), .B1(n18476), .B2(n18162), .ZN(
        n18166) );
  AOI22_X1 U21246 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18164), .B1(
        n18478), .B2(n18163), .ZN(n18165) );
  OAI211_X1 U21247 ( .C1(n18484), .C2(n18190), .A(n18166), .B(n18165), .ZN(
        P3_U2907) );
  NOR2_X2 U21248 ( .A1(n18213), .A2(n18264), .ZN(n18254) );
  INV_X1 U21249 ( .A(n18254), .ZN(n18189) );
  NOR2_X1 U21250 ( .A1(n18213), .A2(n18263), .ZN(n18184) );
  AOI22_X1 U21251 ( .A1(n18435), .A2(n18185), .B1(n18429), .B2(n18184), .ZN(
        n18171) );
  NOR2_X1 U21252 ( .A1(n18530), .A2(n18167), .ZN(n18169) );
  AOI22_X1 U21253 ( .A1(n18434), .A2(n18169), .B1(n18215), .B2(n18168), .ZN(
        n18186) );
  AOI22_X1 U21254 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18186), .B1(
        n18430), .B2(n18208), .ZN(n18170) );
  OAI211_X1 U21255 ( .C1(n18438), .C2(n18189), .A(n18171), .B(n18170), .ZN(
        P3_U2908) );
  AOI22_X1 U21256 ( .A1(n18441), .A2(n18208), .B1(n18439), .B2(n18184), .ZN(
        n18173) );
  AOI22_X1 U21257 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18186), .B1(
        n18440), .B2(n18185), .ZN(n18172) );
  OAI211_X1 U21258 ( .C1(n18444), .C2(n18189), .A(n18173), .B(n18172), .ZN(
        P3_U2909) );
  AOI22_X1 U21259 ( .A1(n18447), .A2(n18208), .B1(n18445), .B2(n18184), .ZN(
        n18175) );
  AOI22_X1 U21260 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18186), .B1(
        n18446), .B2(n18185), .ZN(n18174) );
  OAI211_X1 U21261 ( .C1(n18450), .C2(n18189), .A(n18175), .B(n18174), .ZN(
        P3_U2910) );
  AOI22_X1 U21262 ( .A1(n18452), .A2(n18208), .B1(n18451), .B2(n18184), .ZN(
        n18177) );
  AOI22_X1 U21263 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18186), .B1(
        n18453), .B2(n18185), .ZN(n18176) );
  OAI211_X1 U21264 ( .C1(n18456), .C2(n18189), .A(n18177), .B(n18176), .ZN(
        P3_U2911) );
  AOI22_X1 U21265 ( .A1(n18459), .A2(n18208), .B1(n18457), .B2(n18184), .ZN(
        n18179) );
  AOI22_X1 U21266 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18186), .B1(
        n18458), .B2(n18185), .ZN(n18178) );
  OAI211_X1 U21267 ( .C1(n18462), .C2(n18189), .A(n18179), .B(n18178), .ZN(
        P3_U2912) );
  AOI22_X1 U21268 ( .A1(n18465), .A2(n18185), .B1(n18463), .B2(n18184), .ZN(
        n18181) );
  AOI22_X1 U21269 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18186), .B1(
        n18464), .B2(n18208), .ZN(n18180) );
  OAI211_X1 U21270 ( .C1(n18468), .C2(n18189), .A(n18181), .B(n18180), .ZN(
        P3_U2913) );
  AOI22_X1 U21271 ( .A1(n18470), .A2(n18184), .B1(n18469), .B2(n18185), .ZN(
        n18183) );
  AOI22_X1 U21272 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18186), .B1(
        n18471), .B2(n18208), .ZN(n18182) );
  OAI211_X1 U21273 ( .C1(n18474), .C2(n18189), .A(n18183), .B(n18182), .ZN(
        P3_U2914) );
  AOI22_X1 U21274 ( .A1(n18479), .A2(n18208), .B1(n18476), .B2(n18184), .ZN(
        n18188) );
  AOI22_X1 U21275 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18186), .B1(
        n18478), .B2(n18185), .ZN(n18187) );
  OAI211_X1 U21276 ( .C1(n18484), .C2(n18189), .A(n18188), .B(n18187), .ZN(
        P3_U2915) );
  NOR2_X2 U21277 ( .A1(n18213), .A2(n18294), .ZN(n18288) );
  INV_X1 U21278 ( .A(n18288), .ZN(n18212) );
  NAND2_X1 U21279 ( .A1(n18189), .A2(n18212), .ZN(n18236) );
  NAND2_X1 U21280 ( .A1(n18191), .A2(n18190), .ZN(n18192) );
  OAI221_X1 U21281 ( .B1(n18236), .B2(n18406), .C1(n18236), .C2(n18192), .A(
        n18404), .ZN(n18209) );
  AND2_X1 U21282 ( .A1(n18554), .A2(n18236), .ZN(n18207) );
  AOI22_X1 U21283 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18209), .B1(
        n18429), .B2(n18207), .ZN(n18194) );
  AOI22_X1 U21284 ( .A1(n18430), .A2(n18231), .B1(n18435), .B2(n18208), .ZN(
        n18193) );
  OAI211_X1 U21285 ( .C1(n18438), .C2(n18212), .A(n18194), .B(n18193), .ZN(
        P3_U2916) );
  AOI22_X1 U21286 ( .A1(n18441), .A2(n18231), .B1(n18439), .B2(n18207), .ZN(
        n18196) );
  AOI22_X1 U21287 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18209), .B1(
        n18440), .B2(n18208), .ZN(n18195) );
  OAI211_X1 U21288 ( .C1(n18444), .C2(n18212), .A(n18196), .B(n18195), .ZN(
        P3_U2917) );
  AOI22_X1 U21289 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18209), .B1(
        n18445), .B2(n18207), .ZN(n18198) );
  AOI22_X1 U21290 ( .A1(n18446), .A2(n18208), .B1(n18447), .B2(n18231), .ZN(
        n18197) );
  OAI211_X1 U21291 ( .C1(n18450), .C2(n18212), .A(n18198), .B(n18197), .ZN(
        P3_U2918) );
  AOI22_X1 U21292 ( .A1(n18452), .A2(n18231), .B1(n18451), .B2(n18207), .ZN(
        n18200) );
  AOI22_X1 U21293 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18209), .B1(
        n18453), .B2(n18208), .ZN(n18199) );
  OAI211_X1 U21294 ( .C1(n18456), .C2(n18212), .A(n18200), .B(n18199), .ZN(
        P3_U2919) );
  AOI22_X1 U21295 ( .A1(n18458), .A2(n18208), .B1(n18457), .B2(n18207), .ZN(
        n18202) );
  AOI22_X1 U21296 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18209), .B1(
        n18459), .B2(n18231), .ZN(n18201) );
  OAI211_X1 U21297 ( .C1(n18462), .C2(n18212), .A(n18202), .B(n18201), .ZN(
        P3_U2920) );
  AOI22_X1 U21298 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18209), .B1(
        n18463), .B2(n18207), .ZN(n18204) );
  AOI22_X1 U21299 ( .A1(n18464), .A2(n18231), .B1(n18465), .B2(n18208), .ZN(
        n18203) );
  OAI211_X1 U21300 ( .C1(n18468), .C2(n18212), .A(n18204), .B(n18203), .ZN(
        P3_U2921) );
  AOI22_X1 U21301 ( .A1(n18470), .A2(n18207), .B1(n18469), .B2(n18208), .ZN(
        n18206) );
  AOI22_X1 U21302 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18209), .B1(
        n18471), .B2(n18231), .ZN(n18205) );
  OAI211_X1 U21303 ( .C1(n18474), .C2(n18212), .A(n18206), .B(n18205), .ZN(
        P3_U2922) );
  AOI22_X1 U21304 ( .A1(n18478), .A2(n18208), .B1(n18476), .B2(n18207), .ZN(
        n18211) );
  AOI22_X1 U21305 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18209), .B1(
        n18479), .B2(n18231), .ZN(n18210) );
  OAI211_X1 U21306 ( .C1(n18484), .C2(n18212), .A(n18211), .B(n18210), .ZN(
        P3_U2923) );
  NOR2_X2 U21307 ( .A1(n18529), .A2(n18213), .ZN(n18327) );
  INV_X1 U21308 ( .A(n18327), .ZN(n18235) );
  AOI22_X1 U21309 ( .A1(n18430), .A2(n18254), .B1(n18429), .B2(n18230), .ZN(
        n18217) );
  NAND2_X1 U21310 ( .A1(n18215), .A2(n18214), .ZN(n18232) );
  AOI22_X1 U21311 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18232), .B1(
        n18435), .B2(n18231), .ZN(n18216) );
  OAI211_X1 U21312 ( .C1(n18438), .C2(n18235), .A(n18217), .B(n18216), .ZN(
        P3_U2924) );
  AOI22_X1 U21313 ( .A1(n18441), .A2(n18254), .B1(n18439), .B2(n18230), .ZN(
        n18219) );
  AOI22_X1 U21314 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18232), .B1(
        n18440), .B2(n18231), .ZN(n18218) );
  OAI211_X1 U21315 ( .C1(n18444), .C2(n18235), .A(n18219), .B(n18218), .ZN(
        P3_U2925) );
  AOI22_X1 U21316 ( .A1(n18446), .A2(n18231), .B1(n18445), .B2(n18230), .ZN(
        n18221) );
  AOI22_X1 U21317 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18232), .B1(
        n18447), .B2(n18254), .ZN(n18220) );
  OAI211_X1 U21318 ( .C1(n18450), .C2(n18235), .A(n18221), .B(n18220), .ZN(
        P3_U2926) );
  AOI22_X1 U21319 ( .A1(n18452), .A2(n18254), .B1(n18451), .B2(n18230), .ZN(
        n18223) );
  AOI22_X1 U21320 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18232), .B1(
        n18453), .B2(n18231), .ZN(n18222) );
  OAI211_X1 U21321 ( .C1(n18456), .C2(n18235), .A(n18223), .B(n18222), .ZN(
        P3_U2927) );
  AOI22_X1 U21322 ( .A1(n18459), .A2(n18254), .B1(n18457), .B2(n18230), .ZN(
        n18225) );
  AOI22_X1 U21323 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18232), .B1(
        n18458), .B2(n18231), .ZN(n18224) );
  OAI211_X1 U21324 ( .C1(n18462), .C2(n18235), .A(n18225), .B(n18224), .ZN(
        P3_U2928) );
  AOI22_X1 U21325 ( .A1(n18464), .A2(n18254), .B1(n18463), .B2(n18230), .ZN(
        n18227) );
  AOI22_X1 U21326 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18232), .B1(
        n18465), .B2(n18231), .ZN(n18226) );
  OAI211_X1 U21327 ( .C1(n18468), .C2(n18235), .A(n18227), .B(n18226), .ZN(
        P3_U2929) );
  AOI22_X1 U21328 ( .A1(n18470), .A2(n18230), .B1(n18469), .B2(n18231), .ZN(
        n18229) );
  AOI22_X1 U21329 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18232), .B1(
        n18471), .B2(n18254), .ZN(n18228) );
  OAI211_X1 U21330 ( .C1(n18474), .C2(n18235), .A(n18229), .B(n18228), .ZN(
        P3_U2930) );
  AOI22_X1 U21331 ( .A1(n18478), .A2(n18231), .B1(n18476), .B2(n18230), .ZN(
        n18234) );
  AOI22_X1 U21332 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18232), .B1(
        n18479), .B2(n18254), .ZN(n18233) );
  OAI211_X1 U21333 ( .C1(n18484), .C2(n18235), .A(n18234), .B(n18233), .ZN(
        P3_U2931) );
  NOR2_X2 U21334 ( .A1(n18531), .A2(n18331), .ZN(n18347) );
  INV_X1 U21335 ( .A(n18347), .ZN(n18257) );
  NOR2_X1 U21336 ( .A1(n18327), .A2(n18347), .ZN(n18298) );
  NOR2_X1 U21337 ( .A1(n18400), .A2(n18298), .ZN(n18252) );
  AOI22_X1 U21338 ( .A1(n18435), .A2(n18254), .B1(n18429), .B2(n18252), .ZN(
        n18239) );
  INV_X1 U21339 ( .A(n18298), .ZN(n18237) );
  OAI221_X1 U21340 ( .B1(n18237), .B2(n18406), .C1(n18237), .C2(n18236), .A(
        n18404), .ZN(n18253) );
  AOI22_X1 U21341 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18253), .B1(
        n18430), .B2(n18288), .ZN(n18238) );
  OAI211_X1 U21342 ( .C1(n18438), .C2(n18257), .A(n18239), .B(n18238), .ZN(
        P3_U2932) );
  AOI22_X1 U21343 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18253), .B1(
        n18439), .B2(n18252), .ZN(n18241) );
  AOI22_X1 U21344 ( .A1(n18440), .A2(n18254), .B1(n18441), .B2(n18288), .ZN(
        n18240) );
  OAI211_X1 U21345 ( .C1(n18444), .C2(n18257), .A(n18241), .B(n18240), .ZN(
        P3_U2933) );
  AOI22_X1 U21346 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18253), .B1(
        n18445), .B2(n18252), .ZN(n18243) );
  AOI22_X1 U21347 ( .A1(n18446), .A2(n18254), .B1(n18447), .B2(n18288), .ZN(
        n18242) );
  OAI211_X1 U21348 ( .C1(n18450), .C2(n18257), .A(n18243), .B(n18242), .ZN(
        P3_U2934) );
  AOI22_X1 U21349 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18253), .B1(
        n18451), .B2(n18252), .ZN(n18245) );
  AOI22_X1 U21350 ( .A1(n18452), .A2(n18288), .B1(n18453), .B2(n18254), .ZN(
        n18244) );
  OAI211_X1 U21351 ( .C1(n18456), .C2(n18257), .A(n18245), .B(n18244), .ZN(
        P3_U2935) );
  AOI22_X1 U21352 ( .A1(n18459), .A2(n18288), .B1(n18457), .B2(n18252), .ZN(
        n18247) );
  AOI22_X1 U21353 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18253), .B1(
        n18458), .B2(n18254), .ZN(n18246) );
  OAI211_X1 U21354 ( .C1(n18462), .C2(n18257), .A(n18247), .B(n18246), .ZN(
        P3_U2936) );
  AOI22_X1 U21355 ( .A1(n18464), .A2(n18288), .B1(n18463), .B2(n18252), .ZN(
        n18249) );
  AOI22_X1 U21356 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18253), .B1(
        n18465), .B2(n18254), .ZN(n18248) );
  OAI211_X1 U21357 ( .C1(n18468), .C2(n18257), .A(n18249), .B(n18248), .ZN(
        P3_U2937) );
  AOI22_X1 U21358 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18253), .B1(
        n18470), .B2(n18252), .ZN(n18251) );
  AOI22_X1 U21359 ( .A1(n18471), .A2(n18288), .B1(n18469), .B2(n18254), .ZN(
        n18250) );
  OAI211_X1 U21360 ( .C1(n18474), .C2(n18257), .A(n18251), .B(n18250), .ZN(
        P3_U2938) );
  AOI22_X1 U21361 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18253), .B1(
        n18476), .B2(n18252), .ZN(n18256) );
  AOI22_X1 U21362 ( .A1(n18479), .A2(n18288), .B1(n18478), .B2(n18254), .ZN(
        n18255) );
  OAI211_X1 U21363 ( .C1(n18484), .C2(n18257), .A(n18256), .B(n18255), .ZN(
        P3_U2939) );
  OR2_X1 U21364 ( .A1(n18258), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18261) );
  NAND2_X1 U21365 ( .A1(n18352), .A2(n18530), .ZN(n18259) );
  OAI22_X1 U21366 ( .A1(n18262), .A2(n18261), .B1(n18260), .B2(n18259), .ZN(
        n18292) );
  NOR2_X1 U21367 ( .A1(n18331), .A2(n18263), .ZN(n18287) );
  AOI22_X1 U21368 ( .A1(n18430), .A2(n18327), .B1(n18429), .B2(n18287), .ZN(
        n18266) );
  NOR2_X1 U21369 ( .A1(n18331), .A2(n18264), .ZN(n18372) );
  AOI22_X1 U21370 ( .A1(n18300), .A2(n18372), .B1(n18435), .B2(n18288), .ZN(
        n18265) );
  OAI211_X1 U21371 ( .C1(n18267), .C2(n18292), .A(n18266), .B(n18265), .ZN(
        P3_U2940) );
  AOI22_X1 U21372 ( .A1(n18440), .A2(n18288), .B1(n18439), .B2(n18287), .ZN(
        n18270) );
  INV_X1 U21373 ( .A(n18372), .ZN(n18299) );
  INV_X1 U21374 ( .A(n18299), .ZN(n18368) );
  AOI22_X1 U21375 ( .A1(n18268), .A2(n18368), .B1(n18441), .B2(n18327), .ZN(
        n18269) );
  OAI211_X1 U21376 ( .C1(n18271), .C2(n18292), .A(n18270), .B(n18269), .ZN(
        P3_U2941) );
  AOI22_X1 U21377 ( .A1(n18446), .A2(n18288), .B1(n18445), .B2(n18287), .ZN(
        n18273) );
  AOI22_X1 U21378 ( .A1(n18306), .A2(n18372), .B1(n18447), .B2(n18327), .ZN(
        n18272) );
  OAI211_X1 U21379 ( .C1(n18274), .C2(n18292), .A(n18273), .B(n18272), .ZN(
        P3_U2942) );
  AOI22_X1 U21380 ( .A1(n18453), .A2(n18288), .B1(n18451), .B2(n18287), .ZN(
        n18276) );
  AOI22_X1 U21381 ( .A1(n18452), .A2(n18327), .B1(n18310), .B2(n18368), .ZN(
        n18275) );
  OAI211_X1 U21382 ( .C1(n20910), .C2(n18292), .A(n18276), .B(n18275), .ZN(
        P3_U2943) );
  AOI22_X1 U21383 ( .A1(n18459), .A2(n18327), .B1(n18457), .B2(n18287), .ZN(
        n18279) );
  AOI22_X1 U21384 ( .A1(n18277), .A2(n18372), .B1(n18458), .B2(n18288), .ZN(
        n18278) );
  OAI211_X1 U21385 ( .C1(n18280), .C2(n18292), .A(n18279), .B(n18278), .ZN(
        P3_U2944) );
  AOI22_X1 U21386 ( .A1(n18465), .A2(n18288), .B1(n18463), .B2(n18287), .ZN(
        n18282) );
  AOI22_X1 U21387 ( .A1(n18464), .A2(n18327), .B1(n18316), .B2(n18368), .ZN(
        n18281) );
  OAI211_X1 U21388 ( .C1(n18283), .C2(n18292), .A(n18282), .B(n18281), .ZN(
        P3_U2945) );
  AOI22_X1 U21389 ( .A1(n18471), .A2(n18327), .B1(n18470), .B2(n18287), .ZN(
        n18285) );
  AOI22_X1 U21390 ( .A1(n18320), .A2(n18372), .B1(n18469), .B2(n18288), .ZN(
        n18284) );
  OAI211_X1 U21391 ( .C1(n18286), .C2(n18292), .A(n18285), .B(n18284), .ZN(
        P3_U2946) );
  AOI22_X1 U21392 ( .A1(n18479), .A2(n18327), .B1(n18476), .B2(n18287), .ZN(
        n18291) );
  AOI22_X1 U21393 ( .A1(n18289), .A2(n18372), .B1(n18478), .B2(n18288), .ZN(
        n18290) );
  OAI211_X1 U21394 ( .C1(n18293), .C2(n18292), .A(n18291), .B(n18290), .ZN(
        P3_U2947) );
  NOR2_X1 U21395 ( .A1(n18331), .A2(n18294), .ZN(n18394) );
  CLKBUF_X1 U21396 ( .A(n18394), .Z(n18390) );
  NOR2_X1 U21397 ( .A1(n18368), .A2(n18390), .ZN(n18297) );
  AOI221_X1 U21398 ( .B1(n18298), .B2(n18297), .C1(n18296), .C2(n18297), .A(
        n18295), .ZN(n18324) );
  INV_X1 U21399 ( .A(n18394), .ZN(n18330) );
  AOI21_X1 U21400 ( .B1(n18299), .B2(n18330), .A(n18400), .ZN(n18325) );
  AOI22_X1 U21401 ( .A1(n18430), .A2(n18347), .B1(n18429), .B2(n18325), .ZN(
        n18302) );
  AOI22_X1 U21402 ( .A1(n18300), .A2(n18390), .B1(n18435), .B2(n18327), .ZN(
        n18301) );
  OAI211_X1 U21403 ( .C1(n18324), .C2(n18303), .A(n18302), .B(n18301), .ZN(
        P3_U2948) );
  INV_X1 U21404 ( .A(n18324), .ZN(n18326) );
  AOI22_X1 U21405 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18326), .B1(
        n18439), .B2(n18325), .ZN(n18305) );
  AOI22_X1 U21406 ( .A1(n18440), .A2(n18327), .B1(n18441), .B2(n18347), .ZN(
        n18304) );
  OAI211_X1 U21407 ( .C1(n18444), .C2(n18330), .A(n18305), .B(n18304), .ZN(
        P3_U2949) );
  AOI22_X1 U21408 ( .A1(n18446), .A2(n18327), .B1(n18445), .B2(n18325), .ZN(
        n18308) );
  AOI22_X1 U21409 ( .A1(n18306), .A2(n18390), .B1(n18447), .B2(n18347), .ZN(
        n18307) );
  OAI211_X1 U21410 ( .C1(n18324), .C2(n18309), .A(n18308), .B(n18307), .ZN(
        P3_U2950) );
  AOI22_X1 U21411 ( .A1(n18453), .A2(n18327), .B1(n18451), .B2(n18325), .ZN(
        n18312) );
  AOI22_X1 U21412 ( .A1(n18452), .A2(n18347), .B1(n18310), .B2(n18394), .ZN(
        n18311) );
  OAI211_X1 U21413 ( .C1(n18324), .C2(n18313), .A(n18312), .B(n18311), .ZN(
        P3_U2951) );
  AOI22_X1 U21414 ( .A1(n18458), .A2(n18327), .B1(n18457), .B2(n18325), .ZN(
        n18315) );
  AOI22_X1 U21415 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18326), .B1(
        n18459), .B2(n18347), .ZN(n18314) );
  OAI211_X1 U21416 ( .C1(n18462), .C2(n18330), .A(n18315), .B(n18314), .ZN(
        P3_U2952) );
  AOI22_X1 U21417 ( .A1(n18465), .A2(n18327), .B1(n18463), .B2(n18325), .ZN(
        n18318) );
  AOI22_X1 U21418 ( .A1(n18464), .A2(n18347), .B1(n18316), .B2(n18394), .ZN(
        n18317) );
  OAI211_X1 U21419 ( .C1(n18324), .C2(n18319), .A(n18318), .B(n18317), .ZN(
        P3_U2953) );
  AOI22_X1 U21420 ( .A1(n18470), .A2(n18325), .B1(n18469), .B2(n18327), .ZN(
        n18322) );
  AOI22_X1 U21421 ( .A1(n18471), .A2(n18347), .B1(n18320), .B2(n18390), .ZN(
        n18321) );
  OAI211_X1 U21422 ( .C1(n18324), .C2(n18323), .A(n18322), .B(n18321), .ZN(
        P3_U2954) );
  AOI22_X1 U21423 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18326), .B1(
        n18476), .B2(n18325), .ZN(n18329) );
  AOI22_X1 U21424 ( .A1(n18479), .A2(n18347), .B1(n18478), .B2(n18327), .ZN(
        n18328) );
  OAI211_X1 U21425 ( .C1(n18484), .C2(n18330), .A(n18329), .B(n18328), .ZN(
        P3_U2955) );
  NOR2_X2 U21426 ( .A1(n18529), .A2(n18331), .ZN(n18423) );
  INV_X1 U21427 ( .A(n18423), .ZN(n18403) );
  NOR2_X1 U21428 ( .A1(n18530), .A2(n18331), .ZN(n18377) );
  AND2_X1 U21429 ( .A1(n18554), .A2(n18377), .ZN(n18346) );
  AOI22_X1 U21430 ( .A1(n18430), .A2(n18372), .B1(n18429), .B2(n18346), .ZN(
        n18333) );
  OAI211_X1 U21431 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18434), .A(
        n18432), .B(n18352), .ZN(n18348) );
  AOI22_X1 U21432 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18348), .B1(
        n18435), .B2(n18347), .ZN(n18332) );
  OAI211_X1 U21433 ( .C1(n18438), .C2(n18403), .A(n18333), .B(n18332), .ZN(
        P3_U2956) );
  AOI22_X1 U21434 ( .A1(n18441), .A2(n18372), .B1(n18439), .B2(n18346), .ZN(
        n18335) );
  AOI22_X1 U21435 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18348), .B1(
        n18440), .B2(n18347), .ZN(n18334) );
  OAI211_X1 U21436 ( .C1(n18444), .C2(n18403), .A(n18335), .B(n18334), .ZN(
        P3_U2957) );
  AOI22_X1 U21437 ( .A1(n18447), .A2(n18372), .B1(n18445), .B2(n18346), .ZN(
        n18337) );
  AOI22_X1 U21438 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18348), .B1(
        n18446), .B2(n18347), .ZN(n18336) );
  OAI211_X1 U21439 ( .C1(n18450), .C2(n18403), .A(n18337), .B(n18336), .ZN(
        P3_U2958) );
  AOI22_X1 U21440 ( .A1(n18452), .A2(n18372), .B1(n18451), .B2(n18346), .ZN(
        n18339) );
  AOI22_X1 U21441 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18348), .B1(
        n18453), .B2(n18347), .ZN(n18338) );
  OAI211_X1 U21442 ( .C1(n18456), .C2(n18403), .A(n18339), .B(n18338), .ZN(
        P3_U2959) );
  AOI22_X1 U21443 ( .A1(n18458), .A2(n18347), .B1(n18457), .B2(n18346), .ZN(
        n18341) );
  AOI22_X1 U21444 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18348), .B1(
        n18459), .B2(n18368), .ZN(n18340) );
  OAI211_X1 U21445 ( .C1(n18462), .C2(n18403), .A(n18341), .B(n18340), .ZN(
        P3_U2960) );
  AOI22_X1 U21446 ( .A1(n18465), .A2(n18347), .B1(n18463), .B2(n18346), .ZN(
        n18343) );
  AOI22_X1 U21447 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18348), .B1(
        n18464), .B2(n18368), .ZN(n18342) );
  OAI211_X1 U21448 ( .C1(n18468), .C2(n18403), .A(n18343), .B(n18342), .ZN(
        P3_U2961) );
  AOI22_X1 U21449 ( .A1(n18471), .A2(n18372), .B1(n18470), .B2(n18346), .ZN(
        n18345) );
  AOI22_X1 U21450 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18348), .B1(
        n18469), .B2(n18347), .ZN(n18344) );
  OAI211_X1 U21451 ( .C1(n18474), .C2(n18403), .A(n18345), .B(n18344), .ZN(
        P3_U2962) );
  AOI22_X1 U21452 ( .A1(n18478), .A2(n18347), .B1(n18476), .B2(n18346), .ZN(
        n18350) );
  AOI22_X1 U21453 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18348), .B1(
        n18479), .B2(n18368), .ZN(n18349) );
  OAI211_X1 U21454 ( .C1(n18484), .C2(n18403), .A(n18350), .B(n18349), .ZN(
        P3_U2963) );
  INV_X1 U21455 ( .A(n18433), .ZN(n18376) );
  NOR2_X2 U21456 ( .A1(n18376), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18477) );
  INV_X1 U21457 ( .A(n18477), .ZN(n18402) );
  AOI21_X1 U21458 ( .B1(n18403), .B2(n18402), .A(n18400), .ZN(n18371) );
  AOI22_X1 U21459 ( .A1(n18430), .A2(n18394), .B1(n18429), .B2(n18371), .ZN(
        n18357) );
  NAND3_X1 U21460 ( .A1(n18352), .A2(n18406), .A3(n18351), .ZN(n18353) );
  AOI21_X1 U21461 ( .B1(n18403), .B2(n18353), .A(P3_STATE2_REG_3__SCAN_IN), 
        .ZN(n18355) );
  OAI21_X1 U21462 ( .B1(n18477), .B2(n18355), .A(n18354), .ZN(n18373) );
  AOI22_X1 U21463 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18373), .B1(
        n18435), .B2(n18368), .ZN(n18356) );
  OAI211_X1 U21464 ( .C1(n18438), .C2(n18402), .A(n18357), .B(n18356), .ZN(
        P3_U2964) );
  AOI22_X1 U21465 ( .A1(n18441), .A2(n18390), .B1(n18439), .B2(n18371), .ZN(
        n18359) );
  AOI22_X1 U21466 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18373), .B1(
        n18440), .B2(n18368), .ZN(n18358) );
  OAI211_X1 U21467 ( .C1(n18444), .C2(n18402), .A(n18359), .B(n18358), .ZN(
        P3_U2965) );
  AOI22_X1 U21468 ( .A1(n18447), .A2(n18390), .B1(n18445), .B2(n18371), .ZN(
        n18361) );
  AOI22_X1 U21469 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18373), .B1(
        n18446), .B2(n18368), .ZN(n18360) );
  OAI211_X1 U21470 ( .C1(n18450), .C2(n18402), .A(n18361), .B(n18360), .ZN(
        P3_U2966) );
  AOI22_X1 U21471 ( .A1(n18452), .A2(n18390), .B1(n18451), .B2(n18371), .ZN(
        n18363) );
  AOI22_X1 U21472 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18373), .B1(
        n18453), .B2(n18368), .ZN(n18362) );
  OAI211_X1 U21473 ( .C1(n18456), .C2(n18402), .A(n18363), .B(n18362), .ZN(
        P3_U2967) );
  AOI22_X1 U21474 ( .A1(n18459), .A2(n18394), .B1(n18457), .B2(n18371), .ZN(
        n18365) );
  AOI22_X1 U21475 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18373), .B1(
        n18458), .B2(n18368), .ZN(n18364) );
  OAI211_X1 U21476 ( .C1(n18462), .C2(n18402), .A(n18365), .B(n18364), .ZN(
        P3_U2968) );
  AOI22_X1 U21477 ( .A1(n18464), .A2(n18390), .B1(n18463), .B2(n18371), .ZN(
        n18367) );
  AOI22_X1 U21478 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18373), .B1(
        n18465), .B2(n18368), .ZN(n18366) );
  OAI211_X1 U21479 ( .C1(n18468), .C2(n18402), .A(n18367), .B(n18366), .ZN(
        P3_U2969) );
  AOI22_X1 U21480 ( .A1(n18471), .A2(n18394), .B1(n18470), .B2(n18371), .ZN(
        n18370) );
  AOI22_X1 U21481 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18373), .B1(
        n18469), .B2(n18368), .ZN(n18369) );
  OAI211_X1 U21482 ( .C1(n18474), .C2(n18402), .A(n18370), .B(n18369), .ZN(
        P3_U2970) );
  AOI22_X1 U21483 ( .A1(n18478), .A2(n18372), .B1(n18476), .B2(n18371), .ZN(
        n18375) );
  AOI22_X1 U21484 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18373), .B1(
        n18479), .B2(n18394), .ZN(n18374) );
  OAI211_X1 U21485 ( .C1(n18484), .C2(n18402), .A(n18375), .B(n18374), .ZN(
        P3_U2971) );
  NOR2_X1 U21486 ( .A1(n18400), .A2(n18376), .ZN(n18393) );
  AOI22_X1 U21487 ( .A1(n18430), .A2(n18423), .B1(n18429), .B2(n18393), .ZN(
        n18379) );
  AOI22_X1 U21488 ( .A1(n18434), .A2(n18377), .B1(n18433), .B2(n18432), .ZN(
        n18395) );
  AOI22_X1 U21489 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18395), .B1(
        n18435), .B2(n18394), .ZN(n18378) );
  OAI211_X1 U21490 ( .C1(n18438), .C2(n18398), .A(n18379), .B(n18378), .ZN(
        P3_U2972) );
  AOI22_X1 U21491 ( .A1(n18441), .A2(n18423), .B1(n18439), .B2(n18393), .ZN(
        n18381) );
  AOI22_X1 U21492 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18395), .B1(
        n18440), .B2(n18390), .ZN(n18380) );
  OAI211_X1 U21493 ( .C1(n18398), .C2(n18444), .A(n18381), .B(n18380), .ZN(
        P3_U2973) );
  AOI22_X1 U21494 ( .A1(n18446), .A2(n18394), .B1(n18445), .B2(n18393), .ZN(
        n18383) );
  AOI22_X1 U21495 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18395), .B1(
        n18447), .B2(n18423), .ZN(n18382) );
  OAI211_X1 U21496 ( .C1(n18398), .C2(n18450), .A(n18383), .B(n18382), .ZN(
        P3_U2974) );
  AOI22_X1 U21497 ( .A1(n18452), .A2(n18423), .B1(n18451), .B2(n18393), .ZN(
        n18385) );
  AOI22_X1 U21498 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18395), .B1(
        n18453), .B2(n18394), .ZN(n18384) );
  OAI211_X1 U21499 ( .C1(n18398), .C2(n18456), .A(n18385), .B(n18384), .ZN(
        P3_U2975) );
  AOI22_X1 U21500 ( .A1(n18459), .A2(n18423), .B1(n18457), .B2(n18393), .ZN(
        n18387) );
  AOI22_X1 U21501 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18395), .B1(
        n18458), .B2(n18390), .ZN(n18386) );
  OAI211_X1 U21502 ( .C1(n18398), .C2(n18462), .A(n18387), .B(n18386), .ZN(
        P3_U2976) );
  AOI22_X1 U21503 ( .A1(n18465), .A2(n18390), .B1(n18463), .B2(n18393), .ZN(
        n18389) );
  AOI22_X1 U21504 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18395), .B1(
        n18464), .B2(n18423), .ZN(n18388) );
  OAI211_X1 U21505 ( .C1(n18398), .C2(n18468), .A(n18389), .B(n18388), .ZN(
        P3_U2977) );
  AOI22_X1 U21506 ( .A1(n18470), .A2(n18393), .B1(n18469), .B2(n18390), .ZN(
        n18392) );
  AOI22_X1 U21507 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18395), .B1(
        n18471), .B2(n18423), .ZN(n18391) );
  OAI211_X1 U21508 ( .C1(n18398), .C2(n18474), .A(n18392), .B(n18391), .ZN(
        P3_U2978) );
  AOI22_X1 U21509 ( .A1(n18479), .A2(n18423), .B1(n18476), .B2(n18393), .ZN(
        n18397) );
  AOI22_X1 U21510 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18395), .B1(
        n18478), .B2(n18394), .ZN(n18396) );
  OAI211_X1 U21511 ( .C1(n18398), .C2(n18484), .A(n18397), .B(n18396), .ZN(
        P3_U2979) );
  INV_X1 U21512 ( .A(n18399), .ZN(n18427) );
  NOR2_X1 U21513 ( .A1(n18400), .A2(n18401), .ZN(n18422) );
  AOI22_X1 U21514 ( .A1(n18430), .A2(n18477), .B1(n18429), .B2(n18422), .ZN(
        n18409) );
  INV_X1 U21515 ( .A(n18401), .ZN(n18407) );
  NAND2_X1 U21516 ( .A1(n18403), .A2(n18402), .ZN(n18405) );
  OAI221_X1 U21517 ( .B1(n18407), .B2(n18406), .C1(n18407), .C2(n18405), .A(
        n18404), .ZN(n18424) );
  AOI22_X1 U21518 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18424), .B1(
        n18435), .B2(n18423), .ZN(n18408) );
  OAI211_X1 U21519 ( .C1(n18427), .C2(n18438), .A(n18409), .B(n18408), .ZN(
        P3_U2980) );
  AOI22_X1 U21520 ( .A1(n18441), .A2(n18477), .B1(n18439), .B2(n18422), .ZN(
        n18411) );
  AOI22_X1 U21521 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18424), .B1(
        n18440), .B2(n18423), .ZN(n18410) );
  OAI211_X1 U21522 ( .C1(n18427), .C2(n18444), .A(n18411), .B(n18410), .ZN(
        P3_U2981) );
  AOI22_X1 U21523 ( .A1(n18446), .A2(n18423), .B1(n18445), .B2(n18422), .ZN(
        n18413) );
  AOI22_X1 U21524 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18424), .B1(
        n18447), .B2(n18477), .ZN(n18412) );
  OAI211_X1 U21525 ( .C1(n18427), .C2(n18450), .A(n18413), .B(n18412), .ZN(
        P3_U2982) );
  AOI22_X1 U21526 ( .A1(n18452), .A2(n18477), .B1(n18451), .B2(n18422), .ZN(
        n18415) );
  AOI22_X1 U21527 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18424), .B1(
        n18453), .B2(n18423), .ZN(n18414) );
  OAI211_X1 U21528 ( .C1(n18427), .C2(n18456), .A(n18415), .B(n18414), .ZN(
        P3_U2983) );
  AOI22_X1 U21529 ( .A1(n18458), .A2(n18423), .B1(n18457), .B2(n18422), .ZN(
        n18417) );
  AOI22_X1 U21530 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18424), .B1(
        n18459), .B2(n18477), .ZN(n18416) );
  OAI211_X1 U21531 ( .C1(n18427), .C2(n18462), .A(n18417), .B(n18416), .ZN(
        P3_U2984) );
  AOI22_X1 U21532 ( .A1(n18464), .A2(n18477), .B1(n18463), .B2(n18422), .ZN(
        n18419) );
  AOI22_X1 U21533 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18424), .B1(
        n18465), .B2(n18423), .ZN(n18418) );
  OAI211_X1 U21534 ( .C1(n18427), .C2(n18468), .A(n18419), .B(n18418), .ZN(
        P3_U2985) );
  AOI22_X1 U21535 ( .A1(n18470), .A2(n18422), .B1(n18469), .B2(n18423), .ZN(
        n18421) );
  AOI22_X1 U21536 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18424), .B1(
        n18471), .B2(n18477), .ZN(n18420) );
  OAI211_X1 U21537 ( .C1(n18427), .C2(n18474), .A(n18421), .B(n18420), .ZN(
        P3_U2986) );
  AOI22_X1 U21538 ( .A1(n18478), .A2(n18423), .B1(n18476), .B2(n18422), .ZN(
        n18426) );
  AOI22_X1 U21539 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18424), .B1(
        n18479), .B2(n18477), .ZN(n18425) );
  OAI211_X1 U21540 ( .C1(n18427), .C2(n18484), .A(n18426), .B(n18425), .ZN(
        P3_U2987) );
  INV_X1 U21541 ( .A(n18428), .ZN(n18485) );
  AND2_X1 U21542 ( .A1(n18554), .A2(n18431), .ZN(n18475) );
  AOI22_X1 U21543 ( .A1(n18430), .A2(n18480), .B1(n18429), .B2(n18475), .ZN(
        n18437) );
  AOI22_X1 U21544 ( .A1(n18434), .A2(n18433), .B1(n18432), .B2(n18431), .ZN(
        n18481) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18481), .B1(
        n18435), .B2(n18477), .ZN(n18436) );
  OAI211_X1 U21546 ( .C1(n18485), .C2(n18438), .A(n18437), .B(n18436), .ZN(
        P3_U2988) );
  AOI22_X1 U21547 ( .A1(n18440), .A2(n18477), .B1(n18439), .B2(n18475), .ZN(
        n18443) );
  AOI22_X1 U21548 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18481), .B1(
        n18480), .B2(n18441), .ZN(n18442) );
  OAI211_X1 U21549 ( .C1(n18485), .C2(n18444), .A(n18443), .B(n18442), .ZN(
        P3_U2989) );
  AOI22_X1 U21550 ( .A1(n18446), .A2(n18477), .B1(n18445), .B2(n18475), .ZN(
        n18449) );
  AOI22_X1 U21551 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18481), .B1(
        n18480), .B2(n18447), .ZN(n18448) );
  OAI211_X1 U21552 ( .C1(n18485), .C2(n18450), .A(n18449), .B(n18448), .ZN(
        P3_U2990) );
  AOI22_X1 U21553 ( .A1(n18480), .A2(n18452), .B1(n18451), .B2(n18475), .ZN(
        n18455) );
  AOI22_X1 U21554 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18481), .B1(
        n18453), .B2(n18477), .ZN(n18454) );
  OAI211_X1 U21555 ( .C1(n18485), .C2(n18456), .A(n18455), .B(n18454), .ZN(
        P3_U2991) );
  AOI22_X1 U21556 ( .A1(n18458), .A2(n18477), .B1(n18457), .B2(n18475), .ZN(
        n18461) );
  AOI22_X1 U21557 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18481), .B1(
        n18480), .B2(n18459), .ZN(n18460) );
  OAI211_X1 U21558 ( .C1(n18485), .C2(n18462), .A(n18461), .B(n18460), .ZN(
        P3_U2992) );
  AOI22_X1 U21559 ( .A1(n18480), .A2(n18464), .B1(n18463), .B2(n18475), .ZN(
        n18467) );
  AOI22_X1 U21560 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18481), .B1(
        n18465), .B2(n18477), .ZN(n18466) );
  OAI211_X1 U21561 ( .C1(n18485), .C2(n18468), .A(n18467), .B(n18466), .ZN(
        P3_U2993) );
  AOI22_X1 U21562 ( .A1(n18470), .A2(n18475), .B1(n18469), .B2(n18477), .ZN(
        n18473) );
  AOI22_X1 U21563 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18481), .B1(
        n18480), .B2(n18471), .ZN(n18472) );
  OAI211_X1 U21564 ( .C1(n18485), .C2(n18474), .A(n18473), .B(n18472), .ZN(
        P3_U2994) );
  AOI22_X1 U21565 ( .A1(n18478), .A2(n18477), .B1(n18476), .B2(n18475), .ZN(
        n18483) );
  AOI22_X1 U21566 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18481), .B1(
        n18480), .B2(n18479), .ZN(n18482) );
  OAI211_X1 U21567 ( .C1(n18485), .C2(n18484), .A(n18483), .B(n18482), .ZN(
        P3_U2995) );
  NOR2_X1 U21568 ( .A1(n18497), .A2(n18486), .ZN(n18489) );
  OAI222_X1 U21569 ( .A1(n18492), .A2(n18491), .B1(n18490), .B2(n18489), .C1(
        n18488), .C2(n18487), .ZN(n18696) );
  OAI21_X1 U21570 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(P3_MORE_REG_SCAN_IN), .A(
        n18493), .ZN(n18494) );
  OAI211_X1 U21571 ( .C1(n18523), .C2(n18496), .A(n18495), .B(n18494), .ZN(
        n18544) );
  NOR2_X1 U21572 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18506), .ZN(
        n18527) );
  INV_X1 U21573 ( .A(n18527), .ZN(n18498) );
  NAND2_X1 U21574 ( .A1(n18671), .A2(n18509), .ZN(n18503) );
  AOI22_X1 U21575 ( .A1(n18499), .A2(n18498), .B1(n18497), .B2(n18503), .ZN(
        n18656) );
  NOR2_X1 U21576 ( .A1(n18533), .A2(n18656), .ZN(n18508) );
  AOI21_X1 U21577 ( .B1(n18502), .B2(n18501), .A(n18500), .ZN(n18510) );
  OAI21_X1 U21578 ( .B1(n18504), .B2(n18510), .A(n18503), .ZN(n18505) );
  AOI21_X1 U21579 ( .B1(n18512), .B2(n18506), .A(n18505), .ZN(n18654) );
  NAND2_X1 U21580 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18654), .ZN(
        n18507) );
  OAI22_X1 U21581 ( .A1(n18508), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n18533), .B2(n18507), .ZN(n18542) );
  AND2_X1 U21582 ( .A1(n18509), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n18522) );
  OAI21_X1 U21583 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18511), .A(
        n18510), .ZN(n18521) );
  OAI211_X1 U21584 ( .C1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n18513), .B(n18512), .ZN(
        n18518) );
  NOR2_X1 U21585 ( .A1(n18514), .A2(n18683), .ZN(n18516) );
  OAI211_X1 U21586 ( .C1(n18516), .C2(n18515), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n18671), .ZN(n18517) );
  OAI211_X1 U21587 ( .C1(n18669), .C2(n18519), .A(n18518), .B(n18517), .ZN(
        n18520) );
  AOI21_X1 U21588 ( .B1(n18522), .B2(n18521), .A(n18520), .ZN(n18667) );
  AOI22_X1 U21589 ( .A1(n18533), .A2(n18671), .B1(n18667), .B2(n18523), .ZN(
        n18537) );
  NOR2_X1 U21590 ( .A1(n18525), .A2(n18524), .ZN(n18528) );
  AOI22_X1 U21591 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18526), .B1(
        n18528), .B2(n18683), .ZN(n18679) );
  OAI22_X1 U21592 ( .A1(n18528), .A2(n18672), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18527), .ZN(n18676) );
  AOI222_X1 U21593 ( .A1(n18679), .A2(n18676), .B1(n18679), .B2(n18530), .C1(
        n18676), .C2(n18529), .ZN(n18532) );
  OAI21_X1 U21594 ( .B1(n18533), .B2(n18532), .A(n18531), .ZN(n18536) );
  AND2_X1 U21595 ( .A1(n18537), .A2(n18536), .ZN(n18534) );
  OAI221_X1 U21596 ( .B1(n18537), .B2(n18536), .C1(n18535), .C2(n18534), .A(
        n18539), .ZN(n18541) );
  AOI21_X1 U21597 ( .B1(n18539), .B2(n18538), .A(n18537), .ZN(n18540) );
  AOI222_X1 U21598 ( .A1(n18542), .A2(n18541), .B1(n18542), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18541), .C2(n18540), .ZN(
        n18543) );
  NOR4_X1 U21599 ( .A1(n18545), .A2(n18696), .A3(n18544), .A4(n18543), .ZN(
        n18553) );
  AOI22_X1 U21600 ( .A1(n18703), .A2(n17264), .B1(n18678), .B2(n18708), .ZN(
        n18550) );
  OAI211_X1 U21601 ( .C1(P3_STATE2_REG_1__SCAN_IN), .C2(n18554), .A(
        P3_STATE2_REG_0__SCAN_IN), .B(n18546), .ZN(n18549) );
  OAI211_X1 U21602 ( .C1(n18548), .C2(n18547), .A(n18700), .B(n18553), .ZN(
        n18652) );
  OAI21_X1 U21603 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18697), .A(n18652), 
        .ZN(n18560) );
  OAI22_X1 U21604 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18550), .B1(n18549), 
        .B2(n18560), .ZN(n18551) );
  OAI21_X1 U21605 ( .B1(n18553), .B2(n18552), .A(n18551), .ZN(P3_U2996) );
  NAND2_X1 U21606 ( .A1(n18555), .A2(n18554), .ZN(n18559) );
  AND3_X1 U21607 ( .A1(n18715), .A2(n18703), .A3(n18556), .ZN(n18562) );
  AOI211_X1 U21608 ( .C1(n18703), .C2(n17264), .A(n9662), .B(n18562), .ZN(
        n18558) );
  OAI21_X1 U21609 ( .B1(n18560), .B2(n18559), .A(n18558), .ZN(P3_U2997) );
  OAI21_X1 U21610 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18561), .ZN(n18563) );
  AOI21_X1 U21611 ( .B1(n18564), .B2(n18563), .A(n18562), .ZN(P3_U2998) );
  INV_X1 U21612 ( .A(n18650), .ZN(n18565) );
  AND2_X1 U21613 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18565), .ZN(
        P3_U2999) );
  AND2_X1 U21614 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18565), .ZN(
        P3_U3000) );
  AND2_X1 U21615 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18565), .ZN(
        P3_U3001) );
  AND2_X1 U21616 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18565), .ZN(
        P3_U3002) );
  AND2_X1 U21617 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18565), .ZN(
        P3_U3003) );
  AND2_X1 U21618 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18565), .ZN(
        P3_U3004) );
  AND2_X1 U21619 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18565), .ZN(
        P3_U3005) );
  AND2_X1 U21620 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18565), .ZN(
        P3_U3006) );
  AND2_X1 U21621 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18565), .ZN(
        P3_U3007) );
  AND2_X1 U21622 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18565), .ZN(
        P3_U3008) );
  AND2_X1 U21623 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18565), .ZN(
        P3_U3009) );
  AND2_X1 U21624 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18565), .ZN(
        P3_U3010) );
  AND2_X1 U21625 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18565), .ZN(
        P3_U3011) );
  AND2_X1 U21626 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18565), .ZN(
        P3_U3012) );
  AND2_X1 U21627 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18565), .ZN(
        P3_U3013) );
  INV_X1 U21628 ( .A(P3_DATAWIDTH_REG_16__SCAN_IN), .ZN(n20872) );
  NOR2_X1 U21629 ( .A1(n20872), .A2(n18650), .ZN(P3_U3014) );
  AND2_X1 U21630 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18565), .ZN(
        P3_U3015) );
  AND2_X1 U21631 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18565), .ZN(
        P3_U3016) );
  AND2_X1 U21632 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18565), .ZN(
        P3_U3017) );
  AND2_X1 U21633 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18565), .ZN(
        P3_U3018) );
  AND2_X1 U21634 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18565), .ZN(
        P3_U3019) );
  AND2_X1 U21635 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18565), .ZN(
        P3_U3020) );
  AND2_X1 U21636 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18565), .ZN(P3_U3021) );
  AND2_X1 U21637 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18565), .ZN(P3_U3022) );
  AND2_X1 U21638 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18565), .ZN(P3_U3023) );
  AND2_X1 U21639 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18565), .ZN(P3_U3024) );
  AND2_X1 U21640 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18565), .ZN(P3_U3025) );
  AND2_X1 U21641 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18565), .ZN(P3_U3026) );
  AND2_X1 U21642 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18565), .ZN(P3_U3027) );
  AND2_X1 U21643 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18565), .ZN(P3_U3028) );
  OAI21_X1 U21644 ( .B1(n18566), .B2(n19687), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18567) );
  AOI22_X1 U21645 ( .A1(n18578), .A2(n18580), .B1(n18713), .B2(n18567), .ZN(
        n18568) );
  INV_X1 U21646 ( .A(NA), .ZN(n20697) );
  OR3_X1 U21647 ( .A1(n20697), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n18573) );
  OAI211_X1 U21648 ( .C1(n18697), .C2(n18569), .A(n18568), .B(n18573), .ZN(
        P3_U3029) );
  INV_X1 U21649 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18710) );
  NOR2_X1 U21650 ( .A1(n18580), .A2(n19687), .ZN(n18576) );
  OAI22_X1 U21651 ( .A1(n18710), .A2(n18576), .B1(n19687), .B2(n18569), .ZN(
        n18570) );
  INV_X1 U21652 ( .A(n18570), .ZN(n18572) );
  NAND2_X1 U21653 ( .A1(n18703), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18574) );
  OAI211_X1 U21654 ( .C1(n18572), .C2(n18578), .A(n18574), .B(n18571), .ZN(
        P3_U3030) );
  AOI22_X1 U21655 ( .A1(n18703), .A2(P3_STATE_REG_1__SCAN_IN), .B1(n18578), 
        .B2(n18573), .ZN(n18579) );
  OAI22_X1 U21656 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18574), .ZN(n18575) );
  OAI22_X1 U21657 ( .A1(n18576), .A2(n18575), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18577) );
  OAI22_X1 U21658 ( .A1(n18579), .A2(n18580), .B1(n18578), .B2(n18577), .ZN(
        P3_U3031) );
  OAI222_X1 U21659 ( .A1(n18685), .A2(n9583), .B1(n18581), .B2(n18712), .C1(
        n18582), .C2(n18639), .ZN(P3_U3032) );
  OAI222_X1 U21660 ( .A1(n18639), .A2(n18584), .B1(n18583), .B2(n18712), .C1(
        n18582), .C2(n9583), .ZN(P3_U3033) );
  OAI222_X1 U21661 ( .A1(n18639), .A2(n18587), .B1(n18585), .B2(n18712), .C1(
        n18584), .C2(n9583), .ZN(P3_U3034) );
  INV_X1 U21662 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18590) );
  OAI222_X1 U21663 ( .A1(n18639), .A2(n18590), .B1(n18588), .B2(n18712), .C1(
        n18587), .C2(n9583), .ZN(P3_U3035) );
  OAI222_X1 U21664 ( .A1(n18590), .A2(n9583), .B1(n18589), .B2(n18712), .C1(
        n18591), .C2(n18639), .ZN(P3_U3036) );
  OAI222_X1 U21665 ( .A1(n18639), .A2(n18593), .B1(n18592), .B2(n18712), .C1(
        n18591), .C2(n9583), .ZN(P3_U3037) );
  OAI222_X1 U21666 ( .A1(n18639), .A2(n18595), .B1(n18594), .B2(n18712), .C1(
        n18593), .C2(n9583), .ZN(P3_U3038) );
  OAI222_X1 U21667 ( .A1(n18639), .A2(n18598), .B1(n18596), .B2(n18712), .C1(
        n18595), .C2(n9583), .ZN(P3_U3039) );
  OAI222_X1 U21668 ( .A1(n18598), .A2(n9583), .B1(n18597), .B2(n18712), .C1(
        n18599), .C2(n18639), .ZN(P3_U3040) );
  OAI222_X1 U21669 ( .A1(n18639), .A2(n18601), .B1(n18600), .B2(n18712), .C1(
        n18599), .C2(n9583), .ZN(P3_U3041) );
  OAI222_X1 U21670 ( .A1(n18639), .A2(n18603), .B1(n18602), .B2(n18712), .C1(
        n18601), .C2(n9583), .ZN(P3_U3042) );
  OAI222_X1 U21671 ( .A1(n18639), .A2(n18605), .B1(n18604), .B2(n18712), .C1(
        n18603), .C2(n9583), .ZN(P3_U3043) );
  OAI222_X1 U21672 ( .A1(n18639), .A2(n18608), .B1(n18606), .B2(n18712), .C1(
        n18605), .C2(n9583), .ZN(P3_U3044) );
  OAI222_X1 U21673 ( .A1(n18608), .A2(n9583), .B1(n18607), .B2(n18712), .C1(
        n18609), .C2(n18639), .ZN(P3_U3045) );
  OAI222_X1 U21674 ( .A1(n18639), .A2(n18611), .B1(n18610), .B2(n18712), .C1(
        n18609), .C2(n9583), .ZN(P3_U3046) );
  OAI222_X1 U21675 ( .A1(n18639), .A2(n18614), .B1(n18612), .B2(n18712), .C1(
        n18611), .C2(n9583), .ZN(P3_U3047) );
  OAI222_X1 U21676 ( .A1(n18614), .A2(n9583), .B1(n18613), .B2(n18712), .C1(
        n18615), .C2(n18639), .ZN(P3_U3048) );
  OAI222_X1 U21677 ( .A1(n18639), .A2(n18618), .B1(n18616), .B2(n18712), .C1(
        n18615), .C2(n9583), .ZN(P3_U3049) );
  OAI222_X1 U21678 ( .A1(n18618), .A2(n9583), .B1(n18617), .B2(n18712), .C1(
        n18619), .C2(n18639), .ZN(P3_U3050) );
  OAI222_X1 U21679 ( .A1(n18639), .A2(n18622), .B1(n18620), .B2(n18712), .C1(
        n18619), .C2(n9583), .ZN(P3_U3051) );
  OAI222_X1 U21680 ( .A1(n18622), .A2(n9583), .B1(n18621), .B2(n18712), .C1(
        n18623), .C2(n18639), .ZN(P3_U3052) );
  OAI222_X1 U21681 ( .A1(n18639), .A2(n18626), .B1(n18624), .B2(n18712), .C1(
        n18623), .C2(n9583), .ZN(P3_U3053) );
  OAI222_X1 U21682 ( .A1(n18626), .A2(n9583), .B1(n18625), .B2(n18712), .C1(
        n18627), .C2(n18639), .ZN(P3_U3054) );
  INV_X1 U21683 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18629) );
  OAI222_X1 U21684 ( .A1(n18639), .A2(n18629), .B1(n18628), .B2(n18712), .C1(
        n18627), .C2(n9583), .ZN(P3_U3055) );
  INV_X1 U21685 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18631) );
  OAI222_X1 U21686 ( .A1(n18639), .A2(n18631), .B1(n18630), .B2(n18712), .C1(
        n18629), .C2(n9583), .ZN(P3_U3056) );
  OAI222_X1 U21687 ( .A1(n18639), .A2(n18633), .B1(n18632), .B2(n18712), .C1(
        n18631), .C2(n9583), .ZN(P3_U3057) );
  OAI222_X1 U21688 ( .A1(n18639), .A2(n18636), .B1(n18634), .B2(n18712), .C1(
        n18633), .C2(n9583), .ZN(P3_U3058) );
  OAI222_X1 U21689 ( .A1(n18636), .A2(n9583), .B1(n18635), .B2(n18712), .C1(
        n18637), .C2(n18639), .ZN(P3_U3059) );
  OAI222_X1 U21690 ( .A1(n18639), .A2(n18642), .B1(n18638), .B2(n18712), .C1(
        n18637), .C2(n9583), .ZN(P3_U3060) );
  INV_X1 U21691 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18640) );
  OAI222_X1 U21692 ( .A1(n9583), .A2(n18642), .B1(n18641), .B2(n18712), .C1(
        n18640), .C2(n18639), .ZN(P3_U3061) );
  OAI22_X1 U21693 ( .A1(n18713), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18712), .ZN(n18643) );
  INV_X1 U21694 ( .A(n18643), .ZN(P3_U3274) );
  OAI22_X1 U21695 ( .A1(n18713), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18712), .ZN(n18644) );
  INV_X1 U21696 ( .A(n18644), .ZN(P3_U3275) );
  OAI22_X1 U21697 ( .A1(n18713), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18712), .ZN(n18645) );
  INV_X1 U21698 ( .A(n18645), .ZN(P3_U3276) );
  OAI22_X1 U21699 ( .A1(n18713), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18712), .ZN(n18646) );
  INV_X1 U21700 ( .A(n18646), .ZN(P3_U3277) );
  OAI21_X1 U21701 ( .B1(n18650), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18648), 
        .ZN(n18647) );
  INV_X1 U21702 ( .A(n18647), .ZN(P3_U3280) );
  OAI21_X1 U21703 ( .B1(n18650), .B2(n18649), .A(n18648), .ZN(P3_U3281) );
  OAI221_X1 U21704 ( .B1(n18653), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18653), 
        .C2(n18652), .A(n18651), .ZN(P3_U3282) );
  NOR2_X1 U21705 ( .A1(n18654), .A2(n18666), .ZN(n18655) );
  NOR2_X1 U21706 ( .A1(n18655), .A2(n18684), .ZN(n18660) );
  NOR3_X1 U21707 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18656), .A3(
        n18666), .ZN(n18657) );
  AOI21_X1 U21708 ( .B1(n18678), .B2(n18658), .A(n18657), .ZN(n18659) );
  OAI22_X1 U21709 ( .A1(n18661), .A2(n18660), .B1(n18684), .B2(n18659), .ZN(
        P3_U3285) );
  AOI22_X1 U21710 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n18663), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18662), .ZN(n18674) );
  NOR2_X1 U21711 ( .A1(n18664), .A2(n18680), .ZN(n18673) );
  INV_X1 U21712 ( .A(n18673), .ZN(n18665) );
  OAI22_X1 U21713 ( .A1(n18667), .A2(n18666), .B1(n18674), .B2(n18665), .ZN(
        n18668) );
  AOI21_X1 U21714 ( .B1(n18678), .B2(n18669), .A(n18668), .ZN(n18670) );
  INV_X1 U21715 ( .A(n18684), .ZN(n18681) );
  AOI22_X1 U21716 ( .A1(n18684), .A2(n18671), .B1(n18670), .B2(n18681), .ZN(
        P3_U3288) );
  INV_X1 U21717 ( .A(n18672), .ZN(n18675) );
  AOI222_X1 U21718 ( .A1(n18676), .A2(n18716), .B1(n18678), .B2(n18675), .C1(
        n18674), .C2(n18673), .ZN(n18677) );
  AOI22_X1 U21719 ( .A1(n18684), .A2(n10687), .B1(n18677), .B2(n18681), .ZN(
        P3_U3289) );
  AOI222_X1 U21720 ( .A1(n18680), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18716), 
        .B2(n18679), .C1(n18683), .C2(n18678), .ZN(n18682) );
  AOI22_X1 U21721 ( .A1(n18684), .A2(n18683), .B1(n18682), .B2(n18681), .ZN(
        P3_U3290) );
  AOI21_X1 U21722 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18686) );
  AOI22_X1 U21723 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18686), .B2(n18685), .ZN(n18688) );
  INV_X1 U21724 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18687) );
  AOI22_X1 U21725 ( .A1(n18689), .A2(n18688), .B1(n18687), .B2(n18692), .ZN(
        P3_U3292) );
  INV_X1 U21726 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18693) );
  NOR2_X1 U21727 ( .A1(n18692), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18690) );
  AOI22_X1 U21728 ( .A1(n18693), .A2(n18692), .B1(n18691), .B2(n18690), .ZN(
        P3_U3293) );
  INV_X1 U21729 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18719) );
  OAI22_X1 U21730 ( .A1(n18713), .A2(n18719), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n18712), .ZN(n18694) );
  INV_X1 U21731 ( .A(n18694), .ZN(P3_U3294) );
  MUX2_X1 U21732 ( .A(P3_MORE_REG_SCAN_IN), .B(n18696), .S(n18695), .Z(
        P3_U3295) );
  AOI21_X1 U21733 ( .B1(n17264), .B2(n18697), .A(n18718), .ZN(n18698) );
  OAI21_X1 U21734 ( .B1(n18700), .B2(n18699), .A(n18698), .ZN(n18711) );
  OAI21_X1 U21735 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n18702), .A(n18701), 
        .ZN(n18704) );
  AOI211_X1 U21736 ( .C1(n18717), .C2(n18704), .A(n18703), .B(n18715), .ZN(
        n18706) );
  NOR2_X1 U21737 ( .A1(n18706), .A2(n18705), .ZN(n18707) );
  OAI21_X1 U21738 ( .B1(n18708), .B2(n18707), .A(n18711), .ZN(n18709) );
  OAI21_X1 U21739 ( .B1(n18711), .B2(n18710), .A(n18709), .ZN(P3_U3296) );
  OAI22_X1 U21740 ( .A1(n18713), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18712), .ZN(n18714) );
  INV_X1 U21741 ( .A(n18714), .ZN(P3_U3297) );
  AOI21_X1 U21742 ( .B1(n18716), .B2(n18715), .A(n18718), .ZN(n18722) );
  AOI22_X1 U21743 ( .A1(n18722), .A2(n18719), .B1(n18718), .B2(n18717), .ZN(
        P3_U3298) );
  INV_X1 U21744 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18721) );
  AOI21_X1 U21745 ( .B1(n18722), .B2(n18721), .A(n18720), .ZN(P3_U3299) );
  INV_X1 U21746 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n18728) );
  NAND2_X1 U21747 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19698), .ZN(n19686) );
  NAND2_X1 U21748 ( .A1(n18728), .A2(n18723), .ZN(n19683) );
  OAI21_X1 U21749 ( .B1(n18728), .B2(n19686), .A(n19683), .ZN(n19756) );
  AOI21_X1 U21750 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19756), .ZN(n18724) );
  INV_X1 U21751 ( .A(n18724), .ZN(P2_U2815) );
  INV_X1 U21752 ( .A(n18725), .ZN(n18726) );
  INV_X1 U21753 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18727) );
  OAI22_X1 U21754 ( .A1(n18726), .A2(n18727), .B1(n19666), .B2(n19670), .ZN(
        P2_U2816) );
  AOI21_X1 U21755 ( .B1(P2_STATE_REG_1__SCAN_IN), .B2(n18727), .A(n19691), 
        .ZN(n18730) );
  NAND2_X1 U21756 ( .A1(n18728), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19810) );
  INV_X1 U21757 ( .A(P2_D_C_N_REG_SCAN_IN), .ZN(n18729) );
  OAI22_X1 U21758 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n18730), .B1(n19744), 
        .B2(n18729), .ZN(P2_U2817) );
  OAI21_X1 U21759 ( .B1(n19691), .B2(BS16), .A(n19756), .ZN(n19754) );
  OAI21_X1 U21760 ( .B1(n19756), .B2(n19544), .A(n19754), .ZN(P2_U2818) );
  NOR4_X1 U21761 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18734) );
  NOR4_X1 U21762 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18733) );
  NOR4_X1 U21763 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18732) );
  NOR4_X1 U21764 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18731) );
  NAND4_X1 U21765 ( .A1(n18734), .A2(n18733), .A3(n18732), .A4(n18731), .ZN(
        n18740) );
  NOR4_X1 U21766 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18738) );
  AOI211_X1 U21767 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_14__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18737) );
  NOR4_X1 U21768 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n18736) );
  NOR4_X1 U21769 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18735) );
  NAND4_X1 U21770 ( .A1(n18738), .A2(n18737), .A3(n18736), .A4(n18735), .ZN(
        n18739) );
  NOR2_X1 U21771 ( .A1(n18740), .A2(n18739), .ZN(n18749) );
  INV_X1 U21772 ( .A(n18749), .ZN(n18748) );
  NOR2_X1 U21773 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18748), .ZN(n18743) );
  INV_X1 U21774 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18741) );
  AOI22_X1 U21775 ( .A1(n18743), .A2(n18865), .B1(n18748), .B2(n18741), .ZN(
        P2_U2820) );
  OR3_X1 U21776 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18747) );
  INV_X1 U21777 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18742) );
  AOI22_X1 U21778 ( .A1(n18743), .A2(n18747), .B1(n18748), .B2(n18742), .ZN(
        P2_U2821) );
  INV_X1 U21779 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19755) );
  NAND2_X1 U21780 ( .A1(n18743), .A2(n19755), .ZN(n18746) );
  OAI21_X1 U21781 ( .B1(n19699), .B2(n18865), .A(n18749), .ZN(n18744) );
  OAI21_X1 U21782 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18749), .A(n18744), 
        .ZN(n18745) );
  OAI221_X1 U21783 ( .B1(n18746), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18746), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18745), .ZN(P2_U2822) );
  INV_X1 U21784 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19750) );
  OAI221_X1 U21785 ( .B1(n18749), .B2(n19750), .C1(n18748), .C2(n18747), .A(
        n18746), .ZN(P2_U2823) );
  NOR2_X1 U21786 ( .A1(n18849), .A2(n18750), .ZN(n18751) );
  XOR2_X1 U21787 ( .A(n18752), .B(n18751), .Z(n18762) );
  AOI22_X1 U21788 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18879), .B1(
        P2_REIP_REG_19__SCAN_IN), .B2(n18853), .ZN(n18753) );
  OAI211_X1 U21789 ( .C1(n18864), .C2(n18754), .A(n18753), .B(n18765), .ZN(
        n18755) );
  AOI21_X1 U21790 ( .B1(n18756), .B2(n18786), .A(n18755), .ZN(n18761) );
  OAI22_X1 U21791 ( .A1(n18758), .A2(n18856), .B1(n18757), .B2(n18858), .ZN(
        n18759) );
  INV_X1 U21792 ( .A(n18759), .ZN(n18760) );
  OAI211_X1 U21793 ( .C1(n18863), .C2(n18762), .A(n18761), .B(n18760), .ZN(
        P2_U2836) );
  NAND2_X1 U21794 ( .A1(n9567), .A2(n18777), .ZN(n18763) );
  XOR2_X1 U21795 ( .A(n18764), .B(n18763), .Z(n18776) );
  AOI22_X1 U21796 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18879), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n18853), .ZN(n18766) );
  OAI211_X1 U21797 ( .C1(n18864), .C2(n18767), .A(n18766), .B(n18765), .ZN(
        n18768) );
  AOI21_X1 U21798 ( .B1(n18769), .B2(n18786), .A(n18768), .ZN(n18775) );
  INV_X1 U21799 ( .A(n18770), .ZN(n18771) );
  OAI22_X1 U21800 ( .A1(n18772), .A2(n18856), .B1(n18771), .B2(n18858), .ZN(
        n18773) );
  INV_X1 U21801 ( .A(n18773), .ZN(n18774) );
  OAI211_X1 U21802 ( .C1(n18863), .C2(n18776), .A(n18775), .B(n18774), .ZN(
        P2_U2837) );
  OAI21_X1 U21803 ( .B1(n18778), .B2(n18796), .A(n18777), .ZN(n18789) );
  NAND2_X1 U21804 ( .A1(n18779), .A2(n18874), .ZN(n18784) );
  NAND2_X1 U21805 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n18879), .ZN(
        n18780) );
  OAI211_X1 U21806 ( .C1(n18864), .C2(n18781), .A(n18765), .B(n18780), .ZN(
        n18782) );
  AOI21_X1 U21807 ( .B1(n18853), .B2(P2_REIP_REG_17__SCAN_IN), .A(n18782), 
        .ZN(n18783) );
  NAND2_X1 U21808 ( .A1(n18784), .A2(n18783), .ZN(n18785) );
  AOI21_X1 U21809 ( .B1(n18787), .B2(n18786), .A(n18785), .ZN(n18788) );
  OAI21_X1 U21810 ( .B1(n18790), .B2(n18789), .A(n18788), .ZN(n18791) );
  INV_X1 U21811 ( .A(n18791), .ZN(n18795) );
  INV_X1 U21812 ( .A(n18792), .ZN(n18793) );
  NAND2_X1 U21813 ( .A1(n18869), .A2(n18793), .ZN(n18794) );
  OAI211_X1 U21814 ( .C1(n18835), .C2(n18796), .A(n18795), .B(n18794), .ZN(
        P2_U2838) );
  NOR2_X1 U21815 ( .A1(n18849), .A2(n18797), .ZN(n18799) );
  XOR2_X1 U21816 ( .A(n18799), .B(n18798), .Z(n18807) );
  OAI21_X1 U21817 ( .B1(n18864), .B2(n10632), .A(n18765), .ZN(n18800) );
  AOI21_X1 U21818 ( .B1(n18853), .B2(P2_REIP_REG_15__SCAN_IN), .A(n18800), 
        .ZN(n18801) );
  OAI21_X1 U21819 ( .B1(n18802), .B2(n18871), .A(n18801), .ZN(n18805) );
  OAI22_X1 U21820 ( .A1(n18803), .A2(n18856), .B1(n18937), .B2(n18858), .ZN(
        n18804) );
  AOI211_X1 U21821 ( .C1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n18879), .A(
        n18805), .B(n18804), .ZN(n18806) );
  OAI21_X1 U21822 ( .B1(n18863), .B2(n18807), .A(n18806), .ZN(P2_U2840) );
  INV_X1 U21823 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n20892) );
  OAI21_X1 U21824 ( .B1(n18864), .B2(n18808), .A(n18765), .ZN(n18811) );
  NOR2_X1 U21825 ( .A1(n18809), .A2(n18871), .ZN(n18810) );
  AOI211_X1 U21826 ( .C1(n18853), .C2(P2_REIP_REG_12__SCAN_IN), .A(n18811), 
        .B(n18810), .ZN(n18817) );
  NAND2_X1 U21827 ( .A1(n9567), .A2(n18829), .ZN(n18812) );
  XOR2_X1 U21828 ( .A(n18813), .B(n18812), .Z(n18815) );
  OAI22_X1 U21829 ( .A1(n18944), .A2(n18858), .B1(n18902), .B2(n18856), .ZN(
        n18814) );
  AOI21_X1 U21830 ( .B1(n19673), .B2(n18815), .A(n18814), .ZN(n18816) );
  OAI211_X1 U21831 ( .C1(n20892), .C2(n18821), .A(n18817), .B(n18816), .ZN(
        P2_U2843) );
  INV_X1 U21832 ( .A(n18946), .ZN(n18828) );
  NAND2_X1 U21833 ( .A1(n18818), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n18819) );
  OAI211_X1 U21834 ( .C1(n18821), .C2(n18820), .A(n18819), .B(n18765), .ZN(
        n18824) );
  NOR2_X1 U21835 ( .A1(n18822), .A2(n18856), .ZN(n18823) );
  AOI211_X1 U21836 ( .C1(n18853), .C2(P2_REIP_REG_11__SCAN_IN), .A(n18824), 
        .B(n18823), .ZN(n18825) );
  OAI21_X1 U21837 ( .B1(n18826), .B2(n18871), .A(n18825), .ZN(n18827) );
  AOI21_X1 U21838 ( .B1(n18828), .B2(n18869), .A(n18827), .ZN(n18833) );
  OAI211_X1 U21839 ( .C1(n18831), .C2(n18834), .A(n18830), .B(n18829), .ZN(
        n18832) );
  OAI211_X1 U21840 ( .C1(n18835), .C2(n18834), .A(n18833), .B(n18832), .ZN(
        P2_U2844) );
  NOR2_X1 U21841 ( .A1(n18849), .A2(n18836), .ZN(n18838) );
  XOR2_X1 U21842 ( .A(n18838), .B(n18837), .Z(n18847) );
  INV_X1 U21843 ( .A(n18839), .ZN(n18842) );
  OAI21_X1 U21844 ( .B1(n18864), .B2(n10611), .A(n18765), .ZN(n18840) );
  AOI21_X1 U21845 ( .B1(n18853), .B2(P2_REIP_REG_9__SCAN_IN), .A(n18840), .ZN(
        n18841) );
  OAI21_X1 U21846 ( .B1(n18842), .B2(n18871), .A(n18841), .ZN(n18845) );
  OAI22_X1 U21847 ( .A1(n18843), .A2(n18856), .B1(n18951), .B2(n18858), .ZN(
        n18844) );
  AOI211_X1 U21848 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n18879), .A(
        n18845), .B(n18844), .ZN(n18846) );
  OAI21_X1 U21849 ( .B1(n18863), .B2(n18847), .A(n18846), .ZN(P2_U2846) );
  NOR2_X1 U21850 ( .A1(n18849), .A2(n18848), .ZN(n18850) );
  XOR2_X1 U21851 ( .A(n18851), .B(n18850), .Z(n18862) );
  OAI21_X1 U21852 ( .B1(n18864), .B2(n10602), .A(n18765), .ZN(n18852) );
  AOI21_X1 U21853 ( .B1(n18853), .B2(P2_REIP_REG_7__SCAN_IN), .A(n18852), .ZN(
        n18854) );
  OAI21_X1 U21854 ( .B1(n18855), .B2(n18871), .A(n18854), .ZN(n18860) );
  OAI22_X1 U21855 ( .A1(n18955), .A2(n18858), .B1(n18857), .B2(n18856), .ZN(
        n18859) );
  AOI211_X1 U21856 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n18879), .A(
        n18860), .B(n18859), .ZN(n18861) );
  OAI21_X1 U21857 ( .B1(n18863), .B2(n18862), .A(n18861), .ZN(P2_U2848) );
  OAI22_X1 U21858 ( .A1(n18866), .A2(n18865), .B1(n11161), .B2(n18864), .ZN(
        n18867) );
  AOI21_X1 U21859 ( .B1(n18869), .B2(n18868), .A(n18867), .ZN(n18870) );
  OAI21_X1 U21860 ( .B1(n18872), .B2(n18871), .A(n18870), .ZN(n18873) );
  AOI21_X1 U21861 ( .B1(n18875), .B2(n18874), .A(n18873), .ZN(n18882) );
  AOI22_X1 U21862 ( .A1(n18877), .A2(n19673), .B1(n19334), .B2(n18876), .ZN(
        n18881) );
  OAI21_X1 U21863 ( .B1(n18879), .B2(n18878), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18880) );
  NAND3_X1 U21864 ( .A1(n18882), .A2(n18881), .A3(n18880), .ZN(P2_U2855) );
  AND2_X1 U21865 ( .A1(n18884), .A2(n18883), .ZN(n18885) );
  OR2_X1 U21866 ( .A1(n18885), .A2(n13895), .ZN(n18930) );
  OAI22_X1 U21867 ( .A1(n18930), .A2(n18919), .B1(n20956), .B2(n18886), .ZN(
        n18887) );
  INV_X1 U21868 ( .A(n18887), .ZN(n18888) );
  OAI21_X1 U21869 ( .B1(n20964), .B2(n18889), .A(n18888), .ZN(P2_U2871) );
  XNOR2_X1 U21870 ( .A(n14077), .B(n18890), .ZN(n18892) );
  AOI22_X1 U21871 ( .A1(n18892), .A2(n18891), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n20964), .ZN(n18893) );
  OAI21_X1 U21872 ( .B1(n18894), .B2(n20964), .A(n18893), .ZN(P2_U2873) );
  AND2_X1 U21873 ( .A1(n13410), .A2(n18895), .ZN(n20958) );
  AOI21_X1 U21874 ( .B1(n18903), .B2(n18897), .A(n18896), .ZN(n18898) );
  OR3_X1 U21875 ( .A1(n20958), .A2(n18898), .A3(n18919), .ZN(n18900) );
  NAND2_X1 U21876 ( .A1(n20964), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n18899) );
  AND2_X1 U21877 ( .A1(n18900), .A2(n18899), .ZN(n18901) );
  OAI21_X1 U21878 ( .B1(n18902), .B2(n20964), .A(n18901), .ZN(P2_U2875) );
  AOI211_X1 U21879 ( .C1(n18905), .C2(n18904), .A(n18919), .B(n18903), .ZN(
        n18906) );
  AOI21_X1 U21880 ( .B1(n18907), .B2(n20956), .A(n18906), .ZN(n18908) );
  OAI21_X1 U21881 ( .B1(n20956), .B2(n10614), .A(n18908), .ZN(P2_U2877) );
  AND2_X1 U21882 ( .A1(n13410), .A2(n18909), .ZN(n18911) );
  NAND2_X1 U21883 ( .A1(n18911), .A2(n18910), .ZN(n18913) );
  AOI211_X1 U21884 ( .C1(n18914), .C2(n18913), .A(n18919), .B(n18912), .ZN(
        n18915) );
  AOI21_X1 U21885 ( .B1(P2_EBX_REG_8__SCAN_IN), .B2(n20964), .A(n18915), .ZN(
        n18916) );
  OAI21_X1 U21886 ( .B1(n18917), .B2(n20964), .A(n18916), .ZN(P2_U2879) );
  OAI22_X1 U21887 ( .A1(n18969), .A2(n18919), .B1(n20964), .B2(n18918), .ZN(
        n18920) );
  INV_X1 U21888 ( .A(n18920), .ZN(n18921) );
  OAI21_X1 U21889 ( .B1(n20956), .B2(n18922), .A(n18921), .ZN(P2_U2883) );
  AOI22_X1 U21890 ( .A1(n15811), .A2(n18982), .B1(n18927), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n18924) );
  AOI22_X1 U21891 ( .A1(n18928), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n18981), .ZN(n18923) );
  NAND2_X1 U21892 ( .A1(n18924), .A2(n18923), .ZN(P2_U2888) );
  AOI22_X1 U21893 ( .A1(n18926), .A2(n18925), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n18981), .ZN(n18934) );
  AOI22_X1 U21894 ( .A1(n18928), .A2(BUF1_REG_16__SCAN_IN), .B1(n18927), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n18933) );
  OAI22_X1 U21895 ( .A1(n18930), .A2(n18986), .B1(n18935), .B2(n18929), .ZN(
        n18931) );
  INV_X1 U21896 ( .A(n18931), .ZN(n18932) );
  NAND3_X1 U21897 ( .A1(n18934), .A2(n18933), .A3(n18932), .ZN(P2_U2903) );
  OAI222_X1 U21898 ( .A1(n18937), .A2(n18966), .B1(n13156), .B2(n18956), .C1(
        n18936), .C2(n18990), .ZN(P2_U2904) );
  INV_X1 U21899 ( .A(n18938), .ZN(n18940) );
  AOI22_X1 U21900 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n18981), .B1(n19030), 
        .B2(n18958), .ZN(n18939) );
  OAI21_X1 U21901 ( .B1(n18966), .B2(n18940), .A(n18939), .ZN(P2_U2905) );
  INV_X1 U21902 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19000) );
  OAI222_X1 U21903 ( .A1(n18942), .A2(n18966), .B1(n19000), .B2(n18956), .C1(
        n18990), .C2(n18941), .ZN(P2_U2906) );
  INV_X1 U21904 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19002) );
  OAI222_X1 U21905 ( .A1(n18944), .A2(n18966), .B1(n19002), .B2(n18956), .C1(
        n18990), .C2(n18943), .ZN(P2_U2907) );
  INV_X1 U21906 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19004) );
  OAI222_X1 U21907 ( .A1(n18946), .A2(n18966), .B1(n19004), .B2(n18956), .C1(
        n18990), .C2(n18945), .ZN(P2_U2908) );
  AOI22_X1 U21908 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n18981), .B1(n18947), 
        .B2(n18958), .ZN(n18948) );
  OAI21_X1 U21909 ( .B1(n18966), .B2(n18949), .A(n18948), .ZN(P2_U2909) );
  INV_X1 U21910 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19008) );
  OAI222_X1 U21911 ( .A1(n18951), .A2(n18966), .B1(n19008), .B2(n18956), .C1(
        n18990), .C2(n18950), .ZN(P2_U2910) );
  INV_X1 U21912 ( .A(n18952), .ZN(n18954) );
  INV_X1 U21913 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19010) );
  OAI222_X1 U21914 ( .A1(n18954), .A2(n18966), .B1(n19010), .B2(n18956), .C1(
        n18990), .C2(n18953), .ZN(P2_U2911) );
  OAI222_X1 U21915 ( .A1(n18955), .A2(n18966), .B1(n19012), .B2(n18956), .C1(
        n18990), .C2(n19088), .ZN(P2_U2912) );
  INV_X1 U21916 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19014) );
  OAI222_X1 U21917 ( .A1(n18957), .A2(n18966), .B1(n19014), .B2(n18956), .C1(
        n18990), .C2(n19077), .ZN(P2_U2913) );
  AOI22_X1 U21918 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n18981), .B1(n18959), .B2(
        n18958), .ZN(n18964) );
  AOI21_X1 U21919 ( .B1(n19772), .B2(n19770), .A(n18960), .ZN(n18977) );
  XNOR2_X1 U21920 ( .A(n19761), .B(n18961), .ZN(n18976) );
  NOR2_X1 U21921 ( .A1(n18977), .A2(n18976), .ZN(n18975) );
  AOI21_X1 U21922 ( .B1(n18961), .B2(n19761), .A(n18975), .ZN(n18962) );
  NOR2_X1 U21923 ( .A1(n18962), .A2(n18967), .ZN(n18968) );
  OR3_X1 U21924 ( .A1(n18968), .A2(n18969), .A3(n18986), .ZN(n18963) );
  OAI211_X1 U21925 ( .C1(n18966), .C2(n18965), .A(n18964), .B(n18963), .ZN(
        P2_U2914) );
  AOI22_X1 U21926 ( .A1(n18982), .A2(n18967), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n18981), .ZN(n18973) );
  XOR2_X1 U21927 ( .A(n18969), .B(n18968), .Z(n18971) );
  NAND2_X1 U21928 ( .A1(n18971), .A2(n18970), .ZN(n18972) );
  OAI211_X1 U21929 ( .C1(n18974), .C2(n18990), .A(n18973), .B(n18972), .ZN(
        P2_U2915) );
  AOI22_X1 U21930 ( .A1(n19767), .A2(n18982), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n18981), .ZN(n18980) );
  AOI21_X1 U21931 ( .B1(n18977), .B2(n18976), .A(n18975), .ZN(n18978) );
  OR2_X1 U21932 ( .A1(n18978), .A2(n18986), .ZN(n18979) );
  OAI211_X1 U21933 ( .C1(n19066), .C2(n18990), .A(n18980), .B(n18979), .ZN(
        P2_U2916) );
  AOI22_X1 U21934 ( .A1(n19786), .A2(n18982), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n18981), .ZN(n18989) );
  AOI21_X1 U21935 ( .B1(n18985), .B2(n18984), .A(n18983), .ZN(n18987) );
  OR2_X1 U21936 ( .A1(n18987), .A2(n18986), .ZN(n18988) );
  OAI211_X1 U21937 ( .C1(n19056), .C2(n18990), .A(n18989), .B(n18988), .ZN(
        P2_U2918) );
  NOR2_X1 U21938 ( .A1(n18995), .A2(n18991), .ZN(P2_U2920) );
  INV_X1 U21939 ( .A(n18992), .ZN(n18993) );
  AOI22_X1 U21940 ( .A1(n18993), .A2(P2_EAX_REG_30__SCAN_IN), .B1(
        P2_UWORD_REG_14__SCAN_IN), .B2(n19026), .ZN(n18994) );
  OAI21_X1 U21941 ( .B1(n20866), .B2(n18995), .A(n18994), .ZN(P2_U2921) );
  AOI22_X1 U21942 ( .A1(n19026), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n18996) );
  OAI21_X1 U21943 ( .B1(n13156), .B2(n19028), .A(n18996), .ZN(P2_U2936) );
  INV_X1 U21944 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n18998) );
  AOI22_X1 U21945 ( .A1(n19026), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n18997) );
  OAI21_X1 U21946 ( .B1(n18998), .B2(n19028), .A(n18997), .ZN(P2_U2937) );
  AOI22_X1 U21947 ( .A1(n19026), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n18999) );
  OAI21_X1 U21948 ( .B1(n19000), .B2(n19028), .A(n18999), .ZN(P2_U2938) );
  AOI22_X1 U21949 ( .A1(n19026), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19001) );
  OAI21_X1 U21950 ( .B1(n19002), .B2(n19028), .A(n19001), .ZN(P2_U2939) );
  AOI22_X1 U21951 ( .A1(n19026), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19003) );
  OAI21_X1 U21952 ( .B1(n19004), .B2(n19028), .A(n19003), .ZN(P2_U2940) );
  AOI22_X1 U21953 ( .A1(n19026), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19005) );
  OAI21_X1 U21954 ( .B1(n19006), .B2(n19028), .A(n19005), .ZN(P2_U2941) );
  AOI22_X1 U21955 ( .A1(n19026), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19007) );
  OAI21_X1 U21956 ( .B1(n19008), .B2(n19028), .A(n19007), .ZN(P2_U2942) );
  AOI22_X1 U21957 ( .A1(n19026), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19009) );
  OAI21_X1 U21958 ( .B1(n19010), .B2(n19028), .A(n19009), .ZN(P2_U2943) );
  AOI22_X1 U21959 ( .A1(n19026), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19011) );
  OAI21_X1 U21960 ( .B1(n19012), .B2(n19028), .A(n19011), .ZN(P2_U2944) );
  AOI22_X1 U21961 ( .A1(n19026), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19013) );
  OAI21_X1 U21962 ( .B1(n19014), .B2(n19028), .A(n19013), .ZN(P2_U2945) );
  INV_X1 U21963 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19016) );
  AOI22_X1 U21964 ( .A1(n19026), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19015) );
  OAI21_X1 U21965 ( .B1(n19016), .B2(n19028), .A(n19015), .ZN(P2_U2946) );
  INV_X1 U21966 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19018) );
  AOI22_X1 U21967 ( .A1(n19026), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19017) );
  OAI21_X1 U21968 ( .B1(n19018), .B2(n19028), .A(n19017), .ZN(P2_U2947) );
  INV_X1 U21969 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19020) );
  AOI22_X1 U21970 ( .A1(n19026), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19019) );
  OAI21_X1 U21971 ( .B1(n19020), .B2(n19028), .A(n19019), .ZN(P2_U2948) );
  INV_X1 U21972 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19022) );
  AOI22_X1 U21973 ( .A1(n19026), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19021) );
  OAI21_X1 U21974 ( .B1(n19022), .B2(n19028), .A(n19021), .ZN(P2_U2949) );
  AOI22_X1 U21975 ( .A1(n19026), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19023) );
  OAI21_X1 U21976 ( .B1(n19024), .B2(n19028), .A(n19023), .ZN(P2_U2950) );
  INV_X1 U21977 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19029) );
  AOI22_X1 U21978 ( .A1(n19026), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19025), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19027) );
  OAI21_X1 U21979 ( .B1(n19029), .B2(n19028), .A(n19027), .ZN(P2_U2951) );
  AOI22_X1 U21980 ( .A1(n9582), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n19033), .ZN(n19032) );
  NAND2_X1 U21981 ( .A1(n19031), .A2(n19030), .ZN(n19034) );
  NAND2_X1 U21982 ( .A1(n19032), .A2(n19034), .ZN(P2_U2966) );
  AOI22_X1 U21983 ( .A1(n9582), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_14__SCAN_IN), .B2(n19033), .ZN(n19035) );
  NAND2_X1 U21984 ( .A1(n19035), .A2(n19034), .ZN(P2_U2981) );
  AOI22_X1 U21985 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19038), .B1(n19037), 
        .B2(n19036), .ZN(n19045) );
  AOI222_X1 U21986 ( .A1(n19043), .A2(n13164), .B1(n19042), .B2(n19041), .C1(
        n19040), .C2(n19039), .ZN(n19044) );
  OAI211_X1 U21987 ( .C1(n19047), .C2(n19046), .A(n19045), .B(n19044), .ZN(
        P2_U3010) );
  AOI22_X1 U21988 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19078), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n19079), .ZN(n19520) );
  INV_X1 U21989 ( .A(n19087), .ZN(n19075) );
  NAND2_X1 U21990 ( .A1(n19086), .A2(n19048), .ZN(n19550) );
  OAI22_X1 U21991 ( .A1(n19640), .A2(n19520), .B1(n19075), .B2(n19550), .ZN(
        n19049) );
  INV_X1 U21992 ( .A(n19049), .ZN(n19052) );
  NOR2_X2 U21993 ( .A1(n19549), .A2(n19050), .ZN(n19602) );
  AOI22_X1 U21994 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19079), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19078), .ZN(n19615) );
  INV_X1 U21995 ( .A(n19615), .ZN(n19517) );
  AOI22_X1 U21996 ( .A1(n19602), .A2(n19091), .B1(n19116), .B2(n19517), .ZN(
        n19051) );
  OAI211_X1 U21997 ( .C1(n19094), .C2(n19053), .A(n19052), .B(n19051), .ZN(
        P2_U3048) );
  AOI22_X1 U21998 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19078), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n19079), .ZN(n19524) );
  NAND2_X1 U21999 ( .A1(n19086), .A2(n19054), .ZN(n19559) );
  OAI22_X1 U22000 ( .A1(n19640), .A2(n19524), .B1(n19075), .B2(n19559), .ZN(
        n19055) );
  INV_X1 U22001 ( .A(n19055), .ZN(n19058) );
  NOR2_X2 U22002 ( .A1(n19549), .A2(n19056), .ZN(n19617) );
  INV_X1 U22003 ( .A(n19621), .ZN(n19521) );
  AOI22_X1 U22004 ( .A1(n19617), .A2(n19091), .B1(n19116), .B2(n19521), .ZN(
        n19057) );
  OAI211_X1 U22005 ( .C1(n19094), .C2(n19059), .A(n19058), .B(n19057), .ZN(
        P2_U3049) );
  AOI22_X1 U22006 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19078), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19079), .ZN(n19527) );
  NAND2_X1 U22007 ( .A1(n19086), .A2(n19060), .ZN(n19396) );
  OAI22_X1 U22008 ( .A1(n19640), .A2(n19527), .B1(n19075), .B2(n19396), .ZN(
        n19061) );
  INV_X1 U22009 ( .A(n19061), .ZN(n19064) );
  NOR2_X2 U22010 ( .A1(n19549), .A2(n19062), .ZN(n19623) );
  INV_X1 U22011 ( .A(n19627), .ZN(n19563) );
  AOI22_X1 U22012 ( .A1(n19623), .A2(n19091), .B1(n19116), .B2(n19563), .ZN(
        n19063) );
  OAI211_X1 U22013 ( .C1(n19094), .C2(n11512), .A(n19064), .B(n19063), .ZN(
        P2_U3050) );
  INV_X1 U22014 ( .A(n19633), .ZN(n19567) );
  AND2_X1 U22015 ( .A1(n19086), .A2(n19065), .ZN(n19628) );
  AOI22_X1 U22016 ( .A1(n19659), .A2(n19567), .B1(n19087), .B2(n19628), .ZN(
        n19068) );
  NOR2_X2 U22017 ( .A1(n19549), .A2(n19066), .ZN(n19629) );
  OAI22_X2 U22018 ( .A1(n14458), .A2(n19089), .B1(n14909), .B2(n19090), .ZN(
        n19630) );
  AOI22_X1 U22019 ( .A1(n19629), .A2(n19091), .B1(n19116), .B2(n19630), .ZN(
        n19067) );
  OAI211_X1 U22020 ( .C1(n19094), .C2(n19069), .A(n19068), .B(n19067), .ZN(
        P2_U3051) );
  AOI22_X1 U22021 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19078), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19079), .ZN(n19647) );
  INV_X1 U22022 ( .A(n19647), .ZN(n19579) );
  INV_X1 U22023 ( .A(n19579), .ZN(n19406) );
  NAND2_X1 U22024 ( .A1(n19086), .A2(n19070), .ZN(n19576) );
  OAI22_X1 U22025 ( .A1(n19640), .A2(n19406), .B1(n19075), .B2(n19576), .ZN(
        n19071) );
  INV_X1 U22026 ( .A(n19071), .ZN(n19074) );
  NOR2_X2 U22027 ( .A1(n19549), .A2(n19072), .ZN(n19643) );
  AOI22_X1 U22028 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19079), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19078), .ZN(n19577) );
  INV_X1 U22029 ( .A(n19577), .ZN(n19644) );
  AOI22_X1 U22030 ( .A1(n19643), .A2(n19091), .B1(n19116), .B2(n19644), .ZN(
        n19073) );
  OAI211_X1 U22031 ( .C1(n19094), .C2(n13450), .A(n19074), .B(n19073), .ZN(
        P2_U3053) );
  INV_X1 U22032 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19082) );
  NAND2_X1 U22033 ( .A1(n19086), .A2(n9589), .ZN(n19584) );
  OAI22_X1 U22034 ( .A1(n19640), .A2(n19653), .B1(n19075), .B2(n19584), .ZN(
        n19076) );
  INV_X1 U22035 ( .A(n19076), .ZN(n19081) );
  NOR2_X2 U22036 ( .A1(n19549), .A2(n19077), .ZN(n19649) );
  AOI22_X1 U22037 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19079), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19078), .ZN(n19585) );
  INV_X1 U22038 ( .A(n19585), .ZN(n19650) );
  AOI22_X1 U22039 ( .A1(n19649), .A2(n19091), .B1(n19116), .B2(n19650), .ZN(
        n19080) );
  OAI211_X1 U22040 ( .C1(n19094), .C2(n19082), .A(n19081), .B(n19080), .ZN(
        P2_U3054) );
  OAI22_X1 U22041 ( .A1(n19084), .A2(n19089), .B1(n19083), .B2(n19090), .ZN(
        n19592) );
  AND2_X1 U22042 ( .A1(n19086), .A2(n9586), .ZN(n19655) );
  AOI22_X1 U22043 ( .A1(n19659), .A2(n19592), .B1(n19087), .B2(n19655), .ZN(
        n19093) );
  NOR2_X2 U22044 ( .A1(n19549), .A2(n19088), .ZN(n19656) );
  OAI22_X2 U22045 ( .A1(n14172), .A2(n19090), .B1(n14437), .B2(n19089), .ZN(
        n19658) );
  AOI22_X1 U22046 ( .A1(n19656), .A2(n19091), .B1(n19116), .B2(n19658), .ZN(
        n19092) );
  OAI211_X1 U22047 ( .C1(n19094), .C2(n11533), .A(n19093), .B(n19092), .ZN(
        P2_U3055) );
  NAND2_X1 U22048 ( .A1(n19761), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19764) );
  OR2_X1 U22049 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19160), .ZN(
        n19103) );
  OAI21_X1 U22050 ( .B1(n19764), .B2(n19388), .A(n19103), .ZN(n19099) );
  NAND2_X1 U22051 ( .A1(n19100), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19095) );
  NAND2_X1 U22052 ( .A1(n19095), .A2(n19611), .ZN(n19097) );
  NOR3_X2 U22053 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19797), .A3(
        n19160), .ZN(n19121) );
  INV_X1 U22054 ( .A(n19121), .ZN(n19096) );
  AOI21_X1 U22055 ( .B1(n19097), .B2(n19096), .A(n19549), .ZN(n19098) );
  AND2_X1 U22056 ( .A1(n19099), .A2(n19098), .ZN(n19107) );
  INV_X1 U22057 ( .A(n19759), .ZN(n19763) );
  INV_X1 U22058 ( .A(n19100), .ZN(n19101) );
  OAI21_X1 U22059 ( .B1(n19101), .B2(n19121), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19102) );
  OAI21_X1 U22060 ( .B1(n19103), .B2(n19763), .A(n19102), .ZN(n19122) );
  INV_X1 U22061 ( .A(n19550), .ZN(n19601) );
  AOI22_X1 U22062 ( .A1(n19122), .A2(n19602), .B1(n19601), .B2(n19121), .ZN(
        n19105) );
  NAND2_X1 U22063 ( .A1(n19761), .A2(n19334), .ZN(n19310) );
  INV_X1 U22064 ( .A(n19520), .ZN(n19612) );
  AOI22_X1 U22065 ( .A1(n19147), .A2(n19517), .B1(n19116), .B2(n19612), .ZN(
        n19104) );
  OAI211_X1 U22066 ( .C1(n19107), .C2(n19106), .A(n19105), .B(n19104), .ZN(
        P2_U3056) );
  INV_X1 U22067 ( .A(n19559), .ZN(n19616) );
  AOI22_X1 U22068 ( .A1(n19122), .A2(n19617), .B1(n19616), .B2(n19121), .ZN(
        n19109) );
  INV_X1 U22069 ( .A(n19524), .ZN(n19618) );
  AOI22_X1 U22070 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19123), .B1(
        n19116), .B2(n19618), .ZN(n19108) );
  OAI211_X1 U22071 ( .C1(n19621), .C2(n19156), .A(n19109), .B(n19108), .ZN(
        P2_U3057) );
  INV_X1 U22072 ( .A(n19396), .ZN(n19622) );
  AOI22_X1 U22073 ( .A1(n19122), .A2(n19623), .B1(n19622), .B2(n19121), .ZN(
        n19111) );
  INV_X1 U22074 ( .A(n19527), .ZN(n19624) );
  AOI22_X1 U22075 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19123), .B1(
        n19116), .B2(n19624), .ZN(n19110) );
  OAI211_X1 U22076 ( .C1(n19627), .C2(n19156), .A(n19111), .B(n19110), .ZN(
        P2_U3058) );
  AOI22_X1 U22077 ( .A1(n19122), .A2(n19629), .B1(n19628), .B2(n19121), .ZN(
        n19113) );
  AOI22_X1 U22078 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19123), .B1(
        n19147), .B2(n19630), .ZN(n19112) );
  OAI211_X1 U22079 ( .C1(n19633), .C2(n19126), .A(n19113), .B(n19112), .ZN(
        P2_U3059) );
  AOI22_X1 U22080 ( .A1(n19122), .A2(n19635), .B1(n19634), .B2(n19121), .ZN(
        n19115) );
  AOI22_X1 U22081 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19123), .B1(
        n19116), .B2(n19636), .ZN(n19114) );
  OAI211_X1 U22082 ( .C1(n19641), .C2(n19156), .A(n19115), .B(n19114), .ZN(
        P2_U3060) );
  INV_X1 U22083 ( .A(n19576), .ZN(n19642) );
  AOI22_X1 U22084 ( .A1(n19122), .A2(n19643), .B1(n19642), .B2(n19121), .ZN(
        n19118) );
  AOI22_X1 U22085 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19123), .B1(
        n19116), .B2(n19579), .ZN(n19117) );
  OAI211_X1 U22086 ( .C1(n19577), .C2(n19156), .A(n19118), .B(n19117), .ZN(
        P2_U3061) );
  INV_X1 U22087 ( .A(n19584), .ZN(n19648) );
  AOI22_X1 U22088 ( .A1(n19122), .A2(n19649), .B1(n19648), .B2(n19121), .ZN(
        n19120) );
  AOI22_X1 U22089 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19123), .B1(
        n19147), .B2(n19650), .ZN(n19119) );
  OAI211_X1 U22090 ( .C1(n19653), .C2(n19126), .A(n19120), .B(n19119), .ZN(
        P2_U3062) );
  INV_X1 U22091 ( .A(n19592), .ZN(n19664) );
  AOI22_X1 U22092 ( .A1(n19122), .A2(n19656), .B1(n19655), .B2(n19121), .ZN(
        n19125) );
  AOI22_X1 U22093 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19123), .B1(
        n19147), .B2(n19658), .ZN(n19124) );
  OAI211_X1 U22094 ( .C1(n19664), .C2(n19126), .A(n19125), .B(n19124), .ZN(
        P2_U3063) );
  NOR3_X2 U22095 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19788), .A3(
        n19160), .ZN(n19150) );
  OAI21_X1 U22096 ( .B1(n19129), .B2(n19150), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19128) );
  NOR2_X1 U22097 ( .A1(n19418), .A2(n19160), .ZN(n19130) );
  INV_X1 U22098 ( .A(n19130), .ZN(n19127) );
  NAND2_X1 U22099 ( .A1(n19128), .A2(n19127), .ZN(n19151) );
  AOI22_X1 U22100 ( .A1(n19151), .A2(n19602), .B1(n19601), .B2(n19150), .ZN(
        n19136) );
  AOI21_X1 U22101 ( .B1(n19129), .B2(n19611), .A(n19150), .ZN(n19133) );
  AOI21_X1 U22102 ( .B1(n19194), .B2(n19156), .A(n19544), .ZN(n19131) );
  NOR2_X1 U22103 ( .A1(n19131), .A2(n19130), .ZN(n19132) );
  MUX2_X1 U22104 ( .A(n19133), .B(n19132), .S(n19759), .Z(n19134) );
  INV_X1 U22105 ( .A(n19194), .ZN(n19152) );
  AOI22_X1 U22106 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19153), .B1(
        n19152), .B2(n19517), .ZN(n19135) );
  OAI211_X1 U22107 ( .C1(n19520), .C2(n19156), .A(n19136), .B(n19135), .ZN(
        P2_U3064) );
  AOI22_X1 U22108 ( .A1(n19151), .A2(n19617), .B1(n19616), .B2(n19150), .ZN(
        n19138) );
  AOI22_X1 U22109 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19153), .B1(
        n19147), .B2(n19618), .ZN(n19137) );
  OAI211_X1 U22110 ( .C1(n19621), .C2(n19194), .A(n19138), .B(n19137), .ZN(
        P2_U3065) );
  AOI22_X1 U22111 ( .A1(n19151), .A2(n19623), .B1(n19622), .B2(n19150), .ZN(
        n19140) );
  AOI22_X1 U22112 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19153), .B1(
        n19147), .B2(n19624), .ZN(n19139) );
  OAI211_X1 U22113 ( .C1(n19627), .C2(n19194), .A(n19140), .B(n19139), .ZN(
        P2_U3066) );
  AOI22_X1 U22114 ( .A1(n19151), .A2(n19629), .B1(n19628), .B2(n19150), .ZN(
        n19142) );
  AOI22_X1 U22115 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19153), .B1(
        n19152), .B2(n19630), .ZN(n19141) );
  OAI211_X1 U22116 ( .C1(n19633), .C2(n19156), .A(n19142), .B(n19141), .ZN(
        P2_U3067) );
  AOI22_X1 U22117 ( .A1(n19151), .A2(n19635), .B1(n19634), .B2(n19150), .ZN(
        n19144) );
  AOI22_X1 U22118 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19153), .B1(
        n19152), .B2(n19530), .ZN(n19143) );
  OAI211_X1 U22119 ( .C1(n19533), .C2(n19156), .A(n19144), .B(n19143), .ZN(
        P2_U3068) );
  AOI22_X1 U22120 ( .A1(n19151), .A2(n19643), .B1(n19642), .B2(n19150), .ZN(
        n19146) );
  AOI22_X1 U22121 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19153), .B1(
        n19147), .B2(n19579), .ZN(n19145) );
  OAI211_X1 U22122 ( .C1(n19577), .C2(n19194), .A(n19146), .B(n19145), .ZN(
        P2_U3069) );
  AOI22_X1 U22123 ( .A1(n19151), .A2(n19649), .B1(n19648), .B2(n19150), .ZN(
        n19149) );
  INV_X1 U22124 ( .A(n19653), .ZN(n19587) );
  AOI22_X1 U22125 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19153), .B1(
        n19147), .B2(n19587), .ZN(n19148) );
  OAI211_X1 U22126 ( .C1(n19585), .C2(n19194), .A(n19149), .B(n19148), .ZN(
        P2_U3070) );
  AOI22_X1 U22127 ( .A1(n19151), .A2(n19656), .B1(n19655), .B2(n19150), .ZN(
        n19155) );
  AOI22_X1 U22128 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19153), .B1(
        n19152), .B2(n19658), .ZN(n19154) );
  OAI211_X1 U22129 ( .C1(n19664), .C2(n19156), .A(n19155), .B(n19154), .ZN(
        P2_U3071) );
  INV_X1 U22130 ( .A(n19757), .ZN(n19452) );
  INV_X1 U22131 ( .A(n19157), .ZN(n19446) );
  INV_X1 U22132 ( .A(n19160), .ZN(n19158) );
  NAND2_X1 U22133 ( .A1(n19446), .A2(n19158), .ZN(n19188) );
  OAI22_X1 U22134 ( .A1(n19194), .A2(n19520), .B1(n19188), .B2(n19550), .ZN(
        n19159) );
  INV_X1 U22135 ( .A(n19159), .ZN(n19169) );
  OAI21_X1 U22136 ( .B1(n19764), .B2(n19452), .A(n19759), .ZN(n19167) );
  NOR2_X1 U22137 ( .A1(n19788), .A2(n19160), .ZN(n19162) );
  OAI211_X1 U22138 ( .C1(n11122), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19188), 
        .B(n19763), .ZN(n19161) );
  OAI211_X1 U22139 ( .C1(n19167), .C2(n19162), .A(n19609), .B(n19161), .ZN(
        n19191) );
  INV_X1 U22140 ( .A(n19162), .ZN(n19166) );
  INV_X1 U22141 ( .A(n19188), .ZN(n19163) );
  OAI21_X1 U22142 ( .B1(n19164), .B2(n19163), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19165) );
  OAI21_X1 U22143 ( .B1(n19167), .B2(n19166), .A(n19165), .ZN(n19190) );
  AOI22_X1 U22144 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19191), .B1(
        n19602), .B2(n19190), .ZN(n19168) );
  OAI211_X1 U22145 ( .C1(n19615), .C2(n19235), .A(n19169), .B(n19168), .ZN(
        P2_U3072) );
  OAI22_X1 U22146 ( .A1(n19235), .A2(n19621), .B1(n19188), .B2(n19559), .ZN(
        n19170) );
  INV_X1 U22147 ( .A(n19170), .ZN(n19172) );
  AOI22_X1 U22148 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19191), .B1(
        n19617), .B2(n19190), .ZN(n19171) );
  OAI211_X1 U22149 ( .C1(n19524), .C2(n19194), .A(n19172), .B(n19171), .ZN(
        P2_U3073) );
  OAI22_X1 U22150 ( .A1(n19235), .A2(n19627), .B1(n19188), .B2(n19396), .ZN(
        n19173) );
  INV_X1 U22151 ( .A(n19173), .ZN(n19175) );
  AOI22_X1 U22152 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19191), .B1(
        n19623), .B2(n19190), .ZN(n19174) );
  OAI211_X1 U22153 ( .C1(n19527), .C2(n19194), .A(n19175), .B(n19174), .ZN(
        P2_U3074) );
  INV_X1 U22154 ( .A(n19630), .ZN(n19356) );
  INV_X1 U22155 ( .A(n19628), .ZN(n19355) );
  OAI22_X1 U22156 ( .A1(n19235), .A2(n19356), .B1(n19188), .B2(n19355), .ZN(
        n19176) );
  INV_X1 U22157 ( .A(n19176), .ZN(n19178) );
  AOI22_X1 U22158 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19191), .B1(
        n19629), .B2(n19190), .ZN(n19177) );
  OAI211_X1 U22159 ( .C1(n19633), .C2(n19194), .A(n19178), .B(n19177), .ZN(
        P2_U3075) );
  INV_X1 U22160 ( .A(n19634), .ZN(n19571) );
  OAI22_X1 U22161 ( .A1(n19194), .A2(n19533), .B1(n19571), .B2(n19188), .ZN(
        n19179) );
  INV_X1 U22162 ( .A(n19179), .ZN(n19181) );
  AOI22_X1 U22163 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19191), .B1(
        n19635), .B2(n19190), .ZN(n19180) );
  OAI211_X1 U22164 ( .C1(n19641), .C2(n19235), .A(n19181), .B(n19180), .ZN(
        P2_U3076) );
  OAI22_X1 U22165 ( .A1(n19194), .A2(n19406), .B1(n19188), .B2(n19576), .ZN(
        n19182) );
  INV_X1 U22166 ( .A(n19182), .ZN(n19184) );
  AOI22_X1 U22167 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19191), .B1(
        n19643), .B2(n19190), .ZN(n19183) );
  OAI211_X1 U22168 ( .C1(n19577), .C2(n19235), .A(n19184), .B(n19183), .ZN(
        P2_U3077) );
  OAI22_X1 U22169 ( .A1(n19194), .A2(n19653), .B1(n19188), .B2(n19584), .ZN(
        n19185) );
  INV_X1 U22170 ( .A(n19185), .ZN(n19187) );
  AOI22_X1 U22171 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19191), .B1(
        n19649), .B2(n19190), .ZN(n19186) );
  OAI211_X1 U22172 ( .C1(n19585), .C2(n19235), .A(n19187), .B(n19186), .ZN(
        P2_U3078) );
  INV_X1 U22173 ( .A(n19658), .ZN(n19371) );
  INV_X1 U22174 ( .A(n19655), .ZN(n19370) );
  OAI22_X1 U22175 ( .A1(n19235), .A2(n19371), .B1(n19188), .B2(n19370), .ZN(
        n19189) );
  INV_X1 U22176 ( .A(n19189), .ZN(n19193) );
  AOI22_X1 U22177 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19191), .B1(
        n19656), .B2(n19190), .ZN(n19192) );
  OAI211_X1 U22178 ( .C1(n19664), .C2(n19194), .A(n19193), .B(n19192), .ZN(
        P2_U3079) );
  INV_X1 U22179 ( .A(n19515), .ZN(n19195) );
  NAND3_X1 U22180 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19769), .A3(
        n19788), .ZN(n19243) );
  NOR2_X1 U22181 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19243), .ZN(
        n19204) );
  INV_X1 U22182 ( .A(n19204), .ZN(n19229) );
  OAI22_X1 U22183 ( .A1(n19273), .A2(n19615), .B1(n19229), .B2(n19550), .ZN(
        n19196) );
  INV_X1 U22184 ( .A(n19196), .ZN(n19210) );
  AOI21_X1 U22185 ( .B1(n19197), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19202) );
  AOI21_X1 U22186 ( .B1(n19273), .B2(n19235), .A(n19544), .ZN(n19198) );
  NOR2_X1 U22187 ( .A1(n19198), .A2(n19763), .ZN(n19203) );
  NAND2_X1 U22188 ( .A1(n19200), .A2(n19199), .ZN(n19479) );
  OR2_X1 U22189 ( .A1(n19478), .A2(n19479), .ZN(n19207) );
  NAND2_X1 U22190 ( .A1(n19203), .A2(n19207), .ZN(n19201) );
  OAI211_X1 U22191 ( .C1(n19204), .C2(n19202), .A(n19201), .B(n19609), .ZN(
        n19232) );
  INV_X1 U22192 ( .A(n19203), .ZN(n19208) );
  OAI21_X1 U22193 ( .B1(n19205), .B2(n19204), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19206) );
  AOI22_X1 U22194 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19232), .B1(
        n19602), .B2(n19231), .ZN(n19209) );
  OAI211_X1 U22195 ( .C1(n19520), .C2(n19235), .A(n19210), .B(n19209), .ZN(
        P2_U3080) );
  OAI22_X1 U22196 ( .A1(n19235), .A2(n19524), .B1(n19559), .B2(n19229), .ZN(
        n19211) );
  INV_X1 U22197 ( .A(n19211), .ZN(n19213) );
  AOI22_X1 U22198 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19232), .B1(
        n19617), .B2(n19231), .ZN(n19212) );
  OAI211_X1 U22199 ( .C1(n19621), .C2(n19273), .A(n19213), .B(n19212), .ZN(
        P2_U3081) );
  OAI22_X1 U22200 ( .A1(n19235), .A2(n19527), .B1(n19396), .B2(n19229), .ZN(
        n19214) );
  INV_X1 U22201 ( .A(n19214), .ZN(n19216) );
  AOI22_X1 U22202 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19232), .B1(
        n19623), .B2(n19231), .ZN(n19215) );
  OAI211_X1 U22203 ( .C1(n19627), .C2(n19273), .A(n19216), .B(n19215), .ZN(
        P2_U3082) );
  OAI22_X1 U22204 ( .A1(n19273), .A2(n19356), .B1(n19355), .B2(n19229), .ZN(
        n19217) );
  INV_X1 U22205 ( .A(n19217), .ZN(n19219) );
  AOI22_X1 U22206 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19232), .B1(
        n19629), .B2(n19231), .ZN(n19218) );
  OAI211_X1 U22207 ( .C1(n19633), .C2(n19235), .A(n19219), .B(n19218), .ZN(
        P2_U3083) );
  OAI22_X1 U22208 ( .A1(n19235), .A2(n19533), .B1(n19571), .B2(n19229), .ZN(
        n19220) );
  INV_X1 U22209 ( .A(n19220), .ZN(n19222) );
  AOI22_X1 U22210 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19232), .B1(
        n19635), .B2(n19231), .ZN(n19221) );
  OAI211_X1 U22211 ( .C1(n19641), .C2(n19273), .A(n19222), .B(n19221), .ZN(
        P2_U3084) );
  OAI22_X1 U22212 ( .A1(n19273), .A2(n19577), .B1(n19229), .B2(n19576), .ZN(
        n19223) );
  INV_X1 U22213 ( .A(n19223), .ZN(n19225) );
  AOI22_X1 U22214 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19232), .B1(
        n19643), .B2(n19231), .ZN(n19224) );
  OAI211_X1 U22215 ( .C1(n19647), .C2(n19235), .A(n19225), .B(n19224), .ZN(
        P2_U3085) );
  OAI22_X1 U22216 ( .A1(n19235), .A2(n19653), .B1(n19229), .B2(n19584), .ZN(
        n19226) );
  INV_X1 U22217 ( .A(n19226), .ZN(n19228) );
  AOI22_X1 U22218 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19232), .B1(
        n19649), .B2(n19231), .ZN(n19227) );
  OAI211_X1 U22219 ( .C1(n19585), .C2(n19273), .A(n19228), .B(n19227), .ZN(
        P2_U3086) );
  OAI22_X1 U22220 ( .A1(n19273), .A2(n19371), .B1(n19370), .B2(n19229), .ZN(
        n19230) );
  INV_X1 U22221 ( .A(n19230), .ZN(n19234) );
  AOI22_X1 U22222 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19232), .B1(
        n19656), .B2(n19231), .ZN(n19233) );
  OAI211_X1 U22223 ( .C1(n19664), .C2(n19235), .A(n19234), .B(n19233), .ZN(
        P2_U3087) );
  OR2_X1 U22224 ( .A1(n19764), .A2(n19515), .ZN(n19236) );
  NOR2_X1 U22225 ( .A1(n19797), .A2(n19243), .ZN(n19279) );
  INV_X1 U22226 ( .A(n19279), .ZN(n19267) );
  OAI211_X1 U22227 ( .C1(n11121), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19267), 
        .B(n19763), .ZN(n19237) );
  NAND2_X1 U22228 ( .A1(n19237), .A2(n19609), .ZN(n19238) );
  AOI21_X1 U22229 ( .B1(n19240), .B2(n19243), .A(n19238), .ZN(n19252) );
  OAI22_X1 U22230 ( .A1(n19302), .A2(n19615), .B1(n19550), .B2(n19267), .ZN(
        n19239) );
  INV_X1 U22231 ( .A(n19239), .ZN(n19247) );
  INV_X1 U22232 ( .A(n19240), .ZN(n19244) );
  OAI21_X1 U22233 ( .B1(n19241), .B2(n19279), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19242) );
  OAI21_X1 U22234 ( .B1(n19244), .B2(n19243), .A(n19242), .ZN(n19269) );
  INV_X1 U22235 ( .A(n19273), .ZN(n19245) );
  AOI22_X1 U22236 ( .A1(n19602), .A2(n19269), .B1(n19245), .B2(n19612), .ZN(
        n19246) );
  OAI211_X1 U22237 ( .C1(n19252), .C2(n20829), .A(n19247), .B(n19246), .ZN(
        P2_U3088) );
  OAI22_X1 U22238 ( .A1(n19273), .A2(n19524), .B1(n19559), .B2(n19267), .ZN(
        n19248) );
  INV_X1 U22239 ( .A(n19248), .ZN(n19250) );
  INV_X1 U22240 ( .A(n19302), .ZN(n19294) );
  AOI22_X1 U22241 ( .A1(n19617), .A2(n19269), .B1(n19294), .B2(n19521), .ZN(
        n19249) );
  OAI211_X1 U22242 ( .C1(n19252), .C2(n11096), .A(n19250), .B(n19249), .ZN(
        P2_U3089) );
  OAI22_X1 U22243 ( .A1(n19302), .A2(n19627), .B1(n19396), .B2(n19267), .ZN(
        n19251) );
  INV_X1 U22244 ( .A(n19251), .ZN(n19254) );
  INV_X1 U22245 ( .A(n19252), .ZN(n19270) );
  AOI22_X1 U22246 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19270), .B1(
        n19623), .B2(n19269), .ZN(n19253) );
  OAI211_X1 U22247 ( .C1(n19527), .C2(n19273), .A(n19254), .B(n19253), .ZN(
        P2_U3090) );
  OAI22_X1 U22248 ( .A1(n19302), .A2(n19356), .B1(n19355), .B2(n19267), .ZN(
        n19255) );
  INV_X1 U22249 ( .A(n19255), .ZN(n19257) );
  AOI22_X1 U22250 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19270), .B1(
        n19629), .B2(n19269), .ZN(n19256) );
  OAI211_X1 U22251 ( .C1(n19633), .C2(n19273), .A(n19257), .B(n19256), .ZN(
        P2_U3091) );
  OAI22_X1 U22252 ( .A1(n19302), .A2(n19641), .B1(n19571), .B2(n19267), .ZN(
        n19258) );
  INV_X1 U22253 ( .A(n19258), .ZN(n19260) );
  AOI22_X1 U22254 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19270), .B1(
        n19635), .B2(n19269), .ZN(n19259) );
  OAI211_X1 U22255 ( .C1(n19533), .C2(n19273), .A(n19260), .B(n19259), .ZN(
        P2_U3092) );
  OAI22_X1 U22256 ( .A1(n19273), .A2(n19406), .B1(n19267), .B2(n19576), .ZN(
        n19261) );
  INV_X1 U22257 ( .A(n19261), .ZN(n19263) );
  AOI22_X1 U22258 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19270), .B1(
        n19643), .B2(n19269), .ZN(n19262) );
  OAI211_X1 U22259 ( .C1(n19577), .C2(n19302), .A(n19263), .B(n19262), .ZN(
        P2_U3093) );
  OAI22_X1 U22260 ( .A1(n19302), .A2(n19585), .B1(n19584), .B2(n19267), .ZN(
        n19264) );
  INV_X1 U22261 ( .A(n19264), .ZN(n19266) );
  AOI22_X1 U22262 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19270), .B1(
        n19649), .B2(n19269), .ZN(n19265) );
  OAI211_X1 U22263 ( .C1(n19653), .C2(n19273), .A(n19266), .B(n19265), .ZN(
        P2_U3094) );
  OAI22_X1 U22264 ( .A1(n19302), .A2(n19371), .B1(n19370), .B2(n19267), .ZN(
        n19268) );
  INV_X1 U22265 ( .A(n19268), .ZN(n19272) );
  AOI22_X1 U22266 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19270), .B1(
        n19656), .B2(n19269), .ZN(n19271) );
  OAI211_X1 U22267 ( .C1(n19664), .C2(n19273), .A(n19272), .B(n19271), .ZN(
        P2_U3095) );
  INV_X1 U22268 ( .A(n19274), .ZN(n19275) );
  NOR2_X2 U22269 ( .A1(n19762), .A2(n19275), .ZN(n19324) );
  NOR2_X1 U22270 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19309), .ZN(
        n19297) );
  NOR2_X1 U22271 ( .A1(n19279), .A2(n19297), .ZN(n19276) );
  OR2_X1 U22272 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19276), .ZN(n19277) );
  NOR3_X1 U22273 ( .A1(n11118), .A2(n19297), .A3(n19665), .ZN(n19280) );
  AOI21_X1 U22274 ( .B1(n19665), .B2(n19277), .A(n19280), .ZN(n19298) );
  AOI22_X1 U22275 ( .A1(n19298), .A2(n19602), .B1(n19601), .B2(n19297), .ZN(
        n19283) );
  AOI21_X1 U22276 ( .B1(n19302), .B2(n19333), .A(n19544), .ZN(n19278) );
  AOI221_X1 U22277 ( .B1(n19611), .B2(n19279), .C1(n19611), .C2(n19278), .A(
        n19297), .ZN(n19281) );
  AOI22_X1 U22278 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19299), .B1(
        n19294), .B2(n19612), .ZN(n19282) );
  OAI211_X1 U22279 ( .C1(n19615), .C2(n19333), .A(n19283), .B(n19282), .ZN(
        P2_U3096) );
  AOI22_X1 U22280 ( .A1(n19298), .A2(n19617), .B1(n19616), .B2(n19297), .ZN(
        n19285) );
  AOI22_X1 U22281 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19299), .B1(
        n19324), .B2(n19521), .ZN(n19284) );
  OAI211_X1 U22282 ( .C1(n19524), .C2(n19302), .A(n19285), .B(n19284), .ZN(
        P2_U3097) );
  AOI22_X1 U22283 ( .A1(n19298), .A2(n19623), .B1(n19622), .B2(n19297), .ZN(
        n19287) );
  AOI22_X1 U22284 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19299), .B1(
        n19324), .B2(n19563), .ZN(n19286) );
  OAI211_X1 U22285 ( .C1(n19527), .C2(n19302), .A(n19287), .B(n19286), .ZN(
        P2_U3098) );
  AOI22_X1 U22286 ( .A1(n19298), .A2(n19629), .B1(n19628), .B2(n19297), .ZN(
        n19289) );
  AOI22_X1 U22287 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19299), .B1(
        n19324), .B2(n19630), .ZN(n19288) );
  OAI211_X1 U22288 ( .C1(n19633), .C2(n19302), .A(n19289), .B(n19288), .ZN(
        P2_U3099) );
  AOI22_X1 U22289 ( .A1(n19298), .A2(n19635), .B1(n19634), .B2(n19297), .ZN(
        n19291) );
  AOI22_X1 U22290 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19299), .B1(
        n19324), .B2(n19530), .ZN(n19290) );
  OAI211_X1 U22291 ( .C1(n19533), .C2(n19302), .A(n19291), .B(n19290), .ZN(
        P2_U3100) );
  AOI22_X1 U22292 ( .A1(n19298), .A2(n19643), .B1(n19642), .B2(n19297), .ZN(
        n19293) );
  AOI22_X1 U22293 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19299), .B1(
        n19324), .B2(n19644), .ZN(n19292) );
  OAI211_X1 U22294 ( .C1(n19647), .C2(n19302), .A(n19293), .B(n19292), .ZN(
        P2_U3101) );
  AOI22_X1 U22295 ( .A1(n19298), .A2(n19649), .B1(n19648), .B2(n19297), .ZN(
        n19296) );
  AOI22_X1 U22296 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19299), .B1(
        n19294), .B2(n19587), .ZN(n19295) );
  OAI211_X1 U22297 ( .C1(n19585), .C2(n19333), .A(n19296), .B(n19295), .ZN(
        P2_U3102) );
  AOI22_X1 U22298 ( .A1(n19298), .A2(n19656), .B1(n19655), .B2(n19297), .ZN(
        n19301) );
  AOI22_X1 U22299 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19299), .B1(
        n19324), .B2(n19658), .ZN(n19300) );
  OAI211_X1 U22300 ( .C1(n19664), .C2(n19302), .A(n19301), .B(n19300), .ZN(
        P2_U3103) );
  OAI21_X1 U22301 ( .B1(n19764), .B2(n19762), .A(n19309), .ZN(n19306) );
  NAND2_X1 U22302 ( .A1(n11124), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19303) );
  NAND2_X1 U22303 ( .A1(n19303), .A2(n19611), .ZN(n19304) );
  AOI21_X1 U22304 ( .B1(n19304), .B2(n19340), .A(n19549), .ZN(n19305) );
  INV_X1 U22305 ( .A(n11124), .ZN(n19307) );
  INV_X1 U22306 ( .A(n19340), .ZN(n19343) );
  OAI21_X1 U22307 ( .B1(n19307), .B2(n19343), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19308) );
  OAI21_X1 U22308 ( .B1(n19309), .B2(n19763), .A(n19308), .ZN(n19328) );
  AOI22_X1 U22309 ( .A1(n19328), .A2(n19602), .B1(n19343), .B2(n19601), .ZN(
        n19312) );
  INV_X1 U22310 ( .A(n19377), .ZN(n19329) );
  AOI22_X1 U22311 ( .A1(n19329), .A2(n19517), .B1(n19324), .B2(n19612), .ZN(
        n19311) );
  OAI211_X1 U22312 ( .C1(n19327), .C2(n11626), .A(n19312), .B(n19311), .ZN(
        P2_U3104) );
  AOI22_X1 U22313 ( .A1(n19328), .A2(n19617), .B1(n19343), .B2(n19616), .ZN(
        n19314) );
  AOI22_X1 U22314 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19330), .B1(
        n19324), .B2(n19618), .ZN(n19313) );
  OAI211_X1 U22315 ( .C1(n19621), .C2(n19377), .A(n19314), .B(n19313), .ZN(
        P2_U3105) );
  AOI22_X1 U22316 ( .A1(n19328), .A2(n19623), .B1(n19343), .B2(n19622), .ZN(
        n19316) );
  AOI22_X1 U22317 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19330), .B1(
        n19324), .B2(n19624), .ZN(n19315) );
  OAI211_X1 U22318 ( .C1(n19627), .C2(n19377), .A(n19316), .B(n19315), .ZN(
        P2_U3106) );
  AOI22_X1 U22319 ( .A1(n19328), .A2(n19629), .B1(n19343), .B2(n19628), .ZN(
        n19318) );
  AOI22_X1 U22320 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19330), .B1(
        n19329), .B2(n19630), .ZN(n19317) );
  OAI211_X1 U22321 ( .C1(n19633), .C2(n19333), .A(n19318), .B(n19317), .ZN(
        P2_U3107) );
  AOI22_X1 U22322 ( .A1(n19328), .A2(n19635), .B1(n19343), .B2(n19634), .ZN(
        n19320) );
  AOI22_X1 U22323 ( .A1(n19329), .A2(n19530), .B1(n19324), .B2(n19636), .ZN(
        n19319) );
  OAI211_X1 U22324 ( .C1(n19327), .C2(n19321), .A(n19320), .B(n19319), .ZN(
        P2_U3108) );
  AOI22_X1 U22325 ( .A1(n19328), .A2(n19643), .B1(n19343), .B2(n19642), .ZN(
        n19323) );
  AOI22_X1 U22326 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19330), .B1(
        n19324), .B2(n19579), .ZN(n19322) );
  OAI211_X1 U22327 ( .C1(n19577), .C2(n19377), .A(n19323), .B(n19322), .ZN(
        P2_U3109) );
  AOI22_X1 U22328 ( .A1(n19328), .A2(n19649), .B1(n19343), .B2(n19648), .ZN(
        n19326) );
  AOI22_X1 U22329 ( .A1(n19329), .A2(n19650), .B1(n19324), .B2(n19587), .ZN(
        n19325) );
  OAI211_X1 U22330 ( .C1(n19327), .C2(n11186), .A(n19326), .B(n19325), .ZN(
        P2_U3110) );
  AOI22_X1 U22331 ( .A1(n19328), .A2(n19656), .B1(n19343), .B2(n19655), .ZN(
        n19332) );
  AOI22_X1 U22332 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19330), .B1(
        n19329), .B2(n19658), .ZN(n19331) );
  OAI211_X1 U22333 ( .C1(n19664), .C2(n19333), .A(n19332), .B(n19331), .ZN(
        P2_U3111) );
  NOR2_X1 U22334 ( .A1(n19769), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19447) );
  INV_X1 U22335 ( .A(n19447), .ZN(n19451) );
  NOR2_X1 U22336 ( .A1(n19336), .A2(n19451), .ZN(n19344) );
  INV_X1 U22337 ( .A(n19344), .ZN(n19369) );
  OAI22_X1 U22338 ( .A1(n19416), .A2(n19615), .B1(n19550), .B2(n19369), .ZN(
        n19337) );
  INV_X1 U22339 ( .A(n19337), .ZN(n19348) );
  NAND2_X1 U22340 ( .A1(n19416), .A2(n19377), .ZN(n19338) );
  AOI21_X1 U22341 ( .B1(n19338), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19763), 
        .ZN(n19342) );
  OAI21_X1 U22342 ( .B1(n11134), .B2(n19665), .A(n19611), .ZN(n19339) );
  AOI21_X1 U22343 ( .B1(n19342), .B2(n19340), .A(n19339), .ZN(n19341) );
  OAI21_X1 U22344 ( .B1(n19343), .B2(n19344), .A(n19342), .ZN(n19346) );
  OAI21_X1 U22345 ( .B1(n11134), .B2(n19344), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19345) );
  NAND2_X1 U22346 ( .A1(n19346), .A2(n19345), .ZN(n19373) );
  AOI22_X1 U22347 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19374), .B1(
        n19602), .B2(n19373), .ZN(n19347) );
  OAI211_X1 U22348 ( .C1(n19520), .C2(n19377), .A(n19348), .B(n19347), .ZN(
        P2_U3112) );
  OAI22_X1 U22349 ( .A1(n19377), .A2(n19524), .B1(n19559), .B2(n19369), .ZN(
        n19349) );
  INV_X1 U22350 ( .A(n19349), .ZN(n19351) );
  AOI22_X1 U22351 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19374), .B1(
        n19373), .B2(n19617), .ZN(n19350) );
  OAI211_X1 U22352 ( .C1(n19621), .C2(n19416), .A(n19351), .B(n19350), .ZN(
        P2_U3113) );
  OAI22_X1 U22353 ( .A1(n19377), .A2(n19527), .B1(n19396), .B2(n19369), .ZN(
        n19352) );
  INV_X1 U22354 ( .A(n19352), .ZN(n19354) );
  AOI22_X1 U22355 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19374), .B1(
        n19373), .B2(n19623), .ZN(n19353) );
  OAI211_X1 U22356 ( .C1(n19627), .C2(n19416), .A(n19354), .B(n19353), .ZN(
        P2_U3114) );
  OAI22_X1 U22357 ( .A1(n19416), .A2(n19356), .B1(n19355), .B2(n19369), .ZN(
        n19357) );
  INV_X1 U22358 ( .A(n19357), .ZN(n19359) );
  AOI22_X1 U22359 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19374), .B1(
        n19373), .B2(n19629), .ZN(n19358) );
  OAI211_X1 U22360 ( .C1(n19633), .C2(n19377), .A(n19359), .B(n19358), .ZN(
        P2_U3115) );
  OAI22_X1 U22361 ( .A1(n19416), .A2(n19641), .B1(n19571), .B2(n19369), .ZN(
        n19360) );
  INV_X1 U22362 ( .A(n19360), .ZN(n19362) );
  AOI22_X1 U22363 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19374), .B1(
        n19373), .B2(n19635), .ZN(n19361) );
  OAI211_X1 U22364 ( .C1(n19533), .C2(n19377), .A(n19362), .B(n19361), .ZN(
        P2_U3116) );
  OAI22_X1 U22365 ( .A1(n19377), .A2(n19406), .B1(n19369), .B2(n19576), .ZN(
        n19363) );
  INV_X1 U22366 ( .A(n19363), .ZN(n19365) );
  AOI22_X1 U22367 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19374), .B1(
        n19373), .B2(n19643), .ZN(n19364) );
  OAI211_X1 U22368 ( .C1(n19577), .C2(n19416), .A(n19365), .B(n19364), .ZN(
        P2_U3117) );
  OAI22_X1 U22369 ( .A1(n19416), .A2(n19585), .B1(n19584), .B2(n19369), .ZN(
        n19366) );
  INV_X1 U22370 ( .A(n19366), .ZN(n19368) );
  AOI22_X1 U22371 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19374), .B1(
        n19373), .B2(n19649), .ZN(n19367) );
  OAI211_X1 U22372 ( .C1(n19653), .C2(n19377), .A(n19368), .B(n19367), .ZN(
        P2_U3118) );
  OAI22_X1 U22373 ( .A1(n19416), .A2(n19371), .B1(n19370), .B2(n19369), .ZN(
        n19372) );
  INV_X1 U22374 ( .A(n19372), .ZN(n19376) );
  AOI22_X1 U22375 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19374), .B1(
        n19373), .B2(n19656), .ZN(n19375) );
  OAI211_X1 U22376 ( .C1(n19664), .C2(n19377), .A(n19376), .B(n19375), .ZN(
        P2_U3119) );
  OR2_X1 U22377 ( .A1(n19761), .A2(n19544), .ZN(n19603) );
  OAI21_X1 U22378 ( .B1(n19603), .B2(n19388), .A(n19759), .ZN(n19387) );
  NAND2_X1 U22379 ( .A1(n19447), .A2(n19788), .ZN(n19386) );
  INV_X1 U22380 ( .A(n19386), .ZN(n19378) );
  OR2_X1 U22381 ( .A1(n19387), .A2(n19378), .ZN(n19382) );
  OR2_X1 U22382 ( .A1(n11187), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19380) );
  NOR3_X1 U22383 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19797), .A3(
        n19451), .ZN(n19420) );
  NOR2_X1 U22384 ( .A1(n19759), .A2(n19420), .ZN(n19379) );
  AOI21_X1 U22385 ( .B1(n19380), .B2(n19379), .A(n19549), .ZN(n19381) );
  INV_X1 U22386 ( .A(n19420), .ZN(n19405) );
  OAI22_X1 U22387 ( .A1(n19416), .A2(n19520), .B1(n19550), .B2(n19405), .ZN(
        n19383) );
  INV_X1 U22388 ( .A(n19383), .ZN(n19390) );
  OAI21_X1 U22389 ( .B1(n19384), .B2(n19420), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19385) );
  OAI21_X1 U22390 ( .B1(n19387), .B2(n19386), .A(n19385), .ZN(n19412) );
  AOI22_X1 U22391 ( .A1(n19602), .A2(n19412), .B1(n19436), .B2(n19517), .ZN(
        n19389) );
  OAI211_X1 U22392 ( .C1(n19393), .C2(n19391), .A(n19390), .B(n19389), .ZN(
        P2_U3120) );
  OAI22_X1 U22393 ( .A1(n19416), .A2(n19524), .B1(n19559), .B2(n19405), .ZN(
        n19392) );
  INV_X1 U22394 ( .A(n19392), .ZN(n19395) );
  AOI22_X1 U22395 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19413), .B1(
        n19617), .B2(n19412), .ZN(n19394) );
  OAI211_X1 U22396 ( .C1(n19621), .C2(n19444), .A(n19395), .B(n19394), .ZN(
        P2_U3121) );
  OAI22_X1 U22397 ( .A1(n19416), .A2(n19527), .B1(n19396), .B2(n19405), .ZN(
        n19397) );
  INV_X1 U22398 ( .A(n19397), .ZN(n19399) );
  AOI22_X1 U22399 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19413), .B1(
        n19623), .B2(n19412), .ZN(n19398) );
  OAI211_X1 U22400 ( .C1(n19627), .C2(n19444), .A(n19399), .B(n19398), .ZN(
        P2_U3122) );
  AOI22_X1 U22401 ( .A1(n19436), .A2(n19630), .B1(n19628), .B2(n19420), .ZN(
        n19401) );
  AOI22_X1 U22402 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19413), .B1(
        n19629), .B2(n19412), .ZN(n19400) );
  OAI211_X1 U22403 ( .C1(n19633), .C2(n19416), .A(n19401), .B(n19400), .ZN(
        P2_U3123) );
  OAI22_X1 U22404 ( .A1(n19416), .A2(n19533), .B1(n19571), .B2(n19405), .ZN(
        n19402) );
  INV_X1 U22405 ( .A(n19402), .ZN(n19404) );
  AOI22_X1 U22406 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19413), .B1(
        n19635), .B2(n19412), .ZN(n19403) );
  OAI211_X1 U22407 ( .C1(n19641), .C2(n19444), .A(n19404), .B(n19403), .ZN(
        P2_U3124) );
  OAI22_X1 U22408 ( .A1(n19416), .A2(n19406), .B1(n19576), .B2(n19405), .ZN(
        n19407) );
  INV_X1 U22409 ( .A(n19407), .ZN(n19409) );
  AOI22_X1 U22410 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19413), .B1(
        n19643), .B2(n19412), .ZN(n19408) );
  OAI211_X1 U22411 ( .C1(n19577), .C2(n19444), .A(n19409), .B(n19408), .ZN(
        P2_U3125) );
  AOI22_X1 U22412 ( .A1(n19436), .A2(n19650), .B1(n19648), .B2(n19420), .ZN(
        n19411) );
  AOI22_X1 U22413 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19413), .B1(
        n19649), .B2(n19412), .ZN(n19410) );
  OAI211_X1 U22414 ( .C1(n19653), .C2(n19416), .A(n19411), .B(n19410), .ZN(
        P2_U3126) );
  AOI22_X1 U22415 ( .A1(n19436), .A2(n19658), .B1(n19655), .B2(n19420), .ZN(
        n19415) );
  AOI22_X1 U22416 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19413), .B1(
        n19656), .B2(n19412), .ZN(n19414) );
  OAI211_X1 U22417 ( .C1(n19664), .C2(n19416), .A(n19415), .B(n19414), .ZN(
        P2_U3127) );
  NOR3_X2 U22418 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19788), .A3(
        n19451), .ZN(n19439) );
  OAI21_X1 U22419 ( .B1(n19419), .B2(n19439), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19417) );
  OAI21_X1 U22420 ( .B1(n19451), .B2(n19418), .A(n19417), .ZN(n19440) );
  AOI22_X1 U22421 ( .A1(n19440), .A2(n19602), .B1(n19601), .B2(n19439), .ZN(
        n19425) );
  INV_X1 U22422 ( .A(n19419), .ZN(n19422) );
  AOI221_X1 U22423 ( .B1(n19436), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19466), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19420), .ZN(n19421) );
  AOI211_X1 U22424 ( .C1(n19422), .C2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19421), .ZN(n19423) );
  AOI22_X1 U22425 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19441), .B1(
        n19466), .B2(n19517), .ZN(n19424) );
  OAI211_X1 U22426 ( .C1(n19520), .C2(n19444), .A(n19425), .B(n19424), .ZN(
        P2_U3128) );
  AOI22_X1 U22427 ( .A1(n19440), .A2(n19617), .B1(n19616), .B2(n19439), .ZN(
        n19427) );
  AOI22_X1 U22428 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19441), .B1(
        n19436), .B2(n19618), .ZN(n19426) );
  OAI211_X1 U22429 ( .C1(n19621), .C2(n19477), .A(n19427), .B(n19426), .ZN(
        P2_U3129) );
  AOI22_X1 U22430 ( .A1(n19440), .A2(n19623), .B1(n19622), .B2(n19439), .ZN(
        n19429) );
  AOI22_X1 U22431 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19441), .B1(
        n19436), .B2(n19624), .ZN(n19428) );
  OAI211_X1 U22432 ( .C1(n19627), .C2(n19477), .A(n19429), .B(n19428), .ZN(
        P2_U3130) );
  AOI22_X1 U22433 ( .A1(n19440), .A2(n19629), .B1(n19628), .B2(n19439), .ZN(
        n19431) );
  AOI22_X1 U22434 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19441), .B1(
        n19466), .B2(n19630), .ZN(n19430) );
  OAI211_X1 U22435 ( .C1(n19633), .C2(n19444), .A(n19431), .B(n19430), .ZN(
        P2_U3131) );
  AOI22_X1 U22436 ( .A1(n19440), .A2(n19635), .B1(n19634), .B2(n19439), .ZN(
        n19433) );
  AOI22_X1 U22437 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19441), .B1(
        n19436), .B2(n19636), .ZN(n19432) );
  OAI211_X1 U22438 ( .C1(n19641), .C2(n19477), .A(n19433), .B(n19432), .ZN(
        P2_U3132) );
  AOI22_X1 U22439 ( .A1(n19440), .A2(n19643), .B1(n19642), .B2(n19439), .ZN(
        n19435) );
  AOI22_X1 U22440 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19441), .B1(
        n19466), .B2(n19644), .ZN(n19434) );
  OAI211_X1 U22441 ( .C1(n19647), .C2(n19444), .A(n19435), .B(n19434), .ZN(
        P2_U3133) );
  AOI22_X1 U22442 ( .A1(n19440), .A2(n19649), .B1(n19648), .B2(n19439), .ZN(
        n19438) );
  AOI22_X1 U22443 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19441), .B1(
        n19436), .B2(n19587), .ZN(n19437) );
  OAI211_X1 U22444 ( .C1(n19585), .C2(n19477), .A(n19438), .B(n19437), .ZN(
        P2_U3134) );
  AOI22_X1 U22445 ( .A1(n19440), .A2(n19656), .B1(n19655), .B2(n19439), .ZN(
        n19443) );
  AOI22_X1 U22446 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19441), .B1(
        n19466), .B2(n19658), .ZN(n19442) );
  OAI211_X1 U22447 ( .C1(n19664), .C2(n19444), .A(n19443), .B(n19442), .ZN(
        P2_U3135) );
  NAND2_X1 U22448 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19447), .ZN(
        n19450) );
  NAND2_X1 U22449 ( .A1(n19447), .A2(n19446), .ZN(n19453) );
  INV_X1 U22450 ( .A(n19453), .ZN(n19471) );
  OAI21_X1 U22451 ( .B1(n19448), .B2(n19471), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19449) );
  OAI21_X1 U22452 ( .B1(n19450), .B2(n19763), .A(n19449), .ZN(n19472) );
  AOI22_X1 U22453 ( .A1(n19472), .A2(n19602), .B1(n19601), .B2(n19471), .ZN(
        n19457) );
  OAI22_X1 U22454 ( .A1(n19603), .A2(n19452), .B1(n19788), .B2(n19451), .ZN(
        n19455) );
  OAI211_X1 U22455 ( .C1(n11123), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19453), 
        .B(n19763), .ZN(n19454) );
  NAND3_X1 U22456 ( .A1(n19455), .A2(n19609), .A3(n19454), .ZN(n19474) );
  AOI22_X1 U22457 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19474), .B1(
        n19466), .B2(n19612), .ZN(n19456) );
  OAI211_X1 U22458 ( .C1(n19615), .C2(n19508), .A(n19457), .B(n19456), .ZN(
        P2_U3136) );
  AOI22_X1 U22459 ( .A1(n19472), .A2(n19617), .B1(n19616), .B2(n19471), .ZN(
        n19459) );
  AOI22_X1 U22460 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19474), .B1(
        n19466), .B2(n19618), .ZN(n19458) );
  OAI211_X1 U22461 ( .C1(n19621), .C2(n19508), .A(n19459), .B(n19458), .ZN(
        P2_U3137) );
  AOI22_X1 U22462 ( .A1(n19472), .A2(n19623), .B1(n19622), .B2(n19471), .ZN(
        n19461) );
  AOI22_X1 U22463 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19474), .B1(
        n19466), .B2(n19624), .ZN(n19460) );
  OAI211_X1 U22464 ( .C1(n19627), .C2(n19508), .A(n19461), .B(n19460), .ZN(
        P2_U3138) );
  AOI22_X1 U22465 ( .A1(n19472), .A2(n19629), .B1(n19628), .B2(n19471), .ZN(
        n19463) );
  INV_X1 U22466 ( .A(n19508), .ZN(n19473) );
  AOI22_X1 U22467 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19474), .B1(
        n19473), .B2(n19630), .ZN(n19462) );
  OAI211_X1 U22468 ( .C1(n19633), .C2(n19477), .A(n19463), .B(n19462), .ZN(
        P2_U3139) );
  AOI22_X1 U22469 ( .A1(n19472), .A2(n19635), .B1(n19634), .B2(n19471), .ZN(
        n19465) );
  AOI22_X1 U22470 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19474), .B1(
        n19473), .B2(n19530), .ZN(n19464) );
  OAI211_X1 U22471 ( .C1(n19533), .C2(n19477), .A(n19465), .B(n19464), .ZN(
        P2_U3140) );
  AOI22_X1 U22472 ( .A1(n19472), .A2(n19643), .B1(n19642), .B2(n19471), .ZN(
        n19468) );
  AOI22_X1 U22473 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19474), .B1(
        n19466), .B2(n19579), .ZN(n19467) );
  OAI211_X1 U22474 ( .C1(n19577), .C2(n19508), .A(n19468), .B(n19467), .ZN(
        P2_U3141) );
  AOI22_X1 U22475 ( .A1(n19472), .A2(n19649), .B1(n19648), .B2(n19471), .ZN(
        n19470) );
  AOI22_X1 U22476 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19474), .B1(
        n19473), .B2(n19650), .ZN(n19469) );
  OAI211_X1 U22477 ( .C1(n19653), .C2(n19477), .A(n19470), .B(n19469), .ZN(
        P2_U3142) );
  AOI22_X1 U22478 ( .A1(n19472), .A2(n19656), .B1(n19655), .B2(n19471), .ZN(
        n19476) );
  AOI22_X1 U22479 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19474), .B1(
        n19473), .B2(n19658), .ZN(n19475) );
  OAI211_X1 U22480 ( .C1(n19664), .C2(n19477), .A(n19476), .B(n19475), .ZN(
        P2_U3143) );
  NAND3_X1 U22481 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19788), .ZN(n19511) );
  NOR2_X1 U22482 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19511), .ZN(
        n19502) );
  NOR3_X1 U22483 ( .A1(n11138), .A2(n19502), .A3(n19665), .ZN(n19483) );
  INV_X1 U22484 ( .A(n19478), .ZN(n19480) );
  NOR2_X1 U22485 ( .A1(n19480), .A2(n19479), .ZN(n19487) );
  AOI21_X1 U22486 ( .B1(n19487), .B2(n19611), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19481) );
  NOR2_X1 U22487 ( .A1(n19483), .A2(n19481), .ZN(n19503) );
  AOI22_X1 U22488 ( .A1(n19503), .A2(n19602), .B1(n19601), .B2(n19502), .ZN(
        n19489) );
  AOI21_X1 U22489 ( .B1(n19508), .B2(n19542), .A(n19544), .ZN(n19486) );
  INV_X1 U22490 ( .A(n19502), .ZN(n19484) );
  AOI211_X1 U22491 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19484), .A(n19549), 
        .B(n19483), .ZN(n19485) );
  AOI22_X1 U22492 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19505), .B1(
        n19504), .B2(n19517), .ZN(n19488) );
  OAI211_X1 U22493 ( .C1(n19520), .C2(n19508), .A(n19489), .B(n19488), .ZN(
        P2_U3144) );
  AOI22_X1 U22494 ( .A1(n19503), .A2(n19617), .B1(n19616), .B2(n19502), .ZN(
        n19491) );
  AOI22_X1 U22495 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19505), .B1(
        n19504), .B2(n19521), .ZN(n19490) );
  OAI211_X1 U22496 ( .C1(n19524), .C2(n19508), .A(n19491), .B(n19490), .ZN(
        P2_U3145) );
  AOI22_X1 U22497 ( .A1(n19503), .A2(n19623), .B1(n19622), .B2(n19502), .ZN(
        n19493) );
  AOI22_X1 U22498 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19505), .B1(
        n19504), .B2(n19563), .ZN(n19492) );
  OAI211_X1 U22499 ( .C1(n19527), .C2(n19508), .A(n19493), .B(n19492), .ZN(
        P2_U3146) );
  AOI22_X1 U22500 ( .A1(n19503), .A2(n19629), .B1(n19628), .B2(n19502), .ZN(
        n19495) );
  AOI22_X1 U22501 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19505), .B1(
        n19504), .B2(n19630), .ZN(n19494) );
  OAI211_X1 U22502 ( .C1(n19633), .C2(n19508), .A(n19495), .B(n19494), .ZN(
        P2_U3147) );
  AOI22_X1 U22503 ( .A1(n19503), .A2(n19635), .B1(n19634), .B2(n19502), .ZN(
        n19497) );
  AOI22_X1 U22504 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19505), .B1(
        n19504), .B2(n19530), .ZN(n19496) );
  OAI211_X1 U22505 ( .C1(n19533), .C2(n19508), .A(n19497), .B(n19496), .ZN(
        P2_U3148) );
  AOI22_X1 U22506 ( .A1(n19503), .A2(n19643), .B1(n19642), .B2(n19502), .ZN(
        n19499) );
  AOI22_X1 U22507 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19505), .B1(
        n19504), .B2(n19644), .ZN(n19498) );
  OAI211_X1 U22508 ( .C1(n19647), .C2(n19508), .A(n19499), .B(n19498), .ZN(
        P2_U3149) );
  AOI22_X1 U22509 ( .A1(n19503), .A2(n19649), .B1(n19648), .B2(n19502), .ZN(
        n19501) );
  AOI22_X1 U22510 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19505), .B1(
        n19504), .B2(n19650), .ZN(n19500) );
  OAI211_X1 U22511 ( .C1(n19653), .C2(n19508), .A(n19501), .B(n19500), .ZN(
        P2_U3150) );
  AOI22_X1 U22512 ( .A1(n19503), .A2(n19656), .B1(n19655), .B2(n19502), .ZN(
        n19507) );
  AOI22_X1 U22513 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19505), .B1(
        n19504), .B2(n19658), .ZN(n19506) );
  OAI211_X1 U22514 ( .C1(n19664), .C2(n19508), .A(n19507), .B(n19506), .ZN(
        P2_U3151) );
  NOR2_X1 U22515 ( .A1(n19797), .A2(n19511), .ZN(n19547) );
  INV_X1 U22516 ( .A(n19547), .ZN(n19509) );
  NAND3_X1 U22517 ( .A1(n11086), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19509), 
        .ZN(n19512) );
  OAI21_X1 U22518 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19511), .A(n19665), 
        .ZN(n19510) );
  AOI22_X1 U22519 ( .A1(n19538), .A2(n19602), .B1(n19601), .B2(n19547), .ZN(
        n19519) );
  NOR3_X1 U22520 ( .A1(n19603), .A2(P2_STATE2_REG_3__SCAN_IN), .A3(n19515), 
        .ZN(n19514) );
  AOI21_X1 U22521 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19797), .A(n19511), 
        .ZN(n19513) );
  OAI211_X1 U22522 ( .C1(n19514), .C2(n19513), .A(n19609), .B(n19512), .ZN(
        n19539) );
  NOR2_X2 U22523 ( .A1(n19516), .A2(n19515), .ZN(n19593) );
  AOI22_X1 U22524 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19539), .B1(
        n19593), .B2(n19517), .ZN(n19518) );
  OAI211_X1 U22525 ( .C1(n19520), .C2(n19542), .A(n19519), .B(n19518), .ZN(
        P2_U3152) );
  AOI22_X1 U22526 ( .A1(n19538), .A2(n19617), .B1(n19616), .B2(n19547), .ZN(
        n19523) );
  AOI22_X1 U22527 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19539), .B1(
        n19593), .B2(n19521), .ZN(n19522) );
  OAI211_X1 U22528 ( .C1(n19524), .C2(n19542), .A(n19523), .B(n19522), .ZN(
        P2_U3153) );
  AOI22_X1 U22529 ( .A1(n19538), .A2(n19623), .B1(n19622), .B2(n19547), .ZN(
        n19526) );
  AOI22_X1 U22530 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19539), .B1(
        n19593), .B2(n19563), .ZN(n19525) );
  OAI211_X1 U22531 ( .C1(n19527), .C2(n19542), .A(n19526), .B(n19525), .ZN(
        P2_U3154) );
  AOI22_X1 U22532 ( .A1(n19538), .A2(n19629), .B1(n19628), .B2(n19547), .ZN(
        n19529) );
  AOI22_X1 U22533 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19539), .B1(
        n19593), .B2(n19630), .ZN(n19528) );
  OAI211_X1 U22534 ( .C1(n19633), .C2(n19542), .A(n19529), .B(n19528), .ZN(
        P2_U3155) );
  AOI22_X1 U22535 ( .A1(n19538), .A2(n19635), .B1(n19634), .B2(n19547), .ZN(
        n19532) );
  AOI22_X1 U22536 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19539), .B1(
        n19593), .B2(n19530), .ZN(n19531) );
  OAI211_X1 U22537 ( .C1(n19533), .C2(n19542), .A(n19532), .B(n19531), .ZN(
        P2_U3156) );
  AOI22_X1 U22538 ( .A1(n19538), .A2(n19643), .B1(n19642), .B2(n19547), .ZN(
        n19535) );
  AOI22_X1 U22539 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19539), .B1(
        n19593), .B2(n19644), .ZN(n19534) );
  OAI211_X1 U22540 ( .C1(n19647), .C2(n19542), .A(n19535), .B(n19534), .ZN(
        P2_U3157) );
  AOI22_X1 U22541 ( .A1(n19538), .A2(n19649), .B1(n19648), .B2(n19547), .ZN(
        n19537) );
  AOI22_X1 U22542 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19539), .B1(
        n19593), .B2(n19650), .ZN(n19536) );
  OAI211_X1 U22543 ( .C1(n19653), .C2(n19542), .A(n19537), .B(n19536), .ZN(
        P2_U3158) );
  AOI22_X1 U22544 ( .A1(n19538), .A2(n19656), .B1(n19655), .B2(n19547), .ZN(
        n19541) );
  AOI22_X1 U22545 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19539), .B1(
        n19593), .B2(n19658), .ZN(n19540) );
  OAI211_X1 U22546 ( .C1(n19664), .C2(n19542), .A(n19541), .B(n19540), .ZN(
        P2_U3159) );
  INV_X1 U22547 ( .A(n19593), .ZN(n19545) );
  AOI21_X1 U22548 ( .B1(n19545), .B2(n19663), .A(n19544), .ZN(n19546) );
  NOR2_X1 U22549 ( .A1(n19546), .A2(n19763), .ZN(n19552) );
  NOR2_X1 U22550 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19607), .ZN(
        n19591) );
  NOR2_X1 U22551 ( .A1(n19591), .A2(n19547), .ZN(n19554) );
  AOI211_X1 U22552 ( .C1(n11119), .C2(n19611), .A(n19591), .B(n19759), .ZN(
        n19548) );
  AOI211_X2 U22553 ( .C1(n19552), .C2(n19554), .A(n19549), .B(n19548), .ZN(
        n19598) );
  INV_X1 U22554 ( .A(n19591), .ZN(n19583) );
  OAI22_X1 U22555 ( .A1(n19663), .A2(n19615), .B1(n19550), .B2(n19583), .ZN(
        n19551) );
  INV_X1 U22556 ( .A(n19551), .ZN(n19557) );
  INV_X1 U22557 ( .A(n19552), .ZN(n19555) );
  OAI21_X1 U22558 ( .B1(n11119), .B2(n19591), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19553) );
  AOI22_X1 U22559 ( .A1(n19602), .A2(n19594), .B1(n19593), .B2(n19612), .ZN(
        n19556) );
  OAI211_X1 U22560 ( .C1(n19598), .C2(n19558), .A(n19557), .B(n19556), .ZN(
        P2_U3160) );
  OAI22_X1 U22561 ( .A1(n19663), .A2(n19621), .B1(n19559), .B2(n19583), .ZN(
        n19560) );
  INV_X1 U22562 ( .A(n19560), .ZN(n19562) );
  AOI22_X1 U22563 ( .A1(n19617), .A2(n19594), .B1(n19593), .B2(n19618), .ZN(
        n19561) );
  OAI211_X1 U22564 ( .C1(n19598), .C2(n11108), .A(n19562), .B(n19561), .ZN(
        P2_U3161) );
  INV_X1 U22565 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n19566) );
  AOI22_X1 U22566 ( .A1(n19593), .A2(n19624), .B1(n19622), .B2(n19591), .ZN(
        n19565) );
  AOI22_X1 U22567 ( .A1(n19623), .A2(n19594), .B1(n19637), .B2(n19563), .ZN(
        n19564) );
  OAI211_X1 U22568 ( .C1(n19598), .C2(n19566), .A(n19565), .B(n19564), .ZN(
        P2_U3162) );
  INV_X1 U22569 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n19570) );
  AOI22_X1 U22570 ( .A1(n19593), .A2(n19567), .B1(n19628), .B2(n19591), .ZN(
        n19569) );
  AOI22_X1 U22571 ( .A1(n19629), .A2(n19594), .B1(n19637), .B2(n19630), .ZN(
        n19568) );
  OAI211_X1 U22572 ( .C1(n19598), .C2(n19570), .A(n19569), .B(n19568), .ZN(
        P2_U3163) );
  INV_X1 U22573 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n19575) );
  OAI22_X1 U22574 ( .A1(n19663), .A2(n19641), .B1(n19571), .B2(n19583), .ZN(
        n19572) );
  INV_X1 U22575 ( .A(n19572), .ZN(n19574) );
  AOI22_X1 U22576 ( .A1(n19635), .A2(n19594), .B1(n19593), .B2(n19636), .ZN(
        n19573) );
  OAI211_X1 U22577 ( .C1(n19598), .C2(n19575), .A(n19574), .B(n19573), .ZN(
        P2_U3164) );
  INV_X1 U22578 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n19582) );
  OAI22_X1 U22579 ( .A1(n19663), .A2(n19577), .B1(n19576), .B2(n19583), .ZN(
        n19578) );
  INV_X1 U22580 ( .A(n19578), .ZN(n19581) );
  AOI22_X1 U22581 ( .A1(n19643), .A2(n19594), .B1(n19593), .B2(n19579), .ZN(
        n19580) );
  OAI211_X1 U22582 ( .C1(n19598), .C2(n19582), .A(n19581), .B(n19580), .ZN(
        P2_U3165) );
  INV_X1 U22583 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n19590) );
  OAI22_X1 U22584 ( .A1(n19663), .A2(n19585), .B1(n19584), .B2(n19583), .ZN(
        n19586) );
  INV_X1 U22585 ( .A(n19586), .ZN(n19589) );
  AOI22_X1 U22586 ( .A1(n19649), .A2(n19594), .B1(n19593), .B2(n19587), .ZN(
        n19588) );
  OAI211_X1 U22587 ( .C1(n19598), .C2(n19590), .A(n19589), .B(n19588), .ZN(
        P2_U3166) );
  INV_X1 U22588 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n19597) );
  AOI22_X1 U22589 ( .A1(n19593), .A2(n19592), .B1(n19655), .B2(n19591), .ZN(
        n19596) );
  AOI22_X1 U22590 ( .A1(n19656), .A2(n19594), .B1(n19637), .B2(n19658), .ZN(
        n19595) );
  OAI211_X1 U22591 ( .C1(n19598), .C2(n19597), .A(n19596), .B(n19595), .ZN(
        P2_U3167) );
  NOR3_X1 U22592 ( .A1(n11128), .A2(n19654), .A3(n19665), .ZN(n19606) );
  INV_X1 U22593 ( .A(n19607), .ZN(n19599) );
  AOI21_X1 U22594 ( .B1(n19611), .B2(n19599), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19600) );
  NOR2_X1 U22595 ( .A1(n19606), .A2(n19600), .ZN(n19657) );
  AOI22_X1 U22596 ( .A1(n19657), .A2(n19602), .B1(n19601), .B2(n19654), .ZN(
        n19614) );
  INV_X1 U22597 ( .A(n19603), .ZN(n19605) );
  NAND2_X1 U22598 ( .A1(n19605), .A2(n19604), .ZN(n19608) );
  AOI21_X1 U22599 ( .B1(n19608), .B2(n19607), .A(n19606), .ZN(n19610) );
  OAI211_X1 U22600 ( .C1(n19654), .C2(n19611), .A(n19610), .B(n19609), .ZN(
        n19660) );
  AOI22_X1 U22601 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19660), .B1(
        n19637), .B2(n19612), .ZN(n19613) );
  OAI211_X1 U22602 ( .C1(n19615), .C2(n19640), .A(n19614), .B(n19613), .ZN(
        P2_U3168) );
  AOI22_X1 U22603 ( .A1(n19657), .A2(n19617), .B1(n19616), .B2(n19654), .ZN(
        n19620) );
  AOI22_X1 U22604 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19660), .B1(
        n19637), .B2(n19618), .ZN(n19619) );
  OAI211_X1 U22605 ( .C1(n19621), .C2(n19640), .A(n19620), .B(n19619), .ZN(
        P2_U3169) );
  AOI22_X1 U22606 ( .A1(n19657), .A2(n19623), .B1(n19622), .B2(n19654), .ZN(
        n19626) );
  AOI22_X1 U22607 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19660), .B1(
        n19637), .B2(n19624), .ZN(n19625) );
  OAI211_X1 U22608 ( .C1(n19627), .C2(n19640), .A(n19626), .B(n19625), .ZN(
        P2_U3170) );
  AOI22_X1 U22609 ( .A1(n19657), .A2(n19629), .B1(n19628), .B2(n19654), .ZN(
        n19632) );
  AOI22_X1 U22610 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19660), .B1(
        n19659), .B2(n19630), .ZN(n19631) );
  OAI211_X1 U22611 ( .C1(n19633), .C2(n19663), .A(n19632), .B(n19631), .ZN(
        P2_U3171) );
  AOI22_X1 U22612 ( .A1(n19657), .A2(n19635), .B1(n19634), .B2(n19654), .ZN(
        n19639) );
  AOI22_X1 U22613 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19660), .B1(
        n19637), .B2(n19636), .ZN(n19638) );
  OAI211_X1 U22614 ( .C1(n19641), .C2(n19640), .A(n19639), .B(n19638), .ZN(
        P2_U3172) );
  AOI22_X1 U22615 ( .A1(n19657), .A2(n19643), .B1(n19642), .B2(n19654), .ZN(
        n19646) );
  AOI22_X1 U22616 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19660), .B1(
        n19659), .B2(n19644), .ZN(n19645) );
  OAI211_X1 U22617 ( .C1(n19647), .C2(n19663), .A(n19646), .B(n19645), .ZN(
        P2_U3173) );
  AOI22_X1 U22618 ( .A1(n19657), .A2(n19649), .B1(n19648), .B2(n19654), .ZN(
        n19652) );
  AOI22_X1 U22619 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19660), .B1(
        n19659), .B2(n19650), .ZN(n19651) );
  OAI211_X1 U22620 ( .C1(n19653), .C2(n19663), .A(n19652), .B(n19651), .ZN(
        P2_U3174) );
  AOI22_X1 U22621 ( .A1(n19657), .A2(n19656), .B1(n19655), .B2(n19654), .ZN(
        n19662) );
  AOI22_X1 U22622 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19660), .B1(
        n19659), .B2(n19658), .ZN(n19661) );
  OAI211_X1 U22623 ( .C1(n19664), .C2(n19663), .A(n19662), .B(n19661), .ZN(
        P2_U3175) );
  OAI22_X1 U22624 ( .A1(n19666), .A2(n19690), .B1(n19665), .B2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19675) );
  INV_X1 U22625 ( .A(n19667), .ZN(n19671) );
  AOI211_X1 U22626 ( .C1(n19671), .C2(n19670), .A(n19669), .B(n19668), .ZN(
        n19672) );
  AOI211_X1 U22627 ( .C1(n19675), .C2(n19674), .A(n19673), .B(n19672), .ZN(
        n19676) );
  INV_X1 U22628 ( .A(n19676), .ZN(P2_U3177) );
  INV_X1 U22629 ( .A(n19756), .ZN(n19677) );
  AND2_X1 U22630 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19677), .ZN(
        P2_U3179) );
  AND2_X1 U22631 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19677), .ZN(
        P2_U3180) );
  AND2_X1 U22632 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19677), .ZN(
        P2_U3181) );
  AND2_X1 U22633 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19677), .ZN(
        P2_U3182) );
  AND2_X1 U22634 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19677), .ZN(
        P2_U3183) );
  AND2_X1 U22635 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19677), .ZN(
        P2_U3184) );
  AND2_X1 U22636 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19677), .ZN(
        P2_U3185) );
  AND2_X1 U22637 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19677), .ZN(
        P2_U3186) );
  AND2_X1 U22638 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19677), .ZN(
        P2_U3187) );
  AND2_X1 U22639 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19677), .ZN(
        P2_U3188) );
  AND2_X1 U22640 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19677), .ZN(
        P2_U3189) );
  AND2_X1 U22641 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19677), .ZN(
        P2_U3190) );
  AND2_X1 U22642 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19677), .ZN(
        P2_U3191) );
  AND2_X1 U22643 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19677), .ZN(
        P2_U3192) );
  AND2_X1 U22644 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19677), .ZN(
        P2_U3193) );
  AND2_X1 U22645 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19677), .ZN(
        P2_U3194) );
  AND2_X1 U22646 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19677), .ZN(
        P2_U3195) );
  INV_X1 U22647 ( .A(P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20928) );
  NOR2_X1 U22648 ( .A1(n20928), .A2(n19756), .ZN(P2_U3196) );
  AND2_X1 U22649 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19677), .ZN(
        P2_U3197) );
  AND2_X1 U22650 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19677), .ZN(
        P2_U3198) );
  AND2_X1 U22651 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19677), .ZN(
        P2_U3199) );
  AND2_X1 U22652 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19677), .ZN(
        P2_U3200) );
  AND2_X1 U22653 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19677), .ZN(P2_U3201) );
  AND2_X1 U22654 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19677), .ZN(P2_U3202) );
  AND2_X1 U22655 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19677), .ZN(P2_U3203) );
  AND2_X1 U22656 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19677), .ZN(P2_U3204) );
  AND2_X1 U22657 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19677), .ZN(P2_U3205) );
  AND2_X1 U22658 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19677), .ZN(P2_U3206) );
  AND2_X1 U22659 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19677), .ZN(P2_U3207) );
  AND2_X1 U22660 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19677), .ZN(P2_U3208) );
  NAND2_X1 U22661 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19690), .ZN(n19692) );
  NAND3_X1 U22662 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n19692), .ZN(n19679) );
  AOI211_X1 U22663 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n19687), .A(
        n19691), .B(n19744), .ZN(n19678) );
  NOR2_X1 U22664 ( .A1(n20697), .A2(n19683), .ZN(n19697) );
  AOI211_X1 U22665 ( .C1(n19698), .C2(n19679), .A(n19678), .B(n19697), .ZN(
        n19680) );
  INV_X1 U22666 ( .A(n19680), .ZN(P2_U3209) );
  INV_X1 U22667 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19681) );
  AOI21_X1 U22668 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n19687), .A(n19698), 
        .ZN(n19688) );
  NOR2_X1 U22669 ( .A1(n19681), .A2(n19688), .ZN(n19684) );
  AOI21_X1 U22670 ( .B1(n19684), .B2(n19683), .A(n19682), .ZN(n19685) );
  OAI211_X1 U22671 ( .C1(n19687), .C2(n19686), .A(n19685), .B(n19692), .ZN(
        P2_U3210) );
  AOI21_X1 U22672 ( .B1(n19690), .B2(n19689), .A(n19688), .ZN(n19696) );
  INV_X1 U22673 ( .A(n19691), .ZN(n19693) );
  OAI22_X1 U22674 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19693), .B1(NA), 
        .B2(n19692), .ZN(n19694) );
  OAI211_X1 U22675 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19694), .ZN(n19695) );
  OAI21_X1 U22676 ( .B1(n19697), .B2(n19696), .A(n19695), .ZN(P2_U3211) );
  NAND2_X1 U22677 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19744), .ZN(n19746) );
  CLKBUF_X1 U22678 ( .A(n19746), .Z(n19742) );
  OAI222_X1 U22679 ( .A1(n19749), .A2(n19701), .B1(n19700), .B2(n19744), .C1(
        n19699), .C2(n19742), .ZN(P2_U3212) );
  OAI222_X1 U22680 ( .A1(n19749), .A2(n13657), .B1(n19702), .B2(n19744), .C1(
        n19701), .C2(n19742), .ZN(P2_U3213) );
  OAI222_X1 U22681 ( .A1(n19749), .A2(n10317), .B1(n19703), .B2(n19744), .C1(
        n13657), .C2(n19742), .ZN(P2_U3214) );
  OAI222_X1 U22682 ( .A1(n19742), .A2(n10317), .B1(n19704), .B2(n19744), .C1(
        n13861), .C2(n19749), .ZN(P2_U3215) );
  OAI222_X1 U22683 ( .A1(n19742), .A2(n13861), .B1(n19705), .B2(n19744), .C1(
        n19707), .C2(n19749), .ZN(P2_U3216) );
  OAI222_X1 U22684 ( .A1(n19746), .A2(n19707), .B1(n19706), .B2(n19744), .C1(
        n19709), .C2(n19749), .ZN(P2_U3217) );
  OAI222_X1 U22685 ( .A1(n19746), .A2(n19709), .B1(n19708), .B2(n19744), .C1(
        n10339), .C2(n19749), .ZN(P2_U3218) );
  OAI222_X1 U22686 ( .A1(n19746), .A2(n10339), .B1(n19710), .B2(n19744), .C1(
        n19712), .C2(n19749), .ZN(P2_U3219) );
  OAI222_X1 U22687 ( .A1(n19742), .A2(n19712), .B1(n19711), .B2(n19744), .C1(
        n10365), .C2(n19749), .ZN(P2_U3220) );
  OAI222_X1 U22688 ( .A1(n19746), .A2(n10365), .B1(n19713), .B2(n19744), .C1(
        n19715), .C2(n19749), .ZN(P2_U3221) );
  OAI222_X1 U22689 ( .A1(n19746), .A2(n19715), .B1(n19714), .B2(n19744), .C1(
        n10397), .C2(n19749), .ZN(P2_U3222) );
  OAI222_X1 U22690 ( .A1(n19746), .A2(n10397), .B1(n20831), .B2(n19744), .C1(
        n19716), .C2(n19749), .ZN(P2_U3223) );
  OAI222_X1 U22691 ( .A1(n19749), .A2(n10423), .B1(n20921), .B2(n19744), .C1(
        n19716), .C2(n19742), .ZN(P2_U3224) );
  OAI222_X1 U22692 ( .A1(n19749), .A2(n19717), .B1(n20832), .B2(n19744), .C1(
        n10423), .C2(n19742), .ZN(P2_U3225) );
  OAI222_X1 U22693 ( .A1(n19749), .A2(n19719), .B1(n19718), .B2(n19744), .C1(
        n19717), .C2(n19746), .ZN(P2_U3226) );
  OAI222_X1 U22694 ( .A1(n19749), .A2(n19721), .B1(n19720), .B2(n19744), .C1(
        n19719), .C2(n19746), .ZN(P2_U3227) );
  OAI222_X1 U22695 ( .A1(n19749), .A2(n19723), .B1(n19722), .B2(n19744), .C1(
        n19721), .C2(n19746), .ZN(P2_U3228) );
  OAI222_X1 U22696 ( .A1(n19749), .A2(n19725), .B1(n19724), .B2(n19744), .C1(
        n19723), .C2(n19742), .ZN(P2_U3229) );
  OAI222_X1 U22697 ( .A1(n19749), .A2(n10452), .B1(n19726), .B2(n19744), .C1(
        n19725), .C2(n19742), .ZN(P2_U3230) );
  OAI222_X1 U22698 ( .A1(n19749), .A2(n19728), .B1(n19727), .B2(n19744), .C1(
        n10452), .C2(n19742), .ZN(P2_U3231) );
  OAI222_X1 U22699 ( .A1(n19749), .A2(n19729), .B1(n20924), .B2(n19744), .C1(
        n19728), .C2(n19742), .ZN(P2_U3232) );
  OAI222_X1 U22700 ( .A1(n19749), .A2(n19731), .B1(n19730), .B2(n19744), .C1(
        n19729), .C2(n19742), .ZN(P2_U3233) );
  OAI222_X1 U22701 ( .A1(n19749), .A2(n19733), .B1(n19732), .B2(n19744), .C1(
        n19731), .C2(n19742), .ZN(P2_U3234) );
  OAI222_X1 U22702 ( .A1(n19749), .A2(n19735), .B1(n19734), .B2(n19744), .C1(
        n19733), .C2(n19742), .ZN(P2_U3235) );
  OAI222_X1 U22703 ( .A1(n19749), .A2(n14961), .B1(n19736), .B2(n19744), .C1(
        n19735), .C2(n19742), .ZN(P2_U3236) );
  OAI222_X1 U22704 ( .A1(n19749), .A2(n19739), .B1(n19737), .B2(n19744), .C1(
        n14961), .C2(n19742), .ZN(P2_U3237) );
  OAI222_X1 U22705 ( .A1(n19746), .A2(n19739), .B1(n19738), .B2(n19744), .C1(
        n19740), .C2(n19749), .ZN(P2_U3238) );
  OAI222_X1 U22706 ( .A1(n19749), .A2(n19743), .B1(n19741), .B2(n19744), .C1(
        n19740), .C2(n19742), .ZN(P2_U3239) );
  OAI222_X1 U22707 ( .A1(n19749), .A2(n14146), .B1(n19745), .B2(n19744), .C1(
        n19743), .C2(n19742), .ZN(P2_U3240) );
  INV_X1 U22708 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19748) );
  OAI222_X1 U22709 ( .A1(n19749), .A2(n19748), .B1(n19747), .B2(n19744), .C1(
        n14146), .C2(n19746), .ZN(P2_U3241) );
  AOI22_X1 U22710 ( .A1(n19744), .A2(n19750), .B1(n20925), .B2(n19810), .ZN(
        P2_U3585) );
  MUX2_X1 U22711 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n19810), .Z(P2_U3586) );
  OAI22_X1 U22712 ( .A1(n19810), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19744), .ZN(n19751) );
  INV_X1 U22713 ( .A(n19751), .ZN(P2_U3587) );
  OAI22_X1 U22714 ( .A1(n19810), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19744), .ZN(n19752) );
  INV_X1 U22715 ( .A(n19752), .ZN(P2_U3588) );
  OAI21_X1 U22716 ( .B1(n19756), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19754), 
        .ZN(n19753) );
  INV_X1 U22717 ( .A(n19753), .ZN(P2_U3591) );
  OAI21_X1 U22718 ( .B1(n19756), .B2(n19755), .A(n19754), .ZN(P2_U3592) );
  INV_X1 U22719 ( .A(n19796), .ZN(n19795) );
  AND2_X1 U22720 ( .A1(n19759), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19784) );
  NAND2_X1 U22721 ( .A1(n19757), .A2(n19784), .ZN(n19773) );
  NAND2_X1 U22722 ( .A1(n19782), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19760) );
  AOI21_X1 U22723 ( .B1(n19760), .B2(n19759), .A(n19758), .ZN(n19771) );
  AOI21_X1 U22724 ( .B1(n19773), .B2(n19771), .A(n19761), .ZN(n19766) );
  NOR3_X1 U22725 ( .A1(n19764), .A2(n19763), .A3(n19762), .ZN(n19765) );
  AOI211_X1 U22726 ( .C1(n19767), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19766), 
        .B(n19765), .ZN(n19768) );
  AOI22_X1 U22727 ( .A1(n19795), .A2(n19769), .B1(n19768), .B2(n19796), .ZN(
        P2_U3602) );
  INV_X1 U22728 ( .A(n19770), .ZN(n19777) );
  INV_X1 U22729 ( .A(n19771), .ZN(n19776) );
  NOR2_X1 U22730 ( .A1(n19772), .A2(n19611), .ZN(n19775) );
  INV_X1 U22731 ( .A(n19773), .ZN(n19774) );
  AOI211_X1 U22732 ( .C1(n19777), .C2(n19776), .A(n19775), .B(n19774), .ZN(
        n19778) );
  AOI22_X1 U22733 ( .A1(n19795), .A2(n19779), .B1(n19778), .B2(n19796), .ZN(
        P2_U3603) );
  INV_X1 U22734 ( .A(n19780), .ZN(n19791) );
  AND2_X1 U22735 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19781) );
  NOR2_X1 U22736 ( .A1(n19791), .A2(n19781), .ZN(n19783) );
  MUX2_X1 U22737 ( .A(n19784), .B(n19783), .S(n19782), .Z(n19785) );
  AOI21_X1 U22738 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19786), .A(n19785), 
        .ZN(n19787) );
  AOI22_X1 U22739 ( .A1(n19795), .A2(n19788), .B1(n19787), .B2(n19796), .ZN(
        P2_U3604) );
  NAND3_X1 U22740 ( .A1(n19789), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19790) );
  OAI21_X1 U22741 ( .B1(n19792), .B2(n19791), .A(n19790), .ZN(n19793) );
  AOI21_X1 U22742 ( .B1(n19797), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19793), 
        .ZN(n19794) );
  OAI22_X1 U22743 ( .A1(n19797), .A2(n19796), .B1(n19795), .B2(n19794), .ZN(
        P2_U3605) );
  AOI22_X1 U22744 ( .A1(n19744), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19798), 
        .B2(n19810), .ZN(P2_U3608) );
  AOI22_X1 U22745 ( .A1(n19802), .A2(n19801), .B1(n19800), .B2(n19799), .ZN(
        n19806) );
  INV_X1 U22746 ( .A(n19803), .ZN(n19804) );
  OAI21_X1 U22747 ( .B1(n19806), .B2(n19805), .A(n19804), .ZN(n19808) );
  MUX2_X1 U22748 ( .A(P2_MORE_REG_SCAN_IN), .B(n19808), .S(n19807), .Z(
        P2_U3609) );
  OAI22_X1 U22749 ( .A1(n19810), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19744), .ZN(n19811) );
  INV_X1 U22750 ( .A(n19811), .ZN(P2_U3611) );
  AOI21_X1 U22751 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20702), .A(n19812), 
        .ZN(n19820) );
  INV_X1 U22752 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19813) );
  NAND2_X1 U22753 ( .A1(n19812), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20738) );
  AOI21_X1 U22754 ( .B1(n19820), .B2(n19813), .A(n20795), .ZN(P1_U2802) );
  INV_X1 U22755 ( .A(n19814), .ZN(n19816) );
  OAI21_X1 U22756 ( .B1(n19816), .B2(n19815), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19817) );
  OAI21_X1 U22757 ( .B1(n19818), .B2(n20071), .A(n19817), .ZN(P1_U2803) );
  INV_X1 U22758 ( .A(n20738), .ZN(n20795) );
  INV_X1 U22759 ( .A(n20795), .ZN(n20796) );
  NOR2_X1 U22760 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19821) );
  OAI21_X1 U22761 ( .B1(n19821), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20796), .ZN(
        n19819) );
  OAI21_X1 U22762 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20796), .A(n19819), 
        .ZN(P1_U2804) );
  NOR2_X1 U22763 ( .A1(n20795), .A2(n19820), .ZN(n20755) );
  OAI21_X1 U22764 ( .B1(BS16), .B2(n19821), .A(n20755), .ZN(n20753) );
  OAI21_X1 U22765 ( .B1(n20755), .B2(n20578), .A(n20753), .ZN(P1_U2805) );
  OAI21_X1 U22766 ( .B1(n19824), .B2(n19823), .A(n19822), .ZN(P1_U2806) );
  NOR4_X1 U22767 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19828) );
  NOR4_X1 U22768 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19827) );
  NOR4_X1 U22769 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19826) );
  NOR4_X1 U22770 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19825) );
  NAND4_X1 U22771 ( .A1(n19828), .A2(n19827), .A3(n19826), .A4(n19825), .ZN(
        n19834) );
  NOR4_X1 U22772 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19832) );
  AOI211_X1 U22773 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_11__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19831) );
  NOR4_X1 U22774 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19830) );
  NOR4_X1 U22775 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19829) );
  NAND4_X1 U22776 ( .A1(n19832), .A2(n19831), .A3(n19830), .A4(n19829), .ZN(
        n19833) );
  NOR2_X1 U22777 ( .A1(n19834), .A2(n19833), .ZN(n20782) );
  INV_X1 U22778 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19836) );
  NOR3_X1 U22779 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19837) );
  OAI21_X1 U22780 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19837), .A(n20782), .ZN(
        n19835) );
  OAI21_X1 U22781 ( .B1(n20782), .B2(n19836), .A(n19835), .ZN(P1_U2807) );
  INV_X1 U22782 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20754) );
  AOI21_X1 U22783 ( .B1(n20775), .B2(n20754), .A(n19837), .ZN(n19839) );
  INV_X1 U22784 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19838) );
  INV_X1 U22785 ( .A(n20782), .ZN(n20777) );
  AOI22_X1 U22786 ( .A1(n20782), .A2(n19839), .B1(n19838), .B2(n20777), .ZN(
        P1_U2808) );
  AOI22_X1 U22787 ( .A1(n9561), .A2(n19841), .B1(n19840), .B2(n20713), .ZN(
        n19849) );
  AOI22_X1 U22788 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n19866), .B1(
        n19842), .B2(n19907), .ZN(n19848) );
  AOI21_X1 U22789 ( .B1(n19876), .B2(P1_EBX_REG_9__SCAN_IN), .A(n19854), .ZN(
        n19847) );
  INV_X1 U22790 ( .A(n19843), .ZN(n19845) );
  AOI22_X1 U22791 ( .A1(n19845), .A2(n19870), .B1(P1_REIP_REG_9__SCAN_IN), 
        .B2(n19844), .ZN(n19846) );
  NAND4_X1 U22792 ( .A1(n19849), .A2(n19848), .A3(n19847), .A4(n19846), .ZN(
        P1_U2831) );
  AOI21_X1 U22793 ( .B1(n19882), .B2(n19864), .A(n19850), .ZN(n19874) );
  NAND2_X1 U22794 ( .A1(n19851), .A2(n19870), .ZN(n19861) );
  NOR3_X1 U22795 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19852), .A3(n19864), .ZN(
        n19853) );
  AOI211_X1 U22796 ( .C1(n19866), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n19854), .B(n19853), .ZN(n19860) );
  INV_X1 U22797 ( .A(n19855), .ZN(n19856) );
  AOI22_X1 U22798 ( .A1(n19876), .A2(P1_EBX_REG_7__SCAN_IN), .B1(n19856), .B2(
        n19907), .ZN(n19859) );
  NAND2_X1 U22799 ( .A1(n19857), .A2(n9561), .ZN(n19858) );
  AND4_X1 U22800 ( .A1(n19861), .A2(n19860), .A3(n19859), .A4(n19858), .ZN(
        n19862) );
  OAI21_X1 U22801 ( .B1(n19874), .B2(n20710), .A(n19862), .ZN(P1_U2833) );
  INV_X1 U22802 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n19873) );
  AND3_X1 U22803 ( .A1(n19882), .A2(n19864), .A3(n19863), .ZN(n19865) );
  AOI21_X1 U22804 ( .B1(n19876), .B2(P1_EBX_REG_6__SCAN_IN), .A(n19865), .ZN(
        n19872) );
  AOI22_X1 U22805 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n19866), .B1(
        n9561), .B2(n19912), .ZN(n19867) );
  OAI211_X1 U22806 ( .C1(n19890), .C2(n19868), .A(n19867), .B(n19878), .ZN(
        n19869) );
  AOI21_X1 U22807 ( .B1(n19915), .B2(n19870), .A(n19869), .ZN(n19871) );
  OAI211_X1 U22808 ( .C1(n19874), .C2(n19873), .A(n19872), .B(n19871), .ZN(
        P1_U2834) );
  NOR2_X1 U22809 ( .A1(n19875), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n19883) );
  AOI22_X1 U22810 ( .A1(n19877), .A2(n9561), .B1(n19876), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n19879) );
  OAI211_X1 U22811 ( .C1(n19894), .C2(n19880), .A(n19879), .B(n19878), .ZN(
        n19881) );
  AOI21_X1 U22812 ( .B1(n19883), .B2(n19882), .A(n19881), .ZN(n19889) );
  INV_X1 U22813 ( .A(n19884), .ZN(n19887) );
  AOI22_X1 U22814 ( .A1(n19887), .A2(n19886), .B1(n19885), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n19888) );
  OAI211_X1 U22815 ( .C1(n19891), .C2(n19890), .A(n19889), .B(n19888), .ZN(
        P1_U2835) );
  OAI221_X1 U22816 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(P1_REIP_REG_2__SCAN_IN), 
        .C1(P1_REIP_REG_3__SCAN_IN), .C2(n19893), .A(n19892), .ZN(n19910) );
  OAI22_X1 U22817 ( .A1(n19897), .A2(n19896), .B1(n19895), .B2(n19894), .ZN(
        n19901) );
  NOR2_X1 U22818 ( .A1(n19899), .A2(n19898), .ZN(n19900) );
  AOI211_X1 U22819 ( .C1(n9561), .C2(n20010), .A(n19901), .B(n19900), .ZN(
        n19903) );
  OAI21_X1 U22820 ( .B1(n19905), .B2(n19904), .A(n19903), .ZN(n19906) );
  AOI21_X1 U22821 ( .B1(n19908), .B2(n19907), .A(n19906), .ZN(n19909) );
  OAI21_X1 U22822 ( .B1(n19911), .B2(n19910), .A(n19909), .ZN(P1_U2837) );
  AOI22_X1 U22823 ( .A1(n19915), .A2(n19914), .B1(n19913), .B2(n19912), .ZN(
        n19916) );
  OAI21_X1 U22824 ( .B1(n19918), .B2(n19917), .A(n19916), .ZN(P1_U2866) );
  AOI22_X1 U22825 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n19922), .B1(n19945), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19919) );
  OAI21_X1 U22826 ( .B1(n19921), .B2(n19920), .A(n19919), .ZN(P1_U2921) );
  AOI22_X1 U22827 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n19930), .B1(n19945), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19923) );
  OAI21_X1 U22828 ( .B1(n14006), .B2(n19947), .A(n19923), .ZN(P1_U2922) );
  AOI22_X1 U22829 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n19930), .B1(n19945), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19924) );
  OAI21_X1 U22830 ( .B1(n13998), .B2(n19947), .A(n19924), .ZN(P1_U2923) );
  AOI22_X1 U22831 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n19945), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n19930), .ZN(n19925) );
  OAI21_X1 U22832 ( .B1(n13979), .B2(n19947), .A(n19925), .ZN(P1_U2924) );
  AOI22_X1 U22833 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n19930), .B1(n19945), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19926) );
  OAI21_X1 U22834 ( .B1(n14011), .B2(n19947), .A(n19926), .ZN(P1_U2925) );
  AOI22_X1 U22835 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n19930), .B1(n19934), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19927) );
  OAI21_X1 U22836 ( .B1(n13841), .B2(n19947), .A(n19927), .ZN(P1_U2926) );
  AOI22_X1 U22837 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n19930), .B1(n19934), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19928) );
  OAI21_X1 U22838 ( .B1(n13909), .B2(n19947), .A(n19928), .ZN(P1_U2927) );
  AOI22_X1 U22839 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n19930), .B1(n19934), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19929) );
  OAI21_X1 U22840 ( .B1(n13903), .B2(n19947), .A(n19929), .ZN(P1_U2928) );
  AOI22_X1 U22841 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n19945), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n19930), .ZN(n19931) );
  OAI21_X1 U22842 ( .B1(n12212), .B2(n19947), .A(n19931), .ZN(P1_U2929) );
  AOI22_X1 U22843 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n19930), .B1(n19945), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19932) );
  OAI21_X1 U22844 ( .B1(n19933), .B2(n19947), .A(n19932), .ZN(P1_U2930) );
  AOI22_X1 U22845 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n19930), .B1(n19934), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19935) );
  OAI21_X1 U22846 ( .B1(n19936), .B2(n19947), .A(n19935), .ZN(P1_U2931) );
  AOI22_X1 U22847 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n19930), .B1(n19945), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19937) );
  OAI21_X1 U22848 ( .B1(n19938), .B2(n19947), .A(n19937), .ZN(P1_U2932) );
  AOI22_X1 U22849 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n19930), .B1(n19945), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19939) );
  OAI21_X1 U22850 ( .B1(n19940), .B2(n19947), .A(n19939), .ZN(P1_U2933) );
  AOI22_X1 U22851 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n19930), .B1(n19945), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19941) );
  OAI21_X1 U22852 ( .B1(n19942), .B2(n19947), .A(n19941), .ZN(P1_U2934) );
  AOI22_X1 U22853 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n19930), .B1(n19945), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19943) );
  OAI21_X1 U22854 ( .B1(n19944), .B2(n19947), .A(n19943), .ZN(P1_U2935) );
  AOI22_X1 U22855 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n19930), .B1(n19945), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19946) );
  OAI21_X1 U22856 ( .B1(n19948), .B2(n19947), .A(n19946), .ZN(P1_U2936) );
  AOI22_X1 U22857 ( .A1(n19981), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n19974), .ZN(n19951) );
  INV_X1 U22858 ( .A(n19949), .ZN(n19950) );
  NAND2_X1 U22859 ( .A1(n19966), .A2(n19950), .ZN(n19968) );
  NAND2_X1 U22860 ( .A1(n19951), .A2(n19968), .ZN(P1_U2945) );
  AOI22_X1 U22861 ( .A1(n19981), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n19974), .ZN(n19954) );
  INV_X1 U22862 ( .A(n19952), .ZN(n19953) );
  NAND2_X1 U22863 ( .A1(n19966), .A2(n19953), .ZN(n19970) );
  NAND2_X1 U22864 ( .A1(n19954), .A2(n19970), .ZN(P1_U2946) );
  AOI22_X1 U22865 ( .A1(n19981), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n19974), .ZN(n19957) );
  INV_X1 U22866 ( .A(n19955), .ZN(n19956) );
  NAND2_X1 U22867 ( .A1(n19966), .A2(n19956), .ZN(n19972) );
  NAND2_X1 U22868 ( .A1(n19957), .A2(n19972), .ZN(P1_U2947) );
  AOI22_X1 U22869 ( .A1(n19981), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n19974), .ZN(n19960) );
  INV_X1 U22870 ( .A(n19958), .ZN(n19959) );
  NAND2_X1 U22871 ( .A1(n19966), .A2(n19959), .ZN(n19975) );
  NAND2_X1 U22872 ( .A1(n19960), .A2(n19975), .ZN(P1_U2948) );
  AOI22_X1 U22873 ( .A1(n19981), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n19974), .ZN(n19963) );
  INV_X1 U22874 ( .A(n19961), .ZN(n19962) );
  NAND2_X1 U22875 ( .A1(n19966), .A2(n19962), .ZN(n19979) );
  NAND2_X1 U22876 ( .A1(n19963), .A2(n19979), .ZN(P1_U2950) );
  AOI22_X1 U22877 ( .A1(n19981), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n19974), .ZN(n19967) );
  INV_X1 U22878 ( .A(n19964), .ZN(n19965) );
  NAND2_X1 U22879 ( .A1(n19966), .A2(n19965), .ZN(n19982) );
  NAND2_X1 U22880 ( .A1(n19967), .A2(n19982), .ZN(P1_U2951) );
  AOI22_X1 U22881 ( .A1(n19981), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n19974), .ZN(n19969) );
  NAND2_X1 U22882 ( .A1(n19969), .A2(n19968), .ZN(P1_U2960) );
  AOI22_X1 U22883 ( .A1(n19981), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n19974), .ZN(n19971) );
  NAND2_X1 U22884 ( .A1(n19971), .A2(n19970), .ZN(P1_U2961) );
  AOI22_X1 U22885 ( .A1(n19981), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n19974), .ZN(n19973) );
  NAND2_X1 U22886 ( .A1(n19973), .A2(n19972), .ZN(P1_U2962) );
  AOI22_X1 U22887 ( .A1(n19981), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n19974), .ZN(n19976) );
  NAND2_X1 U22888 ( .A1(n19976), .A2(n19975), .ZN(P1_U2963) );
  AOI22_X1 U22889 ( .A1(n19981), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n19974), .ZN(n19978) );
  NAND2_X1 U22890 ( .A1(n19978), .A2(n19977), .ZN(P1_U2964) );
  AOI22_X1 U22891 ( .A1(n19981), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n19974), .ZN(n19980) );
  NAND2_X1 U22892 ( .A1(n19980), .A2(n19979), .ZN(P1_U2965) );
  AOI22_X1 U22893 ( .A1(n19981), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n19974), .ZN(n19983) );
  NAND2_X1 U22894 ( .A1(n19983), .A2(n19982), .ZN(P1_U2966) );
  AOI22_X1 U22895 ( .A1(n19984), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20053), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n19993) );
  OR2_X1 U22896 ( .A1(n19986), .A2(n19985), .ZN(n19987) );
  NAND2_X1 U22897 ( .A1(n19988), .A2(n19987), .ZN(n19999) );
  INV_X1 U22898 ( .A(n19999), .ZN(n19991) );
  AOI22_X1 U22899 ( .A1(n19991), .A2(n19990), .B1(n13319), .B2(n19989), .ZN(
        n19992) );
  OAI211_X1 U22900 ( .C1(n19995), .C2(n19994), .A(n19993), .B(n19992), .ZN(
        P1_U2995) );
  INV_X1 U22901 ( .A(n20020), .ZN(n19997) );
  AOI21_X1 U22902 ( .B1(n20047), .B2(n19997), .A(n19996), .ZN(n20017) );
  AOI211_X1 U22903 ( .C1(n20009), .C2(n20016), .A(n19998), .B(n20012), .ZN(
        n20007) );
  NOR2_X1 U22904 ( .A1(n19999), .A2(n20050), .ZN(n20006) );
  INV_X1 U22905 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20004) );
  INV_X1 U22906 ( .A(n20000), .ZN(n20002) );
  NAND2_X1 U22907 ( .A1(n20002), .A2(n20001), .ZN(n20003) );
  OAI21_X1 U22908 ( .B1(n20004), .B2(n20035), .A(n20003), .ZN(n20005) );
  NOR3_X1 U22909 ( .A1(n20007), .A2(n20006), .A3(n20005), .ZN(n20008) );
  OAI21_X1 U22910 ( .B1(n20017), .B2(n20009), .A(n20008), .ZN(P1_U3027) );
  AOI22_X1 U22911 ( .A1(n20053), .A2(P1_REIP_REG_3__SCAN_IN), .B1(n20042), 
        .B2(n20010), .ZN(n20015) );
  OAI22_X1 U22912 ( .A1(n20012), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20011), .B2(n20050), .ZN(n20013) );
  INV_X1 U22913 ( .A(n20013), .ZN(n20014) );
  OAI211_X1 U22914 ( .C1(n20017), .C2(n20016), .A(n20015), .B(n20014), .ZN(
        P1_U3028) );
  AOI21_X1 U22915 ( .B1(n20044), .B2(n20018), .A(n20033), .ZN(n20028) );
  NOR2_X1 U22916 ( .A1(n20019), .A2(n20050), .ZN(n20026) );
  NAND2_X1 U22917 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20021) );
  OAI21_X1 U22918 ( .B1(n20029), .B2(n20021), .A(n20020), .ZN(n20022) );
  AOI22_X1 U22919 ( .A1(n20047), .A2(n20022), .B1(n20053), .B2(
        P1_REIP_REG_2__SCAN_IN), .ZN(n20023) );
  OAI21_X1 U22920 ( .B1(n20049), .B2(n20024), .A(n20023), .ZN(n20025) );
  AOI21_X1 U22921 ( .B1(n20026), .B2(n13517), .A(n20025), .ZN(n20027) );
  OAI221_X1 U22922 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20030), .C1(
        n20029), .C2(n20028), .A(n20027), .ZN(P1_U3029) );
  NAND2_X1 U22923 ( .A1(n20032), .A2(n20031), .ZN(n20045) );
  AOI21_X1 U22924 ( .B1(n20047), .B2(n20034), .A(n20033), .ZN(n20056) );
  NOR2_X1 U22925 ( .A1(n20035), .A2(n20775), .ZN(n20040) );
  AND3_X1 U22926 ( .A1(n20038), .A2(n20037), .A3(n20036), .ZN(n20039) );
  AOI211_X1 U22927 ( .C1(n20042), .C2(n20041), .A(n20040), .B(n20039), .ZN(
        n20043) );
  OAI221_X1 U22928 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20045), .C1(
        n20044), .C2(n20056), .A(n20043), .ZN(P1_U3030) );
  NOR3_X1 U22929 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20047), .A3(
        n20046), .ZN(n20057) );
  OAI22_X1 U22930 ( .A1(n20051), .A2(n20050), .B1(n20049), .B2(n20048), .ZN(
        n20052) );
  AOI21_X1 U22931 ( .B1(n20053), .B2(P1_REIP_REG_0__SCAN_IN), .A(n20052), .ZN(
        n20054) );
  OAI221_X1 U22932 ( .B1(n20057), .B2(n20056), .C1(n20057), .C2(n20055), .A(
        n20054), .ZN(P1_U3031) );
  NOR2_X1 U22933 ( .A1(n20058), .A2(n20774), .ZN(P1_U3032) );
  INV_X1 U22934 ( .A(n20426), .ZN(n20359) );
  NAND2_X1 U22935 ( .A1(n20358), .A2(n20359), .ZN(n20235) );
  NAND2_X1 U22936 ( .A1(n20075), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20574) );
  NAND2_X1 U22937 ( .A1(n20112), .A2(n20574), .ZN(n20364) );
  NAND2_X1 U22938 ( .A1(n9569), .A2(n20061), .ZN(n20479) );
  NAND2_X1 U22939 ( .A1(n20624), .A2(n20334), .ZN(n20673) );
  OAI21_X1 U22940 ( .B1(n20147), .B2(n20680), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20062) );
  NAND2_X1 U22941 ( .A1(n20062), .A2(n20632), .ZN(n20077) );
  OR2_X1 U22942 ( .A1(n20357), .A2(n20063), .ZN(n20196) );
  OR2_X1 U22943 ( .A1(n20196), .A2(n20580), .ZN(n20076) );
  INV_X1 U22944 ( .A(n20076), .ZN(n20064) );
  NOR3_X1 U22945 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20129) );
  INV_X1 U22946 ( .A(n20129), .ZN(n20120) );
  NOR2_X1 U22947 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20120), .ZN(
        n20111) );
  OAI22_X1 U22948 ( .A1(n20077), .A2(n20064), .B1(n20111), .B2(n20756), .ZN(
        n20065) );
  AOI211_X2 U22949 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20235), .A(n20364), 
        .B(n20065), .ZN(n20119) );
  INV_X1 U22950 ( .A(n20068), .ZN(n20066) );
  NOR2_X2 U22951 ( .A1(n20067), .A2(n20066), .ZN(n20114) );
  INV_X1 U22952 ( .A(n20636), .ZN(n20431) );
  NOR2_X2 U22953 ( .A1(n20110), .A2(n20072), .ZN(n20622) );
  AOI22_X1 U22954 ( .A1(n20680), .A2(n20431), .B1(n20622), .B2(n20111), .ZN(
        n20079) );
  NAND2_X1 U22955 ( .A1(n20073), .A2(n20112), .ZN(n20440) );
  NOR2_X1 U22956 ( .A1(n20075), .A2(n20074), .ZN(n20428) );
  INV_X1 U22957 ( .A(n20428), .ZN(n20157) );
  OAI22_X1 U22958 ( .A1(n20077), .A2(n20076), .B1(n20157), .B2(n20235), .ZN(
        n20115) );
  AOI22_X1 U22959 ( .A1(DATAI_16_), .A2(n20069), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20114), .ZN(n20506) );
  INV_X1 U22960 ( .A(n20506), .ZN(n20633) );
  AOI22_X1 U22961 ( .A1(n20623), .A2(n20115), .B1(n20147), .B2(n20633), .ZN(
        n20078) );
  OAI211_X1 U22962 ( .C1(n20119), .C2(n20080), .A(n20079), .B(n20078), .ZN(
        P1_U3033) );
  AOI22_X1 U22963 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20114), .B1(DATAI_25_), 
        .B2(n20069), .ZN(n20591) );
  INV_X1 U22964 ( .A(n20591), .ZN(n20639) );
  NOR2_X2 U22965 ( .A1(n20110), .A2(n11957), .ZN(n20637) );
  AOI22_X1 U22966 ( .A1(n20680), .A2(n20639), .B1(n20637), .B2(n20111), .ZN(
        n20083) );
  NAND2_X1 U22967 ( .A1(n20081), .A2(n20112), .ZN(n20443) );
  AOI22_X1 U22968 ( .A1(DATAI_17_), .A2(n20069), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n20114), .ZN(n20642) );
  INV_X1 U22969 ( .A(n20642), .ZN(n20588) );
  AOI22_X1 U22970 ( .A1(n20638), .A2(n20115), .B1(n20147), .B2(n20588), .ZN(
        n20082) );
  OAI211_X1 U22971 ( .C1(n20119), .C2(n20084), .A(n20083), .B(n20082), .ZN(
        P1_U3034) );
  INV_X1 U22972 ( .A(n20648), .ZN(n20444) );
  NOR2_X2 U22973 ( .A1(n20110), .A2(n20085), .ZN(n20643) );
  AOI22_X1 U22974 ( .A1(n20680), .A2(n20444), .B1(n20643), .B2(n20111), .ZN(
        n20088) );
  NAND2_X1 U22975 ( .A1(n20086), .A2(n20112), .ZN(n20447) );
  AOI22_X1 U22976 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20114), .B1(DATAI_18_), 
        .B2(n20069), .ZN(n20166) );
  INV_X1 U22977 ( .A(n20166), .ZN(n20645) );
  AOI22_X1 U22978 ( .A1(n20644), .A2(n20115), .B1(n20147), .B2(n20645), .ZN(
        n20087) );
  OAI211_X1 U22979 ( .C1(n20119), .C2(n20089), .A(n20088), .B(n20087), .ZN(
        P1_U3035) );
  AOI22_X1 U22980 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20114), .B1(DATAI_27_), 
        .B2(n20069), .ZN(n20597) );
  INV_X1 U22981 ( .A(n20597), .ZN(n20651) );
  NOR2_X2 U22982 ( .A1(n20110), .A2(n20090), .ZN(n20649) );
  AOI22_X1 U22983 ( .A1(n20680), .A2(n20651), .B1(n20649), .B2(n20111), .ZN(
        n20093) );
  NAND2_X1 U22984 ( .A1(n20091), .A2(n20112), .ZN(n20450) );
  AOI22_X1 U22985 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20114), .B1(DATAI_19_), 
        .B2(n20069), .ZN(n20654) );
  INV_X1 U22986 ( .A(n20654), .ZN(n20594) );
  AOI22_X1 U22987 ( .A1(n20650), .A2(n20115), .B1(n20147), .B2(n20594), .ZN(
        n20092) );
  OAI211_X1 U22988 ( .C1(n20119), .C2(n20897), .A(n20093), .B(n20092), .ZN(
        P1_U3036) );
  INV_X1 U22989 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n20098) );
  AOI22_X1 U22990 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20114), .B1(DATAI_28_), 
        .B2(n20069), .ZN(n20660) );
  INV_X1 U22991 ( .A(n20660), .ZN(n20555) );
  NOR2_X2 U22992 ( .A1(n20110), .A2(n20094), .ZN(n20655) );
  AOI22_X1 U22993 ( .A1(n20680), .A2(n20555), .B1(n20655), .B2(n20111), .ZN(
        n20097) );
  NAND2_X1 U22994 ( .A1(n20095), .A2(n20112), .ZN(n20453) );
  AOI22_X1 U22995 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20114), .B1(DATAI_20_), 
        .B2(n20069), .ZN(n20559) );
  INV_X1 U22996 ( .A(n20559), .ZN(n20657) );
  AOI22_X1 U22997 ( .A1(n20656), .A2(n20115), .B1(n20147), .B2(n20657), .ZN(
        n20096) );
  OAI211_X1 U22998 ( .C1(n20119), .C2(n20098), .A(n20097), .B(n20096), .ZN(
        P1_U3037) );
  AOI22_X1 U22999 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20114), .B1(DATAI_29_), 
        .B2(n20069), .ZN(n20603) );
  INV_X1 U23000 ( .A(n20603), .ZN(n20663) );
  AOI22_X1 U23001 ( .A1(n20680), .A2(n20663), .B1(n20661), .B2(n20111), .ZN(
        n20102) );
  NAND2_X1 U23002 ( .A1(n20100), .A2(n20112), .ZN(n20456) );
  AOI22_X1 U23003 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20114), .B1(DATAI_21_), 
        .B2(n20069), .ZN(n20666) );
  INV_X1 U23004 ( .A(n20666), .ZN(n20600) );
  AOI22_X1 U23005 ( .A1(n20662), .A2(n20115), .B1(n20147), .B2(n20600), .ZN(
        n20101) );
  OAI211_X1 U23006 ( .C1(n20119), .C2(n20103), .A(n20102), .B(n20101), .ZN(
        P1_U3038) );
  INV_X1 U23007 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20108) );
  AOI22_X1 U23008 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20114), .B1(DATAI_30_), 
        .B2(n20069), .ZN(n20607) );
  INV_X1 U23009 ( .A(n20607), .ZN(n20669) );
  NOR2_X2 U23010 ( .A1(n20110), .A2(n20104), .ZN(n20667) );
  AOI22_X1 U23011 ( .A1(n20680), .A2(n20669), .B1(n20667), .B2(n20111), .ZN(
        n20107) );
  NAND2_X1 U23012 ( .A1(n20105), .A2(n20112), .ZN(n20459) );
  AOI22_X1 U23013 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20114), .B1(DATAI_22_), 
        .B2(n20069), .ZN(n20674) );
  INV_X1 U23014 ( .A(n20674), .ZN(n20604) );
  AOI22_X1 U23015 ( .A1(n20668), .A2(n20115), .B1(n20147), .B2(n20604), .ZN(
        n20106) );
  OAI211_X1 U23016 ( .C1(n20119), .C2(n20108), .A(n20107), .B(n20106), .ZN(
        P1_U3039) );
  AOI22_X1 U23017 ( .A1(DATAI_31_), .A2(n20069), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20114), .ZN(n20685) );
  INV_X1 U23018 ( .A(n20685), .ZN(n20499) );
  NOR2_X2 U23019 ( .A1(n20110), .A2(n20109), .ZN(n20676) );
  AOI22_X1 U23020 ( .A1(n20680), .A2(n20499), .B1(n20676), .B2(n20111), .ZN(
        n20117) );
  NAND2_X1 U23021 ( .A1(n20113), .A2(n20112), .ZN(n20465) );
  AOI22_X1 U23022 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20114), .B1(DATAI_23_), 
        .B2(n20069), .ZN(n20504) );
  INV_X1 U23023 ( .A(n20504), .ZN(n20679) );
  AOI22_X1 U23024 ( .A1(n20678), .A2(n20115), .B1(n20147), .B2(n20679), .ZN(
        n20116) );
  OAI211_X1 U23025 ( .C1(n20119), .C2(n20118), .A(n20117), .B(n20116), .ZN(
        P1_U3040) );
  OR2_X1 U23026 ( .A1(n20196), .A2(n20540), .ZN(n20122) );
  NOR2_X1 U23027 ( .A1(n20773), .A2(n20120), .ZN(n20145) );
  INV_X1 U23028 ( .A(n20145), .ZN(n20121) );
  NAND2_X1 U23029 ( .A1(n20122), .A2(n20121), .ZN(n20125) );
  NAND2_X1 U23030 ( .A1(n20125), .A2(n20618), .ZN(n20124) );
  NAND2_X1 U23031 ( .A1(n20129), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20123) );
  NAND2_X1 U23032 ( .A1(n20124), .A2(n20123), .ZN(n20146) );
  AOI22_X1 U23033 ( .A1(n20623), .A2(n20146), .B1(n20622), .B2(n20145), .ZN(
        n20131) );
  INV_X1 U23034 ( .A(n20207), .ZN(n20127) );
  INV_X1 U23035 ( .A(n20125), .ZN(n20126) );
  OAI21_X1 U23036 ( .B1(n20127), .B2(n20399), .A(n20126), .ZN(n20128) );
  OAI221_X1 U23037 ( .B1(n20632), .B2(n20129), .C1(n20769), .C2(n20128), .A(
        n20629), .ZN(n20148) );
  AOI22_X1 U23038 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20148), .B1(
        n20152), .B2(n20633), .ZN(n20130) );
  OAI211_X1 U23039 ( .C1(n20636), .C2(n20142), .A(n20131), .B(n20130), .ZN(
        P1_U3041) );
  AOI22_X1 U23040 ( .A1(n20638), .A2(n20146), .B1(n20637), .B2(n20145), .ZN(
        n20133) );
  AOI22_X1 U23041 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20148), .B1(
        n20147), .B2(n20639), .ZN(n20132) );
  OAI211_X1 U23042 ( .C1(n20642), .C2(n20187), .A(n20133), .B(n20132), .ZN(
        P1_U3042) );
  AOI22_X1 U23043 ( .A1(n20644), .A2(n20146), .B1(n20643), .B2(n20145), .ZN(
        n20135) );
  AOI22_X1 U23044 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20148), .B1(
        n20152), .B2(n20645), .ZN(n20134) );
  OAI211_X1 U23045 ( .C1(n20648), .C2(n20142), .A(n20135), .B(n20134), .ZN(
        P1_U3043) );
  AOI22_X1 U23046 ( .A1(n20650), .A2(n20146), .B1(n20649), .B2(n20145), .ZN(
        n20137) );
  AOI22_X1 U23047 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20148), .B1(
        n20152), .B2(n20594), .ZN(n20136) );
  OAI211_X1 U23048 ( .C1(n20597), .C2(n20142), .A(n20137), .B(n20136), .ZN(
        P1_U3044) );
  AOI22_X1 U23049 ( .A1(n20656), .A2(n20146), .B1(n20655), .B2(n20145), .ZN(
        n20139) );
  AOI22_X1 U23050 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20148), .B1(
        n20152), .B2(n20657), .ZN(n20138) );
  OAI211_X1 U23051 ( .C1(n20660), .C2(n20142), .A(n20139), .B(n20138), .ZN(
        P1_U3045) );
  AOI22_X1 U23052 ( .A1(n20662), .A2(n20146), .B1(n20661), .B2(n20145), .ZN(
        n20141) );
  AOI22_X1 U23053 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20148), .B1(
        n20152), .B2(n20600), .ZN(n20140) );
  OAI211_X1 U23054 ( .C1(n20603), .C2(n20142), .A(n20141), .B(n20140), .ZN(
        P1_U3046) );
  AOI22_X1 U23055 ( .A1(n20668), .A2(n20146), .B1(n20667), .B2(n20145), .ZN(
        n20144) );
  AOI22_X1 U23056 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20148), .B1(
        n20147), .B2(n20669), .ZN(n20143) );
  OAI211_X1 U23057 ( .C1(n20674), .C2(n20187), .A(n20144), .B(n20143), .ZN(
        P1_U3047) );
  AOI22_X1 U23058 ( .A1(n20678), .A2(n20146), .B1(n20676), .B2(n20145), .ZN(
        n20150) );
  AOI22_X1 U23059 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20148), .B1(
        n20147), .B2(n20499), .ZN(n20149) );
  OAI211_X1 U23060 ( .C1(n20504), .C2(n20187), .A(n20150), .B(n20149), .ZN(
        P1_U3048) );
  NAND2_X1 U23061 ( .A1(n9569), .A2(n12758), .ZN(n20423) );
  INV_X1 U23062 ( .A(n20622), .ZN(n20200) );
  NOR3_X1 U23063 ( .A1(n20429), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20202) );
  NAND2_X1 U23064 ( .A1(n20773), .A2(n20202), .ZN(n20186) );
  OAI22_X1 U23065 ( .A1(n20228), .A2(n20506), .B1(n20200), .B2(n20186), .ZN(
        n20151) );
  INV_X1 U23066 ( .A(n20151), .ZN(n20161) );
  OAI21_X1 U23067 ( .B1(n20223), .B2(n20152), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20153) );
  NAND2_X1 U23068 ( .A1(n20153), .A2(n20618), .ZN(n20159) );
  NOR2_X1 U23069 ( .A1(n20196), .A2(n20571), .ZN(n20155) );
  NOR2_X1 U23070 ( .A1(n20359), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20156) );
  NOR2_X1 U23071 ( .A1(n20156), .A2(n20074), .ZN(n20297) );
  AOI211_X1 U23072 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20186), .A(n20297), 
        .B(n20364), .ZN(n20154) );
  OAI21_X1 U23073 ( .B1(n20159), .B2(n20155), .A(n20154), .ZN(n20190) );
  INV_X1 U23074 ( .A(n20155), .ZN(n20158) );
  INV_X1 U23075 ( .A(n20156), .ZN(n20300) );
  OAI22_X1 U23076 ( .A1(n20159), .A2(n20158), .B1(n20157), .B2(n20300), .ZN(
        n20189) );
  AOI22_X1 U23077 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20190), .B1(
        n20623), .B2(n20189), .ZN(n20160) );
  OAI211_X1 U23078 ( .C1(n20636), .C2(n20187), .A(n20161), .B(n20160), .ZN(
        P1_U3049) );
  INV_X1 U23079 ( .A(n20637), .ZN(n20210) );
  OAI22_X1 U23080 ( .A1(n20228), .A2(n20642), .B1(n20210), .B2(n20186), .ZN(
        n20162) );
  INV_X1 U23081 ( .A(n20162), .ZN(n20164) );
  AOI22_X1 U23082 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20190), .B1(
        n20638), .B2(n20189), .ZN(n20163) );
  OAI211_X1 U23083 ( .C1(n20591), .C2(n20187), .A(n20164), .B(n20163), .ZN(
        P1_U3050) );
  INV_X1 U23084 ( .A(n20643), .ZN(n20165) );
  OAI22_X1 U23085 ( .A1(n20228), .A2(n20166), .B1(n20165), .B2(n20186), .ZN(
        n20167) );
  INV_X1 U23086 ( .A(n20167), .ZN(n20169) );
  AOI22_X1 U23087 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20190), .B1(
        n20644), .B2(n20189), .ZN(n20168) );
  OAI211_X1 U23088 ( .C1(n20648), .C2(n20187), .A(n20169), .B(n20168), .ZN(
        P1_U3051) );
  INV_X1 U23089 ( .A(n20649), .ZN(n20170) );
  OAI22_X1 U23090 ( .A1(n20187), .A2(n20597), .B1(n20170), .B2(n20186), .ZN(
        n20171) );
  INV_X1 U23091 ( .A(n20171), .ZN(n20173) );
  AOI22_X1 U23092 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20190), .B1(
        n20650), .B2(n20189), .ZN(n20172) );
  OAI211_X1 U23093 ( .C1(n20654), .C2(n20228), .A(n20173), .B(n20172), .ZN(
        P1_U3052) );
  INV_X1 U23094 ( .A(n20655), .ZN(n20174) );
  OAI22_X1 U23095 ( .A1(n20187), .A2(n20660), .B1(n20174), .B2(n20186), .ZN(
        n20175) );
  INV_X1 U23096 ( .A(n20175), .ZN(n20177) );
  AOI22_X1 U23097 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20190), .B1(
        n20656), .B2(n20189), .ZN(n20176) );
  OAI211_X1 U23098 ( .C1(n20559), .C2(n20228), .A(n20177), .B(n20176), .ZN(
        P1_U3053) );
  INV_X1 U23099 ( .A(n20661), .ZN(n20178) );
  OAI22_X1 U23100 ( .A1(n20187), .A2(n20603), .B1(n20178), .B2(n20186), .ZN(
        n20179) );
  INV_X1 U23101 ( .A(n20179), .ZN(n20181) );
  AOI22_X1 U23102 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20190), .B1(
        n20662), .B2(n20189), .ZN(n20180) );
  OAI211_X1 U23103 ( .C1(n20666), .C2(n20228), .A(n20181), .B(n20180), .ZN(
        P1_U3054) );
  INV_X1 U23104 ( .A(n20667), .ZN(n20182) );
  OAI22_X1 U23105 ( .A1(n20187), .A2(n20607), .B1(n20182), .B2(n20186), .ZN(
        n20183) );
  INV_X1 U23106 ( .A(n20183), .ZN(n20185) );
  AOI22_X1 U23107 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20190), .B1(
        n20668), .B2(n20189), .ZN(n20184) );
  OAI211_X1 U23108 ( .C1(n20674), .C2(n20228), .A(n20185), .B(n20184), .ZN(
        P1_U3055) );
  INV_X1 U23109 ( .A(n20676), .ZN(n20227) );
  OAI22_X1 U23110 ( .A1(n20187), .A2(n20685), .B1(n20227), .B2(n20186), .ZN(
        n20188) );
  INV_X1 U23111 ( .A(n20188), .ZN(n20192) );
  AOI22_X1 U23112 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20190), .B1(
        n20678), .B2(n20189), .ZN(n20191) );
  OAI211_X1 U23113 ( .C1(n20504), .C2(n20228), .A(n20192), .B(n20191), .ZN(
        P1_U3056) );
  OAI21_X1 U23114 ( .B1(n20207), .B2(n20769), .A(n20193), .ZN(n20204) );
  AND2_X1 U23115 ( .A1(n20195), .A2(n20194), .ZN(n20467) );
  INV_X1 U23116 ( .A(n20467), .ZN(n20614) );
  OR2_X1 U23117 ( .A1(n20196), .A2(n20614), .ZN(n20198) );
  INV_X1 U23118 ( .A(n20197), .ZN(n20469) );
  NAND2_X1 U23119 ( .A1(n20469), .A2(n20507), .ZN(n20226) );
  AND2_X1 U23120 ( .A1(n20198), .A2(n20226), .ZN(n20205) );
  INV_X1 U23121 ( .A(n20205), .ZN(n20199) );
  AOI22_X1 U23122 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20202), .B1(n20204), 
        .B2(n20199), .ZN(n20233) );
  OAI22_X1 U23123 ( .A1(n20228), .A2(n20636), .B1(n20200), .B2(n20226), .ZN(
        n20201) );
  INV_X1 U23124 ( .A(n20201), .ZN(n20209) );
  OAI21_X1 U23125 ( .B1(n20632), .B2(n20202), .A(n20629), .ZN(n20203) );
  AOI21_X1 U23126 ( .B1(n20205), .B2(n20204), .A(n20203), .ZN(n20206) );
  AOI22_X1 U23127 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20230), .B1(
        n20261), .B2(n20633), .ZN(n20208) );
  OAI211_X1 U23128 ( .C1(n20233), .C2(n20440), .A(n20209), .B(n20208), .ZN(
        P1_U3057) );
  OAI22_X1 U23129 ( .A1(n20228), .A2(n20591), .B1(n20210), .B2(n20226), .ZN(
        n20211) );
  INV_X1 U23130 ( .A(n20211), .ZN(n20213) );
  AOI22_X1 U23131 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20230), .B1(
        n20261), .B2(n20588), .ZN(n20212) );
  OAI211_X1 U23132 ( .C1(n20233), .C2(n20443), .A(n20213), .B(n20212), .ZN(
        P1_U3058) );
  INV_X1 U23133 ( .A(n20226), .ZN(n20222) );
  AOI22_X1 U23134 ( .A1(n20261), .A2(n20645), .B1(n20643), .B2(n20222), .ZN(
        n20215) );
  AOI22_X1 U23135 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20230), .B1(
        n20223), .B2(n20444), .ZN(n20214) );
  OAI211_X1 U23136 ( .C1(n20233), .C2(n20447), .A(n20215), .B(n20214), .ZN(
        P1_U3059) );
  AOI22_X1 U23137 ( .A1(n20261), .A2(n20594), .B1(n20649), .B2(n20222), .ZN(
        n20217) );
  AOI22_X1 U23138 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20230), .B1(
        n20223), .B2(n20651), .ZN(n20216) );
  OAI211_X1 U23139 ( .C1(n20233), .C2(n20450), .A(n20217), .B(n20216), .ZN(
        P1_U3060) );
  AOI22_X1 U23140 ( .A1(n20261), .A2(n20657), .B1(n20655), .B2(n20222), .ZN(
        n20219) );
  AOI22_X1 U23141 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20230), .B1(
        n20223), .B2(n20555), .ZN(n20218) );
  OAI211_X1 U23142 ( .C1(n20233), .C2(n20453), .A(n20219), .B(n20218), .ZN(
        P1_U3061) );
  AOI22_X1 U23143 ( .A1(n20261), .A2(n20600), .B1(n20661), .B2(n20222), .ZN(
        n20221) );
  AOI22_X1 U23144 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20230), .B1(
        n20223), .B2(n20663), .ZN(n20220) );
  OAI211_X1 U23145 ( .C1(n20233), .C2(n20456), .A(n20221), .B(n20220), .ZN(
        P1_U3062) );
  AOI22_X1 U23146 ( .A1(n20261), .A2(n20604), .B1(n20667), .B2(n20222), .ZN(
        n20225) );
  AOI22_X1 U23147 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20230), .B1(
        n20223), .B2(n20669), .ZN(n20224) );
  OAI211_X1 U23148 ( .C1(n20233), .C2(n20459), .A(n20225), .B(n20224), .ZN(
        P1_U3063) );
  OAI22_X1 U23149 ( .A1(n20228), .A2(n20685), .B1(n20227), .B2(n20226), .ZN(
        n20229) );
  INV_X1 U23150 ( .A(n20229), .ZN(n20232) );
  AOI22_X1 U23151 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20230), .B1(
        n20261), .B2(n20679), .ZN(n20231) );
  OAI211_X1 U23152 ( .C1(n20233), .C2(n20465), .A(n20232), .B(n20231), .ZN(
        P1_U3064) );
  INV_X1 U23153 ( .A(n20261), .ZN(n20250) );
  NOR2_X1 U23154 ( .A1(n20512), .A2(n20234), .ZN(n20324) );
  NAND3_X1 U23155 ( .A1(n20324), .A2(n20618), .A3(n20571), .ZN(n20239) );
  INV_X1 U23156 ( .A(n20235), .ZN(n20237) );
  INV_X1 U23157 ( .A(n20574), .ZN(n20236) );
  NAND2_X1 U23158 ( .A1(n20237), .A2(n20236), .ZN(n20238) );
  NAND2_X1 U23159 ( .A1(n20239), .A2(n20238), .ZN(n20260) );
  NOR3_X1 U23160 ( .A1(n12676), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20274) );
  INV_X1 U23161 ( .A(n20274), .ZN(n20265) );
  NOR2_X1 U23162 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20265), .ZN(
        n20259) );
  AOI22_X1 U23163 ( .A1(n20623), .A2(n20260), .B1(n20622), .B2(n20259), .ZN(
        n20245) );
  INV_X1 U23164 ( .A(n20324), .ZN(n20241) );
  OAI21_X1 U23165 ( .B1(n20261), .B2(n20287), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20240) );
  OAI21_X1 U23166 ( .B1(n20580), .B2(n20241), .A(n20240), .ZN(n20243) );
  NOR2_X1 U23167 ( .A1(n20428), .A2(n20242), .ZN(n20584) );
  OAI221_X1 U23168 ( .B1(n20259), .B2(n20756), .C1(n20259), .C2(n20243), .A(
        n20584), .ZN(n20262) );
  AOI22_X1 U23169 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20262), .B1(
        n20287), .B2(n20633), .ZN(n20244) );
  OAI211_X1 U23170 ( .C1(n20636), .C2(n20250), .A(n20245), .B(n20244), .ZN(
        P1_U3065) );
  AOI22_X1 U23171 ( .A1(n20638), .A2(n20260), .B1(n20637), .B2(n20259), .ZN(
        n20247) );
  AOI22_X1 U23172 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20262), .B1(
        n20287), .B2(n20588), .ZN(n20246) );
  OAI211_X1 U23173 ( .C1(n20591), .C2(n20250), .A(n20247), .B(n20246), .ZN(
        P1_U3066) );
  AOI22_X1 U23174 ( .A1(n20644), .A2(n20260), .B1(n20643), .B2(n20259), .ZN(
        n20249) );
  AOI22_X1 U23175 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20262), .B1(
        n20287), .B2(n20645), .ZN(n20248) );
  OAI211_X1 U23176 ( .C1(n20648), .C2(n20250), .A(n20249), .B(n20248), .ZN(
        P1_U3067) );
  AOI22_X1 U23177 ( .A1(n20650), .A2(n20260), .B1(n20649), .B2(n20259), .ZN(
        n20252) );
  AOI22_X1 U23178 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20262), .B1(
        n20261), .B2(n20651), .ZN(n20251) );
  OAI211_X1 U23179 ( .C1(n20654), .C2(n20295), .A(n20252), .B(n20251), .ZN(
        P1_U3068) );
  AOI22_X1 U23180 ( .A1(n20656), .A2(n20260), .B1(n20655), .B2(n20259), .ZN(
        n20254) );
  AOI22_X1 U23181 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20262), .B1(
        n20261), .B2(n20555), .ZN(n20253) );
  OAI211_X1 U23182 ( .C1(n20559), .C2(n20295), .A(n20254), .B(n20253), .ZN(
        P1_U3069) );
  AOI22_X1 U23183 ( .A1(n20662), .A2(n20260), .B1(n20661), .B2(n20259), .ZN(
        n20256) );
  AOI22_X1 U23184 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20262), .B1(
        n20261), .B2(n20663), .ZN(n20255) );
  OAI211_X1 U23185 ( .C1(n20666), .C2(n20295), .A(n20256), .B(n20255), .ZN(
        P1_U3070) );
  AOI22_X1 U23186 ( .A1(n20668), .A2(n20260), .B1(n20667), .B2(n20259), .ZN(
        n20258) );
  AOI22_X1 U23187 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20262), .B1(
        n20261), .B2(n20669), .ZN(n20257) );
  OAI211_X1 U23188 ( .C1(n20674), .C2(n20295), .A(n20258), .B(n20257), .ZN(
        P1_U3071) );
  AOI22_X1 U23189 ( .A1(n20678), .A2(n20260), .B1(n20676), .B2(n20259), .ZN(
        n20264) );
  AOI22_X1 U23190 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20262), .B1(
        n20261), .B2(n20499), .ZN(n20263) );
  OAI211_X1 U23191 ( .C1(n20504), .C2(n20295), .A(n20264), .B(n20263), .ZN(
        P1_U3072) );
  INV_X1 U23192 ( .A(n20540), .ZN(n20391) );
  NAND2_X1 U23193 ( .A1(n20324), .A2(n20391), .ZN(n20267) );
  NOR2_X1 U23194 ( .A1(n20773), .A2(n20265), .ZN(n20290) );
  INV_X1 U23195 ( .A(n20290), .ZN(n20266) );
  NAND2_X1 U23196 ( .A1(n20267), .A2(n20266), .ZN(n20270) );
  NAND2_X1 U23197 ( .A1(n20270), .A2(n20618), .ZN(n20269) );
  NAND2_X1 U23198 ( .A1(n20274), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20268) );
  NAND2_X1 U23199 ( .A1(n20269), .A2(n20268), .ZN(n20291) );
  AOI22_X1 U23200 ( .A1(n20623), .A2(n20291), .B1(n20622), .B2(n20290), .ZN(
        n20276) );
  INV_X1 U23201 ( .A(n20270), .ZN(n20271) );
  OAI21_X1 U23202 ( .B1(n20272), .B2(n20399), .A(n20271), .ZN(n20273) );
  OAI221_X1 U23203 ( .B1(n20618), .B2(n20274), .C1(n20769), .C2(n20273), .A(
        n20629), .ZN(n20292) );
  AOI22_X1 U23204 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20292), .B1(
        n20319), .B2(n20633), .ZN(n20275) );
  OAI211_X1 U23205 ( .C1(n20636), .C2(n20295), .A(n20276), .B(n20275), .ZN(
        P1_U3073) );
  AOI22_X1 U23206 ( .A1(n20638), .A2(n20291), .B1(n20637), .B2(n20290), .ZN(
        n20278) );
  AOI22_X1 U23207 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20292), .B1(
        n20287), .B2(n20639), .ZN(n20277) );
  OAI211_X1 U23208 ( .C1(n20642), .C2(n20317), .A(n20278), .B(n20277), .ZN(
        P1_U3074) );
  AOI22_X1 U23209 ( .A1(n20644), .A2(n20291), .B1(n20643), .B2(n20290), .ZN(
        n20280) );
  AOI22_X1 U23210 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20292), .B1(
        n20319), .B2(n20645), .ZN(n20279) );
  OAI211_X1 U23211 ( .C1(n20648), .C2(n20295), .A(n20280), .B(n20279), .ZN(
        P1_U3075) );
  AOI22_X1 U23212 ( .A1(n20650), .A2(n20291), .B1(n20649), .B2(n20290), .ZN(
        n20282) );
  AOI22_X1 U23213 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20292), .B1(
        n20319), .B2(n20594), .ZN(n20281) );
  OAI211_X1 U23214 ( .C1(n20597), .C2(n20295), .A(n20282), .B(n20281), .ZN(
        P1_U3076) );
  AOI22_X1 U23215 ( .A1(n20656), .A2(n20291), .B1(n20655), .B2(n20290), .ZN(
        n20284) );
  AOI22_X1 U23216 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20292), .B1(
        n20319), .B2(n20657), .ZN(n20283) );
  OAI211_X1 U23217 ( .C1(n20660), .C2(n20295), .A(n20284), .B(n20283), .ZN(
        P1_U3077) );
  AOI22_X1 U23218 ( .A1(n20662), .A2(n20291), .B1(n20661), .B2(n20290), .ZN(
        n20286) );
  AOI22_X1 U23219 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20292), .B1(
        n20287), .B2(n20663), .ZN(n20285) );
  OAI211_X1 U23220 ( .C1(n20666), .C2(n20317), .A(n20286), .B(n20285), .ZN(
        P1_U3078) );
  AOI22_X1 U23221 ( .A1(n20668), .A2(n20291), .B1(n20667), .B2(n20290), .ZN(
        n20289) );
  AOI22_X1 U23222 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20292), .B1(
        n20287), .B2(n20669), .ZN(n20288) );
  OAI211_X1 U23223 ( .C1(n20674), .C2(n20317), .A(n20289), .B(n20288), .ZN(
        P1_U3079) );
  AOI22_X1 U23224 ( .A1(n20678), .A2(n20291), .B1(n20676), .B2(n20290), .ZN(
        n20294) );
  AOI22_X1 U23225 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20292), .B1(
        n20319), .B2(n20679), .ZN(n20293) );
  OAI211_X1 U23226 ( .C1(n20685), .C2(n20295), .A(n20294), .B(n20293), .ZN(
        P1_U3080) );
  NOR2_X1 U23227 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20327), .ZN(
        n20318) );
  AOI22_X1 U23228 ( .A1(n20353), .A2(n20633), .B1(n20622), .B2(n20318), .ZN(
        n20304) );
  NAND2_X1 U23229 ( .A1(n20348), .A2(n20317), .ZN(n20296) );
  AOI21_X1 U23230 ( .B1(n20296), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20769), 
        .ZN(n20299) );
  NAND2_X1 U23231 ( .A1(n20324), .A2(n20580), .ZN(n20301) );
  AOI21_X1 U23232 ( .B1(n20299), .B2(n20301), .A(n20297), .ZN(n20298) );
  OAI211_X1 U23233 ( .C1(n20318), .C2(n20756), .A(n20584), .B(n20298), .ZN(
        n20321) );
  INV_X1 U23234 ( .A(n20299), .ZN(n20302) );
  OAI22_X1 U23235 ( .A1(n20302), .A2(n20301), .B1(n20300), .B2(n20574), .ZN(
        n20320) );
  AOI22_X1 U23236 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20321), .B1(
        n20623), .B2(n20320), .ZN(n20303) );
  OAI211_X1 U23237 ( .C1(n20636), .C2(n20317), .A(n20304), .B(n20303), .ZN(
        P1_U3081) );
  AOI22_X1 U23238 ( .A1(n20319), .A2(n20639), .B1(n20637), .B2(n20318), .ZN(
        n20306) );
  AOI22_X1 U23239 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20321), .B1(
        n20638), .B2(n20320), .ZN(n20305) );
  OAI211_X1 U23240 ( .C1(n20642), .C2(n20348), .A(n20306), .B(n20305), .ZN(
        P1_U3082) );
  AOI22_X1 U23241 ( .A1(n20353), .A2(n20645), .B1(n20643), .B2(n20318), .ZN(
        n20308) );
  AOI22_X1 U23242 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20321), .B1(
        n20644), .B2(n20320), .ZN(n20307) );
  OAI211_X1 U23243 ( .C1(n20648), .C2(n20317), .A(n20308), .B(n20307), .ZN(
        P1_U3083) );
  AOI22_X1 U23244 ( .A1(n20353), .A2(n20594), .B1(n20649), .B2(n20318), .ZN(
        n20310) );
  AOI22_X1 U23245 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20321), .B1(
        n20650), .B2(n20320), .ZN(n20309) );
  OAI211_X1 U23246 ( .C1(n20597), .C2(n20317), .A(n20310), .B(n20309), .ZN(
        P1_U3084) );
  AOI22_X1 U23247 ( .A1(n20319), .A2(n20555), .B1(n20655), .B2(n20318), .ZN(
        n20312) );
  AOI22_X1 U23248 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20321), .B1(
        n20656), .B2(n20320), .ZN(n20311) );
  OAI211_X1 U23249 ( .C1(n20559), .C2(n20348), .A(n20312), .B(n20311), .ZN(
        P1_U3085) );
  AOI22_X1 U23250 ( .A1(n20353), .A2(n20600), .B1(n20661), .B2(n20318), .ZN(
        n20314) );
  AOI22_X1 U23251 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20321), .B1(
        n20662), .B2(n20320), .ZN(n20313) );
  OAI211_X1 U23252 ( .C1(n20603), .C2(n20317), .A(n20314), .B(n20313), .ZN(
        P1_U3086) );
  AOI22_X1 U23253 ( .A1(n20353), .A2(n20604), .B1(n20667), .B2(n20318), .ZN(
        n20316) );
  AOI22_X1 U23254 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20321), .B1(
        n20668), .B2(n20320), .ZN(n20315) );
  OAI211_X1 U23255 ( .C1(n20607), .C2(n20317), .A(n20316), .B(n20315), .ZN(
        P1_U3087) );
  AOI22_X1 U23256 ( .A1(n20319), .A2(n20499), .B1(n20676), .B2(n20318), .ZN(
        n20323) );
  AOI22_X1 U23257 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20321), .B1(
        n20678), .B2(n20320), .ZN(n20322) );
  OAI211_X1 U23258 ( .C1(n20504), .C2(n20348), .A(n20323), .B(n20322), .ZN(
        P1_U3088) );
  NAND2_X1 U23259 ( .A1(n20324), .A2(n20467), .ZN(n20326) );
  INV_X1 U23260 ( .A(n20351), .ZN(n20325) );
  NAND2_X1 U23261 ( .A1(n20326), .A2(n20325), .ZN(n20330) );
  NAND2_X1 U23262 ( .A1(n20330), .A2(n20618), .ZN(n20329) );
  INV_X1 U23263 ( .A(n20327), .ZN(n20333) );
  NAND2_X1 U23264 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20333), .ZN(n20328) );
  NAND2_X1 U23265 ( .A1(n20329), .A2(n20328), .ZN(n20352) );
  AOI22_X1 U23266 ( .A1(n20623), .A2(n20352), .B1(n20622), .B2(n20351), .ZN(
        n20337) );
  OR2_X1 U23267 ( .A1(n20331), .A2(n20330), .ZN(n20332) );
  OAI221_X1 U23268 ( .B1(n20632), .B2(n20333), .C1(n20769), .C2(n20332), .A(
        n20629), .ZN(n20354) );
  AOI22_X1 U23269 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20354), .B1(
        n20366), .B2(n20633), .ZN(n20336) );
  OAI211_X1 U23270 ( .C1(n20636), .C2(n20348), .A(n20337), .B(n20336), .ZN(
        P1_U3089) );
  AOI22_X1 U23271 ( .A1(n20638), .A2(n20352), .B1(n20637), .B2(n20351), .ZN(
        n20339) );
  AOI22_X1 U23272 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20354), .B1(
        n20366), .B2(n20588), .ZN(n20338) );
  OAI211_X1 U23273 ( .C1(n20591), .C2(n20348), .A(n20339), .B(n20338), .ZN(
        P1_U3090) );
  AOI22_X1 U23274 ( .A1(n20644), .A2(n20352), .B1(n20643), .B2(n20351), .ZN(
        n20341) );
  AOI22_X1 U23275 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20354), .B1(
        n20366), .B2(n20645), .ZN(n20340) );
  OAI211_X1 U23276 ( .C1(n20648), .C2(n20348), .A(n20341), .B(n20340), .ZN(
        P1_U3091) );
  AOI22_X1 U23277 ( .A1(n20650), .A2(n20352), .B1(n20649), .B2(n20351), .ZN(
        n20343) );
  AOI22_X1 U23278 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20354), .B1(
        n20353), .B2(n20651), .ZN(n20342) );
  OAI211_X1 U23279 ( .C1(n20654), .C2(n20390), .A(n20343), .B(n20342), .ZN(
        P1_U3092) );
  AOI22_X1 U23280 ( .A1(n20656), .A2(n20352), .B1(n20655), .B2(n20351), .ZN(
        n20345) );
  AOI22_X1 U23281 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20354), .B1(
        n20353), .B2(n20555), .ZN(n20344) );
  OAI211_X1 U23282 ( .C1(n20559), .C2(n20390), .A(n20345), .B(n20344), .ZN(
        P1_U3093) );
  AOI22_X1 U23283 ( .A1(n20662), .A2(n20352), .B1(n20661), .B2(n20351), .ZN(
        n20347) );
  AOI22_X1 U23284 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20354), .B1(
        n20366), .B2(n20600), .ZN(n20346) );
  OAI211_X1 U23285 ( .C1(n20603), .C2(n20348), .A(n20347), .B(n20346), .ZN(
        P1_U3094) );
  AOI22_X1 U23286 ( .A1(n20668), .A2(n20352), .B1(n20667), .B2(n20351), .ZN(
        n20350) );
  AOI22_X1 U23287 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20354), .B1(
        n20353), .B2(n20669), .ZN(n20349) );
  OAI211_X1 U23288 ( .C1(n20674), .C2(n20390), .A(n20350), .B(n20349), .ZN(
        P1_U3095) );
  AOI22_X1 U23289 ( .A1(n20678), .A2(n20352), .B1(n20676), .B2(n20351), .ZN(
        n20356) );
  AOI22_X1 U23290 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20354), .B1(
        n20353), .B2(n20499), .ZN(n20355) );
  OAI211_X1 U23291 ( .C1(n20504), .C2(n20390), .A(n20356), .B(n20355), .ZN(
        P1_U3096) );
  AND2_X1 U23292 ( .A1(n20512), .A2(n20357), .ZN(n20468) );
  NOR3_X1 U23293 ( .A1(n20507), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20401) );
  INV_X1 U23294 ( .A(n20401), .ZN(n20392) );
  NOR2_X1 U23295 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20392), .ZN(
        n20384) );
  AOI21_X1 U23296 ( .B1(n20468), .B2(n20571), .A(n20384), .ZN(n20367) );
  OR2_X1 U23297 ( .A1(n20367), .A2(n20769), .ZN(n20363) );
  INV_X1 U23298 ( .A(n20358), .ZN(n20360) );
  NAND2_X1 U23299 ( .A1(n20360), .A2(n20359), .ZN(n20515) );
  INV_X1 U23300 ( .A(n20515), .ZN(n20361) );
  NAND2_X1 U23301 ( .A1(n20361), .A2(n20428), .ZN(n20362) );
  NAND2_X1 U23302 ( .A1(n20363), .A2(n20362), .ZN(n20385) );
  AOI22_X1 U23303 ( .A1(n20623), .A2(n20385), .B1(n20622), .B2(n20384), .ZN(
        n20371) );
  INV_X1 U23304 ( .A(n20364), .ZN(n20433) );
  OAI21_X1 U23305 ( .B1(n20386), .B2(n20366), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20368) );
  NAND2_X1 U23306 ( .A1(n20368), .A2(n20367), .ZN(n20369) );
  AOI22_X1 U23307 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20387), .B1(
        n20386), .B2(n20633), .ZN(n20370) );
  OAI211_X1 U23308 ( .C1(n20636), .C2(n20390), .A(n20371), .B(n20370), .ZN(
        P1_U3097) );
  AOI22_X1 U23309 ( .A1(n20638), .A2(n20385), .B1(n20637), .B2(n20384), .ZN(
        n20373) );
  AOI22_X1 U23310 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20387), .B1(
        n20386), .B2(n20588), .ZN(n20372) );
  OAI211_X1 U23311 ( .C1(n20591), .C2(n20390), .A(n20373), .B(n20372), .ZN(
        P1_U3098) );
  AOI22_X1 U23312 ( .A1(n20644), .A2(n20385), .B1(n20643), .B2(n20384), .ZN(
        n20375) );
  AOI22_X1 U23313 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20387), .B1(
        n20386), .B2(n20645), .ZN(n20374) );
  OAI211_X1 U23314 ( .C1(n20648), .C2(n20390), .A(n20375), .B(n20374), .ZN(
        P1_U3099) );
  AOI22_X1 U23315 ( .A1(n20650), .A2(n20385), .B1(n20649), .B2(n20384), .ZN(
        n20377) );
  AOI22_X1 U23316 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20387), .B1(
        n20386), .B2(n20594), .ZN(n20376) );
  OAI211_X1 U23317 ( .C1(n20597), .C2(n20390), .A(n20377), .B(n20376), .ZN(
        P1_U3100) );
  AOI22_X1 U23318 ( .A1(n20656), .A2(n20385), .B1(n20655), .B2(n20384), .ZN(
        n20379) );
  AOI22_X1 U23319 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20387), .B1(
        n20386), .B2(n20657), .ZN(n20378) );
  OAI211_X1 U23320 ( .C1(n20660), .C2(n20390), .A(n20379), .B(n20378), .ZN(
        P1_U3101) );
  AOI22_X1 U23321 ( .A1(n20662), .A2(n20385), .B1(n20661), .B2(n20384), .ZN(
        n20381) );
  AOI22_X1 U23322 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20387), .B1(
        n20386), .B2(n20600), .ZN(n20380) );
  OAI211_X1 U23323 ( .C1(n20603), .C2(n20390), .A(n20381), .B(n20380), .ZN(
        P1_U3102) );
  AOI22_X1 U23324 ( .A1(n20668), .A2(n20385), .B1(n20667), .B2(n20384), .ZN(
        n20383) );
  AOI22_X1 U23325 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20387), .B1(
        n20386), .B2(n20604), .ZN(n20382) );
  OAI211_X1 U23326 ( .C1(n20607), .C2(n20390), .A(n20383), .B(n20382), .ZN(
        P1_U3103) );
  AOI22_X1 U23327 ( .A1(n20678), .A2(n20385), .B1(n20676), .B2(n20384), .ZN(
        n20389) );
  AOI22_X1 U23328 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20387), .B1(
        n20386), .B2(n20679), .ZN(n20388) );
  OAI211_X1 U23329 ( .C1(n20685), .C2(n20390), .A(n20389), .B(n20388), .ZN(
        P1_U3104) );
  NAND2_X1 U23330 ( .A1(n20468), .A2(n20391), .ZN(n20394) );
  NOR2_X1 U23331 ( .A1(n20773), .A2(n20392), .ZN(n20417) );
  INV_X1 U23332 ( .A(n20417), .ZN(n20393) );
  NAND2_X1 U23333 ( .A1(n20394), .A2(n20393), .ZN(n20397) );
  NAND2_X1 U23334 ( .A1(n20397), .A2(n20618), .ZN(n20396) );
  NAND2_X1 U23335 ( .A1(n20401), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20395) );
  NAND2_X1 U23336 ( .A1(n20396), .A2(n20395), .ZN(n20418) );
  AOI22_X1 U23337 ( .A1(n20623), .A2(n20418), .B1(n20622), .B2(n20417), .ZN(
        n20404) );
  INV_X1 U23338 ( .A(n20397), .ZN(n20398) );
  OAI21_X1 U23339 ( .B1(n20480), .B2(n20399), .A(n20398), .ZN(n20400) );
  OAI221_X1 U23340 ( .B1(n20618), .B2(n20401), .C1(n20769), .C2(n20400), .A(
        n20629), .ZN(n20419) );
  NOR2_X2 U23341 ( .A1(n20480), .A2(n20402), .ZN(n20461) );
  AOI22_X1 U23342 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20419), .B1(
        n20461), .B2(n20633), .ZN(n20403) );
  OAI211_X1 U23343 ( .C1(n20636), .C2(n20422), .A(n20404), .B(n20403), .ZN(
        P1_U3105) );
  AOI22_X1 U23344 ( .A1(n20638), .A2(n20418), .B1(n20637), .B2(n20417), .ZN(
        n20406) );
  AOI22_X1 U23345 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20419), .B1(
        n20461), .B2(n20588), .ZN(n20405) );
  OAI211_X1 U23346 ( .C1(n20591), .C2(n20422), .A(n20406), .B(n20405), .ZN(
        P1_U3106) );
  AOI22_X1 U23347 ( .A1(n20644), .A2(n20418), .B1(n20643), .B2(n20417), .ZN(
        n20408) );
  AOI22_X1 U23348 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20419), .B1(
        n20461), .B2(n20645), .ZN(n20407) );
  OAI211_X1 U23349 ( .C1(n20648), .C2(n20422), .A(n20408), .B(n20407), .ZN(
        P1_U3107) );
  AOI22_X1 U23350 ( .A1(n20650), .A2(n20418), .B1(n20649), .B2(n20417), .ZN(
        n20410) );
  AOI22_X1 U23351 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20419), .B1(
        n20461), .B2(n20594), .ZN(n20409) );
  OAI211_X1 U23352 ( .C1(n20597), .C2(n20422), .A(n20410), .B(n20409), .ZN(
        P1_U3108) );
  AOI22_X1 U23353 ( .A1(n20656), .A2(n20418), .B1(n20655), .B2(n20417), .ZN(
        n20412) );
  AOI22_X1 U23354 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20419), .B1(
        n20461), .B2(n20657), .ZN(n20411) );
  OAI211_X1 U23355 ( .C1(n20660), .C2(n20422), .A(n20412), .B(n20411), .ZN(
        P1_U3109) );
  AOI22_X1 U23356 ( .A1(n20662), .A2(n20418), .B1(n20661), .B2(n20417), .ZN(
        n20414) );
  AOI22_X1 U23357 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20419), .B1(
        n20461), .B2(n20600), .ZN(n20413) );
  OAI211_X1 U23358 ( .C1(n20603), .C2(n20422), .A(n20414), .B(n20413), .ZN(
        P1_U3110) );
  AOI22_X1 U23359 ( .A1(n20668), .A2(n20418), .B1(n20667), .B2(n20417), .ZN(
        n20416) );
  AOI22_X1 U23360 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20419), .B1(
        n20461), .B2(n20604), .ZN(n20415) );
  OAI211_X1 U23361 ( .C1(n20607), .C2(n20422), .A(n20416), .B(n20415), .ZN(
        P1_U3111) );
  AOI22_X1 U23362 ( .A1(n20678), .A2(n20418), .B1(n20676), .B2(n20417), .ZN(
        n20421) );
  AOI22_X1 U23363 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20419), .B1(
        n20461), .B2(n20679), .ZN(n20420) );
  OAI211_X1 U23364 ( .C1(n20685), .C2(n20422), .A(n20421), .B(n20420), .ZN(
        P1_U3112) );
  INV_X1 U23365 ( .A(n20461), .ZN(n20424) );
  AOI21_X1 U23366 ( .B1(n20424), .B2(n20496), .A(n20578), .ZN(n20425) );
  NOR2_X1 U23367 ( .A1(n20425), .A2(n20769), .ZN(n20436) );
  AND2_X1 U23368 ( .A1(n20468), .A2(n20580), .ZN(n20432) );
  NAND2_X1 U23369 ( .A1(n20426), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20573) );
  INV_X1 U23370 ( .A(n20573), .ZN(n20427) );
  AOI22_X1 U23371 ( .A1(n20436), .A2(n20432), .B1(n20428), .B2(n20427), .ZN(
        n20466) );
  NOR3_X1 U23372 ( .A1(n20507), .A2(n20429), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20478) );
  INV_X1 U23373 ( .A(n20478), .ZN(n20430) );
  NOR2_X1 U23374 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20430), .ZN(
        n20460) );
  AOI22_X1 U23375 ( .A1(n20461), .A2(n20431), .B1(n20622), .B2(n20460), .ZN(
        n20439) );
  INV_X1 U23376 ( .A(n20432), .ZN(n20435) );
  NAND2_X1 U23377 ( .A1(n20573), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20583) );
  OAI211_X1 U23378 ( .C1(n20756), .C2(n20460), .A(n20583), .B(n20433), .ZN(
        n20434) );
  AOI21_X1 U23379 ( .B1(n20436), .B2(n20435), .A(n20434), .ZN(n20437) );
  AOI22_X1 U23380 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20462), .B1(
        n20500), .B2(n20633), .ZN(n20438) );
  OAI211_X1 U23381 ( .C1(n20466), .C2(n20440), .A(n20439), .B(n20438), .ZN(
        P1_U3113) );
  AOI22_X1 U23382 ( .A1(n20461), .A2(n20639), .B1(n20637), .B2(n20460), .ZN(
        n20442) );
  AOI22_X1 U23383 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20462), .B1(
        n20500), .B2(n20588), .ZN(n20441) );
  OAI211_X1 U23384 ( .C1(n20466), .C2(n20443), .A(n20442), .B(n20441), .ZN(
        P1_U3114) );
  AOI22_X1 U23385 ( .A1(n20461), .A2(n20444), .B1(n20643), .B2(n20460), .ZN(
        n20446) );
  AOI22_X1 U23386 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20462), .B1(
        n20500), .B2(n20645), .ZN(n20445) );
  OAI211_X1 U23387 ( .C1(n20466), .C2(n20447), .A(n20446), .B(n20445), .ZN(
        P1_U3115) );
  AOI22_X1 U23388 ( .A1(n20461), .A2(n20651), .B1(n20649), .B2(n20460), .ZN(
        n20449) );
  AOI22_X1 U23389 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20462), .B1(
        n20500), .B2(n20594), .ZN(n20448) );
  OAI211_X1 U23390 ( .C1(n20466), .C2(n20450), .A(n20449), .B(n20448), .ZN(
        P1_U3116) );
  AOI22_X1 U23391 ( .A1(n20461), .A2(n20555), .B1(n20655), .B2(n20460), .ZN(
        n20452) );
  AOI22_X1 U23392 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20462), .B1(
        n20500), .B2(n20657), .ZN(n20451) );
  OAI211_X1 U23393 ( .C1(n20466), .C2(n20453), .A(n20452), .B(n20451), .ZN(
        P1_U3117) );
  AOI22_X1 U23394 ( .A1(n20461), .A2(n20663), .B1(n20661), .B2(n20460), .ZN(
        n20455) );
  AOI22_X1 U23395 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20462), .B1(
        n20500), .B2(n20600), .ZN(n20454) );
  OAI211_X1 U23396 ( .C1(n20466), .C2(n20456), .A(n20455), .B(n20454), .ZN(
        P1_U3118) );
  AOI22_X1 U23397 ( .A1(n20461), .A2(n20669), .B1(n20667), .B2(n20460), .ZN(
        n20458) );
  AOI22_X1 U23398 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20462), .B1(
        n20500), .B2(n20604), .ZN(n20457) );
  OAI211_X1 U23399 ( .C1(n20466), .C2(n20459), .A(n20458), .B(n20457), .ZN(
        P1_U3119) );
  AOI22_X1 U23400 ( .A1(n20461), .A2(n20499), .B1(n20676), .B2(n20460), .ZN(
        n20464) );
  AOI22_X1 U23401 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20462), .B1(
        n20500), .B2(n20679), .ZN(n20463) );
  OAI211_X1 U23402 ( .C1(n20466), .C2(n20465), .A(n20464), .B(n20463), .ZN(
        P1_U3120) );
  NAND2_X1 U23403 ( .A1(n20468), .A2(n20467), .ZN(n20470) );
  NAND2_X1 U23404 ( .A1(n20469), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20474) );
  NAND2_X1 U23405 ( .A1(n20470), .A2(n20474), .ZN(n20471) );
  NAND2_X1 U23406 ( .A1(n20471), .A2(n20618), .ZN(n20473) );
  NAND2_X1 U23407 ( .A1(n20478), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20472) );
  NAND2_X1 U23408 ( .A1(n20473), .A2(n20472), .ZN(n20498) );
  INV_X1 U23409 ( .A(n20474), .ZN(n20497) );
  AOI22_X1 U23410 ( .A1(n20623), .A2(n20498), .B1(n20622), .B2(n20497), .ZN(
        n20482) );
  INV_X1 U23411 ( .A(n20475), .ZN(n20476) );
  NOR2_X1 U23412 ( .A1(n20480), .A2(n20476), .ZN(n20477) );
  OAI21_X1 U23413 ( .B1(n20478), .B2(n20477), .A(n20629), .ZN(n20501) );
  INV_X1 U23414 ( .A(n20537), .ZN(n20493) );
  AOI22_X1 U23415 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20501), .B1(
        n20493), .B2(n20633), .ZN(n20481) );
  OAI211_X1 U23416 ( .C1(n20636), .C2(n20496), .A(n20482), .B(n20481), .ZN(
        P1_U3121) );
  AOI22_X1 U23417 ( .A1(n20638), .A2(n20498), .B1(n20637), .B2(n20497), .ZN(
        n20484) );
  AOI22_X1 U23418 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20501), .B1(
        n20500), .B2(n20639), .ZN(n20483) );
  OAI211_X1 U23419 ( .C1(n20642), .C2(n20537), .A(n20484), .B(n20483), .ZN(
        P1_U3122) );
  AOI22_X1 U23420 ( .A1(n20644), .A2(n20498), .B1(n20643), .B2(n20497), .ZN(
        n20486) );
  AOI22_X1 U23421 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20501), .B1(
        n20493), .B2(n20645), .ZN(n20485) );
  OAI211_X1 U23422 ( .C1(n20648), .C2(n20496), .A(n20486), .B(n20485), .ZN(
        P1_U3123) );
  AOI22_X1 U23423 ( .A1(n20650), .A2(n20498), .B1(n20649), .B2(n20497), .ZN(
        n20488) );
  AOI22_X1 U23424 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20501), .B1(
        n20500), .B2(n20651), .ZN(n20487) );
  OAI211_X1 U23425 ( .C1(n20654), .C2(n20537), .A(n20488), .B(n20487), .ZN(
        P1_U3124) );
  AOI22_X1 U23426 ( .A1(n20656), .A2(n20498), .B1(n20655), .B2(n20497), .ZN(
        n20490) );
  AOI22_X1 U23427 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20501), .B1(
        n20493), .B2(n20657), .ZN(n20489) );
  OAI211_X1 U23428 ( .C1(n20660), .C2(n20496), .A(n20490), .B(n20489), .ZN(
        P1_U3125) );
  AOI22_X1 U23429 ( .A1(n20662), .A2(n20498), .B1(n20661), .B2(n20497), .ZN(
        n20492) );
  AOI22_X1 U23430 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20501), .B1(
        n20500), .B2(n20663), .ZN(n20491) );
  OAI211_X1 U23431 ( .C1(n20666), .C2(n20537), .A(n20492), .B(n20491), .ZN(
        P1_U3126) );
  AOI22_X1 U23432 ( .A1(n20668), .A2(n20498), .B1(n20667), .B2(n20497), .ZN(
        n20495) );
  AOI22_X1 U23433 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20501), .B1(
        n20493), .B2(n20604), .ZN(n20494) );
  OAI211_X1 U23434 ( .C1(n20607), .C2(n20496), .A(n20495), .B(n20494), .ZN(
        P1_U3127) );
  AOI22_X1 U23435 ( .A1(n20678), .A2(n20498), .B1(n20676), .B2(n20497), .ZN(
        n20503) );
  AOI22_X1 U23436 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20501), .B1(
        n20500), .B2(n20499), .ZN(n20502) );
  OAI211_X1 U23437 ( .C1(n20504), .C2(n20537), .A(n20503), .B(n20502), .ZN(
        P1_U3128) );
  NAND2_X1 U23438 ( .A1(n20624), .A2(n20505), .ZN(n20570) );
  OR2_X1 U23439 ( .A1(n20570), .A2(n20506), .ZN(n20509) );
  NOR3_X1 U23440 ( .A1(n12676), .A2(n20507), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20545) );
  INV_X1 U23441 ( .A(n20545), .ZN(n20538) );
  NOR2_X1 U23442 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20538), .ZN(
        n20532) );
  NAND2_X1 U23443 ( .A1(n20622), .A2(n20532), .ZN(n20508) );
  AND2_X1 U23444 ( .A1(n20509), .A2(n20508), .ZN(n20519) );
  NAND2_X1 U23445 ( .A1(n20537), .A2(n20570), .ZN(n20510) );
  AOI21_X1 U23446 ( .B1(n20510), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20769), 
        .ZN(n20514) );
  OR2_X1 U23447 ( .A1(n20512), .A2(n20511), .ZN(n20615) );
  OR2_X1 U23448 ( .A1(n20615), .A2(n20580), .ZN(n20516) );
  AOI22_X1 U23449 ( .A1(n20514), .A2(n20516), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20515), .ZN(n20513) );
  OAI211_X1 U23450 ( .C1(n20532), .C2(n20756), .A(n20584), .B(n20513), .ZN(
        n20534) );
  INV_X1 U23451 ( .A(n20514), .ZN(n20517) );
  AOI22_X1 U23452 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20534), .B1(
        n20623), .B2(n20533), .ZN(n20518) );
  OAI211_X1 U23453 ( .C1(n20636), .C2(n20537), .A(n20519), .B(n20518), .ZN(
        P1_U3129) );
  INV_X1 U23454 ( .A(n20570), .ZN(n20556) );
  AOI22_X1 U23455 ( .A1(n20556), .A2(n20588), .B1(n20637), .B2(n20532), .ZN(
        n20521) );
  AOI22_X1 U23456 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20534), .B1(
        n20638), .B2(n20533), .ZN(n20520) );
  OAI211_X1 U23457 ( .C1(n20591), .C2(n20537), .A(n20521), .B(n20520), .ZN(
        P1_U3130) );
  AOI22_X1 U23458 ( .A1(n20556), .A2(n20645), .B1(n20643), .B2(n20532), .ZN(
        n20523) );
  AOI22_X1 U23459 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20534), .B1(
        n20644), .B2(n20533), .ZN(n20522) );
  OAI211_X1 U23460 ( .C1(n20648), .C2(n20537), .A(n20523), .B(n20522), .ZN(
        P1_U3131) );
  AOI22_X1 U23461 ( .A1(n20556), .A2(n20594), .B1(n20649), .B2(n20532), .ZN(
        n20525) );
  AOI22_X1 U23462 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20534), .B1(
        n20650), .B2(n20533), .ZN(n20524) );
  OAI211_X1 U23463 ( .C1(n20597), .C2(n20537), .A(n20525), .B(n20524), .ZN(
        P1_U3132) );
  AOI22_X1 U23464 ( .A1(n20556), .A2(n20657), .B1(n20655), .B2(n20532), .ZN(
        n20527) );
  AOI22_X1 U23465 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20534), .B1(
        n20656), .B2(n20533), .ZN(n20526) );
  OAI211_X1 U23466 ( .C1(n20660), .C2(n20537), .A(n20527), .B(n20526), .ZN(
        P1_U3133) );
  AOI22_X1 U23467 ( .A1(n20556), .A2(n20600), .B1(n20661), .B2(n20532), .ZN(
        n20529) );
  AOI22_X1 U23468 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20534), .B1(
        n20662), .B2(n20533), .ZN(n20528) );
  OAI211_X1 U23469 ( .C1(n20603), .C2(n20537), .A(n20529), .B(n20528), .ZN(
        P1_U3134) );
  AOI22_X1 U23470 ( .A1(n20556), .A2(n20604), .B1(n20667), .B2(n20532), .ZN(
        n20531) );
  AOI22_X1 U23471 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20534), .B1(
        n20668), .B2(n20533), .ZN(n20530) );
  OAI211_X1 U23472 ( .C1(n20607), .C2(n20537), .A(n20531), .B(n20530), .ZN(
        P1_U3135) );
  AOI22_X1 U23473 ( .A1(n20556), .A2(n20679), .B1(n20676), .B2(n20532), .ZN(
        n20536) );
  AOI22_X1 U23474 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20534), .B1(
        n20678), .B2(n20533), .ZN(n20535) );
  OAI211_X1 U23475 ( .C1(n20685), .C2(n20537), .A(n20536), .B(n20535), .ZN(
        P1_U3136) );
  NOR2_X1 U23476 ( .A1(n20773), .A2(n20538), .ZN(n20564) );
  INV_X1 U23477 ( .A(n20564), .ZN(n20539) );
  OAI21_X1 U23478 ( .B1(n20615), .B2(n20540), .A(n20539), .ZN(n20541) );
  NAND2_X1 U23479 ( .A1(n20541), .A2(n20632), .ZN(n20543) );
  NAND2_X1 U23480 ( .A1(n20545), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20542) );
  NAND2_X1 U23481 ( .A1(n20543), .A2(n20542), .ZN(n20565) );
  AOI22_X1 U23482 ( .A1(n20623), .A2(n20565), .B1(n20622), .B2(n20564), .ZN(
        n20548) );
  OAI21_X1 U23483 ( .B1(n20545), .B2(n20544), .A(n20629), .ZN(n20567) );
  NAND2_X1 U23484 ( .A1(n20624), .A2(n20546), .ZN(n20613) );
  INV_X1 U23485 ( .A(n20613), .ZN(n20566) );
  AOI22_X1 U23486 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20567), .B1(
        n20566), .B2(n20633), .ZN(n20547) );
  OAI211_X1 U23487 ( .C1(n20636), .C2(n20570), .A(n20548), .B(n20547), .ZN(
        P1_U3137) );
  AOI22_X1 U23488 ( .A1(n20638), .A2(n20565), .B1(n20637), .B2(n20564), .ZN(
        n20550) );
  AOI22_X1 U23489 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20567), .B1(
        n20566), .B2(n20588), .ZN(n20549) );
  OAI211_X1 U23490 ( .C1(n20591), .C2(n20570), .A(n20550), .B(n20549), .ZN(
        P1_U3138) );
  AOI22_X1 U23491 ( .A1(n20644), .A2(n20565), .B1(n20643), .B2(n20564), .ZN(
        n20552) );
  AOI22_X1 U23492 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20567), .B1(
        n20566), .B2(n20645), .ZN(n20551) );
  OAI211_X1 U23493 ( .C1(n20648), .C2(n20570), .A(n20552), .B(n20551), .ZN(
        P1_U3139) );
  AOI22_X1 U23494 ( .A1(n20650), .A2(n20565), .B1(n20649), .B2(n20564), .ZN(
        n20554) );
  AOI22_X1 U23495 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20567), .B1(
        n20566), .B2(n20594), .ZN(n20553) );
  OAI211_X1 U23496 ( .C1(n20597), .C2(n20570), .A(n20554), .B(n20553), .ZN(
        P1_U3140) );
  AOI22_X1 U23497 ( .A1(n20656), .A2(n20565), .B1(n20655), .B2(n20564), .ZN(
        n20558) );
  AOI22_X1 U23498 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20567), .B1(
        n20556), .B2(n20555), .ZN(n20557) );
  OAI211_X1 U23499 ( .C1(n20559), .C2(n20613), .A(n20558), .B(n20557), .ZN(
        P1_U3141) );
  AOI22_X1 U23500 ( .A1(n20662), .A2(n20565), .B1(n20661), .B2(n20564), .ZN(
        n20561) );
  AOI22_X1 U23501 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20567), .B1(
        n20566), .B2(n20600), .ZN(n20560) );
  OAI211_X1 U23502 ( .C1(n20603), .C2(n20570), .A(n20561), .B(n20560), .ZN(
        P1_U3142) );
  AOI22_X1 U23503 ( .A1(n20668), .A2(n20565), .B1(n20667), .B2(n20564), .ZN(
        n20563) );
  AOI22_X1 U23504 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20567), .B1(
        n20566), .B2(n20604), .ZN(n20562) );
  OAI211_X1 U23505 ( .C1(n20607), .C2(n20570), .A(n20563), .B(n20562), .ZN(
        P1_U3143) );
  AOI22_X1 U23506 ( .A1(n20678), .A2(n20565), .B1(n20676), .B2(n20564), .ZN(
        n20569) );
  AOI22_X1 U23507 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20567), .B1(
        n20566), .B2(n20679), .ZN(n20568) );
  OAI211_X1 U23508 ( .C1(n20685), .C2(n20570), .A(n20569), .B(n20568), .ZN(
        P1_U3144) );
  OR2_X1 U23509 ( .A1(n20571), .A2(n20769), .ZN(n20572) );
  OR2_X1 U23510 ( .A1(n20615), .A2(n20572), .ZN(n20576) );
  OR2_X1 U23511 ( .A1(n20574), .A2(n20573), .ZN(n20575) );
  NAND2_X1 U23512 ( .A1(n20576), .A2(n20575), .ZN(n20609) );
  NOR2_X1 U23513 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20619), .ZN(
        n20608) );
  AOI22_X1 U23514 ( .A1(n20623), .A2(n20609), .B1(n20622), .B2(n20608), .ZN(
        n20587) );
  INV_X1 U23515 ( .A(n20615), .ZN(n20581) );
  NAND2_X1 U23516 ( .A1(n20624), .A2(n20577), .ZN(n20684) );
  AOI21_X1 U23517 ( .B1(n20684), .B2(n20613), .A(n20578), .ZN(n20579) );
  AOI21_X1 U23518 ( .B1(n20581), .B2(n20580), .A(n20579), .ZN(n20582) );
  NOR2_X1 U23519 ( .A1(n20582), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20585) );
  OAI211_X1 U23520 ( .C1(n20608), .C2(n20585), .A(n20584), .B(n20583), .ZN(
        n20610) );
  AOI22_X1 U23521 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20610), .B1(
        n20670), .B2(n20633), .ZN(n20586) );
  OAI211_X1 U23522 ( .C1(n20636), .C2(n20613), .A(n20587), .B(n20586), .ZN(
        P1_U3145) );
  AOI22_X1 U23523 ( .A1(n20638), .A2(n20609), .B1(n20637), .B2(n20608), .ZN(
        n20590) );
  AOI22_X1 U23524 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20610), .B1(
        n20670), .B2(n20588), .ZN(n20589) );
  OAI211_X1 U23525 ( .C1(n20591), .C2(n20613), .A(n20590), .B(n20589), .ZN(
        P1_U3146) );
  AOI22_X1 U23526 ( .A1(n20644), .A2(n20609), .B1(n20643), .B2(n20608), .ZN(
        n20593) );
  AOI22_X1 U23527 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20610), .B1(
        n20670), .B2(n20645), .ZN(n20592) );
  OAI211_X1 U23528 ( .C1(n20648), .C2(n20613), .A(n20593), .B(n20592), .ZN(
        P1_U3147) );
  AOI22_X1 U23529 ( .A1(n20650), .A2(n20609), .B1(n20649), .B2(n20608), .ZN(
        n20596) );
  AOI22_X1 U23530 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20610), .B1(
        n20670), .B2(n20594), .ZN(n20595) );
  OAI211_X1 U23531 ( .C1(n20597), .C2(n20613), .A(n20596), .B(n20595), .ZN(
        P1_U3148) );
  AOI22_X1 U23532 ( .A1(n20656), .A2(n20609), .B1(n20655), .B2(n20608), .ZN(
        n20599) );
  AOI22_X1 U23533 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20610), .B1(
        n20670), .B2(n20657), .ZN(n20598) );
  OAI211_X1 U23534 ( .C1(n20660), .C2(n20613), .A(n20599), .B(n20598), .ZN(
        P1_U3149) );
  AOI22_X1 U23535 ( .A1(n20662), .A2(n20609), .B1(n20661), .B2(n20608), .ZN(
        n20602) );
  AOI22_X1 U23536 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20610), .B1(
        n20670), .B2(n20600), .ZN(n20601) );
  OAI211_X1 U23537 ( .C1(n20603), .C2(n20613), .A(n20602), .B(n20601), .ZN(
        P1_U3150) );
  AOI22_X1 U23538 ( .A1(n20668), .A2(n20609), .B1(n20667), .B2(n20608), .ZN(
        n20606) );
  AOI22_X1 U23539 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20610), .B1(
        n20670), .B2(n20604), .ZN(n20605) );
  OAI211_X1 U23540 ( .C1(n20607), .C2(n20613), .A(n20606), .B(n20605), .ZN(
        P1_U3151) );
  AOI22_X1 U23541 ( .A1(n20678), .A2(n20609), .B1(n20676), .B2(n20608), .ZN(
        n20612) );
  AOI22_X1 U23542 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20610), .B1(
        n20670), .B2(n20679), .ZN(n20611) );
  OAI211_X1 U23543 ( .C1(n20685), .C2(n20613), .A(n20612), .B(n20611), .ZN(
        P1_U3152) );
  OR2_X1 U23544 ( .A1(n20615), .A2(n20614), .ZN(n20617) );
  INV_X1 U23545 ( .A(n20675), .ZN(n20616) );
  NAND2_X1 U23546 ( .A1(n20617), .A2(n20616), .ZN(n20625) );
  NAND2_X1 U23547 ( .A1(n20625), .A2(n20618), .ZN(n20621) );
  NAND2_X1 U23548 ( .A1(n20631), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20620) );
  NAND2_X1 U23549 ( .A1(n20621), .A2(n20620), .ZN(n20677) );
  AOI22_X1 U23550 ( .A1(n20623), .A2(n20677), .B1(n20622), .B2(n20675), .ZN(
        n20635) );
  INV_X1 U23551 ( .A(n20624), .ZN(n20628) );
  INV_X1 U23552 ( .A(n20625), .ZN(n20626) );
  OAI21_X1 U23553 ( .B1(n20628), .B2(n20627), .A(n20626), .ZN(n20630) );
  OAI221_X1 U23554 ( .B1(n20632), .B2(n20631), .C1(n20769), .C2(n20630), .A(
        n20629), .ZN(n20681) );
  AOI22_X1 U23555 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20681), .B1(
        n20680), .B2(n20633), .ZN(n20634) );
  OAI211_X1 U23556 ( .C1(n20636), .C2(n20684), .A(n20635), .B(n20634), .ZN(
        P1_U3153) );
  AOI22_X1 U23557 ( .A1(n20638), .A2(n20677), .B1(n20637), .B2(n20675), .ZN(
        n20641) );
  AOI22_X1 U23558 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20681), .B1(
        n20670), .B2(n20639), .ZN(n20640) );
  OAI211_X1 U23559 ( .C1(n20642), .C2(n20673), .A(n20641), .B(n20640), .ZN(
        P1_U3154) );
  AOI22_X1 U23560 ( .A1(n20644), .A2(n20677), .B1(n20643), .B2(n20675), .ZN(
        n20647) );
  AOI22_X1 U23561 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20681), .B1(
        n20680), .B2(n20645), .ZN(n20646) );
  OAI211_X1 U23562 ( .C1(n20648), .C2(n20684), .A(n20647), .B(n20646), .ZN(
        P1_U3155) );
  AOI22_X1 U23563 ( .A1(n20650), .A2(n20677), .B1(n20649), .B2(n20675), .ZN(
        n20653) );
  AOI22_X1 U23564 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20681), .B1(
        n20670), .B2(n20651), .ZN(n20652) );
  OAI211_X1 U23565 ( .C1(n20654), .C2(n20673), .A(n20653), .B(n20652), .ZN(
        P1_U3156) );
  AOI22_X1 U23566 ( .A1(n20656), .A2(n20677), .B1(n20655), .B2(n20675), .ZN(
        n20659) );
  AOI22_X1 U23567 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20681), .B1(
        n20680), .B2(n20657), .ZN(n20658) );
  OAI211_X1 U23568 ( .C1(n20660), .C2(n20684), .A(n20659), .B(n20658), .ZN(
        P1_U3157) );
  AOI22_X1 U23569 ( .A1(n20662), .A2(n20677), .B1(n20661), .B2(n20675), .ZN(
        n20665) );
  AOI22_X1 U23570 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20681), .B1(
        n20670), .B2(n20663), .ZN(n20664) );
  OAI211_X1 U23571 ( .C1(n20666), .C2(n20673), .A(n20665), .B(n20664), .ZN(
        P1_U3158) );
  AOI22_X1 U23572 ( .A1(n20668), .A2(n20677), .B1(n20667), .B2(n20675), .ZN(
        n20672) );
  AOI22_X1 U23573 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20681), .B1(
        n20670), .B2(n20669), .ZN(n20671) );
  OAI211_X1 U23574 ( .C1(n20674), .C2(n20673), .A(n20672), .B(n20671), .ZN(
        P1_U3159) );
  AOI22_X1 U23575 ( .A1(n20678), .A2(n20677), .B1(n20676), .B2(n20675), .ZN(
        n20683) );
  AOI22_X1 U23576 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20681), .B1(
        n20680), .B2(n20679), .ZN(n20682) );
  OAI211_X1 U23577 ( .C1(n20685), .C2(n20684), .A(n20683), .B(n20682), .ZN(
        P1_U3160) );
  NAND3_X1 U23578 ( .A1(n20687), .A2(n20686), .A3(n9989), .ZN(P1_U3163) );
  INV_X1 U23579 ( .A(n20755), .ZN(n20688) );
  AND2_X1 U23580 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20688), .ZN(
        P1_U3164) );
  AND2_X1 U23581 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20688), .ZN(
        P1_U3165) );
  AND2_X1 U23582 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20688), .ZN(
        P1_U3166) );
  AND2_X1 U23583 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20688), .ZN(
        P1_U3167) );
  AND2_X1 U23584 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20688), .ZN(
        P1_U3168) );
  AND2_X1 U23585 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20688), .ZN(
        P1_U3169) );
  AND2_X1 U23586 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20688), .ZN(
        P1_U3170) );
  AND2_X1 U23587 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20688), .ZN(
        P1_U3171) );
  AND2_X1 U23588 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20688), .ZN(
        P1_U3172) );
  AND2_X1 U23589 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20688), .ZN(
        P1_U3173) );
  AND2_X1 U23590 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20688), .ZN(
        P1_U3174) );
  AND2_X1 U23591 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20688), .ZN(
        P1_U3175) );
  AND2_X1 U23592 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20688), .ZN(
        P1_U3176) );
  AND2_X1 U23593 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20688), .ZN(
        P1_U3177) );
  AND2_X1 U23594 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20688), .ZN(
        P1_U3178) );
  AND2_X1 U23595 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20688), .ZN(
        P1_U3179) );
  AND2_X1 U23596 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20688), .ZN(
        P1_U3180) );
  AND2_X1 U23597 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20688), .ZN(
        P1_U3181) );
  AND2_X1 U23598 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20688), .ZN(
        P1_U3182) );
  AND2_X1 U23599 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20688), .ZN(
        P1_U3183) );
  AND2_X1 U23600 ( .A1(n20688), .A2(P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(
        P1_U3184) );
  AND2_X1 U23601 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20688), .ZN(
        P1_U3185) );
  AND2_X1 U23602 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20688), .ZN(P1_U3186) );
  AND2_X1 U23603 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20688), .ZN(P1_U3187) );
  AND2_X1 U23604 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20688), .ZN(P1_U3188) );
  AND2_X1 U23605 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20688), .ZN(P1_U3189) );
  AND2_X1 U23606 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20688), .ZN(P1_U3190) );
  AND2_X1 U23607 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20688), .ZN(P1_U3191) );
  AND2_X1 U23608 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20688), .ZN(P1_U3192) );
  AND2_X1 U23609 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20688), .ZN(P1_U3193) );
  INV_X1 U23610 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20701) );
  OAI21_X1 U23611 ( .B1(n20701), .B2(n20786), .A(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20696) );
  INV_X1 U23612 ( .A(n20696), .ZN(n20692) );
  OAI21_X1 U23613 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20697), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20689) );
  AOI211_X1 U23614 ( .C1(HOLD), .C2(P1_STATE_REG_1__SCAN_IN), .A(n20690), .B(
        n20689), .ZN(n20691) );
  OAI22_X1 U23615 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20692), .B1(n20795), 
        .B2(n20691), .ZN(P1_U3194) );
  NAND4_X1 U23616 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20693), .A3(
        P1_REQUESTPENDING_REG_SCAN_IN), .A4(n20697), .ZN(n20700) );
  NAND2_X1 U23617 ( .A1(n20693), .A2(n20697), .ZN(n20694) );
  OAI221_X1 U23618 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(
        P1_STATE_REG_1__SCAN_IN), .C1(P1_REQUESTPENDING_REG_SCAN_IN), .C2(
        n20694), .A(n20702), .ZN(n20695) );
  NAND3_X1 U23619 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(HOLD), .A3(n20695), .ZN(
        n20699) );
  OAI211_X1 U23620 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n20697), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20696), .ZN(n20698) );
  OAI211_X1 U23621 ( .C1(n20701), .C2(n20700), .A(n20699), .B(n20698), .ZN(
        P1_U3196) );
  OR2_X1 U23622 ( .A1(n20738), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20746) );
  INV_X1 U23623 ( .A(n20746), .ZN(n20740) );
  OR2_X1 U23624 ( .A1(n20702), .A2(n20796), .ZN(n20742) );
  INV_X1 U23625 ( .A(n20742), .ZN(n20744) );
  AOI222_X1 U23626 ( .A1(n20740), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20738), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n20744), .ZN(n20703) );
  INV_X1 U23627 ( .A(n20703), .ZN(P1_U3197) );
  AOI22_X1 U23628 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n20796), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n20740), .ZN(n20704) );
  OAI21_X1 U23629 ( .B1(n13077), .B2(n20742), .A(n20704), .ZN(P1_U3198) );
  AOI222_X1 U23630 ( .A1(n20744), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n20738), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20740), .ZN(n20705) );
  INV_X1 U23631 ( .A(n20705), .ZN(P1_U3199) );
  AOI222_X1 U23632 ( .A1(n20744), .A2(P1_REIP_REG_4__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20738), .C1(P1_REIP_REG_5__SCAN_IN), 
        .C2(n20740), .ZN(n20706) );
  INV_X1 U23633 ( .A(n20706), .ZN(P1_U3200) );
  AOI222_X1 U23634 ( .A1(n20744), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20738), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20740), .ZN(n20707) );
  INV_X1 U23635 ( .A(n20707), .ZN(P1_U3201) );
  AOI222_X1 U23636 ( .A1(n20744), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20738), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20740), .ZN(n20708) );
  INV_X1 U23637 ( .A(n20708), .ZN(P1_U3202) );
  INV_X1 U23638 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20709) );
  INV_X1 U23639 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20711) );
  OAI222_X1 U23640 ( .A1(n20742), .A2(n20710), .B1(n20709), .B2(n20795), .C1(
        n20711), .C2(n20746), .ZN(P1_U3203) );
  INV_X1 U23641 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20712) );
  OAI222_X1 U23642 ( .A1(n20746), .A2(n20713), .B1(n20712), .B2(n20795), .C1(
        n20711), .C2(n20742), .ZN(P1_U3204) );
  AOI222_X1 U23643 ( .A1(n20744), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20738), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20740), .ZN(n20714) );
  INV_X1 U23644 ( .A(n20714), .ZN(P1_U3205) );
  AOI222_X1 U23645 ( .A1(n20740), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20738), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20744), .ZN(n20715) );
  INV_X1 U23646 ( .A(n20715), .ZN(P1_U3206) );
  AOI222_X1 U23647 ( .A1(n20744), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20738), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20740), .ZN(n20716) );
  INV_X1 U23648 ( .A(n20716), .ZN(P1_U3207) );
  INV_X1 U23649 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20869) );
  OAI222_X1 U23650 ( .A1(n20742), .A2(n20718), .B1(n20869), .B2(n20795), .C1(
        n20717), .C2(n20746), .ZN(P1_U3208) );
  AOI222_X1 U23651 ( .A1(n20744), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20738), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20740), .ZN(n20719) );
  INV_X1 U23652 ( .A(n20719), .ZN(P1_U3209) );
  AOI222_X1 U23653 ( .A1(n20740), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20738), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20744), .ZN(n20720) );
  INV_X1 U23654 ( .A(n20720), .ZN(P1_U3210) );
  AOI222_X1 U23655 ( .A1(n20744), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20796), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20740), .ZN(n20721) );
  INV_X1 U23656 ( .A(n20721), .ZN(P1_U3211) );
  AOI22_X1 U23657 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20796), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20740), .ZN(n20722) );
  OAI21_X1 U23658 ( .B1(n20723), .B2(n20742), .A(n20722), .ZN(P1_U3212) );
  AOI22_X1 U23659 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20796), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20744), .ZN(n20724) );
  OAI21_X1 U23660 ( .B1(n20725), .B2(n20746), .A(n20724), .ZN(P1_U3213) );
  AOI222_X1 U23661 ( .A1(n20744), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20738), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20740), .ZN(n20726) );
  INV_X1 U23662 ( .A(n20726), .ZN(P1_U3214) );
  AOI222_X1 U23663 ( .A1(n20744), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20738), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n20740), .ZN(n20727) );
  INV_X1 U23664 ( .A(n20727), .ZN(P1_U3215) );
  AOI222_X1 U23665 ( .A1(n20744), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20738), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20740), .ZN(n20728) );
  INV_X1 U23666 ( .A(n20728), .ZN(P1_U3216) );
  AOI222_X1 U23667 ( .A1(n20744), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20738), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n20740), .ZN(n20729) );
  INV_X1 U23668 ( .A(n20729), .ZN(P1_U3217) );
  AOI22_X1 U23669 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20796), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20740), .ZN(n20730) );
  OAI21_X1 U23670 ( .B1(n20731), .B2(n20742), .A(n20730), .ZN(P1_U3218) );
  AOI22_X1 U23671 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n20796), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20744), .ZN(n20732) );
  OAI21_X1 U23672 ( .B1(n20733), .B2(n20746), .A(n20732), .ZN(P1_U3219) );
  AOI222_X1 U23673 ( .A1(n20744), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20738), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20740), .ZN(n20734) );
  INV_X1 U23674 ( .A(n20734), .ZN(P1_U3220) );
  AOI222_X1 U23675 ( .A1(n20744), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20738), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20740), .ZN(n20735) );
  INV_X1 U23676 ( .A(n20735), .ZN(P1_U3221) );
  AOI222_X1 U23677 ( .A1(n20744), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20738), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20740), .ZN(n20736) );
  INV_X1 U23678 ( .A(n20736), .ZN(P1_U3222) );
  AOI222_X1 U23679 ( .A1(n20744), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20738), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20740), .ZN(n20737) );
  INV_X1 U23680 ( .A(n20737), .ZN(P1_U3223) );
  AOI222_X1 U23681 ( .A1(n20744), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20738), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20740), .ZN(n20739) );
  INV_X1 U23682 ( .A(n20739), .ZN(P1_U3224) );
  AOI22_X1 U23683 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20740), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20796), .ZN(n20741) );
  OAI21_X1 U23684 ( .B1(n20743), .B2(n20742), .A(n20741), .ZN(P1_U3225) );
  AOI22_X1 U23685 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20744), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20796), .ZN(n20745) );
  OAI21_X1 U23686 ( .B1(n20747), .B2(n20746), .A(n20745), .ZN(P1_U3226) );
  OAI22_X1 U23687 ( .A1(n20796), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20795), .ZN(n20748) );
  INV_X1 U23688 ( .A(n20748), .ZN(P1_U3458) );
  OAI22_X1 U23689 ( .A1(n20796), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20795), .ZN(n20749) );
  INV_X1 U23690 ( .A(n20749), .ZN(P1_U3459) );
  OAI22_X1 U23691 ( .A1(n20796), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20795), .ZN(n20750) );
  INV_X1 U23692 ( .A(n20750), .ZN(P1_U3460) );
  OAI22_X1 U23693 ( .A1(n20796), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20795), .ZN(n20751) );
  INV_X1 U23694 ( .A(n20751), .ZN(P1_U3461) );
  OAI21_X1 U23695 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20755), .A(n20753), 
        .ZN(n20752) );
  INV_X1 U23696 ( .A(n20752), .ZN(P1_U3464) );
  OAI21_X1 U23697 ( .B1(n20755), .B2(n20754), .A(n20753), .ZN(P1_U3465) );
  AOI21_X1 U23698 ( .B1(n20757), .B2(n20756), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n20759) );
  OAI22_X1 U23699 ( .A1(n20760), .A2(n20759), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20758), .ZN(n20762) );
  AOI22_X1 U23700 ( .A1(n20763), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20762), .B2(n20761), .ZN(n20764) );
  OAI21_X1 U23701 ( .B1(n20766), .B2(n20765), .A(n20764), .ZN(P1_U3474) );
  OAI22_X1 U23702 ( .A1(n12758), .A2(n20769), .B1(n20768), .B2(n20767), .ZN(
        n20770) );
  OAI21_X1 U23703 ( .B1(n20771), .B2(n20770), .A(n20774), .ZN(n20772) );
  OAI21_X1 U23704 ( .B1(n20774), .B2(n20773), .A(n20772), .ZN(P1_U3478) );
  AOI21_X1 U23705 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20776) );
  AOI22_X1 U23706 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20776), .B2(n20775), .ZN(n20779) );
  INV_X1 U23707 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20778) );
  AOI22_X1 U23708 ( .A1(n20782), .A2(n20779), .B1(n20778), .B2(n20777), .ZN(
        P1_U3481) );
  INV_X1 U23709 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20781) );
  OAI21_X1 U23710 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20782), .ZN(n20780) );
  OAI21_X1 U23711 ( .B1(n20782), .B2(n20781), .A(n20780), .ZN(P1_U3482) );
  AOI22_X1 U23712 ( .A1(n20795), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20783), 
        .B2(n20796), .ZN(P1_U3483) );
  AOI211_X1 U23713 ( .C1(n19930), .C2(n20786), .A(n20785), .B(n20784), .ZN(
        n20794) );
  INV_X1 U23714 ( .A(n20787), .ZN(n20788) );
  OAI211_X1 U23715 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20789), .A(n20788), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20791) );
  AOI21_X1 U23716 ( .B1(n20791), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n20790), 
        .ZN(n20793) );
  NAND2_X1 U23717 ( .A1(n20794), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20792) );
  OAI21_X1 U23718 ( .B1(n20794), .B2(n20793), .A(n20792), .ZN(P1_U3485) );
  OAI22_X1 U23719 ( .A1(n20796), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n20795), .ZN(n20797) );
  INV_X1 U23720 ( .A(n20797), .ZN(P1_U3486) );
  INV_X1 U23721 ( .A(keyinput55), .ZN(n20824) );
  NAND3_X1 U23722 ( .A1(keyinput50), .A2(keyinput27), .A3(keyinput4), .ZN(
        n20801) );
  INV_X1 U23723 ( .A(keyinput17), .ZN(n20894) );
  NAND4_X1 U23724 ( .A1(keyinput62), .A2(keyinput43), .A3(keyinput19), .A4(
        n20894), .ZN(n20800) );
  INV_X1 U23725 ( .A(keyinput48), .ZN(n20889) );
  NOR4_X1 U23726 ( .A1(keyinput35), .A2(keyinput22), .A3(keyinput36), .A4(
        n20889), .ZN(n20798) );
  NAND4_X1 U23727 ( .A1(keyinput16), .A2(keyinput13), .A3(keyinput63), .A4(
        n20798), .ZN(n20799) );
  NOR4_X1 U23728 ( .A1(keyinput53), .A2(n20801), .A3(n20800), .A4(n20799), 
        .ZN(n20822) );
  NAND2_X1 U23729 ( .A1(keyinput20), .A2(keyinput5), .ZN(n20807) );
  NOR2_X1 U23730 ( .A1(keyinput12), .A2(keyinput15), .ZN(n20805) );
  NAND3_X1 U23731 ( .A1(keyinput25), .A2(keyinput45), .A3(keyinput42), .ZN(
        n20803) );
  NAND3_X1 U23732 ( .A1(keyinput52), .A2(keyinput3), .A3(keyinput30), .ZN(
        n20802) );
  NOR4_X1 U23733 ( .A1(keyinput59), .A2(keyinput40), .A3(n20803), .A4(n20802), 
        .ZN(n20804) );
  NAND4_X1 U23734 ( .A1(keyinput31), .A2(keyinput28), .A3(n20805), .A4(n20804), 
        .ZN(n20806) );
  NOR4_X1 U23735 ( .A1(keyinput23), .A2(keyinput47), .A3(n20807), .A4(n20806), 
        .ZN(n20821) );
  NOR2_X1 U23736 ( .A1(keyinput9), .A2(keyinput18), .ZN(n20808) );
  NAND3_X1 U23737 ( .A1(keyinput0), .A2(keyinput7), .A3(n20808), .ZN(n20813)
         );
  NAND3_X1 U23738 ( .A1(keyinput24), .A2(keyinput26), .A3(keyinput46), .ZN(
        n20812) );
  NOR3_X1 U23739 ( .A1(keyinput60), .A2(keyinput11), .A3(keyinput1), .ZN(
        n20810) );
  INV_X1 U23740 ( .A(keyinput57), .ZN(n20834) );
  NOR3_X1 U23741 ( .A1(keyinput61), .A2(keyinput21), .A3(n20834), .ZN(n20809)
         );
  NAND4_X1 U23742 ( .A1(keyinput41), .A2(n20810), .A3(keyinput10), .A4(n20809), 
        .ZN(n20811) );
  NOR4_X1 U23743 ( .A1(keyinput58), .A2(n20813), .A3(n20812), .A4(n20811), 
        .ZN(n20820) );
  INV_X1 U23744 ( .A(keyinput49), .ZN(n20862) );
  NAND3_X1 U23745 ( .A1(keyinput2), .A2(keyinput38), .A3(n20862), .ZN(n20818)
         );
  NAND4_X1 U23746 ( .A1(keyinput51), .A2(keyinput34), .A3(keyinput44), .A4(
        keyinput39), .ZN(n20817) );
  NOR3_X1 U23747 ( .A1(keyinput8), .A2(keyinput29), .A3(keyinput33), .ZN(
        n20815) );
  NOR3_X1 U23748 ( .A1(keyinput6), .A2(keyinput14), .A3(keyinput56), .ZN(
        n20814) );
  NAND4_X1 U23749 ( .A1(keyinput37), .A2(n20815), .A3(keyinput54), .A4(n20814), 
        .ZN(n20816) );
  NOR4_X1 U23750 ( .A1(keyinput32), .A2(n20818), .A3(n20817), .A4(n20816), 
        .ZN(n20819) );
  NAND4_X1 U23751 ( .A1(n20822), .A2(n20821), .A3(n20820), .A4(n20819), .ZN(
        n20823) );
  AOI21_X1 U23752 ( .B1(n20824), .B2(n20823), .A(P2_DATAWIDTH_REG_14__SCAN_IN), 
        .ZN(n20955) );
  INV_X1 U23753 ( .A(keyinput46), .ZN(n20826) );
  OAI22_X1 U23754 ( .A1(n14411), .A2(keyinput61), .B1(n20826), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n20825) );
  AOI221_X1 U23755 ( .B1(n14411), .B2(keyinput61), .C1(
        P1_DATAO_REG_12__SCAN_IN), .C2(n20826), .A(n20825), .ZN(n20839) );
  OAI22_X1 U23756 ( .A1(n20829), .A2(keyinput58), .B1(n20828), .B2(keyinput26), 
        .ZN(n20827) );
  AOI221_X1 U23757 ( .B1(n20829), .B2(keyinput58), .C1(keyinput26), .C2(n20828), .A(n20827), .ZN(n20838) );
  OAI22_X1 U23758 ( .A1(n20832), .A2(keyinput21), .B1(n20831), .B2(keyinput37), 
        .ZN(n20830) );
  AOI221_X1 U23759 ( .B1(n20832), .B2(keyinput21), .C1(keyinput37), .C2(n20831), .A(n20830), .ZN(n20837) );
  INV_X1 U23760 ( .A(DATAI_9_), .ZN(n20835) );
  OAI22_X1 U23761 ( .A1(n20835), .A2(keyinput10), .B1(n20834), .B2(
        P1_DATAO_REG_31__SCAN_IN), .ZN(n20833) );
  AOI221_X1 U23762 ( .B1(n20835), .B2(keyinput10), .C1(
        P1_DATAO_REG_31__SCAN_IN), .C2(n20834), .A(n20833), .ZN(n20836) );
  NAND4_X1 U23763 ( .A1(n20839), .A2(n20838), .A3(n20837), .A4(n20836), .ZN(
        n20954) );
  OAI22_X1 U23764 ( .A1(n11626), .A2(keyinput11), .B1(n11453), .B2(keyinput0), 
        .ZN(n20840) );
  AOI221_X1 U23765 ( .B1(n11626), .B2(keyinput11), .C1(keyinput0), .C2(n11453), 
        .A(n20840), .ZN(n20852) );
  INV_X1 U23766 ( .A(keyinput1), .ZN(n20842) );
  OAI22_X1 U23767 ( .A1(n14875), .A2(keyinput60), .B1(n20842), .B2(
        P3_DATAO_REG_23__SCAN_IN), .ZN(n20841) );
  AOI221_X1 U23768 ( .B1(n14875), .B2(keyinput60), .C1(
        P3_DATAO_REG_23__SCAN_IN), .C2(n20842), .A(n20841), .ZN(n20851) );
  INV_X1 U23769 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n20845) );
  OAI22_X1 U23770 ( .A1(n20845), .A2(keyinput18), .B1(n20844), .B2(keyinput24), 
        .ZN(n20843) );
  AOI221_X1 U23771 ( .B1(n20845), .B2(keyinput18), .C1(keyinput24), .C2(n20844), .A(n20843), .ZN(n20850) );
  INV_X1 U23772 ( .A(keyinput7), .ZN(n20847) );
  OAI22_X1 U23773 ( .A1(keyinput9), .A2(n20848), .B1(n20847), .B2(
        P3_UWORD_REG_11__SCAN_IN), .ZN(n20846) );
  AOI221_X1 U23774 ( .B1(n20848), .B2(keyinput9), .C1(n20847), .C2(
        P3_UWORD_REG_11__SCAN_IN), .A(n20846), .ZN(n20849) );
  NAND4_X1 U23775 ( .A1(n20852), .A2(n20851), .A3(n20850), .A4(n20849), .ZN(
        n20953) );
  INV_X1 U23776 ( .A(keyinput56), .ZN(n20855) );
  INV_X1 U23777 ( .A(keyinput38), .ZN(n20854) );
  AOI22_X1 U23778 ( .A1(n20855), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(
        P1_DATAWIDTH_REG_11__SCAN_IN), .B2(n20854), .ZN(n20853) );
  OAI221_X1 U23779 ( .B1(n20855), .B2(P1_UWORD_REG_11__SCAN_IN), .C1(n20854), 
        .C2(P1_DATAWIDTH_REG_11__SCAN_IN), .A(n20853), .ZN(n20886) );
  INV_X1 U23780 ( .A(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n20857) );
  AOI22_X1 U23781 ( .A1(n20858), .A2(keyinput6), .B1(n20857), .B2(keyinput14), 
        .ZN(n20856) );
  OAI221_X1 U23782 ( .B1(n20858), .B2(keyinput6), .C1(n20857), .C2(keyinput14), 
        .A(n20856), .ZN(n20885) );
  INV_X1 U23783 ( .A(keyinput32), .ZN(n20865) );
  AOI22_X1 U23784 ( .A1(n20860), .A2(keyinput2), .B1(n15666), .B2(keyinput51), 
        .ZN(n20859) );
  OAI221_X1 U23785 ( .B1(n20860), .B2(keyinput2), .C1(n15666), .C2(keyinput51), 
        .A(n20859), .ZN(n20861) );
  AOI221_X1 U23786 ( .B1(keyinput49), .B2(n20863), .C1(n20862), .C2(
        P3_EBX_REG_6__SCAN_IN), .A(n20861), .ZN(n20864) );
  OAI221_X1 U23787 ( .B1(keyinput32), .B2(n20866), .C1(n20865), .C2(
        P2_DATAO_REG_30__SCAN_IN), .A(n20864), .ZN(n20884) );
  OAI22_X1 U23788 ( .A1(n20869), .A2(keyinput29), .B1(n20868), .B2(keyinput54), 
        .ZN(n20867) );
  AOI221_X1 U23789 ( .B1(n20869), .B2(keyinput29), .C1(keyinput54), .C2(n20868), .A(n20867), .ZN(n20882) );
  INV_X1 U23790 ( .A(keyinput33), .ZN(n20871) );
  OAI22_X1 U23791 ( .A1(keyinput8), .A2(n20872), .B1(n20871), .B2(
        P1_ADS_N_REG_SCAN_IN), .ZN(n20870) );
  AOI221_X1 U23792 ( .B1(n20872), .B2(keyinput8), .C1(n20871), .C2(
        P1_ADS_N_REG_SCAN_IN), .A(n20870), .ZN(n20881) );
  OAI22_X1 U23793 ( .A1(n20875), .A2(keyinput63), .B1(n20874), .B2(keyinput39), 
        .ZN(n20873) );
  AOI221_X1 U23794 ( .B1(n20875), .B2(keyinput63), .C1(keyinput39), .C2(n20874), .A(n20873), .ZN(n20880) );
  INV_X1 U23795 ( .A(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n20878) );
  INV_X1 U23796 ( .A(keyinput34), .ZN(n20877) );
  OAI22_X1 U23797 ( .A1(n20878), .A2(keyinput44), .B1(n20877), .B2(
        P3_EAX_REG_20__SCAN_IN), .ZN(n20876) );
  AOI221_X1 U23798 ( .B1(n20878), .B2(keyinput44), .C1(P3_EAX_REG_20__SCAN_IN), 
        .C2(n20877), .A(n20876), .ZN(n20879) );
  NAND4_X1 U23799 ( .A1(n20882), .A2(n20881), .A3(n20880), .A4(n20879), .ZN(
        n20883) );
  NOR4_X1 U23800 ( .A1(n20886), .A2(n20885), .A3(n20884), .A4(n20883), .ZN(
        n20951) );
  INV_X1 U23801 ( .A(keyinput22), .ZN(n20888) );
  AOI22_X1 U23802 ( .A1(n20889), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n20888), .ZN(n20887) );
  OAI221_X1 U23803 ( .B1(n20889), .B2(P3_UWORD_REG_13__SCAN_IN), .C1(n20888), 
        .C2(P1_DATAO_REG_7__SCAN_IN), .A(n20887), .ZN(n20902) );
  AOI22_X1 U23804 ( .A1(n20892), .A2(keyinput36), .B1(keyinput62), .B2(n20891), 
        .ZN(n20890) );
  OAI221_X1 U23805 ( .B1(n20892), .B2(keyinput36), .C1(n20891), .C2(keyinput62), .A(n20890), .ZN(n20901) );
  AOI22_X1 U23806 ( .A1(n20895), .A2(keyinput43), .B1(P3_LWORD_REG_10__SCAN_IN), .B2(n20894), .ZN(n20893) );
  OAI221_X1 U23807 ( .B1(n20895), .B2(keyinput43), .C1(n20894), .C2(
        P3_LWORD_REG_10__SCAN_IN), .A(n20893), .ZN(n20900) );
  AOI22_X1 U23808 ( .A1(n20898), .A2(keyinput19), .B1(n20897), .B2(keyinput20), 
        .ZN(n20896) );
  OAI221_X1 U23809 ( .B1(n20898), .B2(keyinput19), .C1(n20897), .C2(keyinput20), .A(n20896), .ZN(n20899) );
  NOR4_X1 U23810 ( .A1(n20902), .A2(n20901), .A3(n20900), .A4(n20899), .ZN(
        n20950) );
  INV_X1 U23811 ( .A(keyinput23), .ZN(n20905) );
  INV_X1 U23812 ( .A(keyinput5), .ZN(n20904) );
  AOI22_X1 U23813 ( .A1(n20905), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(
        P3_ADDRESS_REG_20__SCAN_IN), .B2(n20904), .ZN(n20903) );
  OAI221_X1 U23814 ( .B1(n20905), .B2(P3_READREQUEST_REG_SCAN_IN), .C1(n20904), 
        .C2(P3_ADDRESS_REG_20__SCAN_IN), .A(n20903), .ZN(n20916) );
  INV_X1 U23815 ( .A(keyinput59), .ZN(n20907) );
  AOI22_X1 U23816 ( .A1(n10143), .A2(keyinput47), .B1(P3_FLUSH_REG_SCAN_IN), 
        .B2(n20907), .ZN(n20906) );
  OAI221_X1 U23817 ( .B1(n10143), .B2(keyinput47), .C1(n20907), .C2(
        P3_FLUSH_REG_SCAN_IN), .A(n20906), .ZN(n20915) );
  AOI22_X1 U23818 ( .A1(n20910), .A2(keyinput25), .B1(keyinput45), .B2(n20909), 
        .ZN(n20908) );
  OAI221_X1 U23819 ( .B1(n20910), .B2(keyinput25), .C1(n20909), .C2(keyinput45), .A(n20908), .ZN(n20914) );
  INV_X1 U23820 ( .A(keyinput31), .ZN(n20912) );
  AOI22_X1 U23821 ( .A1(n12824), .A2(keyinput42), .B1(P2_DATAO_REG_25__SCAN_IN), .B2(n20912), .ZN(n20911) );
  OAI221_X1 U23822 ( .B1(n12824), .B2(keyinput42), .C1(n20912), .C2(
        P2_DATAO_REG_25__SCAN_IN), .A(n20911), .ZN(n20913) );
  NOR4_X1 U23823 ( .A1(n20916), .A2(n20915), .A3(n20914), .A4(n20913), .ZN(
        n20949) );
  INV_X1 U23824 ( .A(keyinput50), .ZN(n20918) );
  AOI22_X1 U23825 ( .A1(n11737), .A2(keyinput13), .B1(P1_DATAO_REG_29__SCAN_IN), .B2(n20918), .ZN(n20917) );
  OAI221_X1 U23826 ( .B1(n11737), .B2(keyinput13), .C1(n20918), .C2(
        P1_DATAO_REG_29__SCAN_IN), .A(n20917), .ZN(n20947) );
  AOI22_X1 U23827 ( .A1(n20921), .A2(keyinput53), .B1(keyinput27), .B2(n20920), 
        .ZN(n20919) );
  OAI221_X1 U23828 ( .B1(n20921), .B2(keyinput53), .C1(n20920), .C2(keyinput27), .A(n20919), .ZN(n20946) );
  OAI22_X1 U23829 ( .A1(n20924), .A2(keyinput4), .B1(n20923), .B2(keyinput35), 
        .ZN(n20922) );
  AOI221_X1 U23830 ( .B1(n20924), .B2(keyinput4), .C1(keyinput35), .C2(n20923), 
        .A(n20922), .ZN(n20927) );
  XOR2_X1 U23831 ( .A(keyinput16), .B(n20925), .Z(n20926) );
  OAI211_X1 U23832 ( .C1(keyinput55), .C2(n20928), .A(n20927), .B(n20926), 
        .ZN(n20945) );
  INV_X1 U23833 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20931) );
  INV_X1 U23834 ( .A(keyinput12), .ZN(n20930) );
  OAI22_X1 U23835 ( .A1(n20931), .A2(keyinput28), .B1(n20930), .B2(DATAI_15_), 
        .ZN(n20929) );
  AOI221_X1 U23836 ( .B1(n20931), .B2(keyinput28), .C1(DATAI_15_), .C2(n20930), 
        .A(n20929), .ZN(n20943) );
  INV_X1 U23837 ( .A(keyinput52), .ZN(n20933) );
  OAI22_X1 U23838 ( .A1(keyinput15), .A2(n20934), .B1(n20933), .B2(
        P3_ADDRESS_REG_29__SCAN_IN), .ZN(n20932) );
  AOI221_X1 U23839 ( .B1(n20934), .B2(keyinput15), .C1(n20933), .C2(
        P3_ADDRESS_REG_29__SCAN_IN), .A(n20932), .ZN(n20942) );
  OAI22_X1 U23840 ( .A1(n20937), .A2(keyinput3), .B1(n20936), .B2(keyinput40), 
        .ZN(n20935) );
  AOI221_X1 U23841 ( .B1(n20937), .B2(keyinput3), .C1(keyinput40), .C2(n20936), 
        .A(n20935), .ZN(n20941) );
  INV_X1 U23842 ( .A(keyinput30), .ZN(n20939) );
  OAI22_X1 U23843 ( .A1(n10632), .A2(keyinput41), .B1(n20939), .B2(
        P3_EAX_REG_26__SCAN_IN), .ZN(n20938) );
  AOI221_X1 U23844 ( .B1(n10632), .B2(keyinput41), .C1(P3_EAX_REG_26__SCAN_IN), 
        .C2(n20939), .A(n20938), .ZN(n20940) );
  NAND4_X1 U23845 ( .A1(n20943), .A2(n20942), .A3(n20941), .A4(n20940), .ZN(
        n20944) );
  NOR4_X1 U23846 ( .A1(n20947), .A2(n20946), .A3(n20945), .A4(n20944), .ZN(
        n20948) );
  NAND4_X1 U23847 ( .A1(n20951), .A2(n20950), .A3(n20949), .A4(n20948), .ZN(
        n20952) );
  NOR4_X1 U23848 ( .A1(n20955), .A2(n20954), .A3(n20953), .A4(n20952), .ZN(
        n20966) );
  AND2_X1 U23849 ( .A1(n20957), .A2(n20956), .ZN(n20963) );
  INV_X1 U23850 ( .A(n20958), .ZN(n20960) );
  INV_X1 U23851 ( .A(n14077), .ZN(n20959) );
  AOI211_X1 U23852 ( .C1(n20961), .C2(n20960), .A(n18919), .B(n20959), .ZN(
        n20962) );
  AOI211_X1 U23853 ( .C1(P2_EBX_REG_13__SCAN_IN), .C2(n20964), .A(n20963), .B(
        n20962), .ZN(n20965) );
  XNOR2_X1 U23854 ( .A(n20966), .B(n20965), .ZN(P2_U2874) );
  XNOR2_X1 U11009 ( .A(n12785), .B(n20009), .ZN(n19985) );
  CLKBUF_X1 U11024 ( .A(n12113), .Z(n13588) );
  CLKBUF_X1 U11068 ( .A(n11120), .Z(n19129) );
  CLKBUF_X1 U11070 ( .A(n10814), .Z(n16756) );
  CLKBUF_X1 U11073 ( .A(n15414), .Z(n9577) );
  XOR2_X1 U11085 ( .A(n17189), .B(n10781), .Z(n10769) );
  CLKBUF_X1 U11106 ( .A(n13595), .Z(n9569) );
  CLKBUF_X1 U11108 ( .A(n13600), .Z(n20059) );
  CLKBUF_X3 U11110 ( .A(n13685), .Z(n9567) );
  OR3_X2 U11115 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n10699), .ZN(n10740) );
  NOR2_X2 U11128 ( .A1(n14059), .A2(n18515), .ZN(n18513) );
  CLKBUF_X1 U11137 ( .A(n12867), .Z(n14520) );
  CLKBUF_X1 U11139 ( .A(n9593), .Z(n15388) );
  CLKBUF_X1 U11145 ( .A(n10745), .Z(n17014) );
  CLKBUF_X1 U11159 ( .A(n17294), .Z(n17319) );
  NAND2_X2 U11924 ( .A1(n17907), .A2(n18514), .ZN(n17926) );
  CLKBUF_X1 U11999 ( .A(n17696), .Z(n9594) );
  INV_X2 U12098 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10687) );
endmodule

